magic
tech sky130A
timestamp 1616095553
<< nwell >>
rect 3450 8500 4058 8650
rect 7814 8513 8422 8663
rect 12191 8525 12799 8675
rect 16555 8538 17163 8688
rect 401 8346 1009 8496
rect 1199 8162 1807 8312
rect 2653 8272 3261 8422
rect 4765 8359 5373 8509
rect 3451 8088 4059 8238
rect 5563 8175 6171 8325
rect 7017 8285 7625 8435
rect 9142 8371 9750 8521
rect 7815 8101 8423 8251
rect 9940 8187 10548 8337
rect 11394 8297 12002 8447
rect 13506 8384 14114 8534
rect 12192 8113 12800 8263
rect 14304 8200 14912 8350
rect 15758 8310 16366 8460
rect 16556 8126 17164 8276
rect 402 7934 1010 8084
rect 2554 7862 3162 8012
rect 4766 7947 5374 8097
rect 6918 7875 7526 8025
rect 9143 7959 9751 8109
rect 11295 7887 11903 8037
rect 13507 7972 14115 8122
rect 15659 7900 16267 8050
rect 1281 7554 1889 7704
rect 3433 7482 4041 7632
rect 5645 7567 6253 7717
rect 7797 7495 8405 7645
rect 10022 7579 10630 7729
rect 12174 7507 12782 7657
rect 14386 7592 14994 7742
rect 16538 7520 17146 7670
rect 384 7328 992 7478
rect 1182 7144 1790 7294
rect 2636 7254 3244 7404
rect 4748 7341 5356 7491
rect 3434 7070 4042 7220
rect 5546 7157 6154 7307
rect 7000 7267 7608 7417
rect 9125 7353 9733 7503
rect 7798 7083 8406 7233
rect 9923 7169 10531 7319
rect 11377 7279 11985 7429
rect 13489 7366 14097 7516
rect 12175 7095 12783 7245
rect 14287 7182 14895 7332
rect 15741 7292 16349 7442
rect 16539 7108 17147 7258
rect 385 6916 993 7066
rect 2471 6846 3079 6996
rect 4749 6929 5357 7079
rect 6835 6859 7443 7009
rect 9126 6941 9734 7091
rect 11212 6871 11820 7021
rect 13490 6954 14098 7104
rect 15576 6884 16184 7034
rect 1327 6534 1935 6684
rect 3413 6464 4021 6614
rect 5691 6547 6299 6697
rect 7777 6477 8385 6627
rect 10068 6559 10676 6709
rect 12154 6489 12762 6639
rect 14432 6572 15040 6722
rect 16518 6502 17126 6652
rect 364 6310 972 6460
rect 1162 6126 1770 6276
rect 2616 6236 3224 6386
rect 4728 6323 5336 6473
rect 3414 6052 4022 6202
rect 5526 6139 6134 6289
rect 6980 6249 7588 6399
rect 9105 6335 9713 6485
rect 7778 6065 8386 6215
rect 9903 6151 10511 6301
rect 11357 6261 11965 6411
rect 13469 6348 14077 6498
rect 12155 6077 12763 6227
rect 14267 6164 14875 6314
rect 15721 6274 16329 6424
rect 16519 6090 17127 6240
rect 365 5898 973 6048
rect 2517 5826 3125 5976
rect 4729 5911 5337 6061
rect 6881 5839 7489 5989
rect 9106 5923 9714 6073
rect 11258 5851 11866 6001
rect 13470 5936 14078 6086
rect 15622 5864 16230 6014
rect 1244 5518 1852 5668
rect 3396 5446 4004 5596
rect 5608 5531 6216 5681
rect 7760 5459 8368 5609
rect 9985 5543 10593 5693
rect 12137 5471 12745 5621
rect 14349 5556 14957 5706
rect 16501 5484 17109 5634
rect 347 5292 955 5442
rect 1145 5108 1753 5258
rect 2599 5218 3207 5368
rect 4711 5305 5319 5455
rect 3397 5034 4005 5184
rect 5509 5121 6117 5271
rect 6963 5231 7571 5381
rect 9088 5317 9696 5467
rect 7761 5047 8369 5197
rect 9886 5133 10494 5283
rect 11340 5243 11948 5393
rect 13452 5330 14060 5480
rect 12138 5059 12746 5209
rect 14250 5146 14858 5296
rect 15704 5256 16312 5406
rect 16502 5072 17110 5222
rect 348 4880 956 5030
rect 2295 4812 2903 4962
rect 4712 4893 5320 5043
rect 6659 4825 7267 4975
rect 9089 4905 9697 5055
rect 11036 4837 11644 4987
rect 13453 4918 14061 5068
rect 15400 4850 16008 5000
rect 1430 4496 2038 4646
rect 3377 4428 3985 4578
rect 5794 4509 6402 4659
rect 7741 4441 8349 4591
rect 10171 4521 10779 4671
rect 12118 4453 12726 4603
rect 14535 4534 15143 4684
rect 16482 4466 17090 4616
rect 328 4274 936 4424
rect 1126 4090 1734 4240
rect 2580 4200 3188 4350
rect 4692 4287 5300 4437
rect 3378 4016 3986 4166
rect 5490 4103 6098 4253
rect 6944 4213 7552 4363
rect 9069 4299 9677 4449
rect 7742 4029 8350 4179
rect 9867 4115 10475 4265
rect 11321 4225 11929 4375
rect 13433 4312 14041 4462
rect 12119 4041 12727 4191
rect 14231 4128 14839 4278
rect 15685 4238 16293 4388
rect 16483 4054 17091 4204
rect 329 3862 937 4012
rect 2481 3790 3089 3940
rect 4693 3875 5301 4025
rect 6845 3803 7453 3953
rect 9070 3887 9678 4037
rect 11222 3815 11830 3965
rect 13434 3900 14042 4050
rect 15586 3828 16194 3978
rect 1208 3482 1816 3632
rect 3360 3410 3968 3560
rect 5572 3495 6180 3645
rect 7724 3423 8332 3573
rect 9949 3507 10557 3657
rect 12101 3435 12709 3585
rect 14313 3520 14921 3670
rect 16465 3448 17073 3598
rect 311 3256 919 3406
rect 1109 3072 1717 3222
rect 2563 3182 3171 3332
rect 4675 3269 5283 3419
rect 3361 2998 3969 3148
rect 5473 3085 6081 3235
rect 6927 3195 7535 3345
rect 9052 3281 9660 3431
rect 7725 3011 8333 3161
rect 9850 3097 10458 3247
rect 11304 3207 11912 3357
rect 13416 3294 14024 3444
rect 12102 3023 12710 3173
rect 14214 3110 14822 3260
rect 15668 3220 16276 3370
rect 16466 3036 17074 3186
rect 312 2844 920 2994
rect 2398 2774 3006 2924
rect 4676 2857 5284 3007
rect 6762 2787 7370 2937
rect 9053 2869 9661 3019
rect 11139 2799 11747 2949
rect 13417 2882 14025 3032
rect 15503 2812 16111 2962
rect 1254 2462 1862 2612
rect 3340 2392 3948 2542
rect 5618 2475 6226 2625
rect 7704 2405 8312 2555
rect 9995 2487 10603 2637
rect 12081 2417 12689 2567
rect 14359 2500 14967 2650
rect 16445 2430 17053 2580
rect 291 2238 899 2388
rect 1089 2054 1697 2204
rect 2543 2164 3151 2314
rect 4655 2251 5263 2401
rect 3341 1980 3949 2130
rect 5453 2067 6061 2217
rect 6907 2177 7515 2327
rect 9032 2263 9640 2413
rect 7705 1993 8313 2143
rect 9830 2079 10438 2229
rect 11284 2189 11892 2339
rect 13396 2276 14004 2426
rect 12082 2005 12690 2155
rect 14194 2092 14802 2242
rect 15648 2202 16256 2352
rect 16446 2018 17054 2168
rect 292 1826 900 1976
rect 2444 1754 3052 1904
rect 4656 1839 5264 1989
rect 6808 1767 7416 1917
rect 9033 1851 9641 2001
rect 11185 1779 11793 1929
rect 13397 1864 14005 2014
rect 15549 1792 16157 1942
rect 1171 1446 1779 1596
rect 3323 1374 3931 1524
rect 5535 1459 6143 1609
rect 7687 1387 8295 1537
rect 9912 1471 10520 1621
rect 12064 1399 12672 1549
rect 14276 1484 14884 1634
rect 16428 1412 17036 1562
rect 274 1220 882 1370
rect 1072 1036 1680 1186
rect 2526 1146 3134 1296
rect 4638 1233 5246 1383
rect 3324 962 3932 1112
rect 5436 1049 6044 1199
rect 6890 1159 7498 1309
rect 9015 1245 9623 1395
rect 7688 975 8296 1125
rect 9813 1061 10421 1211
rect 11267 1171 11875 1321
rect 13379 1258 13987 1408
rect 12065 987 12673 1137
rect 14177 1074 14785 1224
rect 15631 1184 16239 1334
rect 16429 1000 17037 1150
rect 275 808 883 958
rect 4639 821 5247 971
rect 9016 833 9624 983
rect 13380 846 13988 996
rect 1488 232 2096 382
rect 3977 158 4585 308
rect 5852 245 6460 395
rect 8425 182 9033 332
rect 10229 257 10837 407
rect 12718 183 13326 333
rect 14593 270 15201 420
<< nmos >>
rect 3518 8709 3568 8751
rect 3726 8709 3776 8751
rect 3944 8709 3994 8751
rect 7882 8722 7932 8764
rect 8090 8722 8140 8764
rect 8308 8722 8358 8764
rect 12259 8734 12309 8776
rect 12467 8734 12517 8776
rect 12685 8734 12735 8776
rect 2721 8481 2771 8523
rect 2929 8481 2979 8523
rect 3147 8481 3197 8523
rect 16623 8747 16673 8789
rect 16831 8747 16881 8789
rect 17049 8747 17099 8789
rect 7085 8494 7135 8536
rect 7293 8494 7343 8536
rect 7511 8494 7561 8536
rect 11462 8506 11512 8548
rect 11670 8506 11720 8548
rect 11888 8506 11938 8548
rect 15826 8519 15876 8561
rect 16034 8519 16084 8561
rect 16252 8519 16302 8561
rect 465 8245 515 8287
rect 683 8245 733 8287
rect 891 8245 941 8287
rect 3519 8297 3569 8339
rect 3727 8297 3777 8339
rect 3945 8297 3995 8339
rect 4829 8258 4879 8300
rect 5047 8258 5097 8300
rect 5255 8258 5305 8300
rect 7883 8310 7933 8352
rect 8091 8310 8141 8352
rect 8309 8310 8359 8352
rect 9206 8270 9256 8312
rect 9424 8270 9474 8312
rect 9632 8270 9682 8312
rect 12260 8322 12310 8364
rect 12468 8322 12518 8364
rect 12686 8322 12736 8364
rect 1263 8061 1313 8103
rect 1481 8061 1531 8103
rect 1689 8061 1739 8103
rect 2622 8071 2672 8113
rect 2830 8071 2880 8113
rect 3048 8071 3098 8113
rect 13570 8283 13620 8325
rect 13788 8283 13838 8325
rect 13996 8283 14046 8325
rect 16624 8335 16674 8377
rect 16832 8335 16882 8377
rect 17050 8335 17100 8377
rect 5627 8074 5677 8116
rect 5845 8074 5895 8116
rect 6053 8074 6103 8116
rect 6986 8084 7036 8126
rect 7194 8084 7244 8126
rect 7412 8084 7462 8126
rect 10004 8086 10054 8128
rect 10222 8086 10272 8128
rect 10430 8086 10480 8128
rect 11363 8096 11413 8138
rect 11571 8096 11621 8138
rect 11789 8096 11839 8138
rect 466 7833 516 7875
rect 684 7833 734 7875
rect 892 7833 942 7875
rect 14368 8099 14418 8141
rect 14586 8099 14636 8141
rect 14794 8099 14844 8141
rect 15727 8109 15777 8151
rect 15935 8109 15985 8151
rect 16153 8109 16203 8151
rect 4830 7846 4880 7888
rect 5048 7846 5098 7888
rect 5256 7846 5306 7888
rect 9207 7858 9257 7900
rect 9425 7858 9475 7900
rect 9633 7858 9683 7900
rect 13571 7871 13621 7913
rect 13789 7871 13839 7913
rect 13997 7871 14047 7913
rect 3501 7691 3551 7733
rect 3709 7691 3759 7733
rect 3927 7691 3977 7733
rect 7865 7704 7915 7746
rect 8073 7704 8123 7746
rect 8291 7704 8341 7746
rect 12242 7716 12292 7758
rect 12450 7716 12500 7758
rect 12668 7716 12718 7758
rect 1345 7453 1395 7495
rect 1563 7453 1613 7495
rect 1771 7453 1821 7495
rect 2704 7463 2754 7505
rect 2912 7463 2962 7505
rect 3130 7463 3180 7505
rect 16606 7729 16656 7771
rect 16814 7729 16864 7771
rect 17032 7729 17082 7771
rect 5709 7466 5759 7508
rect 5927 7466 5977 7508
rect 6135 7466 6185 7508
rect 7068 7476 7118 7518
rect 7276 7476 7326 7518
rect 7494 7476 7544 7518
rect 10086 7478 10136 7520
rect 10304 7478 10354 7520
rect 10512 7478 10562 7520
rect 11445 7488 11495 7530
rect 11653 7488 11703 7530
rect 11871 7488 11921 7530
rect 448 7227 498 7269
rect 666 7227 716 7269
rect 874 7227 924 7269
rect 3502 7279 3552 7321
rect 3710 7279 3760 7321
rect 3928 7279 3978 7321
rect 14450 7491 14500 7533
rect 14668 7491 14718 7533
rect 14876 7491 14926 7533
rect 15809 7501 15859 7543
rect 16017 7501 16067 7543
rect 16235 7501 16285 7543
rect 4812 7240 4862 7282
rect 5030 7240 5080 7282
rect 5238 7240 5288 7282
rect 7866 7292 7916 7334
rect 8074 7292 8124 7334
rect 8292 7292 8342 7334
rect 9189 7252 9239 7294
rect 9407 7252 9457 7294
rect 9615 7252 9665 7294
rect 12243 7304 12293 7346
rect 12451 7304 12501 7346
rect 12669 7304 12719 7346
rect 1246 7043 1296 7085
rect 1464 7043 1514 7085
rect 1672 7043 1722 7085
rect 2539 7055 2589 7097
rect 2747 7055 2797 7097
rect 2965 7055 3015 7097
rect 13553 7265 13603 7307
rect 13771 7265 13821 7307
rect 13979 7265 14029 7307
rect 16607 7317 16657 7359
rect 16815 7317 16865 7359
rect 17033 7317 17083 7359
rect 5610 7056 5660 7098
rect 5828 7056 5878 7098
rect 6036 7056 6086 7098
rect 6903 7068 6953 7110
rect 7111 7068 7161 7110
rect 7329 7068 7379 7110
rect 9987 7068 10037 7110
rect 10205 7068 10255 7110
rect 10413 7068 10463 7110
rect 11280 7080 11330 7122
rect 11488 7080 11538 7122
rect 11706 7080 11756 7122
rect 449 6815 499 6857
rect 667 6815 717 6857
rect 875 6815 925 6857
rect 14351 7081 14401 7123
rect 14569 7081 14619 7123
rect 14777 7081 14827 7123
rect 15644 7093 15694 7135
rect 15852 7093 15902 7135
rect 16070 7093 16120 7135
rect 4813 6828 4863 6870
rect 5031 6828 5081 6870
rect 5239 6828 5289 6870
rect 9190 6840 9240 6882
rect 9408 6840 9458 6882
rect 9616 6840 9666 6882
rect 13554 6853 13604 6895
rect 13772 6853 13822 6895
rect 13980 6853 14030 6895
rect 3481 6673 3531 6715
rect 3689 6673 3739 6715
rect 3907 6673 3957 6715
rect 7845 6686 7895 6728
rect 8053 6686 8103 6728
rect 8271 6686 8321 6728
rect 12222 6698 12272 6740
rect 12430 6698 12480 6740
rect 12648 6698 12698 6740
rect 1391 6433 1441 6475
rect 1609 6433 1659 6475
rect 1817 6433 1867 6475
rect 2684 6445 2734 6487
rect 2892 6445 2942 6487
rect 3110 6445 3160 6487
rect 16586 6711 16636 6753
rect 16794 6711 16844 6753
rect 17012 6711 17062 6753
rect 5755 6446 5805 6488
rect 5973 6446 6023 6488
rect 6181 6446 6231 6488
rect 7048 6458 7098 6500
rect 7256 6458 7306 6500
rect 7474 6458 7524 6500
rect 10132 6458 10182 6500
rect 10350 6458 10400 6500
rect 10558 6458 10608 6500
rect 11425 6470 11475 6512
rect 11633 6470 11683 6512
rect 11851 6470 11901 6512
rect 428 6209 478 6251
rect 646 6209 696 6251
rect 854 6209 904 6251
rect 3482 6261 3532 6303
rect 3690 6261 3740 6303
rect 3908 6261 3958 6303
rect 14496 6471 14546 6513
rect 14714 6471 14764 6513
rect 14922 6471 14972 6513
rect 15789 6483 15839 6525
rect 15997 6483 16047 6525
rect 16215 6483 16265 6525
rect 4792 6222 4842 6264
rect 5010 6222 5060 6264
rect 5218 6222 5268 6264
rect 7846 6274 7896 6316
rect 8054 6274 8104 6316
rect 8272 6274 8322 6316
rect 9169 6234 9219 6276
rect 9387 6234 9437 6276
rect 9595 6234 9645 6276
rect 12223 6286 12273 6328
rect 12431 6286 12481 6328
rect 12649 6286 12699 6328
rect 1226 6025 1276 6067
rect 1444 6025 1494 6067
rect 1652 6025 1702 6067
rect 2585 6035 2635 6077
rect 2793 6035 2843 6077
rect 3011 6035 3061 6077
rect 13533 6247 13583 6289
rect 13751 6247 13801 6289
rect 13959 6247 14009 6289
rect 16587 6299 16637 6341
rect 16795 6299 16845 6341
rect 17013 6299 17063 6341
rect 5590 6038 5640 6080
rect 5808 6038 5858 6080
rect 6016 6038 6066 6080
rect 6949 6048 6999 6090
rect 7157 6048 7207 6090
rect 7375 6048 7425 6090
rect 9967 6050 10017 6092
rect 10185 6050 10235 6092
rect 10393 6050 10443 6092
rect 11326 6060 11376 6102
rect 11534 6060 11584 6102
rect 11752 6060 11802 6102
rect 429 5797 479 5839
rect 647 5797 697 5839
rect 855 5797 905 5839
rect 14331 6063 14381 6105
rect 14549 6063 14599 6105
rect 14757 6063 14807 6105
rect 15690 6073 15740 6115
rect 15898 6073 15948 6115
rect 16116 6073 16166 6115
rect 4793 5810 4843 5852
rect 5011 5810 5061 5852
rect 5219 5810 5269 5852
rect 9170 5822 9220 5864
rect 9388 5822 9438 5864
rect 9596 5822 9646 5864
rect 13534 5835 13584 5877
rect 13752 5835 13802 5877
rect 13960 5835 14010 5877
rect 3464 5655 3514 5697
rect 3672 5655 3722 5697
rect 3890 5655 3940 5697
rect 7828 5668 7878 5710
rect 8036 5668 8086 5710
rect 8254 5668 8304 5710
rect 12205 5680 12255 5722
rect 12413 5680 12463 5722
rect 12631 5680 12681 5722
rect 1308 5417 1358 5459
rect 1526 5417 1576 5459
rect 1734 5417 1784 5459
rect 2667 5427 2717 5469
rect 2875 5427 2925 5469
rect 3093 5427 3143 5469
rect 16569 5693 16619 5735
rect 16777 5693 16827 5735
rect 16995 5693 17045 5735
rect 5672 5430 5722 5472
rect 5890 5430 5940 5472
rect 6098 5430 6148 5472
rect 7031 5440 7081 5482
rect 7239 5440 7289 5482
rect 7457 5440 7507 5482
rect 10049 5442 10099 5484
rect 10267 5442 10317 5484
rect 10475 5442 10525 5484
rect 11408 5452 11458 5494
rect 11616 5452 11666 5494
rect 11834 5452 11884 5494
rect 411 5191 461 5233
rect 629 5191 679 5233
rect 837 5191 887 5233
rect 3465 5243 3515 5285
rect 3673 5243 3723 5285
rect 3891 5243 3941 5285
rect 14413 5455 14463 5497
rect 14631 5455 14681 5497
rect 14839 5455 14889 5497
rect 15772 5465 15822 5507
rect 15980 5465 16030 5507
rect 16198 5465 16248 5507
rect 4775 5204 4825 5246
rect 4993 5204 5043 5246
rect 5201 5204 5251 5246
rect 7829 5256 7879 5298
rect 8037 5256 8087 5298
rect 8255 5256 8305 5298
rect 9152 5216 9202 5258
rect 9370 5216 9420 5258
rect 9578 5216 9628 5258
rect 12206 5268 12256 5310
rect 12414 5268 12464 5310
rect 12632 5268 12682 5310
rect 1209 5007 1259 5049
rect 1427 5007 1477 5049
rect 1635 5007 1685 5049
rect 2363 5021 2413 5063
rect 2571 5021 2621 5063
rect 2789 5021 2839 5063
rect 13516 5229 13566 5271
rect 13734 5229 13784 5271
rect 13942 5229 13992 5271
rect 16570 5281 16620 5323
rect 16778 5281 16828 5323
rect 16996 5281 17046 5323
rect 5573 5020 5623 5062
rect 5791 5020 5841 5062
rect 5999 5020 6049 5062
rect 6727 5034 6777 5076
rect 6935 5034 6985 5076
rect 7153 5034 7203 5076
rect 9950 5032 10000 5074
rect 10168 5032 10218 5074
rect 10376 5032 10426 5074
rect 11104 5046 11154 5088
rect 11312 5046 11362 5088
rect 11530 5046 11580 5088
rect 412 4779 462 4821
rect 630 4779 680 4821
rect 838 4779 888 4821
rect 14314 5045 14364 5087
rect 14532 5045 14582 5087
rect 14740 5045 14790 5087
rect 15468 5059 15518 5101
rect 15676 5059 15726 5101
rect 15894 5059 15944 5101
rect 4776 4792 4826 4834
rect 4994 4792 5044 4834
rect 5202 4792 5252 4834
rect 9153 4804 9203 4846
rect 9371 4804 9421 4846
rect 9579 4804 9629 4846
rect 13517 4817 13567 4859
rect 13735 4817 13785 4859
rect 13943 4817 13993 4859
rect 3445 4637 3495 4679
rect 3653 4637 3703 4679
rect 3871 4637 3921 4679
rect 7809 4650 7859 4692
rect 8017 4650 8067 4692
rect 8235 4650 8285 4692
rect 12186 4662 12236 4704
rect 12394 4662 12444 4704
rect 12612 4662 12662 4704
rect 1494 4395 1544 4437
rect 1712 4395 1762 4437
rect 1920 4395 1970 4437
rect 2648 4409 2698 4451
rect 2856 4409 2906 4451
rect 3074 4409 3124 4451
rect 16550 4675 16600 4717
rect 16758 4675 16808 4717
rect 16976 4675 17026 4717
rect 5858 4408 5908 4450
rect 6076 4408 6126 4450
rect 6284 4408 6334 4450
rect 7012 4422 7062 4464
rect 7220 4422 7270 4464
rect 7438 4422 7488 4464
rect 10235 4420 10285 4462
rect 10453 4420 10503 4462
rect 10661 4420 10711 4462
rect 11389 4434 11439 4476
rect 11597 4434 11647 4476
rect 11815 4434 11865 4476
rect 392 4173 442 4215
rect 610 4173 660 4215
rect 818 4173 868 4215
rect 3446 4225 3496 4267
rect 3654 4225 3704 4267
rect 3872 4225 3922 4267
rect 14599 4433 14649 4475
rect 14817 4433 14867 4475
rect 15025 4433 15075 4475
rect 15753 4447 15803 4489
rect 15961 4447 16011 4489
rect 16179 4447 16229 4489
rect 4756 4186 4806 4228
rect 4974 4186 5024 4228
rect 5182 4186 5232 4228
rect 7810 4238 7860 4280
rect 8018 4238 8068 4280
rect 8236 4238 8286 4280
rect 9133 4198 9183 4240
rect 9351 4198 9401 4240
rect 9559 4198 9609 4240
rect 12187 4250 12237 4292
rect 12395 4250 12445 4292
rect 12613 4250 12663 4292
rect 1190 3989 1240 4031
rect 1408 3989 1458 4031
rect 1616 3989 1666 4031
rect 2549 3999 2599 4041
rect 2757 3999 2807 4041
rect 2975 3999 3025 4041
rect 13497 4211 13547 4253
rect 13715 4211 13765 4253
rect 13923 4211 13973 4253
rect 16551 4263 16601 4305
rect 16759 4263 16809 4305
rect 16977 4263 17027 4305
rect 5554 4002 5604 4044
rect 5772 4002 5822 4044
rect 5980 4002 6030 4044
rect 6913 4012 6963 4054
rect 7121 4012 7171 4054
rect 7339 4012 7389 4054
rect 9931 4014 9981 4056
rect 10149 4014 10199 4056
rect 10357 4014 10407 4056
rect 11290 4024 11340 4066
rect 11498 4024 11548 4066
rect 11716 4024 11766 4066
rect 393 3761 443 3803
rect 611 3761 661 3803
rect 819 3761 869 3803
rect 14295 4027 14345 4069
rect 14513 4027 14563 4069
rect 14721 4027 14771 4069
rect 15654 4037 15704 4079
rect 15862 4037 15912 4079
rect 16080 4037 16130 4079
rect 4757 3774 4807 3816
rect 4975 3774 5025 3816
rect 5183 3774 5233 3816
rect 9134 3786 9184 3828
rect 9352 3786 9402 3828
rect 9560 3786 9610 3828
rect 13498 3799 13548 3841
rect 13716 3799 13766 3841
rect 13924 3799 13974 3841
rect 3428 3619 3478 3661
rect 3636 3619 3686 3661
rect 3854 3619 3904 3661
rect 7792 3632 7842 3674
rect 8000 3632 8050 3674
rect 8218 3632 8268 3674
rect 12169 3644 12219 3686
rect 12377 3644 12427 3686
rect 12595 3644 12645 3686
rect 1272 3381 1322 3423
rect 1490 3381 1540 3423
rect 1698 3381 1748 3423
rect 2631 3391 2681 3433
rect 2839 3391 2889 3433
rect 3057 3391 3107 3433
rect 16533 3657 16583 3699
rect 16741 3657 16791 3699
rect 16959 3657 17009 3699
rect 5636 3394 5686 3436
rect 5854 3394 5904 3436
rect 6062 3394 6112 3436
rect 6995 3404 7045 3446
rect 7203 3404 7253 3446
rect 7421 3404 7471 3446
rect 10013 3406 10063 3448
rect 10231 3406 10281 3448
rect 10439 3406 10489 3448
rect 11372 3416 11422 3458
rect 11580 3416 11630 3458
rect 11798 3416 11848 3458
rect 375 3155 425 3197
rect 593 3155 643 3197
rect 801 3155 851 3197
rect 3429 3207 3479 3249
rect 3637 3207 3687 3249
rect 3855 3207 3905 3249
rect 14377 3419 14427 3461
rect 14595 3419 14645 3461
rect 14803 3419 14853 3461
rect 15736 3429 15786 3471
rect 15944 3429 15994 3471
rect 16162 3429 16212 3471
rect 4739 3168 4789 3210
rect 4957 3168 5007 3210
rect 5165 3168 5215 3210
rect 7793 3220 7843 3262
rect 8001 3220 8051 3262
rect 8219 3220 8269 3262
rect 9116 3180 9166 3222
rect 9334 3180 9384 3222
rect 9542 3180 9592 3222
rect 12170 3232 12220 3274
rect 12378 3232 12428 3274
rect 12596 3232 12646 3274
rect 1173 2971 1223 3013
rect 1391 2971 1441 3013
rect 1599 2971 1649 3013
rect 2466 2983 2516 3025
rect 2674 2983 2724 3025
rect 2892 2983 2942 3025
rect 13480 3193 13530 3235
rect 13698 3193 13748 3235
rect 13906 3193 13956 3235
rect 16534 3245 16584 3287
rect 16742 3245 16792 3287
rect 16960 3245 17010 3287
rect 5537 2984 5587 3026
rect 5755 2984 5805 3026
rect 5963 2984 6013 3026
rect 6830 2996 6880 3038
rect 7038 2996 7088 3038
rect 7256 2996 7306 3038
rect 9914 2996 9964 3038
rect 10132 2996 10182 3038
rect 10340 2996 10390 3038
rect 11207 3008 11257 3050
rect 11415 3008 11465 3050
rect 11633 3008 11683 3050
rect 376 2743 426 2785
rect 594 2743 644 2785
rect 802 2743 852 2785
rect 14278 3009 14328 3051
rect 14496 3009 14546 3051
rect 14704 3009 14754 3051
rect 15571 3021 15621 3063
rect 15779 3021 15829 3063
rect 15997 3021 16047 3063
rect 4740 2756 4790 2798
rect 4958 2756 5008 2798
rect 5166 2756 5216 2798
rect 9117 2768 9167 2810
rect 9335 2768 9385 2810
rect 9543 2768 9593 2810
rect 13481 2781 13531 2823
rect 13699 2781 13749 2823
rect 13907 2781 13957 2823
rect 3408 2601 3458 2643
rect 3616 2601 3666 2643
rect 3834 2601 3884 2643
rect 7772 2614 7822 2656
rect 7980 2614 8030 2656
rect 8198 2614 8248 2656
rect 12149 2626 12199 2668
rect 12357 2626 12407 2668
rect 12575 2626 12625 2668
rect 1318 2361 1368 2403
rect 1536 2361 1586 2403
rect 1744 2361 1794 2403
rect 2611 2373 2661 2415
rect 2819 2373 2869 2415
rect 3037 2373 3087 2415
rect 16513 2639 16563 2681
rect 16721 2639 16771 2681
rect 16939 2639 16989 2681
rect 5682 2374 5732 2416
rect 5900 2374 5950 2416
rect 6108 2374 6158 2416
rect 6975 2386 7025 2428
rect 7183 2386 7233 2428
rect 7401 2386 7451 2428
rect 10059 2386 10109 2428
rect 10277 2386 10327 2428
rect 10485 2386 10535 2428
rect 11352 2398 11402 2440
rect 11560 2398 11610 2440
rect 11778 2398 11828 2440
rect 355 2137 405 2179
rect 573 2137 623 2179
rect 781 2137 831 2179
rect 3409 2189 3459 2231
rect 3617 2189 3667 2231
rect 3835 2189 3885 2231
rect 14423 2399 14473 2441
rect 14641 2399 14691 2441
rect 14849 2399 14899 2441
rect 15716 2411 15766 2453
rect 15924 2411 15974 2453
rect 16142 2411 16192 2453
rect 4719 2150 4769 2192
rect 4937 2150 4987 2192
rect 5145 2150 5195 2192
rect 7773 2202 7823 2244
rect 7981 2202 8031 2244
rect 8199 2202 8249 2244
rect 9096 2162 9146 2204
rect 9314 2162 9364 2204
rect 9522 2162 9572 2204
rect 12150 2214 12200 2256
rect 12358 2214 12408 2256
rect 12576 2214 12626 2256
rect 1153 1953 1203 1995
rect 1371 1953 1421 1995
rect 1579 1953 1629 1995
rect 2512 1963 2562 2005
rect 2720 1963 2770 2005
rect 2938 1963 2988 2005
rect 13460 2175 13510 2217
rect 13678 2175 13728 2217
rect 13886 2175 13936 2217
rect 16514 2227 16564 2269
rect 16722 2227 16772 2269
rect 16940 2227 16990 2269
rect 5517 1966 5567 2008
rect 5735 1966 5785 2008
rect 5943 1966 5993 2008
rect 6876 1976 6926 2018
rect 7084 1976 7134 2018
rect 7302 1976 7352 2018
rect 9894 1978 9944 2020
rect 10112 1978 10162 2020
rect 10320 1978 10370 2020
rect 11253 1988 11303 2030
rect 11461 1988 11511 2030
rect 11679 1988 11729 2030
rect 356 1725 406 1767
rect 574 1725 624 1767
rect 782 1725 832 1767
rect 14258 1991 14308 2033
rect 14476 1991 14526 2033
rect 14684 1991 14734 2033
rect 15617 2001 15667 2043
rect 15825 2001 15875 2043
rect 16043 2001 16093 2043
rect 4720 1738 4770 1780
rect 4938 1738 4988 1780
rect 5146 1738 5196 1780
rect 9097 1750 9147 1792
rect 9315 1750 9365 1792
rect 9523 1750 9573 1792
rect 13461 1763 13511 1805
rect 13679 1763 13729 1805
rect 13887 1763 13937 1805
rect 3391 1583 3441 1625
rect 3599 1583 3649 1625
rect 3817 1583 3867 1625
rect 7755 1596 7805 1638
rect 7963 1596 8013 1638
rect 8181 1596 8231 1638
rect 12132 1608 12182 1650
rect 12340 1608 12390 1650
rect 12558 1608 12608 1650
rect 1235 1345 1285 1387
rect 1453 1345 1503 1387
rect 1661 1345 1711 1387
rect 2594 1355 2644 1397
rect 2802 1355 2852 1397
rect 3020 1355 3070 1397
rect 16496 1621 16546 1663
rect 16704 1621 16754 1663
rect 16922 1621 16972 1663
rect 5599 1358 5649 1400
rect 5817 1358 5867 1400
rect 6025 1358 6075 1400
rect 6958 1368 7008 1410
rect 7166 1368 7216 1410
rect 7384 1368 7434 1410
rect 9976 1370 10026 1412
rect 10194 1370 10244 1412
rect 10402 1370 10452 1412
rect 11335 1380 11385 1422
rect 11543 1380 11593 1422
rect 11761 1380 11811 1422
rect 338 1119 388 1161
rect 556 1119 606 1161
rect 764 1119 814 1161
rect 3392 1171 3442 1213
rect 3600 1171 3650 1213
rect 3818 1171 3868 1213
rect 14340 1383 14390 1425
rect 14558 1383 14608 1425
rect 14766 1383 14816 1425
rect 15699 1393 15749 1435
rect 15907 1393 15957 1435
rect 16125 1393 16175 1435
rect 4702 1132 4752 1174
rect 4920 1132 4970 1174
rect 5128 1132 5178 1174
rect 7756 1184 7806 1226
rect 7964 1184 8014 1226
rect 8182 1184 8232 1226
rect 9079 1144 9129 1186
rect 9297 1144 9347 1186
rect 9505 1144 9555 1186
rect 12133 1196 12183 1238
rect 12341 1196 12391 1238
rect 12559 1196 12609 1238
rect 13443 1157 13493 1199
rect 13661 1157 13711 1199
rect 13869 1157 13919 1199
rect 16497 1209 16547 1251
rect 16705 1209 16755 1251
rect 16923 1209 16973 1251
rect 1136 935 1186 977
rect 1354 935 1404 977
rect 1562 935 1612 977
rect 5500 948 5550 990
rect 5718 948 5768 990
rect 5926 948 5976 990
rect 9877 960 9927 1002
rect 10095 960 10145 1002
rect 10303 960 10353 1002
rect 339 707 389 749
rect 557 707 607 749
rect 765 707 815 749
rect 14241 973 14291 1015
rect 14459 973 14509 1015
rect 14667 973 14717 1015
rect 4703 720 4753 762
rect 4921 720 4971 762
rect 5129 720 5179 762
rect 9080 732 9130 774
rect 9298 732 9348 774
rect 9506 732 9556 774
rect 13444 745 13494 787
rect 13662 745 13712 787
rect 13870 745 13920 787
rect 1552 131 1602 173
rect 1770 131 1820 173
rect 1978 131 2028 173
rect 5916 144 5966 186
rect 6134 144 6184 186
rect 6342 144 6392 186
rect 10293 156 10343 198
rect 10511 156 10561 198
rect 10719 156 10769 198
rect 14657 169 14707 211
rect 14875 169 14925 211
rect 15083 169 15133 211
rect 4041 57 4091 99
rect 4259 57 4309 99
rect 4467 57 4517 99
rect 8489 81 8539 123
rect 8707 81 8757 123
rect 8915 81 8965 123
rect 12782 82 12832 124
rect 13000 82 13050 124
rect 13208 82 13258 124
<< pmos >>
rect 3518 8532 3568 8632
rect 3726 8532 3776 8632
rect 3944 8532 3994 8632
rect 7882 8545 7932 8645
rect 8090 8545 8140 8645
rect 8308 8545 8358 8645
rect 12259 8557 12309 8657
rect 12467 8557 12517 8657
rect 12685 8557 12735 8657
rect 16623 8570 16673 8670
rect 16831 8570 16881 8670
rect 17049 8570 17099 8670
rect 465 8364 515 8464
rect 683 8364 733 8464
rect 891 8364 941 8464
rect 2721 8304 2771 8404
rect 2929 8304 2979 8404
rect 3147 8304 3197 8404
rect 4829 8377 4879 8477
rect 5047 8377 5097 8477
rect 5255 8377 5305 8477
rect 1263 8180 1313 8280
rect 1481 8180 1531 8280
rect 1689 8180 1739 8280
rect 7085 8317 7135 8417
rect 7293 8317 7343 8417
rect 7511 8317 7561 8417
rect 9206 8389 9256 8489
rect 9424 8389 9474 8489
rect 9632 8389 9682 8489
rect 3519 8120 3569 8220
rect 3727 8120 3777 8220
rect 3945 8120 3995 8220
rect 5627 8193 5677 8293
rect 5845 8193 5895 8293
rect 6053 8193 6103 8293
rect 11462 8329 11512 8429
rect 11670 8329 11720 8429
rect 11888 8329 11938 8429
rect 13570 8402 13620 8502
rect 13788 8402 13838 8502
rect 13996 8402 14046 8502
rect 7883 8133 7933 8233
rect 8091 8133 8141 8233
rect 8309 8133 8359 8233
rect 10004 8205 10054 8305
rect 10222 8205 10272 8305
rect 10430 8205 10480 8305
rect 15826 8342 15876 8442
rect 16034 8342 16084 8442
rect 16252 8342 16302 8442
rect 466 7952 516 8052
rect 684 7952 734 8052
rect 892 7952 942 8052
rect 12260 8145 12310 8245
rect 12468 8145 12518 8245
rect 12686 8145 12736 8245
rect 14368 8218 14418 8318
rect 14586 8218 14636 8318
rect 14794 8218 14844 8318
rect 2622 7894 2672 7994
rect 2830 7894 2880 7994
rect 3048 7894 3098 7994
rect 4830 7965 4880 8065
rect 5048 7965 5098 8065
rect 5256 7965 5306 8065
rect 16624 8158 16674 8258
rect 16832 8158 16882 8258
rect 17050 8158 17100 8258
rect 6986 7907 7036 8007
rect 7194 7907 7244 8007
rect 7412 7907 7462 8007
rect 9207 7977 9257 8077
rect 9425 7977 9475 8077
rect 9633 7977 9683 8077
rect 11363 7919 11413 8019
rect 11571 7919 11621 8019
rect 11789 7919 11839 8019
rect 13571 7990 13621 8090
rect 13789 7990 13839 8090
rect 13997 7990 14047 8090
rect 15727 7932 15777 8032
rect 15935 7932 15985 8032
rect 16153 7932 16203 8032
rect 1345 7572 1395 7672
rect 1563 7572 1613 7672
rect 1771 7572 1821 7672
rect 3501 7514 3551 7614
rect 3709 7514 3759 7614
rect 3927 7514 3977 7614
rect 5709 7585 5759 7685
rect 5927 7585 5977 7685
rect 6135 7585 6185 7685
rect 7865 7527 7915 7627
rect 8073 7527 8123 7627
rect 8291 7527 8341 7627
rect 10086 7597 10136 7697
rect 10304 7597 10354 7697
rect 10512 7597 10562 7697
rect 448 7346 498 7446
rect 666 7346 716 7446
rect 874 7346 924 7446
rect 12242 7539 12292 7639
rect 12450 7539 12500 7639
rect 12668 7539 12718 7639
rect 14450 7610 14500 7710
rect 14668 7610 14718 7710
rect 14876 7610 14926 7710
rect 2704 7286 2754 7386
rect 2912 7286 2962 7386
rect 3130 7286 3180 7386
rect 4812 7359 4862 7459
rect 5030 7359 5080 7459
rect 5238 7359 5288 7459
rect 16606 7552 16656 7652
rect 16814 7552 16864 7652
rect 17032 7552 17082 7652
rect 1246 7162 1296 7262
rect 1464 7162 1514 7262
rect 1672 7162 1722 7262
rect 7068 7299 7118 7399
rect 7276 7299 7326 7399
rect 7494 7299 7544 7399
rect 9189 7371 9239 7471
rect 9407 7371 9457 7471
rect 9615 7371 9665 7471
rect 3502 7102 3552 7202
rect 3710 7102 3760 7202
rect 3928 7102 3978 7202
rect 5610 7175 5660 7275
rect 5828 7175 5878 7275
rect 6036 7175 6086 7275
rect 11445 7311 11495 7411
rect 11653 7311 11703 7411
rect 11871 7311 11921 7411
rect 13553 7384 13603 7484
rect 13771 7384 13821 7484
rect 13979 7384 14029 7484
rect 7866 7115 7916 7215
rect 8074 7115 8124 7215
rect 8292 7115 8342 7215
rect 9987 7187 10037 7287
rect 10205 7187 10255 7287
rect 10413 7187 10463 7287
rect 15809 7324 15859 7424
rect 16017 7324 16067 7424
rect 16235 7324 16285 7424
rect 449 6934 499 7034
rect 667 6934 717 7034
rect 875 6934 925 7034
rect 12243 7127 12293 7227
rect 12451 7127 12501 7227
rect 12669 7127 12719 7227
rect 14351 7200 14401 7300
rect 14569 7200 14619 7300
rect 14777 7200 14827 7300
rect 2539 6878 2589 6978
rect 2747 6878 2797 6978
rect 2965 6878 3015 6978
rect 4813 6947 4863 7047
rect 5031 6947 5081 7047
rect 5239 6947 5289 7047
rect 16607 7140 16657 7240
rect 16815 7140 16865 7240
rect 17033 7140 17083 7240
rect 6903 6891 6953 6991
rect 7111 6891 7161 6991
rect 7329 6891 7379 6991
rect 9190 6959 9240 7059
rect 9408 6959 9458 7059
rect 9616 6959 9666 7059
rect 11280 6903 11330 7003
rect 11488 6903 11538 7003
rect 11706 6903 11756 7003
rect 13554 6972 13604 7072
rect 13772 6972 13822 7072
rect 13980 6972 14030 7072
rect 15644 6916 15694 7016
rect 15852 6916 15902 7016
rect 16070 6916 16120 7016
rect 1391 6552 1441 6652
rect 1609 6552 1659 6652
rect 1817 6552 1867 6652
rect 3481 6496 3531 6596
rect 3689 6496 3739 6596
rect 3907 6496 3957 6596
rect 5755 6565 5805 6665
rect 5973 6565 6023 6665
rect 6181 6565 6231 6665
rect 7845 6509 7895 6609
rect 8053 6509 8103 6609
rect 8271 6509 8321 6609
rect 10132 6577 10182 6677
rect 10350 6577 10400 6677
rect 10558 6577 10608 6677
rect 428 6328 478 6428
rect 646 6328 696 6428
rect 854 6328 904 6428
rect 12222 6521 12272 6621
rect 12430 6521 12480 6621
rect 12648 6521 12698 6621
rect 14496 6590 14546 6690
rect 14714 6590 14764 6690
rect 14922 6590 14972 6690
rect 2684 6268 2734 6368
rect 2892 6268 2942 6368
rect 3110 6268 3160 6368
rect 4792 6341 4842 6441
rect 5010 6341 5060 6441
rect 5218 6341 5268 6441
rect 16586 6534 16636 6634
rect 16794 6534 16844 6634
rect 17012 6534 17062 6634
rect 1226 6144 1276 6244
rect 1444 6144 1494 6244
rect 1652 6144 1702 6244
rect 7048 6281 7098 6381
rect 7256 6281 7306 6381
rect 7474 6281 7524 6381
rect 9169 6353 9219 6453
rect 9387 6353 9437 6453
rect 9595 6353 9645 6453
rect 3482 6084 3532 6184
rect 3690 6084 3740 6184
rect 3908 6084 3958 6184
rect 5590 6157 5640 6257
rect 5808 6157 5858 6257
rect 6016 6157 6066 6257
rect 11425 6293 11475 6393
rect 11633 6293 11683 6393
rect 11851 6293 11901 6393
rect 13533 6366 13583 6466
rect 13751 6366 13801 6466
rect 13959 6366 14009 6466
rect 7846 6097 7896 6197
rect 8054 6097 8104 6197
rect 8272 6097 8322 6197
rect 9967 6169 10017 6269
rect 10185 6169 10235 6269
rect 10393 6169 10443 6269
rect 15789 6306 15839 6406
rect 15997 6306 16047 6406
rect 16215 6306 16265 6406
rect 429 5916 479 6016
rect 647 5916 697 6016
rect 855 5916 905 6016
rect 12223 6109 12273 6209
rect 12431 6109 12481 6209
rect 12649 6109 12699 6209
rect 14331 6182 14381 6282
rect 14549 6182 14599 6282
rect 14757 6182 14807 6282
rect 2585 5858 2635 5958
rect 2793 5858 2843 5958
rect 3011 5858 3061 5958
rect 4793 5929 4843 6029
rect 5011 5929 5061 6029
rect 5219 5929 5269 6029
rect 16587 6122 16637 6222
rect 16795 6122 16845 6222
rect 17013 6122 17063 6222
rect 6949 5871 6999 5971
rect 7157 5871 7207 5971
rect 7375 5871 7425 5971
rect 9170 5941 9220 6041
rect 9388 5941 9438 6041
rect 9596 5941 9646 6041
rect 11326 5883 11376 5983
rect 11534 5883 11584 5983
rect 11752 5883 11802 5983
rect 13534 5954 13584 6054
rect 13752 5954 13802 6054
rect 13960 5954 14010 6054
rect 15690 5896 15740 5996
rect 15898 5896 15948 5996
rect 16116 5896 16166 5996
rect 1308 5536 1358 5636
rect 1526 5536 1576 5636
rect 1734 5536 1784 5636
rect 3464 5478 3514 5578
rect 3672 5478 3722 5578
rect 3890 5478 3940 5578
rect 5672 5549 5722 5649
rect 5890 5549 5940 5649
rect 6098 5549 6148 5649
rect 7828 5491 7878 5591
rect 8036 5491 8086 5591
rect 8254 5491 8304 5591
rect 10049 5561 10099 5661
rect 10267 5561 10317 5661
rect 10475 5561 10525 5661
rect 411 5310 461 5410
rect 629 5310 679 5410
rect 837 5310 887 5410
rect 12205 5503 12255 5603
rect 12413 5503 12463 5603
rect 12631 5503 12681 5603
rect 14413 5574 14463 5674
rect 14631 5574 14681 5674
rect 14839 5574 14889 5674
rect 2667 5250 2717 5350
rect 2875 5250 2925 5350
rect 3093 5250 3143 5350
rect 4775 5323 4825 5423
rect 4993 5323 5043 5423
rect 5201 5323 5251 5423
rect 16569 5516 16619 5616
rect 16777 5516 16827 5616
rect 16995 5516 17045 5616
rect 1209 5126 1259 5226
rect 1427 5126 1477 5226
rect 1635 5126 1685 5226
rect 7031 5263 7081 5363
rect 7239 5263 7289 5363
rect 7457 5263 7507 5363
rect 9152 5335 9202 5435
rect 9370 5335 9420 5435
rect 9578 5335 9628 5435
rect 3465 5066 3515 5166
rect 3673 5066 3723 5166
rect 3891 5066 3941 5166
rect 5573 5139 5623 5239
rect 5791 5139 5841 5239
rect 5999 5139 6049 5239
rect 11408 5275 11458 5375
rect 11616 5275 11666 5375
rect 11834 5275 11884 5375
rect 13516 5348 13566 5448
rect 13734 5348 13784 5448
rect 13942 5348 13992 5448
rect 7829 5079 7879 5179
rect 8037 5079 8087 5179
rect 8255 5079 8305 5179
rect 9950 5151 10000 5251
rect 10168 5151 10218 5251
rect 10376 5151 10426 5251
rect 15772 5288 15822 5388
rect 15980 5288 16030 5388
rect 16198 5288 16248 5388
rect 412 4898 462 4998
rect 630 4898 680 4998
rect 838 4898 888 4998
rect 12206 5091 12256 5191
rect 12414 5091 12464 5191
rect 12632 5091 12682 5191
rect 14314 5164 14364 5264
rect 14532 5164 14582 5264
rect 14740 5164 14790 5264
rect 2363 4844 2413 4944
rect 2571 4844 2621 4944
rect 2789 4844 2839 4944
rect 4776 4911 4826 5011
rect 4994 4911 5044 5011
rect 5202 4911 5252 5011
rect 16570 5104 16620 5204
rect 16778 5104 16828 5204
rect 16996 5104 17046 5204
rect 6727 4857 6777 4957
rect 6935 4857 6985 4957
rect 7153 4857 7203 4957
rect 9153 4923 9203 5023
rect 9371 4923 9421 5023
rect 9579 4923 9629 5023
rect 11104 4869 11154 4969
rect 11312 4869 11362 4969
rect 11530 4869 11580 4969
rect 13517 4936 13567 5036
rect 13735 4936 13785 5036
rect 13943 4936 13993 5036
rect 15468 4882 15518 4982
rect 15676 4882 15726 4982
rect 15894 4882 15944 4982
rect 1494 4514 1544 4614
rect 1712 4514 1762 4614
rect 1920 4514 1970 4614
rect 3445 4460 3495 4560
rect 3653 4460 3703 4560
rect 3871 4460 3921 4560
rect 5858 4527 5908 4627
rect 6076 4527 6126 4627
rect 6284 4527 6334 4627
rect 7809 4473 7859 4573
rect 8017 4473 8067 4573
rect 8235 4473 8285 4573
rect 10235 4539 10285 4639
rect 10453 4539 10503 4639
rect 10661 4539 10711 4639
rect 392 4292 442 4392
rect 610 4292 660 4392
rect 818 4292 868 4392
rect 12186 4485 12236 4585
rect 12394 4485 12444 4585
rect 12612 4485 12662 4585
rect 14599 4552 14649 4652
rect 14817 4552 14867 4652
rect 15025 4552 15075 4652
rect 2648 4232 2698 4332
rect 2856 4232 2906 4332
rect 3074 4232 3124 4332
rect 4756 4305 4806 4405
rect 4974 4305 5024 4405
rect 5182 4305 5232 4405
rect 16550 4498 16600 4598
rect 16758 4498 16808 4598
rect 16976 4498 17026 4598
rect 1190 4108 1240 4208
rect 1408 4108 1458 4208
rect 1616 4108 1666 4208
rect 7012 4245 7062 4345
rect 7220 4245 7270 4345
rect 7438 4245 7488 4345
rect 9133 4317 9183 4417
rect 9351 4317 9401 4417
rect 9559 4317 9609 4417
rect 3446 4048 3496 4148
rect 3654 4048 3704 4148
rect 3872 4048 3922 4148
rect 5554 4121 5604 4221
rect 5772 4121 5822 4221
rect 5980 4121 6030 4221
rect 11389 4257 11439 4357
rect 11597 4257 11647 4357
rect 11815 4257 11865 4357
rect 13497 4330 13547 4430
rect 13715 4330 13765 4430
rect 13923 4330 13973 4430
rect 7810 4061 7860 4161
rect 8018 4061 8068 4161
rect 8236 4061 8286 4161
rect 9931 4133 9981 4233
rect 10149 4133 10199 4233
rect 10357 4133 10407 4233
rect 15753 4270 15803 4370
rect 15961 4270 16011 4370
rect 16179 4270 16229 4370
rect 393 3880 443 3980
rect 611 3880 661 3980
rect 819 3880 869 3980
rect 12187 4073 12237 4173
rect 12395 4073 12445 4173
rect 12613 4073 12663 4173
rect 14295 4146 14345 4246
rect 14513 4146 14563 4246
rect 14721 4146 14771 4246
rect 2549 3822 2599 3922
rect 2757 3822 2807 3922
rect 2975 3822 3025 3922
rect 4757 3893 4807 3993
rect 4975 3893 5025 3993
rect 5183 3893 5233 3993
rect 16551 4086 16601 4186
rect 16759 4086 16809 4186
rect 16977 4086 17027 4186
rect 6913 3835 6963 3935
rect 7121 3835 7171 3935
rect 7339 3835 7389 3935
rect 9134 3905 9184 4005
rect 9352 3905 9402 4005
rect 9560 3905 9610 4005
rect 11290 3847 11340 3947
rect 11498 3847 11548 3947
rect 11716 3847 11766 3947
rect 13498 3918 13548 4018
rect 13716 3918 13766 4018
rect 13924 3918 13974 4018
rect 15654 3860 15704 3960
rect 15862 3860 15912 3960
rect 16080 3860 16130 3960
rect 1272 3500 1322 3600
rect 1490 3500 1540 3600
rect 1698 3500 1748 3600
rect 3428 3442 3478 3542
rect 3636 3442 3686 3542
rect 3854 3442 3904 3542
rect 5636 3513 5686 3613
rect 5854 3513 5904 3613
rect 6062 3513 6112 3613
rect 7792 3455 7842 3555
rect 8000 3455 8050 3555
rect 8218 3455 8268 3555
rect 10013 3525 10063 3625
rect 10231 3525 10281 3625
rect 10439 3525 10489 3625
rect 375 3274 425 3374
rect 593 3274 643 3374
rect 801 3274 851 3374
rect 12169 3467 12219 3567
rect 12377 3467 12427 3567
rect 12595 3467 12645 3567
rect 14377 3538 14427 3638
rect 14595 3538 14645 3638
rect 14803 3538 14853 3638
rect 2631 3214 2681 3314
rect 2839 3214 2889 3314
rect 3057 3214 3107 3314
rect 4739 3287 4789 3387
rect 4957 3287 5007 3387
rect 5165 3287 5215 3387
rect 16533 3480 16583 3580
rect 16741 3480 16791 3580
rect 16959 3480 17009 3580
rect 1173 3090 1223 3190
rect 1391 3090 1441 3190
rect 1599 3090 1649 3190
rect 6995 3227 7045 3327
rect 7203 3227 7253 3327
rect 7421 3227 7471 3327
rect 9116 3299 9166 3399
rect 9334 3299 9384 3399
rect 9542 3299 9592 3399
rect 3429 3030 3479 3130
rect 3637 3030 3687 3130
rect 3855 3030 3905 3130
rect 5537 3103 5587 3203
rect 5755 3103 5805 3203
rect 5963 3103 6013 3203
rect 11372 3239 11422 3339
rect 11580 3239 11630 3339
rect 11798 3239 11848 3339
rect 13480 3312 13530 3412
rect 13698 3312 13748 3412
rect 13906 3312 13956 3412
rect 7793 3043 7843 3143
rect 8001 3043 8051 3143
rect 8219 3043 8269 3143
rect 9914 3115 9964 3215
rect 10132 3115 10182 3215
rect 10340 3115 10390 3215
rect 15736 3252 15786 3352
rect 15944 3252 15994 3352
rect 16162 3252 16212 3352
rect 376 2862 426 2962
rect 594 2862 644 2962
rect 802 2862 852 2962
rect 12170 3055 12220 3155
rect 12378 3055 12428 3155
rect 12596 3055 12646 3155
rect 14278 3128 14328 3228
rect 14496 3128 14546 3228
rect 14704 3128 14754 3228
rect 2466 2806 2516 2906
rect 2674 2806 2724 2906
rect 2892 2806 2942 2906
rect 4740 2875 4790 2975
rect 4958 2875 5008 2975
rect 5166 2875 5216 2975
rect 16534 3068 16584 3168
rect 16742 3068 16792 3168
rect 16960 3068 17010 3168
rect 6830 2819 6880 2919
rect 7038 2819 7088 2919
rect 7256 2819 7306 2919
rect 9117 2887 9167 2987
rect 9335 2887 9385 2987
rect 9543 2887 9593 2987
rect 11207 2831 11257 2931
rect 11415 2831 11465 2931
rect 11633 2831 11683 2931
rect 13481 2900 13531 3000
rect 13699 2900 13749 3000
rect 13907 2900 13957 3000
rect 15571 2844 15621 2944
rect 15779 2844 15829 2944
rect 15997 2844 16047 2944
rect 1318 2480 1368 2580
rect 1536 2480 1586 2580
rect 1744 2480 1794 2580
rect 3408 2424 3458 2524
rect 3616 2424 3666 2524
rect 3834 2424 3884 2524
rect 5682 2493 5732 2593
rect 5900 2493 5950 2593
rect 6108 2493 6158 2593
rect 7772 2437 7822 2537
rect 7980 2437 8030 2537
rect 8198 2437 8248 2537
rect 10059 2505 10109 2605
rect 10277 2505 10327 2605
rect 10485 2505 10535 2605
rect 355 2256 405 2356
rect 573 2256 623 2356
rect 781 2256 831 2356
rect 12149 2449 12199 2549
rect 12357 2449 12407 2549
rect 12575 2449 12625 2549
rect 14423 2518 14473 2618
rect 14641 2518 14691 2618
rect 14849 2518 14899 2618
rect 2611 2196 2661 2296
rect 2819 2196 2869 2296
rect 3037 2196 3087 2296
rect 4719 2269 4769 2369
rect 4937 2269 4987 2369
rect 5145 2269 5195 2369
rect 16513 2462 16563 2562
rect 16721 2462 16771 2562
rect 16939 2462 16989 2562
rect 1153 2072 1203 2172
rect 1371 2072 1421 2172
rect 1579 2072 1629 2172
rect 6975 2209 7025 2309
rect 7183 2209 7233 2309
rect 7401 2209 7451 2309
rect 9096 2281 9146 2381
rect 9314 2281 9364 2381
rect 9522 2281 9572 2381
rect 3409 2012 3459 2112
rect 3617 2012 3667 2112
rect 3835 2012 3885 2112
rect 5517 2085 5567 2185
rect 5735 2085 5785 2185
rect 5943 2085 5993 2185
rect 11352 2221 11402 2321
rect 11560 2221 11610 2321
rect 11778 2221 11828 2321
rect 13460 2294 13510 2394
rect 13678 2294 13728 2394
rect 13886 2294 13936 2394
rect 7773 2025 7823 2125
rect 7981 2025 8031 2125
rect 8199 2025 8249 2125
rect 9894 2097 9944 2197
rect 10112 2097 10162 2197
rect 10320 2097 10370 2197
rect 15716 2234 15766 2334
rect 15924 2234 15974 2334
rect 16142 2234 16192 2334
rect 356 1844 406 1944
rect 574 1844 624 1944
rect 782 1844 832 1944
rect 12150 2037 12200 2137
rect 12358 2037 12408 2137
rect 12576 2037 12626 2137
rect 14258 2110 14308 2210
rect 14476 2110 14526 2210
rect 14684 2110 14734 2210
rect 2512 1786 2562 1886
rect 2720 1786 2770 1886
rect 2938 1786 2988 1886
rect 4720 1857 4770 1957
rect 4938 1857 4988 1957
rect 5146 1857 5196 1957
rect 16514 2050 16564 2150
rect 16722 2050 16772 2150
rect 16940 2050 16990 2150
rect 6876 1799 6926 1899
rect 7084 1799 7134 1899
rect 7302 1799 7352 1899
rect 9097 1869 9147 1969
rect 9315 1869 9365 1969
rect 9523 1869 9573 1969
rect 11253 1811 11303 1911
rect 11461 1811 11511 1911
rect 11679 1811 11729 1911
rect 13461 1882 13511 1982
rect 13679 1882 13729 1982
rect 13887 1882 13937 1982
rect 15617 1824 15667 1924
rect 15825 1824 15875 1924
rect 16043 1824 16093 1924
rect 1235 1464 1285 1564
rect 1453 1464 1503 1564
rect 1661 1464 1711 1564
rect 3391 1406 3441 1506
rect 3599 1406 3649 1506
rect 3817 1406 3867 1506
rect 5599 1477 5649 1577
rect 5817 1477 5867 1577
rect 6025 1477 6075 1577
rect 7755 1419 7805 1519
rect 7963 1419 8013 1519
rect 8181 1419 8231 1519
rect 9976 1489 10026 1589
rect 10194 1489 10244 1589
rect 10402 1489 10452 1589
rect 338 1238 388 1338
rect 556 1238 606 1338
rect 764 1238 814 1338
rect 12132 1431 12182 1531
rect 12340 1431 12390 1531
rect 12558 1431 12608 1531
rect 14340 1502 14390 1602
rect 14558 1502 14608 1602
rect 14766 1502 14816 1602
rect 2594 1178 2644 1278
rect 2802 1178 2852 1278
rect 3020 1178 3070 1278
rect 4702 1251 4752 1351
rect 4920 1251 4970 1351
rect 5128 1251 5178 1351
rect 16496 1444 16546 1544
rect 16704 1444 16754 1544
rect 16922 1444 16972 1544
rect 1136 1054 1186 1154
rect 1354 1054 1404 1154
rect 1562 1054 1612 1154
rect 6958 1191 7008 1291
rect 7166 1191 7216 1291
rect 7384 1191 7434 1291
rect 9079 1263 9129 1363
rect 9297 1263 9347 1363
rect 9505 1263 9555 1363
rect 3392 994 3442 1094
rect 3600 994 3650 1094
rect 3818 994 3868 1094
rect 5500 1067 5550 1167
rect 5718 1067 5768 1167
rect 5926 1067 5976 1167
rect 11335 1203 11385 1303
rect 11543 1203 11593 1303
rect 11761 1203 11811 1303
rect 13443 1276 13493 1376
rect 13661 1276 13711 1376
rect 13869 1276 13919 1376
rect 7756 1007 7806 1107
rect 7964 1007 8014 1107
rect 8182 1007 8232 1107
rect 9877 1079 9927 1179
rect 10095 1079 10145 1179
rect 10303 1079 10353 1179
rect 15699 1216 15749 1316
rect 15907 1216 15957 1316
rect 16125 1216 16175 1316
rect 12133 1019 12183 1119
rect 12341 1019 12391 1119
rect 12559 1019 12609 1119
rect 14241 1092 14291 1192
rect 14459 1092 14509 1192
rect 14667 1092 14717 1192
rect 16497 1032 16547 1132
rect 16705 1032 16755 1132
rect 16923 1032 16973 1132
rect 339 826 389 926
rect 557 826 607 926
rect 765 826 815 926
rect 4703 839 4753 939
rect 4921 839 4971 939
rect 5129 839 5179 939
rect 9080 851 9130 951
rect 9298 851 9348 951
rect 9506 851 9556 951
rect 13444 864 13494 964
rect 13662 864 13712 964
rect 13870 864 13920 964
rect 1552 250 1602 350
rect 1770 250 1820 350
rect 1978 250 2028 350
rect 4041 176 4091 276
rect 4259 176 4309 276
rect 4467 176 4517 276
rect 5916 263 5966 363
rect 6134 263 6184 363
rect 6342 263 6392 363
rect 8489 200 8539 300
rect 8707 200 8757 300
rect 8915 200 8965 300
rect 10293 275 10343 375
rect 10511 275 10561 375
rect 10719 275 10769 375
rect 12782 201 12832 301
rect 13000 201 13050 301
rect 13208 201 13258 301
rect 14657 288 14707 388
rect 14875 288 14925 388
rect 15083 288 15133 388
<< ndiff >>
rect 3469 8739 3518 8751
rect 3469 8719 3480 8739
rect 3500 8719 3518 8739
rect 3469 8709 3518 8719
rect 3568 8735 3612 8751
rect 3568 8715 3583 8735
rect 3603 8715 3612 8735
rect 3568 8709 3612 8715
rect 3682 8735 3726 8751
rect 3682 8715 3691 8735
rect 3711 8715 3726 8735
rect 3682 8709 3726 8715
rect 3776 8739 3825 8751
rect 3776 8719 3794 8739
rect 3814 8719 3825 8739
rect 3776 8709 3825 8719
rect 3900 8735 3944 8751
rect 3900 8715 3909 8735
rect 3929 8715 3944 8735
rect 3900 8709 3944 8715
rect 3994 8739 4043 8751
rect 3994 8719 4012 8739
rect 4032 8719 4043 8739
rect 3994 8709 4043 8719
rect 7833 8752 7882 8764
rect 7833 8732 7844 8752
rect 7864 8732 7882 8752
rect 7833 8722 7882 8732
rect 7932 8748 7976 8764
rect 7932 8728 7947 8748
rect 7967 8728 7976 8748
rect 7932 8722 7976 8728
rect 8046 8748 8090 8764
rect 8046 8728 8055 8748
rect 8075 8728 8090 8748
rect 8046 8722 8090 8728
rect 8140 8752 8189 8764
rect 8140 8732 8158 8752
rect 8178 8732 8189 8752
rect 8140 8722 8189 8732
rect 8264 8748 8308 8764
rect 8264 8728 8273 8748
rect 8293 8728 8308 8748
rect 8264 8722 8308 8728
rect 8358 8752 8407 8764
rect 8358 8732 8376 8752
rect 8396 8732 8407 8752
rect 8358 8722 8407 8732
rect 12210 8764 12259 8776
rect 12210 8744 12221 8764
rect 12241 8744 12259 8764
rect 12210 8734 12259 8744
rect 12309 8760 12353 8776
rect 12309 8740 12324 8760
rect 12344 8740 12353 8760
rect 12309 8734 12353 8740
rect 12423 8760 12467 8776
rect 12423 8740 12432 8760
rect 12452 8740 12467 8760
rect 12423 8734 12467 8740
rect 12517 8764 12566 8776
rect 12517 8744 12535 8764
rect 12555 8744 12566 8764
rect 12517 8734 12566 8744
rect 12641 8760 12685 8776
rect 12641 8740 12650 8760
rect 12670 8740 12685 8760
rect 12641 8734 12685 8740
rect 12735 8764 12784 8776
rect 12735 8744 12753 8764
rect 12773 8744 12784 8764
rect 12735 8734 12784 8744
rect 16574 8777 16623 8789
rect 2672 8511 2721 8523
rect 2672 8491 2683 8511
rect 2703 8491 2721 8511
rect 2672 8481 2721 8491
rect 2771 8507 2815 8523
rect 2771 8487 2786 8507
rect 2806 8487 2815 8507
rect 2771 8481 2815 8487
rect 2885 8507 2929 8523
rect 2885 8487 2894 8507
rect 2914 8487 2929 8507
rect 2885 8481 2929 8487
rect 2979 8511 3028 8523
rect 2979 8491 2997 8511
rect 3017 8491 3028 8511
rect 2979 8481 3028 8491
rect 3103 8507 3147 8523
rect 3103 8487 3112 8507
rect 3132 8487 3147 8507
rect 3103 8481 3147 8487
rect 3197 8511 3246 8523
rect 16574 8757 16585 8777
rect 16605 8757 16623 8777
rect 16574 8747 16623 8757
rect 16673 8773 16717 8789
rect 16673 8753 16688 8773
rect 16708 8753 16717 8773
rect 16673 8747 16717 8753
rect 16787 8773 16831 8789
rect 16787 8753 16796 8773
rect 16816 8753 16831 8773
rect 16787 8747 16831 8753
rect 16881 8777 16930 8789
rect 16881 8757 16899 8777
rect 16919 8757 16930 8777
rect 16881 8747 16930 8757
rect 17005 8773 17049 8789
rect 17005 8753 17014 8773
rect 17034 8753 17049 8773
rect 17005 8747 17049 8753
rect 17099 8777 17148 8789
rect 17099 8757 17117 8777
rect 17137 8757 17148 8777
rect 17099 8747 17148 8757
rect 3197 8491 3215 8511
rect 3235 8491 3246 8511
rect 3197 8481 3246 8491
rect 7036 8524 7085 8536
rect 7036 8504 7047 8524
rect 7067 8504 7085 8524
rect 7036 8494 7085 8504
rect 7135 8520 7179 8536
rect 7135 8500 7150 8520
rect 7170 8500 7179 8520
rect 7135 8494 7179 8500
rect 7249 8520 7293 8536
rect 7249 8500 7258 8520
rect 7278 8500 7293 8520
rect 7249 8494 7293 8500
rect 7343 8524 7392 8536
rect 7343 8504 7361 8524
rect 7381 8504 7392 8524
rect 7343 8494 7392 8504
rect 7467 8520 7511 8536
rect 7467 8500 7476 8520
rect 7496 8500 7511 8520
rect 7467 8494 7511 8500
rect 7561 8524 7610 8536
rect 7561 8504 7579 8524
rect 7599 8504 7610 8524
rect 7561 8494 7610 8504
rect 11413 8536 11462 8548
rect 11413 8516 11424 8536
rect 11444 8516 11462 8536
rect 11413 8506 11462 8516
rect 11512 8532 11556 8548
rect 11512 8512 11527 8532
rect 11547 8512 11556 8532
rect 11512 8506 11556 8512
rect 11626 8532 11670 8548
rect 11626 8512 11635 8532
rect 11655 8512 11670 8532
rect 11626 8506 11670 8512
rect 11720 8536 11769 8548
rect 11720 8516 11738 8536
rect 11758 8516 11769 8536
rect 11720 8506 11769 8516
rect 11844 8532 11888 8548
rect 11844 8512 11853 8532
rect 11873 8512 11888 8532
rect 11844 8506 11888 8512
rect 11938 8536 11987 8548
rect 11938 8516 11956 8536
rect 11976 8516 11987 8536
rect 11938 8506 11987 8516
rect 15777 8549 15826 8561
rect 15777 8529 15788 8549
rect 15808 8529 15826 8549
rect 15777 8519 15826 8529
rect 15876 8545 15920 8561
rect 15876 8525 15891 8545
rect 15911 8525 15920 8545
rect 15876 8519 15920 8525
rect 15990 8545 16034 8561
rect 15990 8525 15999 8545
rect 16019 8525 16034 8545
rect 15990 8519 16034 8525
rect 16084 8549 16133 8561
rect 16084 8529 16102 8549
rect 16122 8529 16133 8549
rect 16084 8519 16133 8529
rect 16208 8545 16252 8561
rect 16208 8525 16217 8545
rect 16237 8525 16252 8545
rect 16208 8519 16252 8525
rect 16302 8549 16351 8561
rect 16302 8529 16320 8549
rect 16340 8529 16351 8549
rect 16302 8519 16351 8529
rect 3470 8327 3519 8339
rect 3470 8307 3481 8327
rect 3501 8307 3519 8327
rect 416 8277 465 8287
rect 416 8257 427 8277
rect 447 8257 465 8277
rect 416 8245 465 8257
rect 515 8281 559 8287
rect 515 8261 530 8281
rect 550 8261 559 8281
rect 515 8245 559 8261
rect 634 8277 683 8287
rect 634 8257 645 8277
rect 665 8257 683 8277
rect 634 8245 683 8257
rect 733 8281 777 8287
rect 733 8261 748 8281
rect 768 8261 777 8281
rect 733 8245 777 8261
rect 847 8281 891 8287
rect 847 8261 856 8281
rect 876 8261 891 8281
rect 847 8245 891 8261
rect 941 8277 990 8287
rect 3470 8297 3519 8307
rect 3569 8323 3613 8339
rect 3569 8303 3584 8323
rect 3604 8303 3613 8323
rect 3569 8297 3613 8303
rect 3683 8323 3727 8339
rect 3683 8303 3692 8323
rect 3712 8303 3727 8323
rect 3683 8297 3727 8303
rect 3777 8327 3826 8339
rect 3777 8307 3795 8327
rect 3815 8307 3826 8327
rect 3777 8297 3826 8307
rect 3901 8323 3945 8339
rect 3901 8303 3910 8323
rect 3930 8303 3945 8323
rect 3901 8297 3945 8303
rect 3995 8327 4044 8339
rect 3995 8307 4013 8327
rect 4033 8307 4044 8327
rect 3995 8297 4044 8307
rect 941 8257 959 8277
rect 979 8257 990 8277
rect 941 8245 990 8257
rect 7834 8340 7883 8352
rect 7834 8320 7845 8340
rect 7865 8320 7883 8340
rect 4780 8290 4829 8300
rect 4780 8270 4791 8290
rect 4811 8270 4829 8290
rect 4780 8258 4829 8270
rect 4879 8294 4923 8300
rect 4879 8274 4894 8294
rect 4914 8274 4923 8294
rect 4879 8258 4923 8274
rect 4998 8290 5047 8300
rect 4998 8270 5009 8290
rect 5029 8270 5047 8290
rect 4998 8258 5047 8270
rect 5097 8294 5141 8300
rect 5097 8274 5112 8294
rect 5132 8274 5141 8294
rect 5097 8258 5141 8274
rect 5211 8294 5255 8300
rect 5211 8274 5220 8294
rect 5240 8274 5255 8294
rect 5211 8258 5255 8274
rect 5305 8290 5354 8300
rect 7834 8310 7883 8320
rect 7933 8336 7977 8352
rect 7933 8316 7948 8336
rect 7968 8316 7977 8336
rect 7933 8310 7977 8316
rect 8047 8336 8091 8352
rect 8047 8316 8056 8336
rect 8076 8316 8091 8336
rect 8047 8310 8091 8316
rect 8141 8340 8190 8352
rect 8141 8320 8159 8340
rect 8179 8320 8190 8340
rect 8141 8310 8190 8320
rect 8265 8336 8309 8352
rect 8265 8316 8274 8336
rect 8294 8316 8309 8336
rect 8265 8310 8309 8316
rect 8359 8340 8408 8352
rect 8359 8320 8377 8340
rect 8397 8320 8408 8340
rect 8359 8310 8408 8320
rect 5305 8270 5323 8290
rect 5343 8270 5354 8290
rect 5305 8258 5354 8270
rect 12211 8352 12260 8364
rect 12211 8332 12222 8352
rect 12242 8332 12260 8352
rect 9157 8302 9206 8312
rect 9157 8282 9168 8302
rect 9188 8282 9206 8302
rect 9157 8270 9206 8282
rect 9256 8306 9300 8312
rect 9256 8286 9271 8306
rect 9291 8286 9300 8306
rect 9256 8270 9300 8286
rect 9375 8302 9424 8312
rect 9375 8282 9386 8302
rect 9406 8282 9424 8302
rect 9375 8270 9424 8282
rect 9474 8306 9518 8312
rect 9474 8286 9489 8306
rect 9509 8286 9518 8306
rect 9474 8270 9518 8286
rect 9588 8306 9632 8312
rect 9588 8286 9597 8306
rect 9617 8286 9632 8306
rect 9588 8270 9632 8286
rect 9682 8302 9731 8312
rect 12211 8322 12260 8332
rect 12310 8348 12354 8364
rect 12310 8328 12325 8348
rect 12345 8328 12354 8348
rect 12310 8322 12354 8328
rect 12424 8348 12468 8364
rect 12424 8328 12433 8348
rect 12453 8328 12468 8348
rect 12424 8322 12468 8328
rect 12518 8352 12567 8364
rect 12518 8332 12536 8352
rect 12556 8332 12567 8352
rect 12518 8322 12567 8332
rect 12642 8348 12686 8364
rect 12642 8328 12651 8348
rect 12671 8328 12686 8348
rect 12642 8322 12686 8328
rect 12736 8352 12785 8364
rect 12736 8332 12754 8352
rect 12774 8332 12785 8352
rect 12736 8322 12785 8332
rect 9682 8282 9700 8302
rect 9720 8282 9731 8302
rect 9682 8270 9731 8282
rect 1214 8093 1263 8103
rect 1214 8073 1225 8093
rect 1245 8073 1263 8093
rect 1214 8061 1263 8073
rect 1313 8097 1357 8103
rect 1313 8077 1328 8097
rect 1348 8077 1357 8097
rect 1313 8061 1357 8077
rect 1432 8093 1481 8103
rect 1432 8073 1443 8093
rect 1463 8073 1481 8093
rect 1432 8061 1481 8073
rect 1531 8097 1575 8103
rect 1531 8077 1546 8097
rect 1566 8077 1575 8097
rect 1531 8061 1575 8077
rect 1645 8097 1689 8103
rect 1645 8077 1654 8097
rect 1674 8077 1689 8097
rect 1645 8061 1689 8077
rect 1739 8093 1788 8103
rect 1739 8073 1757 8093
rect 1777 8073 1788 8093
rect 1739 8061 1788 8073
rect 2573 8101 2622 8113
rect 2573 8081 2584 8101
rect 2604 8081 2622 8101
rect 2573 8071 2622 8081
rect 2672 8097 2716 8113
rect 2672 8077 2687 8097
rect 2707 8077 2716 8097
rect 2672 8071 2716 8077
rect 2786 8097 2830 8113
rect 2786 8077 2795 8097
rect 2815 8077 2830 8097
rect 2786 8071 2830 8077
rect 2880 8101 2929 8113
rect 2880 8081 2898 8101
rect 2918 8081 2929 8101
rect 2880 8071 2929 8081
rect 3004 8097 3048 8113
rect 3004 8077 3013 8097
rect 3033 8077 3048 8097
rect 3004 8071 3048 8077
rect 3098 8101 3147 8113
rect 16575 8365 16624 8377
rect 16575 8345 16586 8365
rect 16606 8345 16624 8365
rect 13521 8315 13570 8325
rect 13521 8295 13532 8315
rect 13552 8295 13570 8315
rect 13521 8283 13570 8295
rect 13620 8319 13664 8325
rect 13620 8299 13635 8319
rect 13655 8299 13664 8319
rect 13620 8283 13664 8299
rect 13739 8315 13788 8325
rect 13739 8295 13750 8315
rect 13770 8295 13788 8315
rect 13739 8283 13788 8295
rect 13838 8319 13882 8325
rect 13838 8299 13853 8319
rect 13873 8299 13882 8319
rect 13838 8283 13882 8299
rect 13952 8319 13996 8325
rect 13952 8299 13961 8319
rect 13981 8299 13996 8319
rect 13952 8283 13996 8299
rect 14046 8315 14095 8325
rect 16575 8335 16624 8345
rect 16674 8361 16718 8377
rect 16674 8341 16689 8361
rect 16709 8341 16718 8361
rect 16674 8335 16718 8341
rect 16788 8361 16832 8377
rect 16788 8341 16797 8361
rect 16817 8341 16832 8361
rect 16788 8335 16832 8341
rect 16882 8365 16931 8377
rect 16882 8345 16900 8365
rect 16920 8345 16931 8365
rect 16882 8335 16931 8345
rect 17006 8361 17050 8377
rect 17006 8341 17015 8361
rect 17035 8341 17050 8361
rect 17006 8335 17050 8341
rect 17100 8365 17149 8377
rect 17100 8345 17118 8365
rect 17138 8345 17149 8365
rect 17100 8335 17149 8345
rect 14046 8295 14064 8315
rect 14084 8295 14095 8315
rect 14046 8283 14095 8295
rect 3098 8081 3116 8101
rect 3136 8081 3147 8101
rect 3098 8071 3147 8081
rect 5578 8106 5627 8116
rect 5578 8086 5589 8106
rect 5609 8086 5627 8106
rect 5578 8074 5627 8086
rect 5677 8110 5721 8116
rect 5677 8090 5692 8110
rect 5712 8090 5721 8110
rect 5677 8074 5721 8090
rect 5796 8106 5845 8116
rect 5796 8086 5807 8106
rect 5827 8086 5845 8106
rect 5796 8074 5845 8086
rect 5895 8110 5939 8116
rect 5895 8090 5910 8110
rect 5930 8090 5939 8110
rect 5895 8074 5939 8090
rect 6009 8110 6053 8116
rect 6009 8090 6018 8110
rect 6038 8090 6053 8110
rect 6009 8074 6053 8090
rect 6103 8106 6152 8116
rect 6103 8086 6121 8106
rect 6141 8086 6152 8106
rect 6103 8074 6152 8086
rect 6937 8114 6986 8126
rect 6937 8094 6948 8114
rect 6968 8094 6986 8114
rect 6937 8084 6986 8094
rect 7036 8110 7080 8126
rect 7036 8090 7051 8110
rect 7071 8090 7080 8110
rect 7036 8084 7080 8090
rect 7150 8110 7194 8126
rect 7150 8090 7159 8110
rect 7179 8090 7194 8110
rect 7150 8084 7194 8090
rect 7244 8114 7293 8126
rect 7244 8094 7262 8114
rect 7282 8094 7293 8114
rect 7244 8084 7293 8094
rect 7368 8110 7412 8126
rect 7368 8090 7377 8110
rect 7397 8090 7412 8110
rect 7368 8084 7412 8090
rect 7462 8114 7511 8126
rect 7462 8094 7480 8114
rect 7500 8094 7511 8114
rect 7462 8084 7511 8094
rect 9955 8118 10004 8128
rect 9955 8098 9966 8118
rect 9986 8098 10004 8118
rect 9955 8086 10004 8098
rect 10054 8122 10098 8128
rect 10054 8102 10069 8122
rect 10089 8102 10098 8122
rect 10054 8086 10098 8102
rect 10173 8118 10222 8128
rect 10173 8098 10184 8118
rect 10204 8098 10222 8118
rect 10173 8086 10222 8098
rect 10272 8122 10316 8128
rect 10272 8102 10287 8122
rect 10307 8102 10316 8122
rect 10272 8086 10316 8102
rect 10386 8122 10430 8128
rect 10386 8102 10395 8122
rect 10415 8102 10430 8122
rect 10386 8086 10430 8102
rect 10480 8118 10529 8128
rect 10480 8098 10498 8118
rect 10518 8098 10529 8118
rect 10480 8086 10529 8098
rect 11314 8126 11363 8138
rect 11314 8106 11325 8126
rect 11345 8106 11363 8126
rect 11314 8096 11363 8106
rect 11413 8122 11457 8138
rect 11413 8102 11428 8122
rect 11448 8102 11457 8122
rect 11413 8096 11457 8102
rect 11527 8122 11571 8138
rect 11527 8102 11536 8122
rect 11556 8102 11571 8122
rect 11527 8096 11571 8102
rect 11621 8126 11670 8138
rect 11621 8106 11639 8126
rect 11659 8106 11670 8126
rect 11621 8096 11670 8106
rect 11745 8122 11789 8138
rect 11745 8102 11754 8122
rect 11774 8102 11789 8122
rect 11745 8096 11789 8102
rect 11839 8126 11888 8138
rect 11839 8106 11857 8126
rect 11877 8106 11888 8126
rect 11839 8096 11888 8106
rect 14319 8131 14368 8141
rect 14319 8111 14330 8131
rect 14350 8111 14368 8131
rect 417 7865 466 7875
rect 417 7845 428 7865
rect 448 7845 466 7865
rect 417 7833 466 7845
rect 516 7869 560 7875
rect 516 7849 531 7869
rect 551 7849 560 7869
rect 516 7833 560 7849
rect 635 7865 684 7875
rect 635 7845 646 7865
rect 666 7845 684 7865
rect 635 7833 684 7845
rect 734 7869 778 7875
rect 734 7849 749 7869
rect 769 7849 778 7869
rect 734 7833 778 7849
rect 848 7869 892 7875
rect 848 7849 857 7869
rect 877 7849 892 7869
rect 848 7833 892 7849
rect 942 7865 991 7875
rect 942 7845 960 7865
rect 980 7845 991 7865
rect 14319 8099 14368 8111
rect 14418 8135 14462 8141
rect 14418 8115 14433 8135
rect 14453 8115 14462 8135
rect 14418 8099 14462 8115
rect 14537 8131 14586 8141
rect 14537 8111 14548 8131
rect 14568 8111 14586 8131
rect 14537 8099 14586 8111
rect 14636 8135 14680 8141
rect 14636 8115 14651 8135
rect 14671 8115 14680 8135
rect 14636 8099 14680 8115
rect 14750 8135 14794 8141
rect 14750 8115 14759 8135
rect 14779 8115 14794 8135
rect 14750 8099 14794 8115
rect 14844 8131 14893 8141
rect 14844 8111 14862 8131
rect 14882 8111 14893 8131
rect 14844 8099 14893 8111
rect 15678 8139 15727 8151
rect 15678 8119 15689 8139
rect 15709 8119 15727 8139
rect 15678 8109 15727 8119
rect 15777 8135 15821 8151
rect 15777 8115 15792 8135
rect 15812 8115 15821 8135
rect 15777 8109 15821 8115
rect 15891 8135 15935 8151
rect 15891 8115 15900 8135
rect 15920 8115 15935 8135
rect 15891 8109 15935 8115
rect 15985 8139 16034 8151
rect 15985 8119 16003 8139
rect 16023 8119 16034 8139
rect 15985 8109 16034 8119
rect 16109 8135 16153 8151
rect 16109 8115 16118 8135
rect 16138 8115 16153 8135
rect 16109 8109 16153 8115
rect 16203 8139 16252 8151
rect 16203 8119 16221 8139
rect 16241 8119 16252 8139
rect 16203 8109 16252 8119
rect 942 7833 991 7845
rect 4781 7878 4830 7888
rect 4781 7858 4792 7878
rect 4812 7858 4830 7878
rect 4781 7846 4830 7858
rect 4880 7882 4924 7888
rect 4880 7862 4895 7882
rect 4915 7862 4924 7882
rect 4880 7846 4924 7862
rect 4999 7878 5048 7888
rect 4999 7858 5010 7878
rect 5030 7858 5048 7878
rect 4999 7846 5048 7858
rect 5098 7882 5142 7888
rect 5098 7862 5113 7882
rect 5133 7862 5142 7882
rect 5098 7846 5142 7862
rect 5212 7882 5256 7888
rect 5212 7862 5221 7882
rect 5241 7862 5256 7882
rect 5212 7846 5256 7862
rect 5306 7878 5355 7888
rect 5306 7858 5324 7878
rect 5344 7858 5355 7878
rect 5306 7846 5355 7858
rect 9158 7890 9207 7900
rect 9158 7870 9169 7890
rect 9189 7870 9207 7890
rect 9158 7858 9207 7870
rect 9257 7894 9301 7900
rect 9257 7874 9272 7894
rect 9292 7874 9301 7894
rect 9257 7858 9301 7874
rect 9376 7890 9425 7900
rect 9376 7870 9387 7890
rect 9407 7870 9425 7890
rect 9376 7858 9425 7870
rect 9475 7894 9519 7900
rect 9475 7874 9490 7894
rect 9510 7874 9519 7894
rect 9475 7858 9519 7874
rect 9589 7894 9633 7900
rect 9589 7874 9598 7894
rect 9618 7874 9633 7894
rect 9589 7858 9633 7874
rect 9683 7890 9732 7900
rect 9683 7870 9701 7890
rect 9721 7870 9732 7890
rect 9683 7858 9732 7870
rect 13522 7903 13571 7913
rect 13522 7883 13533 7903
rect 13553 7883 13571 7903
rect 13522 7871 13571 7883
rect 13621 7907 13665 7913
rect 13621 7887 13636 7907
rect 13656 7887 13665 7907
rect 13621 7871 13665 7887
rect 13740 7903 13789 7913
rect 13740 7883 13751 7903
rect 13771 7883 13789 7903
rect 13740 7871 13789 7883
rect 13839 7907 13883 7913
rect 13839 7887 13854 7907
rect 13874 7887 13883 7907
rect 13839 7871 13883 7887
rect 13953 7907 13997 7913
rect 13953 7887 13962 7907
rect 13982 7887 13997 7907
rect 13953 7871 13997 7887
rect 14047 7903 14096 7913
rect 14047 7883 14065 7903
rect 14085 7883 14096 7903
rect 14047 7871 14096 7883
rect 3452 7721 3501 7733
rect 3452 7701 3463 7721
rect 3483 7701 3501 7721
rect 3452 7691 3501 7701
rect 3551 7717 3595 7733
rect 3551 7697 3566 7717
rect 3586 7697 3595 7717
rect 3551 7691 3595 7697
rect 3665 7717 3709 7733
rect 3665 7697 3674 7717
rect 3694 7697 3709 7717
rect 3665 7691 3709 7697
rect 3759 7721 3808 7733
rect 3759 7701 3777 7721
rect 3797 7701 3808 7721
rect 3759 7691 3808 7701
rect 3883 7717 3927 7733
rect 3883 7697 3892 7717
rect 3912 7697 3927 7717
rect 3883 7691 3927 7697
rect 3977 7721 4026 7733
rect 3977 7701 3995 7721
rect 4015 7701 4026 7721
rect 3977 7691 4026 7701
rect 7816 7734 7865 7746
rect 7816 7714 7827 7734
rect 7847 7714 7865 7734
rect 7816 7704 7865 7714
rect 7915 7730 7959 7746
rect 7915 7710 7930 7730
rect 7950 7710 7959 7730
rect 7915 7704 7959 7710
rect 8029 7730 8073 7746
rect 8029 7710 8038 7730
rect 8058 7710 8073 7730
rect 8029 7704 8073 7710
rect 8123 7734 8172 7746
rect 8123 7714 8141 7734
rect 8161 7714 8172 7734
rect 8123 7704 8172 7714
rect 8247 7730 8291 7746
rect 8247 7710 8256 7730
rect 8276 7710 8291 7730
rect 8247 7704 8291 7710
rect 8341 7734 8390 7746
rect 8341 7714 8359 7734
rect 8379 7714 8390 7734
rect 8341 7704 8390 7714
rect 12193 7746 12242 7758
rect 12193 7726 12204 7746
rect 12224 7726 12242 7746
rect 12193 7716 12242 7726
rect 12292 7742 12336 7758
rect 12292 7722 12307 7742
rect 12327 7722 12336 7742
rect 12292 7716 12336 7722
rect 12406 7742 12450 7758
rect 12406 7722 12415 7742
rect 12435 7722 12450 7742
rect 12406 7716 12450 7722
rect 12500 7746 12549 7758
rect 12500 7726 12518 7746
rect 12538 7726 12549 7746
rect 12500 7716 12549 7726
rect 12624 7742 12668 7758
rect 12624 7722 12633 7742
rect 12653 7722 12668 7742
rect 12624 7716 12668 7722
rect 12718 7746 12767 7758
rect 12718 7726 12736 7746
rect 12756 7726 12767 7746
rect 12718 7716 12767 7726
rect 16557 7759 16606 7771
rect 1296 7485 1345 7495
rect 1296 7465 1307 7485
rect 1327 7465 1345 7485
rect 1296 7453 1345 7465
rect 1395 7489 1439 7495
rect 1395 7469 1410 7489
rect 1430 7469 1439 7489
rect 1395 7453 1439 7469
rect 1514 7485 1563 7495
rect 1514 7465 1525 7485
rect 1545 7465 1563 7485
rect 1514 7453 1563 7465
rect 1613 7489 1657 7495
rect 1613 7469 1628 7489
rect 1648 7469 1657 7489
rect 1613 7453 1657 7469
rect 1727 7489 1771 7495
rect 1727 7469 1736 7489
rect 1756 7469 1771 7489
rect 1727 7453 1771 7469
rect 1821 7485 1870 7495
rect 1821 7465 1839 7485
rect 1859 7465 1870 7485
rect 1821 7453 1870 7465
rect 2655 7493 2704 7505
rect 2655 7473 2666 7493
rect 2686 7473 2704 7493
rect 2655 7463 2704 7473
rect 2754 7489 2798 7505
rect 2754 7469 2769 7489
rect 2789 7469 2798 7489
rect 2754 7463 2798 7469
rect 2868 7489 2912 7505
rect 2868 7469 2877 7489
rect 2897 7469 2912 7489
rect 2868 7463 2912 7469
rect 2962 7493 3011 7505
rect 2962 7473 2980 7493
rect 3000 7473 3011 7493
rect 2962 7463 3011 7473
rect 3086 7489 3130 7505
rect 3086 7469 3095 7489
rect 3115 7469 3130 7489
rect 3086 7463 3130 7469
rect 3180 7493 3229 7505
rect 16557 7739 16568 7759
rect 16588 7739 16606 7759
rect 16557 7729 16606 7739
rect 16656 7755 16700 7771
rect 16656 7735 16671 7755
rect 16691 7735 16700 7755
rect 16656 7729 16700 7735
rect 16770 7755 16814 7771
rect 16770 7735 16779 7755
rect 16799 7735 16814 7755
rect 16770 7729 16814 7735
rect 16864 7759 16913 7771
rect 16864 7739 16882 7759
rect 16902 7739 16913 7759
rect 16864 7729 16913 7739
rect 16988 7755 17032 7771
rect 16988 7735 16997 7755
rect 17017 7735 17032 7755
rect 16988 7729 17032 7735
rect 17082 7759 17131 7771
rect 17082 7739 17100 7759
rect 17120 7739 17131 7759
rect 17082 7729 17131 7739
rect 3180 7473 3198 7493
rect 3218 7473 3229 7493
rect 3180 7463 3229 7473
rect 5660 7498 5709 7508
rect 5660 7478 5671 7498
rect 5691 7478 5709 7498
rect 5660 7466 5709 7478
rect 5759 7502 5803 7508
rect 5759 7482 5774 7502
rect 5794 7482 5803 7502
rect 5759 7466 5803 7482
rect 5878 7498 5927 7508
rect 5878 7478 5889 7498
rect 5909 7478 5927 7498
rect 5878 7466 5927 7478
rect 5977 7502 6021 7508
rect 5977 7482 5992 7502
rect 6012 7482 6021 7502
rect 5977 7466 6021 7482
rect 6091 7502 6135 7508
rect 6091 7482 6100 7502
rect 6120 7482 6135 7502
rect 6091 7466 6135 7482
rect 6185 7498 6234 7508
rect 6185 7478 6203 7498
rect 6223 7478 6234 7498
rect 6185 7466 6234 7478
rect 7019 7506 7068 7518
rect 7019 7486 7030 7506
rect 7050 7486 7068 7506
rect 7019 7476 7068 7486
rect 7118 7502 7162 7518
rect 7118 7482 7133 7502
rect 7153 7482 7162 7502
rect 7118 7476 7162 7482
rect 7232 7502 7276 7518
rect 7232 7482 7241 7502
rect 7261 7482 7276 7502
rect 7232 7476 7276 7482
rect 7326 7506 7375 7518
rect 7326 7486 7344 7506
rect 7364 7486 7375 7506
rect 7326 7476 7375 7486
rect 7450 7502 7494 7518
rect 7450 7482 7459 7502
rect 7479 7482 7494 7502
rect 7450 7476 7494 7482
rect 7544 7506 7593 7518
rect 7544 7486 7562 7506
rect 7582 7486 7593 7506
rect 7544 7476 7593 7486
rect 10037 7510 10086 7520
rect 10037 7490 10048 7510
rect 10068 7490 10086 7510
rect 10037 7478 10086 7490
rect 10136 7514 10180 7520
rect 10136 7494 10151 7514
rect 10171 7494 10180 7514
rect 10136 7478 10180 7494
rect 10255 7510 10304 7520
rect 10255 7490 10266 7510
rect 10286 7490 10304 7510
rect 10255 7478 10304 7490
rect 10354 7514 10398 7520
rect 10354 7494 10369 7514
rect 10389 7494 10398 7514
rect 10354 7478 10398 7494
rect 10468 7514 10512 7520
rect 10468 7494 10477 7514
rect 10497 7494 10512 7514
rect 10468 7478 10512 7494
rect 10562 7510 10611 7520
rect 10562 7490 10580 7510
rect 10600 7490 10611 7510
rect 10562 7478 10611 7490
rect 11396 7518 11445 7530
rect 11396 7498 11407 7518
rect 11427 7498 11445 7518
rect 11396 7488 11445 7498
rect 11495 7514 11539 7530
rect 11495 7494 11510 7514
rect 11530 7494 11539 7514
rect 11495 7488 11539 7494
rect 11609 7514 11653 7530
rect 11609 7494 11618 7514
rect 11638 7494 11653 7514
rect 11609 7488 11653 7494
rect 11703 7518 11752 7530
rect 11703 7498 11721 7518
rect 11741 7498 11752 7518
rect 11703 7488 11752 7498
rect 11827 7514 11871 7530
rect 11827 7494 11836 7514
rect 11856 7494 11871 7514
rect 11827 7488 11871 7494
rect 11921 7518 11970 7530
rect 11921 7498 11939 7518
rect 11959 7498 11970 7518
rect 11921 7488 11970 7498
rect 14401 7523 14450 7533
rect 14401 7503 14412 7523
rect 14432 7503 14450 7523
rect 3453 7309 3502 7321
rect 3453 7289 3464 7309
rect 3484 7289 3502 7309
rect 399 7259 448 7269
rect 399 7239 410 7259
rect 430 7239 448 7259
rect 399 7227 448 7239
rect 498 7263 542 7269
rect 498 7243 513 7263
rect 533 7243 542 7263
rect 498 7227 542 7243
rect 617 7259 666 7269
rect 617 7239 628 7259
rect 648 7239 666 7259
rect 617 7227 666 7239
rect 716 7263 760 7269
rect 716 7243 731 7263
rect 751 7243 760 7263
rect 716 7227 760 7243
rect 830 7263 874 7269
rect 830 7243 839 7263
rect 859 7243 874 7263
rect 830 7227 874 7243
rect 924 7259 973 7269
rect 3453 7279 3502 7289
rect 3552 7305 3596 7321
rect 3552 7285 3567 7305
rect 3587 7285 3596 7305
rect 3552 7279 3596 7285
rect 3666 7305 3710 7321
rect 3666 7285 3675 7305
rect 3695 7285 3710 7305
rect 3666 7279 3710 7285
rect 3760 7309 3809 7321
rect 3760 7289 3778 7309
rect 3798 7289 3809 7309
rect 3760 7279 3809 7289
rect 3884 7305 3928 7321
rect 3884 7285 3893 7305
rect 3913 7285 3928 7305
rect 3884 7279 3928 7285
rect 3978 7309 4027 7321
rect 3978 7289 3996 7309
rect 4016 7289 4027 7309
rect 3978 7279 4027 7289
rect 924 7239 942 7259
rect 962 7239 973 7259
rect 924 7227 973 7239
rect 14401 7491 14450 7503
rect 14500 7527 14544 7533
rect 14500 7507 14515 7527
rect 14535 7507 14544 7527
rect 14500 7491 14544 7507
rect 14619 7523 14668 7533
rect 14619 7503 14630 7523
rect 14650 7503 14668 7523
rect 14619 7491 14668 7503
rect 14718 7527 14762 7533
rect 14718 7507 14733 7527
rect 14753 7507 14762 7527
rect 14718 7491 14762 7507
rect 14832 7527 14876 7533
rect 14832 7507 14841 7527
rect 14861 7507 14876 7527
rect 14832 7491 14876 7507
rect 14926 7523 14975 7533
rect 14926 7503 14944 7523
rect 14964 7503 14975 7523
rect 14926 7491 14975 7503
rect 15760 7531 15809 7543
rect 15760 7511 15771 7531
rect 15791 7511 15809 7531
rect 15760 7501 15809 7511
rect 15859 7527 15903 7543
rect 15859 7507 15874 7527
rect 15894 7507 15903 7527
rect 15859 7501 15903 7507
rect 15973 7527 16017 7543
rect 15973 7507 15982 7527
rect 16002 7507 16017 7527
rect 15973 7501 16017 7507
rect 16067 7531 16116 7543
rect 16067 7511 16085 7531
rect 16105 7511 16116 7531
rect 16067 7501 16116 7511
rect 16191 7527 16235 7543
rect 16191 7507 16200 7527
rect 16220 7507 16235 7527
rect 16191 7501 16235 7507
rect 16285 7531 16334 7543
rect 16285 7511 16303 7531
rect 16323 7511 16334 7531
rect 16285 7501 16334 7511
rect 7817 7322 7866 7334
rect 7817 7302 7828 7322
rect 7848 7302 7866 7322
rect 4763 7272 4812 7282
rect 4763 7252 4774 7272
rect 4794 7252 4812 7272
rect 4763 7240 4812 7252
rect 4862 7276 4906 7282
rect 4862 7256 4877 7276
rect 4897 7256 4906 7276
rect 4862 7240 4906 7256
rect 4981 7272 5030 7282
rect 4981 7252 4992 7272
rect 5012 7252 5030 7272
rect 4981 7240 5030 7252
rect 5080 7276 5124 7282
rect 5080 7256 5095 7276
rect 5115 7256 5124 7276
rect 5080 7240 5124 7256
rect 5194 7276 5238 7282
rect 5194 7256 5203 7276
rect 5223 7256 5238 7276
rect 5194 7240 5238 7256
rect 5288 7272 5337 7282
rect 7817 7292 7866 7302
rect 7916 7318 7960 7334
rect 7916 7298 7931 7318
rect 7951 7298 7960 7318
rect 7916 7292 7960 7298
rect 8030 7318 8074 7334
rect 8030 7298 8039 7318
rect 8059 7298 8074 7318
rect 8030 7292 8074 7298
rect 8124 7322 8173 7334
rect 8124 7302 8142 7322
rect 8162 7302 8173 7322
rect 8124 7292 8173 7302
rect 8248 7318 8292 7334
rect 8248 7298 8257 7318
rect 8277 7298 8292 7318
rect 8248 7292 8292 7298
rect 8342 7322 8391 7334
rect 8342 7302 8360 7322
rect 8380 7302 8391 7322
rect 8342 7292 8391 7302
rect 5288 7252 5306 7272
rect 5326 7252 5337 7272
rect 5288 7240 5337 7252
rect 12194 7334 12243 7346
rect 12194 7314 12205 7334
rect 12225 7314 12243 7334
rect 9140 7284 9189 7294
rect 9140 7264 9151 7284
rect 9171 7264 9189 7284
rect 9140 7252 9189 7264
rect 9239 7288 9283 7294
rect 9239 7268 9254 7288
rect 9274 7268 9283 7288
rect 9239 7252 9283 7268
rect 9358 7284 9407 7294
rect 9358 7264 9369 7284
rect 9389 7264 9407 7284
rect 9358 7252 9407 7264
rect 9457 7288 9501 7294
rect 9457 7268 9472 7288
rect 9492 7268 9501 7288
rect 9457 7252 9501 7268
rect 9571 7288 9615 7294
rect 9571 7268 9580 7288
rect 9600 7268 9615 7288
rect 9571 7252 9615 7268
rect 9665 7284 9714 7294
rect 12194 7304 12243 7314
rect 12293 7330 12337 7346
rect 12293 7310 12308 7330
rect 12328 7310 12337 7330
rect 12293 7304 12337 7310
rect 12407 7330 12451 7346
rect 12407 7310 12416 7330
rect 12436 7310 12451 7330
rect 12407 7304 12451 7310
rect 12501 7334 12550 7346
rect 12501 7314 12519 7334
rect 12539 7314 12550 7334
rect 12501 7304 12550 7314
rect 12625 7330 12669 7346
rect 12625 7310 12634 7330
rect 12654 7310 12669 7330
rect 12625 7304 12669 7310
rect 12719 7334 12768 7346
rect 12719 7314 12737 7334
rect 12757 7314 12768 7334
rect 12719 7304 12768 7314
rect 9665 7264 9683 7284
rect 9703 7264 9714 7284
rect 9665 7252 9714 7264
rect 2490 7085 2539 7097
rect 1197 7075 1246 7085
rect 1197 7055 1208 7075
rect 1228 7055 1246 7075
rect 1197 7043 1246 7055
rect 1296 7079 1340 7085
rect 1296 7059 1311 7079
rect 1331 7059 1340 7079
rect 1296 7043 1340 7059
rect 1415 7075 1464 7085
rect 1415 7055 1426 7075
rect 1446 7055 1464 7075
rect 1415 7043 1464 7055
rect 1514 7079 1558 7085
rect 1514 7059 1529 7079
rect 1549 7059 1558 7079
rect 1514 7043 1558 7059
rect 1628 7079 1672 7085
rect 1628 7059 1637 7079
rect 1657 7059 1672 7079
rect 1628 7043 1672 7059
rect 1722 7075 1771 7085
rect 1722 7055 1740 7075
rect 1760 7055 1771 7075
rect 2490 7065 2501 7085
rect 2521 7065 2539 7085
rect 2490 7055 2539 7065
rect 2589 7081 2633 7097
rect 2589 7061 2604 7081
rect 2624 7061 2633 7081
rect 2589 7055 2633 7061
rect 2703 7081 2747 7097
rect 2703 7061 2712 7081
rect 2732 7061 2747 7081
rect 2703 7055 2747 7061
rect 2797 7085 2846 7097
rect 2797 7065 2815 7085
rect 2835 7065 2846 7085
rect 2797 7055 2846 7065
rect 2921 7081 2965 7097
rect 2921 7061 2930 7081
rect 2950 7061 2965 7081
rect 2921 7055 2965 7061
rect 3015 7085 3064 7097
rect 16558 7347 16607 7359
rect 16558 7327 16569 7347
rect 16589 7327 16607 7347
rect 13504 7297 13553 7307
rect 13504 7277 13515 7297
rect 13535 7277 13553 7297
rect 13504 7265 13553 7277
rect 13603 7301 13647 7307
rect 13603 7281 13618 7301
rect 13638 7281 13647 7301
rect 13603 7265 13647 7281
rect 13722 7297 13771 7307
rect 13722 7277 13733 7297
rect 13753 7277 13771 7297
rect 13722 7265 13771 7277
rect 13821 7301 13865 7307
rect 13821 7281 13836 7301
rect 13856 7281 13865 7301
rect 13821 7265 13865 7281
rect 13935 7301 13979 7307
rect 13935 7281 13944 7301
rect 13964 7281 13979 7301
rect 13935 7265 13979 7281
rect 14029 7297 14078 7307
rect 16558 7317 16607 7327
rect 16657 7343 16701 7359
rect 16657 7323 16672 7343
rect 16692 7323 16701 7343
rect 16657 7317 16701 7323
rect 16771 7343 16815 7359
rect 16771 7323 16780 7343
rect 16800 7323 16815 7343
rect 16771 7317 16815 7323
rect 16865 7347 16914 7359
rect 16865 7327 16883 7347
rect 16903 7327 16914 7347
rect 16865 7317 16914 7327
rect 16989 7343 17033 7359
rect 16989 7323 16998 7343
rect 17018 7323 17033 7343
rect 16989 7317 17033 7323
rect 17083 7347 17132 7359
rect 17083 7327 17101 7347
rect 17121 7327 17132 7347
rect 17083 7317 17132 7327
rect 14029 7277 14047 7297
rect 14067 7277 14078 7297
rect 14029 7265 14078 7277
rect 6854 7098 6903 7110
rect 3015 7065 3033 7085
rect 3053 7065 3064 7085
rect 3015 7055 3064 7065
rect 1722 7043 1771 7055
rect 5561 7088 5610 7098
rect 5561 7068 5572 7088
rect 5592 7068 5610 7088
rect 5561 7056 5610 7068
rect 5660 7092 5704 7098
rect 5660 7072 5675 7092
rect 5695 7072 5704 7092
rect 5660 7056 5704 7072
rect 5779 7088 5828 7098
rect 5779 7068 5790 7088
rect 5810 7068 5828 7088
rect 5779 7056 5828 7068
rect 5878 7092 5922 7098
rect 5878 7072 5893 7092
rect 5913 7072 5922 7092
rect 5878 7056 5922 7072
rect 5992 7092 6036 7098
rect 5992 7072 6001 7092
rect 6021 7072 6036 7092
rect 5992 7056 6036 7072
rect 6086 7088 6135 7098
rect 6086 7068 6104 7088
rect 6124 7068 6135 7088
rect 6854 7078 6865 7098
rect 6885 7078 6903 7098
rect 6854 7068 6903 7078
rect 6953 7094 6997 7110
rect 6953 7074 6968 7094
rect 6988 7074 6997 7094
rect 6953 7068 6997 7074
rect 7067 7094 7111 7110
rect 7067 7074 7076 7094
rect 7096 7074 7111 7094
rect 7067 7068 7111 7074
rect 7161 7098 7210 7110
rect 7161 7078 7179 7098
rect 7199 7078 7210 7098
rect 7161 7068 7210 7078
rect 7285 7094 7329 7110
rect 7285 7074 7294 7094
rect 7314 7074 7329 7094
rect 7285 7068 7329 7074
rect 7379 7098 7428 7110
rect 11231 7110 11280 7122
rect 7379 7078 7397 7098
rect 7417 7078 7428 7098
rect 7379 7068 7428 7078
rect 6086 7056 6135 7068
rect 9938 7100 9987 7110
rect 9938 7080 9949 7100
rect 9969 7080 9987 7100
rect 9938 7068 9987 7080
rect 10037 7104 10081 7110
rect 10037 7084 10052 7104
rect 10072 7084 10081 7104
rect 10037 7068 10081 7084
rect 10156 7100 10205 7110
rect 10156 7080 10167 7100
rect 10187 7080 10205 7100
rect 10156 7068 10205 7080
rect 10255 7104 10299 7110
rect 10255 7084 10270 7104
rect 10290 7084 10299 7104
rect 10255 7068 10299 7084
rect 10369 7104 10413 7110
rect 10369 7084 10378 7104
rect 10398 7084 10413 7104
rect 10369 7068 10413 7084
rect 10463 7100 10512 7110
rect 10463 7080 10481 7100
rect 10501 7080 10512 7100
rect 11231 7090 11242 7110
rect 11262 7090 11280 7110
rect 11231 7080 11280 7090
rect 11330 7106 11374 7122
rect 11330 7086 11345 7106
rect 11365 7086 11374 7106
rect 11330 7080 11374 7086
rect 11444 7106 11488 7122
rect 11444 7086 11453 7106
rect 11473 7086 11488 7106
rect 11444 7080 11488 7086
rect 11538 7110 11587 7122
rect 11538 7090 11556 7110
rect 11576 7090 11587 7110
rect 11538 7080 11587 7090
rect 11662 7106 11706 7122
rect 11662 7086 11671 7106
rect 11691 7086 11706 7106
rect 11662 7080 11706 7086
rect 11756 7110 11805 7122
rect 15595 7123 15644 7135
rect 11756 7090 11774 7110
rect 11794 7090 11805 7110
rect 11756 7080 11805 7090
rect 10463 7068 10512 7080
rect 400 6847 449 6857
rect 400 6827 411 6847
rect 431 6827 449 6847
rect 400 6815 449 6827
rect 499 6851 543 6857
rect 499 6831 514 6851
rect 534 6831 543 6851
rect 499 6815 543 6831
rect 618 6847 667 6857
rect 618 6827 629 6847
rect 649 6827 667 6847
rect 618 6815 667 6827
rect 717 6851 761 6857
rect 717 6831 732 6851
rect 752 6831 761 6851
rect 717 6815 761 6831
rect 831 6851 875 6857
rect 831 6831 840 6851
rect 860 6831 875 6851
rect 831 6815 875 6831
rect 925 6847 974 6857
rect 925 6827 943 6847
rect 963 6827 974 6847
rect 14302 7113 14351 7123
rect 14302 7093 14313 7113
rect 14333 7093 14351 7113
rect 14302 7081 14351 7093
rect 14401 7117 14445 7123
rect 14401 7097 14416 7117
rect 14436 7097 14445 7117
rect 14401 7081 14445 7097
rect 14520 7113 14569 7123
rect 14520 7093 14531 7113
rect 14551 7093 14569 7113
rect 14520 7081 14569 7093
rect 14619 7117 14663 7123
rect 14619 7097 14634 7117
rect 14654 7097 14663 7117
rect 14619 7081 14663 7097
rect 14733 7117 14777 7123
rect 14733 7097 14742 7117
rect 14762 7097 14777 7117
rect 14733 7081 14777 7097
rect 14827 7113 14876 7123
rect 14827 7093 14845 7113
rect 14865 7093 14876 7113
rect 15595 7103 15606 7123
rect 15626 7103 15644 7123
rect 15595 7093 15644 7103
rect 15694 7119 15738 7135
rect 15694 7099 15709 7119
rect 15729 7099 15738 7119
rect 15694 7093 15738 7099
rect 15808 7119 15852 7135
rect 15808 7099 15817 7119
rect 15837 7099 15852 7119
rect 15808 7093 15852 7099
rect 15902 7123 15951 7135
rect 15902 7103 15920 7123
rect 15940 7103 15951 7123
rect 15902 7093 15951 7103
rect 16026 7119 16070 7135
rect 16026 7099 16035 7119
rect 16055 7099 16070 7119
rect 16026 7093 16070 7099
rect 16120 7123 16169 7135
rect 16120 7103 16138 7123
rect 16158 7103 16169 7123
rect 16120 7093 16169 7103
rect 14827 7081 14876 7093
rect 925 6815 974 6827
rect 4764 6860 4813 6870
rect 4764 6840 4775 6860
rect 4795 6840 4813 6860
rect 4764 6828 4813 6840
rect 4863 6864 4907 6870
rect 4863 6844 4878 6864
rect 4898 6844 4907 6864
rect 4863 6828 4907 6844
rect 4982 6860 5031 6870
rect 4982 6840 4993 6860
rect 5013 6840 5031 6860
rect 4982 6828 5031 6840
rect 5081 6864 5125 6870
rect 5081 6844 5096 6864
rect 5116 6844 5125 6864
rect 5081 6828 5125 6844
rect 5195 6864 5239 6870
rect 5195 6844 5204 6864
rect 5224 6844 5239 6864
rect 5195 6828 5239 6844
rect 5289 6860 5338 6870
rect 5289 6840 5307 6860
rect 5327 6840 5338 6860
rect 5289 6828 5338 6840
rect 9141 6872 9190 6882
rect 9141 6852 9152 6872
rect 9172 6852 9190 6872
rect 9141 6840 9190 6852
rect 9240 6876 9284 6882
rect 9240 6856 9255 6876
rect 9275 6856 9284 6876
rect 9240 6840 9284 6856
rect 9359 6872 9408 6882
rect 9359 6852 9370 6872
rect 9390 6852 9408 6872
rect 9359 6840 9408 6852
rect 9458 6876 9502 6882
rect 9458 6856 9473 6876
rect 9493 6856 9502 6876
rect 9458 6840 9502 6856
rect 9572 6876 9616 6882
rect 9572 6856 9581 6876
rect 9601 6856 9616 6876
rect 9572 6840 9616 6856
rect 9666 6872 9715 6882
rect 9666 6852 9684 6872
rect 9704 6852 9715 6872
rect 9666 6840 9715 6852
rect 13505 6885 13554 6895
rect 13505 6865 13516 6885
rect 13536 6865 13554 6885
rect 13505 6853 13554 6865
rect 13604 6889 13648 6895
rect 13604 6869 13619 6889
rect 13639 6869 13648 6889
rect 13604 6853 13648 6869
rect 13723 6885 13772 6895
rect 13723 6865 13734 6885
rect 13754 6865 13772 6885
rect 13723 6853 13772 6865
rect 13822 6889 13866 6895
rect 13822 6869 13837 6889
rect 13857 6869 13866 6889
rect 13822 6853 13866 6869
rect 13936 6889 13980 6895
rect 13936 6869 13945 6889
rect 13965 6869 13980 6889
rect 13936 6853 13980 6869
rect 14030 6885 14079 6895
rect 14030 6865 14048 6885
rect 14068 6865 14079 6885
rect 14030 6853 14079 6865
rect 3432 6703 3481 6715
rect 3432 6683 3443 6703
rect 3463 6683 3481 6703
rect 3432 6673 3481 6683
rect 3531 6699 3575 6715
rect 3531 6679 3546 6699
rect 3566 6679 3575 6699
rect 3531 6673 3575 6679
rect 3645 6699 3689 6715
rect 3645 6679 3654 6699
rect 3674 6679 3689 6699
rect 3645 6673 3689 6679
rect 3739 6703 3788 6715
rect 3739 6683 3757 6703
rect 3777 6683 3788 6703
rect 3739 6673 3788 6683
rect 3863 6699 3907 6715
rect 3863 6679 3872 6699
rect 3892 6679 3907 6699
rect 3863 6673 3907 6679
rect 3957 6703 4006 6715
rect 3957 6683 3975 6703
rect 3995 6683 4006 6703
rect 3957 6673 4006 6683
rect 7796 6716 7845 6728
rect 7796 6696 7807 6716
rect 7827 6696 7845 6716
rect 7796 6686 7845 6696
rect 7895 6712 7939 6728
rect 7895 6692 7910 6712
rect 7930 6692 7939 6712
rect 7895 6686 7939 6692
rect 8009 6712 8053 6728
rect 8009 6692 8018 6712
rect 8038 6692 8053 6712
rect 8009 6686 8053 6692
rect 8103 6716 8152 6728
rect 8103 6696 8121 6716
rect 8141 6696 8152 6716
rect 8103 6686 8152 6696
rect 8227 6712 8271 6728
rect 8227 6692 8236 6712
rect 8256 6692 8271 6712
rect 8227 6686 8271 6692
rect 8321 6716 8370 6728
rect 8321 6696 8339 6716
rect 8359 6696 8370 6716
rect 8321 6686 8370 6696
rect 12173 6728 12222 6740
rect 12173 6708 12184 6728
rect 12204 6708 12222 6728
rect 12173 6698 12222 6708
rect 12272 6724 12316 6740
rect 12272 6704 12287 6724
rect 12307 6704 12316 6724
rect 12272 6698 12316 6704
rect 12386 6724 12430 6740
rect 12386 6704 12395 6724
rect 12415 6704 12430 6724
rect 12386 6698 12430 6704
rect 12480 6728 12529 6740
rect 12480 6708 12498 6728
rect 12518 6708 12529 6728
rect 12480 6698 12529 6708
rect 12604 6724 12648 6740
rect 12604 6704 12613 6724
rect 12633 6704 12648 6724
rect 12604 6698 12648 6704
rect 12698 6728 12747 6740
rect 12698 6708 12716 6728
rect 12736 6708 12747 6728
rect 12698 6698 12747 6708
rect 16537 6741 16586 6753
rect 2635 6475 2684 6487
rect 1342 6465 1391 6475
rect 1342 6445 1353 6465
rect 1373 6445 1391 6465
rect 1342 6433 1391 6445
rect 1441 6469 1485 6475
rect 1441 6449 1456 6469
rect 1476 6449 1485 6469
rect 1441 6433 1485 6449
rect 1560 6465 1609 6475
rect 1560 6445 1571 6465
rect 1591 6445 1609 6465
rect 1560 6433 1609 6445
rect 1659 6469 1703 6475
rect 1659 6449 1674 6469
rect 1694 6449 1703 6469
rect 1659 6433 1703 6449
rect 1773 6469 1817 6475
rect 1773 6449 1782 6469
rect 1802 6449 1817 6469
rect 1773 6433 1817 6449
rect 1867 6465 1916 6475
rect 1867 6445 1885 6465
rect 1905 6445 1916 6465
rect 2635 6455 2646 6475
rect 2666 6455 2684 6475
rect 2635 6445 2684 6455
rect 2734 6471 2778 6487
rect 2734 6451 2749 6471
rect 2769 6451 2778 6471
rect 2734 6445 2778 6451
rect 2848 6471 2892 6487
rect 2848 6451 2857 6471
rect 2877 6451 2892 6471
rect 2848 6445 2892 6451
rect 2942 6475 2991 6487
rect 2942 6455 2960 6475
rect 2980 6455 2991 6475
rect 2942 6445 2991 6455
rect 3066 6471 3110 6487
rect 3066 6451 3075 6471
rect 3095 6451 3110 6471
rect 3066 6445 3110 6451
rect 3160 6475 3209 6487
rect 3160 6455 3178 6475
rect 3198 6455 3209 6475
rect 3160 6445 3209 6455
rect 16537 6721 16548 6741
rect 16568 6721 16586 6741
rect 16537 6711 16586 6721
rect 16636 6737 16680 6753
rect 16636 6717 16651 6737
rect 16671 6717 16680 6737
rect 16636 6711 16680 6717
rect 16750 6737 16794 6753
rect 16750 6717 16759 6737
rect 16779 6717 16794 6737
rect 16750 6711 16794 6717
rect 16844 6741 16893 6753
rect 16844 6721 16862 6741
rect 16882 6721 16893 6741
rect 16844 6711 16893 6721
rect 16968 6737 17012 6753
rect 16968 6717 16977 6737
rect 16997 6717 17012 6737
rect 16968 6711 17012 6717
rect 17062 6741 17111 6753
rect 17062 6721 17080 6741
rect 17100 6721 17111 6741
rect 17062 6711 17111 6721
rect 6999 6488 7048 6500
rect 5706 6478 5755 6488
rect 5706 6458 5717 6478
rect 5737 6458 5755 6478
rect 1867 6433 1916 6445
rect 5706 6446 5755 6458
rect 5805 6482 5849 6488
rect 5805 6462 5820 6482
rect 5840 6462 5849 6482
rect 5805 6446 5849 6462
rect 5924 6478 5973 6488
rect 5924 6458 5935 6478
rect 5955 6458 5973 6478
rect 5924 6446 5973 6458
rect 6023 6482 6067 6488
rect 6023 6462 6038 6482
rect 6058 6462 6067 6482
rect 6023 6446 6067 6462
rect 6137 6482 6181 6488
rect 6137 6462 6146 6482
rect 6166 6462 6181 6482
rect 6137 6446 6181 6462
rect 6231 6478 6280 6488
rect 6231 6458 6249 6478
rect 6269 6458 6280 6478
rect 6999 6468 7010 6488
rect 7030 6468 7048 6488
rect 6999 6458 7048 6468
rect 7098 6484 7142 6500
rect 7098 6464 7113 6484
rect 7133 6464 7142 6484
rect 7098 6458 7142 6464
rect 7212 6484 7256 6500
rect 7212 6464 7221 6484
rect 7241 6464 7256 6484
rect 7212 6458 7256 6464
rect 7306 6488 7355 6500
rect 7306 6468 7324 6488
rect 7344 6468 7355 6488
rect 7306 6458 7355 6468
rect 7430 6484 7474 6500
rect 7430 6464 7439 6484
rect 7459 6464 7474 6484
rect 7430 6458 7474 6464
rect 7524 6488 7573 6500
rect 7524 6468 7542 6488
rect 7562 6468 7573 6488
rect 7524 6458 7573 6468
rect 11376 6500 11425 6512
rect 10083 6490 10132 6500
rect 10083 6470 10094 6490
rect 10114 6470 10132 6490
rect 6231 6446 6280 6458
rect 10083 6458 10132 6470
rect 10182 6494 10226 6500
rect 10182 6474 10197 6494
rect 10217 6474 10226 6494
rect 10182 6458 10226 6474
rect 10301 6490 10350 6500
rect 10301 6470 10312 6490
rect 10332 6470 10350 6490
rect 10301 6458 10350 6470
rect 10400 6494 10444 6500
rect 10400 6474 10415 6494
rect 10435 6474 10444 6494
rect 10400 6458 10444 6474
rect 10514 6494 10558 6500
rect 10514 6474 10523 6494
rect 10543 6474 10558 6494
rect 10514 6458 10558 6474
rect 10608 6490 10657 6500
rect 10608 6470 10626 6490
rect 10646 6470 10657 6490
rect 11376 6480 11387 6500
rect 11407 6480 11425 6500
rect 11376 6470 11425 6480
rect 11475 6496 11519 6512
rect 11475 6476 11490 6496
rect 11510 6476 11519 6496
rect 11475 6470 11519 6476
rect 11589 6496 11633 6512
rect 11589 6476 11598 6496
rect 11618 6476 11633 6496
rect 11589 6470 11633 6476
rect 11683 6500 11732 6512
rect 11683 6480 11701 6500
rect 11721 6480 11732 6500
rect 11683 6470 11732 6480
rect 11807 6496 11851 6512
rect 11807 6476 11816 6496
rect 11836 6476 11851 6496
rect 11807 6470 11851 6476
rect 11901 6500 11950 6512
rect 11901 6480 11919 6500
rect 11939 6480 11950 6500
rect 11901 6470 11950 6480
rect 15740 6513 15789 6525
rect 14447 6503 14496 6513
rect 14447 6483 14458 6503
rect 14478 6483 14496 6503
rect 10608 6458 10657 6470
rect 3433 6291 3482 6303
rect 3433 6271 3444 6291
rect 3464 6271 3482 6291
rect 379 6241 428 6251
rect 379 6221 390 6241
rect 410 6221 428 6241
rect 379 6209 428 6221
rect 478 6245 522 6251
rect 478 6225 493 6245
rect 513 6225 522 6245
rect 478 6209 522 6225
rect 597 6241 646 6251
rect 597 6221 608 6241
rect 628 6221 646 6241
rect 597 6209 646 6221
rect 696 6245 740 6251
rect 696 6225 711 6245
rect 731 6225 740 6245
rect 696 6209 740 6225
rect 810 6245 854 6251
rect 810 6225 819 6245
rect 839 6225 854 6245
rect 810 6209 854 6225
rect 904 6241 953 6251
rect 3433 6261 3482 6271
rect 3532 6287 3576 6303
rect 3532 6267 3547 6287
rect 3567 6267 3576 6287
rect 3532 6261 3576 6267
rect 3646 6287 3690 6303
rect 3646 6267 3655 6287
rect 3675 6267 3690 6287
rect 3646 6261 3690 6267
rect 3740 6291 3789 6303
rect 3740 6271 3758 6291
rect 3778 6271 3789 6291
rect 3740 6261 3789 6271
rect 3864 6287 3908 6303
rect 3864 6267 3873 6287
rect 3893 6267 3908 6287
rect 3864 6261 3908 6267
rect 3958 6291 4007 6303
rect 3958 6271 3976 6291
rect 3996 6271 4007 6291
rect 3958 6261 4007 6271
rect 904 6221 922 6241
rect 942 6221 953 6241
rect 904 6209 953 6221
rect 14447 6471 14496 6483
rect 14546 6507 14590 6513
rect 14546 6487 14561 6507
rect 14581 6487 14590 6507
rect 14546 6471 14590 6487
rect 14665 6503 14714 6513
rect 14665 6483 14676 6503
rect 14696 6483 14714 6503
rect 14665 6471 14714 6483
rect 14764 6507 14808 6513
rect 14764 6487 14779 6507
rect 14799 6487 14808 6507
rect 14764 6471 14808 6487
rect 14878 6507 14922 6513
rect 14878 6487 14887 6507
rect 14907 6487 14922 6507
rect 14878 6471 14922 6487
rect 14972 6503 15021 6513
rect 14972 6483 14990 6503
rect 15010 6483 15021 6503
rect 15740 6493 15751 6513
rect 15771 6493 15789 6513
rect 15740 6483 15789 6493
rect 15839 6509 15883 6525
rect 15839 6489 15854 6509
rect 15874 6489 15883 6509
rect 15839 6483 15883 6489
rect 15953 6509 15997 6525
rect 15953 6489 15962 6509
rect 15982 6489 15997 6509
rect 15953 6483 15997 6489
rect 16047 6513 16096 6525
rect 16047 6493 16065 6513
rect 16085 6493 16096 6513
rect 16047 6483 16096 6493
rect 16171 6509 16215 6525
rect 16171 6489 16180 6509
rect 16200 6489 16215 6509
rect 16171 6483 16215 6489
rect 16265 6513 16314 6525
rect 16265 6493 16283 6513
rect 16303 6493 16314 6513
rect 16265 6483 16314 6493
rect 14972 6471 15021 6483
rect 7797 6304 7846 6316
rect 7797 6284 7808 6304
rect 7828 6284 7846 6304
rect 4743 6254 4792 6264
rect 4743 6234 4754 6254
rect 4774 6234 4792 6254
rect 4743 6222 4792 6234
rect 4842 6258 4886 6264
rect 4842 6238 4857 6258
rect 4877 6238 4886 6258
rect 4842 6222 4886 6238
rect 4961 6254 5010 6264
rect 4961 6234 4972 6254
rect 4992 6234 5010 6254
rect 4961 6222 5010 6234
rect 5060 6258 5104 6264
rect 5060 6238 5075 6258
rect 5095 6238 5104 6258
rect 5060 6222 5104 6238
rect 5174 6258 5218 6264
rect 5174 6238 5183 6258
rect 5203 6238 5218 6258
rect 5174 6222 5218 6238
rect 5268 6254 5317 6264
rect 7797 6274 7846 6284
rect 7896 6300 7940 6316
rect 7896 6280 7911 6300
rect 7931 6280 7940 6300
rect 7896 6274 7940 6280
rect 8010 6300 8054 6316
rect 8010 6280 8019 6300
rect 8039 6280 8054 6300
rect 8010 6274 8054 6280
rect 8104 6304 8153 6316
rect 8104 6284 8122 6304
rect 8142 6284 8153 6304
rect 8104 6274 8153 6284
rect 8228 6300 8272 6316
rect 8228 6280 8237 6300
rect 8257 6280 8272 6300
rect 8228 6274 8272 6280
rect 8322 6304 8371 6316
rect 8322 6284 8340 6304
rect 8360 6284 8371 6304
rect 8322 6274 8371 6284
rect 5268 6234 5286 6254
rect 5306 6234 5317 6254
rect 5268 6222 5317 6234
rect 12174 6316 12223 6328
rect 12174 6296 12185 6316
rect 12205 6296 12223 6316
rect 9120 6266 9169 6276
rect 9120 6246 9131 6266
rect 9151 6246 9169 6266
rect 9120 6234 9169 6246
rect 9219 6270 9263 6276
rect 9219 6250 9234 6270
rect 9254 6250 9263 6270
rect 9219 6234 9263 6250
rect 9338 6266 9387 6276
rect 9338 6246 9349 6266
rect 9369 6246 9387 6266
rect 9338 6234 9387 6246
rect 9437 6270 9481 6276
rect 9437 6250 9452 6270
rect 9472 6250 9481 6270
rect 9437 6234 9481 6250
rect 9551 6270 9595 6276
rect 9551 6250 9560 6270
rect 9580 6250 9595 6270
rect 9551 6234 9595 6250
rect 9645 6266 9694 6276
rect 12174 6286 12223 6296
rect 12273 6312 12317 6328
rect 12273 6292 12288 6312
rect 12308 6292 12317 6312
rect 12273 6286 12317 6292
rect 12387 6312 12431 6328
rect 12387 6292 12396 6312
rect 12416 6292 12431 6312
rect 12387 6286 12431 6292
rect 12481 6316 12530 6328
rect 12481 6296 12499 6316
rect 12519 6296 12530 6316
rect 12481 6286 12530 6296
rect 12605 6312 12649 6328
rect 12605 6292 12614 6312
rect 12634 6292 12649 6312
rect 12605 6286 12649 6292
rect 12699 6316 12748 6328
rect 12699 6296 12717 6316
rect 12737 6296 12748 6316
rect 12699 6286 12748 6296
rect 9645 6246 9663 6266
rect 9683 6246 9694 6266
rect 9645 6234 9694 6246
rect 1177 6057 1226 6067
rect 1177 6037 1188 6057
rect 1208 6037 1226 6057
rect 1177 6025 1226 6037
rect 1276 6061 1320 6067
rect 1276 6041 1291 6061
rect 1311 6041 1320 6061
rect 1276 6025 1320 6041
rect 1395 6057 1444 6067
rect 1395 6037 1406 6057
rect 1426 6037 1444 6057
rect 1395 6025 1444 6037
rect 1494 6061 1538 6067
rect 1494 6041 1509 6061
rect 1529 6041 1538 6061
rect 1494 6025 1538 6041
rect 1608 6061 1652 6067
rect 1608 6041 1617 6061
rect 1637 6041 1652 6061
rect 1608 6025 1652 6041
rect 1702 6057 1751 6067
rect 1702 6037 1720 6057
rect 1740 6037 1751 6057
rect 1702 6025 1751 6037
rect 2536 6065 2585 6077
rect 2536 6045 2547 6065
rect 2567 6045 2585 6065
rect 2536 6035 2585 6045
rect 2635 6061 2679 6077
rect 2635 6041 2650 6061
rect 2670 6041 2679 6061
rect 2635 6035 2679 6041
rect 2749 6061 2793 6077
rect 2749 6041 2758 6061
rect 2778 6041 2793 6061
rect 2749 6035 2793 6041
rect 2843 6065 2892 6077
rect 2843 6045 2861 6065
rect 2881 6045 2892 6065
rect 2843 6035 2892 6045
rect 2967 6061 3011 6077
rect 2967 6041 2976 6061
rect 2996 6041 3011 6061
rect 2967 6035 3011 6041
rect 3061 6065 3110 6077
rect 16538 6329 16587 6341
rect 16538 6309 16549 6329
rect 16569 6309 16587 6329
rect 13484 6279 13533 6289
rect 13484 6259 13495 6279
rect 13515 6259 13533 6279
rect 13484 6247 13533 6259
rect 13583 6283 13627 6289
rect 13583 6263 13598 6283
rect 13618 6263 13627 6283
rect 13583 6247 13627 6263
rect 13702 6279 13751 6289
rect 13702 6259 13713 6279
rect 13733 6259 13751 6279
rect 13702 6247 13751 6259
rect 13801 6283 13845 6289
rect 13801 6263 13816 6283
rect 13836 6263 13845 6283
rect 13801 6247 13845 6263
rect 13915 6283 13959 6289
rect 13915 6263 13924 6283
rect 13944 6263 13959 6283
rect 13915 6247 13959 6263
rect 14009 6279 14058 6289
rect 16538 6299 16587 6309
rect 16637 6325 16681 6341
rect 16637 6305 16652 6325
rect 16672 6305 16681 6325
rect 16637 6299 16681 6305
rect 16751 6325 16795 6341
rect 16751 6305 16760 6325
rect 16780 6305 16795 6325
rect 16751 6299 16795 6305
rect 16845 6329 16894 6341
rect 16845 6309 16863 6329
rect 16883 6309 16894 6329
rect 16845 6299 16894 6309
rect 16969 6325 17013 6341
rect 16969 6305 16978 6325
rect 16998 6305 17013 6325
rect 16969 6299 17013 6305
rect 17063 6329 17112 6341
rect 17063 6309 17081 6329
rect 17101 6309 17112 6329
rect 17063 6299 17112 6309
rect 14009 6259 14027 6279
rect 14047 6259 14058 6279
rect 14009 6247 14058 6259
rect 3061 6045 3079 6065
rect 3099 6045 3110 6065
rect 3061 6035 3110 6045
rect 5541 6070 5590 6080
rect 5541 6050 5552 6070
rect 5572 6050 5590 6070
rect 5541 6038 5590 6050
rect 5640 6074 5684 6080
rect 5640 6054 5655 6074
rect 5675 6054 5684 6074
rect 5640 6038 5684 6054
rect 5759 6070 5808 6080
rect 5759 6050 5770 6070
rect 5790 6050 5808 6070
rect 5759 6038 5808 6050
rect 5858 6074 5902 6080
rect 5858 6054 5873 6074
rect 5893 6054 5902 6074
rect 5858 6038 5902 6054
rect 5972 6074 6016 6080
rect 5972 6054 5981 6074
rect 6001 6054 6016 6074
rect 5972 6038 6016 6054
rect 6066 6070 6115 6080
rect 6066 6050 6084 6070
rect 6104 6050 6115 6070
rect 6066 6038 6115 6050
rect 6900 6078 6949 6090
rect 6900 6058 6911 6078
rect 6931 6058 6949 6078
rect 6900 6048 6949 6058
rect 6999 6074 7043 6090
rect 6999 6054 7014 6074
rect 7034 6054 7043 6074
rect 6999 6048 7043 6054
rect 7113 6074 7157 6090
rect 7113 6054 7122 6074
rect 7142 6054 7157 6074
rect 7113 6048 7157 6054
rect 7207 6078 7256 6090
rect 7207 6058 7225 6078
rect 7245 6058 7256 6078
rect 7207 6048 7256 6058
rect 7331 6074 7375 6090
rect 7331 6054 7340 6074
rect 7360 6054 7375 6074
rect 7331 6048 7375 6054
rect 7425 6078 7474 6090
rect 7425 6058 7443 6078
rect 7463 6058 7474 6078
rect 7425 6048 7474 6058
rect 9918 6082 9967 6092
rect 9918 6062 9929 6082
rect 9949 6062 9967 6082
rect 9918 6050 9967 6062
rect 10017 6086 10061 6092
rect 10017 6066 10032 6086
rect 10052 6066 10061 6086
rect 10017 6050 10061 6066
rect 10136 6082 10185 6092
rect 10136 6062 10147 6082
rect 10167 6062 10185 6082
rect 10136 6050 10185 6062
rect 10235 6086 10279 6092
rect 10235 6066 10250 6086
rect 10270 6066 10279 6086
rect 10235 6050 10279 6066
rect 10349 6086 10393 6092
rect 10349 6066 10358 6086
rect 10378 6066 10393 6086
rect 10349 6050 10393 6066
rect 10443 6082 10492 6092
rect 10443 6062 10461 6082
rect 10481 6062 10492 6082
rect 10443 6050 10492 6062
rect 11277 6090 11326 6102
rect 11277 6070 11288 6090
rect 11308 6070 11326 6090
rect 11277 6060 11326 6070
rect 11376 6086 11420 6102
rect 11376 6066 11391 6086
rect 11411 6066 11420 6086
rect 11376 6060 11420 6066
rect 11490 6086 11534 6102
rect 11490 6066 11499 6086
rect 11519 6066 11534 6086
rect 11490 6060 11534 6066
rect 11584 6090 11633 6102
rect 11584 6070 11602 6090
rect 11622 6070 11633 6090
rect 11584 6060 11633 6070
rect 11708 6086 11752 6102
rect 11708 6066 11717 6086
rect 11737 6066 11752 6086
rect 11708 6060 11752 6066
rect 11802 6090 11851 6102
rect 11802 6070 11820 6090
rect 11840 6070 11851 6090
rect 11802 6060 11851 6070
rect 14282 6095 14331 6105
rect 14282 6075 14293 6095
rect 14313 6075 14331 6095
rect 380 5829 429 5839
rect 380 5809 391 5829
rect 411 5809 429 5829
rect 380 5797 429 5809
rect 479 5833 523 5839
rect 479 5813 494 5833
rect 514 5813 523 5833
rect 479 5797 523 5813
rect 598 5829 647 5839
rect 598 5809 609 5829
rect 629 5809 647 5829
rect 598 5797 647 5809
rect 697 5833 741 5839
rect 697 5813 712 5833
rect 732 5813 741 5833
rect 697 5797 741 5813
rect 811 5833 855 5839
rect 811 5813 820 5833
rect 840 5813 855 5833
rect 811 5797 855 5813
rect 905 5829 954 5839
rect 905 5809 923 5829
rect 943 5809 954 5829
rect 14282 6063 14331 6075
rect 14381 6099 14425 6105
rect 14381 6079 14396 6099
rect 14416 6079 14425 6099
rect 14381 6063 14425 6079
rect 14500 6095 14549 6105
rect 14500 6075 14511 6095
rect 14531 6075 14549 6095
rect 14500 6063 14549 6075
rect 14599 6099 14643 6105
rect 14599 6079 14614 6099
rect 14634 6079 14643 6099
rect 14599 6063 14643 6079
rect 14713 6099 14757 6105
rect 14713 6079 14722 6099
rect 14742 6079 14757 6099
rect 14713 6063 14757 6079
rect 14807 6095 14856 6105
rect 14807 6075 14825 6095
rect 14845 6075 14856 6095
rect 14807 6063 14856 6075
rect 15641 6103 15690 6115
rect 15641 6083 15652 6103
rect 15672 6083 15690 6103
rect 15641 6073 15690 6083
rect 15740 6099 15784 6115
rect 15740 6079 15755 6099
rect 15775 6079 15784 6099
rect 15740 6073 15784 6079
rect 15854 6099 15898 6115
rect 15854 6079 15863 6099
rect 15883 6079 15898 6099
rect 15854 6073 15898 6079
rect 15948 6103 15997 6115
rect 15948 6083 15966 6103
rect 15986 6083 15997 6103
rect 15948 6073 15997 6083
rect 16072 6099 16116 6115
rect 16072 6079 16081 6099
rect 16101 6079 16116 6099
rect 16072 6073 16116 6079
rect 16166 6103 16215 6115
rect 16166 6083 16184 6103
rect 16204 6083 16215 6103
rect 16166 6073 16215 6083
rect 905 5797 954 5809
rect 4744 5842 4793 5852
rect 4744 5822 4755 5842
rect 4775 5822 4793 5842
rect 4744 5810 4793 5822
rect 4843 5846 4887 5852
rect 4843 5826 4858 5846
rect 4878 5826 4887 5846
rect 4843 5810 4887 5826
rect 4962 5842 5011 5852
rect 4962 5822 4973 5842
rect 4993 5822 5011 5842
rect 4962 5810 5011 5822
rect 5061 5846 5105 5852
rect 5061 5826 5076 5846
rect 5096 5826 5105 5846
rect 5061 5810 5105 5826
rect 5175 5846 5219 5852
rect 5175 5826 5184 5846
rect 5204 5826 5219 5846
rect 5175 5810 5219 5826
rect 5269 5842 5318 5852
rect 5269 5822 5287 5842
rect 5307 5822 5318 5842
rect 5269 5810 5318 5822
rect 9121 5854 9170 5864
rect 9121 5834 9132 5854
rect 9152 5834 9170 5854
rect 9121 5822 9170 5834
rect 9220 5858 9264 5864
rect 9220 5838 9235 5858
rect 9255 5838 9264 5858
rect 9220 5822 9264 5838
rect 9339 5854 9388 5864
rect 9339 5834 9350 5854
rect 9370 5834 9388 5854
rect 9339 5822 9388 5834
rect 9438 5858 9482 5864
rect 9438 5838 9453 5858
rect 9473 5838 9482 5858
rect 9438 5822 9482 5838
rect 9552 5858 9596 5864
rect 9552 5838 9561 5858
rect 9581 5838 9596 5858
rect 9552 5822 9596 5838
rect 9646 5854 9695 5864
rect 9646 5834 9664 5854
rect 9684 5834 9695 5854
rect 9646 5822 9695 5834
rect 13485 5867 13534 5877
rect 13485 5847 13496 5867
rect 13516 5847 13534 5867
rect 13485 5835 13534 5847
rect 13584 5871 13628 5877
rect 13584 5851 13599 5871
rect 13619 5851 13628 5871
rect 13584 5835 13628 5851
rect 13703 5867 13752 5877
rect 13703 5847 13714 5867
rect 13734 5847 13752 5867
rect 13703 5835 13752 5847
rect 13802 5871 13846 5877
rect 13802 5851 13817 5871
rect 13837 5851 13846 5871
rect 13802 5835 13846 5851
rect 13916 5871 13960 5877
rect 13916 5851 13925 5871
rect 13945 5851 13960 5871
rect 13916 5835 13960 5851
rect 14010 5867 14059 5877
rect 14010 5847 14028 5867
rect 14048 5847 14059 5867
rect 14010 5835 14059 5847
rect 3415 5685 3464 5697
rect 3415 5665 3426 5685
rect 3446 5665 3464 5685
rect 3415 5655 3464 5665
rect 3514 5681 3558 5697
rect 3514 5661 3529 5681
rect 3549 5661 3558 5681
rect 3514 5655 3558 5661
rect 3628 5681 3672 5697
rect 3628 5661 3637 5681
rect 3657 5661 3672 5681
rect 3628 5655 3672 5661
rect 3722 5685 3771 5697
rect 3722 5665 3740 5685
rect 3760 5665 3771 5685
rect 3722 5655 3771 5665
rect 3846 5681 3890 5697
rect 3846 5661 3855 5681
rect 3875 5661 3890 5681
rect 3846 5655 3890 5661
rect 3940 5685 3989 5697
rect 3940 5665 3958 5685
rect 3978 5665 3989 5685
rect 3940 5655 3989 5665
rect 7779 5698 7828 5710
rect 7779 5678 7790 5698
rect 7810 5678 7828 5698
rect 7779 5668 7828 5678
rect 7878 5694 7922 5710
rect 7878 5674 7893 5694
rect 7913 5674 7922 5694
rect 7878 5668 7922 5674
rect 7992 5694 8036 5710
rect 7992 5674 8001 5694
rect 8021 5674 8036 5694
rect 7992 5668 8036 5674
rect 8086 5698 8135 5710
rect 8086 5678 8104 5698
rect 8124 5678 8135 5698
rect 8086 5668 8135 5678
rect 8210 5694 8254 5710
rect 8210 5674 8219 5694
rect 8239 5674 8254 5694
rect 8210 5668 8254 5674
rect 8304 5698 8353 5710
rect 8304 5678 8322 5698
rect 8342 5678 8353 5698
rect 8304 5668 8353 5678
rect 12156 5710 12205 5722
rect 12156 5690 12167 5710
rect 12187 5690 12205 5710
rect 12156 5680 12205 5690
rect 12255 5706 12299 5722
rect 12255 5686 12270 5706
rect 12290 5686 12299 5706
rect 12255 5680 12299 5686
rect 12369 5706 12413 5722
rect 12369 5686 12378 5706
rect 12398 5686 12413 5706
rect 12369 5680 12413 5686
rect 12463 5710 12512 5722
rect 12463 5690 12481 5710
rect 12501 5690 12512 5710
rect 12463 5680 12512 5690
rect 12587 5706 12631 5722
rect 12587 5686 12596 5706
rect 12616 5686 12631 5706
rect 12587 5680 12631 5686
rect 12681 5710 12730 5722
rect 12681 5690 12699 5710
rect 12719 5690 12730 5710
rect 12681 5680 12730 5690
rect 16520 5723 16569 5735
rect 1259 5449 1308 5459
rect 1259 5429 1270 5449
rect 1290 5429 1308 5449
rect 1259 5417 1308 5429
rect 1358 5453 1402 5459
rect 1358 5433 1373 5453
rect 1393 5433 1402 5453
rect 1358 5417 1402 5433
rect 1477 5449 1526 5459
rect 1477 5429 1488 5449
rect 1508 5429 1526 5449
rect 1477 5417 1526 5429
rect 1576 5453 1620 5459
rect 1576 5433 1591 5453
rect 1611 5433 1620 5453
rect 1576 5417 1620 5433
rect 1690 5453 1734 5459
rect 1690 5433 1699 5453
rect 1719 5433 1734 5453
rect 1690 5417 1734 5433
rect 1784 5449 1833 5459
rect 1784 5429 1802 5449
rect 1822 5429 1833 5449
rect 1784 5417 1833 5429
rect 2618 5457 2667 5469
rect 2618 5437 2629 5457
rect 2649 5437 2667 5457
rect 2618 5427 2667 5437
rect 2717 5453 2761 5469
rect 2717 5433 2732 5453
rect 2752 5433 2761 5453
rect 2717 5427 2761 5433
rect 2831 5453 2875 5469
rect 2831 5433 2840 5453
rect 2860 5433 2875 5453
rect 2831 5427 2875 5433
rect 2925 5457 2974 5469
rect 2925 5437 2943 5457
rect 2963 5437 2974 5457
rect 2925 5427 2974 5437
rect 3049 5453 3093 5469
rect 3049 5433 3058 5453
rect 3078 5433 3093 5453
rect 3049 5427 3093 5433
rect 3143 5457 3192 5469
rect 16520 5703 16531 5723
rect 16551 5703 16569 5723
rect 16520 5693 16569 5703
rect 16619 5719 16663 5735
rect 16619 5699 16634 5719
rect 16654 5699 16663 5719
rect 16619 5693 16663 5699
rect 16733 5719 16777 5735
rect 16733 5699 16742 5719
rect 16762 5699 16777 5719
rect 16733 5693 16777 5699
rect 16827 5723 16876 5735
rect 16827 5703 16845 5723
rect 16865 5703 16876 5723
rect 16827 5693 16876 5703
rect 16951 5719 16995 5735
rect 16951 5699 16960 5719
rect 16980 5699 16995 5719
rect 16951 5693 16995 5699
rect 17045 5723 17094 5735
rect 17045 5703 17063 5723
rect 17083 5703 17094 5723
rect 17045 5693 17094 5703
rect 3143 5437 3161 5457
rect 3181 5437 3192 5457
rect 3143 5427 3192 5437
rect 5623 5462 5672 5472
rect 5623 5442 5634 5462
rect 5654 5442 5672 5462
rect 5623 5430 5672 5442
rect 5722 5466 5766 5472
rect 5722 5446 5737 5466
rect 5757 5446 5766 5466
rect 5722 5430 5766 5446
rect 5841 5462 5890 5472
rect 5841 5442 5852 5462
rect 5872 5442 5890 5462
rect 5841 5430 5890 5442
rect 5940 5466 5984 5472
rect 5940 5446 5955 5466
rect 5975 5446 5984 5466
rect 5940 5430 5984 5446
rect 6054 5466 6098 5472
rect 6054 5446 6063 5466
rect 6083 5446 6098 5466
rect 6054 5430 6098 5446
rect 6148 5462 6197 5472
rect 6148 5442 6166 5462
rect 6186 5442 6197 5462
rect 6148 5430 6197 5442
rect 6982 5470 7031 5482
rect 6982 5450 6993 5470
rect 7013 5450 7031 5470
rect 6982 5440 7031 5450
rect 7081 5466 7125 5482
rect 7081 5446 7096 5466
rect 7116 5446 7125 5466
rect 7081 5440 7125 5446
rect 7195 5466 7239 5482
rect 7195 5446 7204 5466
rect 7224 5446 7239 5466
rect 7195 5440 7239 5446
rect 7289 5470 7338 5482
rect 7289 5450 7307 5470
rect 7327 5450 7338 5470
rect 7289 5440 7338 5450
rect 7413 5466 7457 5482
rect 7413 5446 7422 5466
rect 7442 5446 7457 5466
rect 7413 5440 7457 5446
rect 7507 5470 7556 5482
rect 7507 5450 7525 5470
rect 7545 5450 7556 5470
rect 7507 5440 7556 5450
rect 10000 5474 10049 5484
rect 10000 5454 10011 5474
rect 10031 5454 10049 5474
rect 10000 5442 10049 5454
rect 10099 5478 10143 5484
rect 10099 5458 10114 5478
rect 10134 5458 10143 5478
rect 10099 5442 10143 5458
rect 10218 5474 10267 5484
rect 10218 5454 10229 5474
rect 10249 5454 10267 5474
rect 10218 5442 10267 5454
rect 10317 5478 10361 5484
rect 10317 5458 10332 5478
rect 10352 5458 10361 5478
rect 10317 5442 10361 5458
rect 10431 5478 10475 5484
rect 10431 5458 10440 5478
rect 10460 5458 10475 5478
rect 10431 5442 10475 5458
rect 10525 5474 10574 5484
rect 10525 5454 10543 5474
rect 10563 5454 10574 5474
rect 10525 5442 10574 5454
rect 11359 5482 11408 5494
rect 11359 5462 11370 5482
rect 11390 5462 11408 5482
rect 11359 5452 11408 5462
rect 11458 5478 11502 5494
rect 11458 5458 11473 5478
rect 11493 5458 11502 5478
rect 11458 5452 11502 5458
rect 11572 5478 11616 5494
rect 11572 5458 11581 5478
rect 11601 5458 11616 5478
rect 11572 5452 11616 5458
rect 11666 5482 11715 5494
rect 11666 5462 11684 5482
rect 11704 5462 11715 5482
rect 11666 5452 11715 5462
rect 11790 5478 11834 5494
rect 11790 5458 11799 5478
rect 11819 5458 11834 5478
rect 11790 5452 11834 5458
rect 11884 5482 11933 5494
rect 11884 5462 11902 5482
rect 11922 5462 11933 5482
rect 11884 5452 11933 5462
rect 14364 5487 14413 5497
rect 14364 5467 14375 5487
rect 14395 5467 14413 5487
rect 3416 5273 3465 5285
rect 3416 5253 3427 5273
rect 3447 5253 3465 5273
rect 362 5223 411 5233
rect 362 5203 373 5223
rect 393 5203 411 5223
rect 362 5191 411 5203
rect 461 5227 505 5233
rect 461 5207 476 5227
rect 496 5207 505 5227
rect 461 5191 505 5207
rect 580 5223 629 5233
rect 580 5203 591 5223
rect 611 5203 629 5223
rect 580 5191 629 5203
rect 679 5227 723 5233
rect 679 5207 694 5227
rect 714 5207 723 5227
rect 679 5191 723 5207
rect 793 5227 837 5233
rect 793 5207 802 5227
rect 822 5207 837 5227
rect 793 5191 837 5207
rect 887 5223 936 5233
rect 3416 5243 3465 5253
rect 3515 5269 3559 5285
rect 3515 5249 3530 5269
rect 3550 5249 3559 5269
rect 3515 5243 3559 5249
rect 3629 5269 3673 5285
rect 3629 5249 3638 5269
rect 3658 5249 3673 5269
rect 3629 5243 3673 5249
rect 3723 5273 3772 5285
rect 3723 5253 3741 5273
rect 3761 5253 3772 5273
rect 3723 5243 3772 5253
rect 3847 5269 3891 5285
rect 3847 5249 3856 5269
rect 3876 5249 3891 5269
rect 3847 5243 3891 5249
rect 3941 5273 3990 5285
rect 3941 5253 3959 5273
rect 3979 5253 3990 5273
rect 3941 5243 3990 5253
rect 887 5203 905 5223
rect 925 5203 936 5223
rect 887 5191 936 5203
rect 14364 5455 14413 5467
rect 14463 5491 14507 5497
rect 14463 5471 14478 5491
rect 14498 5471 14507 5491
rect 14463 5455 14507 5471
rect 14582 5487 14631 5497
rect 14582 5467 14593 5487
rect 14613 5467 14631 5487
rect 14582 5455 14631 5467
rect 14681 5491 14725 5497
rect 14681 5471 14696 5491
rect 14716 5471 14725 5491
rect 14681 5455 14725 5471
rect 14795 5491 14839 5497
rect 14795 5471 14804 5491
rect 14824 5471 14839 5491
rect 14795 5455 14839 5471
rect 14889 5487 14938 5497
rect 14889 5467 14907 5487
rect 14927 5467 14938 5487
rect 14889 5455 14938 5467
rect 15723 5495 15772 5507
rect 15723 5475 15734 5495
rect 15754 5475 15772 5495
rect 15723 5465 15772 5475
rect 15822 5491 15866 5507
rect 15822 5471 15837 5491
rect 15857 5471 15866 5491
rect 15822 5465 15866 5471
rect 15936 5491 15980 5507
rect 15936 5471 15945 5491
rect 15965 5471 15980 5491
rect 15936 5465 15980 5471
rect 16030 5495 16079 5507
rect 16030 5475 16048 5495
rect 16068 5475 16079 5495
rect 16030 5465 16079 5475
rect 16154 5491 16198 5507
rect 16154 5471 16163 5491
rect 16183 5471 16198 5491
rect 16154 5465 16198 5471
rect 16248 5495 16297 5507
rect 16248 5475 16266 5495
rect 16286 5475 16297 5495
rect 16248 5465 16297 5475
rect 7780 5286 7829 5298
rect 7780 5266 7791 5286
rect 7811 5266 7829 5286
rect 4726 5236 4775 5246
rect 4726 5216 4737 5236
rect 4757 5216 4775 5236
rect 4726 5204 4775 5216
rect 4825 5240 4869 5246
rect 4825 5220 4840 5240
rect 4860 5220 4869 5240
rect 4825 5204 4869 5220
rect 4944 5236 4993 5246
rect 4944 5216 4955 5236
rect 4975 5216 4993 5236
rect 4944 5204 4993 5216
rect 5043 5240 5087 5246
rect 5043 5220 5058 5240
rect 5078 5220 5087 5240
rect 5043 5204 5087 5220
rect 5157 5240 5201 5246
rect 5157 5220 5166 5240
rect 5186 5220 5201 5240
rect 5157 5204 5201 5220
rect 5251 5236 5300 5246
rect 7780 5256 7829 5266
rect 7879 5282 7923 5298
rect 7879 5262 7894 5282
rect 7914 5262 7923 5282
rect 7879 5256 7923 5262
rect 7993 5282 8037 5298
rect 7993 5262 8002 5282
rect 8022 5262 8037 5282
rect 7993 5256 8037 5262
rect 8087 5286 8136 5298
rect 8087 5266 8105 5286
rect 8125 5266 8136 5286
rect 8087 5256 8136 5266
rect 8211 5282 8255 5298
rect 8211 5262 8220 5282
rect 8240 5262 8255 5282
rect 8211 5256 8255 5262
rect 8305 5286 8354 5298
rect 8305 5266 8323 5286
rect 8343 5266 8354 5286
rect 8305 5256 8354 5266
rect 5251 5216 5269 5236
rect 5289 5216 5300 5236
rect 5251 5204 5300 5216
rect 12157 5298 12206 5310
rect 12157 5278 12168 5298
rect 12188 5278 12206 5298
rect 9103 5248 9152 5258
rect 9103 5228 9114 5248
rect 9134 5228 9152 5248
rect 9103 5216 9152 5228
rect 9202 5252 9246 5258
rect 9202 5232 9217 5252
rect 9237 5232 9246 5252
rect 9202 5216 9246 5232
rect 9321 5248 9370 5258
rect 9321 5228 9332 5248
rect 9352 5228 9370 5248
rect 9321 5216 9370 5228
rect 9420 5252 9464 5258
rect 9420 5232 9435 5252
rect 9455 5232 9464 5252
rect 9420 5216 9464 5232
rect 9534 5252 9578 5258
rect 9534 5232 9543 5252
rect 9563 5232 9578 5252
rect 9534 5216 9578 5232
rect 9628 5248 9677 5258
rect 12157 5268 12206 5278
rect 12256 5294 12300 5310
rect 12256 5274 12271 5294
rect 12291 5274 12300 5294
rect 12256 5268 12300 5274
rect 12370 5294 12414 5310
rect 12370 5274 12379 5294
rect 12399 5274 12414 5294
rect 12370 5268 12414 5274
rect 12464 5298 12513 5310
rect 12464 5278 12482 5298
rect 12502 5278 12513 5298
rect 12464 5268 12513 5278
rect 12588 5294 12632 5310
rect 12588 5274 12597 5294
rect 12617 5274 12632 5294
rect 12588 5268 12632 5274
rect 12682 5298 12731 5310
rect 12682 5278 12700 5298
rect 12720 5278 12731 5298
rect 12682 5268 12731 5278
rect 9628 5228 9646 5248
rect 9666 5228 9677 5248
rect 9628 5216 9677 5228
rect 2314 5051 2363 5063
rect 1160 5039 1209 5049
rect 1160 5019 1171 5039
rect 1191 5019 1209 5039
rect 1160 5007 1209 5019
rect 1259 5043 1303 5049
rect 1259 5023 1274 5043
rect 1294 5023 1303 5043
rect 1259 5007 1303 5023
rect 1378 5039 1427 5049
rect 1378 5019 1389 5039
rect 1409 5019 1427 5039
rect 1378 5007 1427 5019
rect 1477 5043 1521 5049
rect 1477 5023 1492 5043
rect 1512 5023 1521 5043
rect 1477 5007 1521 5023
rect 1591 5043 1635 5049
rect 1591 5023 1600 5043
rect 1620 5023 1635 5043
rect 1591 5007 1635 5023
rect 1685 5039 1734 5049
rect 1685 5019 1703 5039
rect 1723 5019 1734 5039
rect 2314 5031 2325 5051
rect 2345 5031 2363 5051
rect 2314 5021 2363 5031
rect 2413 5047 2457 5063
rect 2413 5027 2428 5047
rect 2448 5027 2457 5047
rect 2413 5021 2457 5027
rect 2527 5047 2571 5063
rect 2527 5027 2536 5047
rect 2556 5027 2571 5047
rect 2527 5021 2571 5027
rect 2621 5051 2670 5063
rect 2621 5031 2639 5051
rect 2659 5031 2670 5051
rect 2621 5021 2670 5031
rect 2745 5047 2789 5063
rect 2745 5027 2754 5047
rect 2774 5027 2789 5047
rect 2745 5021 2789 5027
rect 2839 5051 2888 5063
rect 16521 5311 16570 5323
rect 16521 5291 16532 5311
rect 16552 5291 16570 5311
rect 13467 5261 13516 5271
rect 13467 5241 13478 5261
rect 13498 5241 13516 5261
rect 13467 5229 13516 5241
rect 13566 5265 13610 5271
rect 13566 5245 13581 5265
rect 13601 5245 13610 5265
rect 13566 5229 13610 5245
rect 13685 5261 13734 5271
rect 13685 5241 13696 5261
rect 13716 5241 13734 5261
rect 13685 5229 13734 5241
rect 13784 5265 13828 5271
rect 13784 5245 13799 5265
rect 13819 5245 13828 5265
rect 13784 5229 13828 5245
rect 13898 5265 13942 5271
rect 13898 5245 13907 5265
rect 13927 5245 13942 5265
rect 13898 5229 13942 5245
rect 13992 5261 14041 5271
rect 16521 5281 16570 5291
rect 16620 5307 16664 5323
rect 16620 5287 16635 5307
rect 16655 5287 16664 5307
rect 16620 5281 16664 5287
rect 16734 5307 16778 5323
rect 16734 5287 16743 5307
rect 16763 5287 16778 5307
rect 16734 5281 16778 5287
rect 16828 5311 16877 5323
rect 16828 5291 16846 5311
rect 16866 5291 16877 5311
rect 16828 5281 16877 5291
rect 16952 5307 16996 5323
rect 16952 5287 16961 5307
rect 16981 5287 16996 5307
rect 16952 5281 16996 5287
rect 17046 5311 17095 5323
rect 17046 5291 17064 5311
rect 17084 5291 17095 5311
rect 17046 5281 17095 5291
rect 13992 5241 14010 5261
rect 14030 5241 14041 5261
rect 13992 5229 14041 5241
rect 6678 5064 6727 5076
rect 2839 5031 2857 5051
rect 2877 5031 2888 5051
rect 2839 5021 2888 5031
rect 1685 5007 1734 5019
rect 5524 5052 5573 5062
rect 5524 5032 5535 5052
rect 5555 5032 5573 5052
rect 5524 5020 5573 5032
rect 5623 5056 5667 5062
rect 5623 5036 5638 5056
rect 5658 5036 5667 5056
rect 5623 5020 5667 5036
rect 5742 5052 5791 5062
rect 5742 5032 5753 5052
rect 5773 5032 5791 5052
rect 5742 5020 5791 5032
rect 5841 5056 5885 5062
rect 5841 5036 5856 5056
rect 5876 5036 5885 5056
rect 5841 5020 5885 5036
rect 5955 5056 5999 5062
rect 5955 5036 5964 5056
rect 5984 5036 5999 5056
rect 5955 5020 5999 5036
rect 6049 5052 6098 5062
rect 6049 5032 6067 5052
rect 6087 5032 6098 5052
rect 6678 5044 6689 5064
rect 6709 5044 6727 5064
rect 6678 5034 6727 5044
rect 6777 5060 6821 5076
rect 6777 5040 6792 5060
rect 6812 5040 6821 5060
rect 6777 5034 6821 5040
rect 6891 5060 6935 5076
rect 6891 5040 6900 5060
rect 6920 5040 6935 5060
rect 6891 5034 6935 5040
rect 6985 5064 7034 5076
rect 6985 5044 7003 5064
rect 7023 5044 7034 5064
rect 6985 5034 7034 5044
rect 7109 5060 7153 5076
rect 7109 5040 7118 5060
rect 7138 5040 7153 5060
rect 7109 5034 7153 5040
rect 7203 5064 7252 5076
rect 11055 5076 11104 5088
rect 7203 5044 7221 5064
rect 7241 5044 7252 5064
rect 7203 5034 7252 5044
rect 6049 5020 6098 5032
rect 9901 5064 9950 5074
rect 9901 5044 9912 5064
rect 9932 5044 9950 5064
rect 9901 5032 9950 5044
rect 10000 5068 10044 5074
rect 10000 5048 10015 5068
rect 10035 5048 10044 5068
rect 10000 5032 10044 5048
rect 10119 5064 10168 5074
rect 10119 5044 10130 5064
rect 10150 5044 10168 5064
rect 10119 5032 10168 5044
rect 10218 5068 10262 5074
rect 10218 5048 10233 5068
rect 10253 5048 10262 5068
rect 10218 5032 10262 5048
rect 10332 5068 10376 5074
rect 10332 5048 10341 5068
rect 10361 5048 10376 5068
rect 10332 5032 10376 5048
rect 10426 5064 10475 5074
rect 10426 5044 10444 5064
rect 10464 5044 10475 5064
rect 11055 5056 11066 5076
rect 11086 5056 11104 5076
rect 11055 5046 11104 5056
rect 11154 5072 11198 5088
rect 11154 5052 11169 5072
rect 11189 5052 11198 5072
rect 11154 5046 11198 5052
rect 11268 5072 11312 5088
rect 11268 5052 11277 5072
rect 11297 5052 11312 5072
rect 11268 5046 11312 5052
rect 11362 5076 11411 5088
rect 11362 5056 11380 5076
rect 11400 5056 11411 5076
rect 11362 5046 11411 5056
rect 11486 5072 11530 5088
rect 11486 5052 11495 5072
rect 11515 5052 11530 5072
rect 11486 5046 11530 5052
rect 11580 5076 11629 5088
rect 15419 5089 15468 5101
rect 11580 5056 11598 5076
rect 11618 5056 11629 5076
rect 11580 5046 11629 5056
rect 10426 5032 10475 5044
rect 363 4811 412 4821
rect 363 4791 374 4811
rect 394 4791 412 4811
rect 363 4779 412 4791
rect 462 4815 506 4821
rect 462 4795 477 4815
rect 497 4795 506 4815
rect 462 4779 506 4795
rect 581 4811 630 4821
rect 581 4791 592 4811
rect 612 4791 630 4811
rect 581 4779 630 4791
rect 680 4815 724 4821
rect 680 4795 695 4815
rect 715 4795 724 4815
rect 680 4779 724 4795
rect 794 4815 838 4821
rect 794 4795 803 4815
rect 823 4795 838 4815
rect 794 4779 838 4795
rect 888 4811 937 4821
rect 888 4791 906 4811
rect 926 4791 937 4811
rect 14265 5077 14314 5087
rect 14265 5057 14276 5077
rect 14296 5057 14314 5077
rect 14265 5045 14314 5057
rect 14364 5081 14408 5087
rect 14364 5061 14379 5081
rect 14399 5061 14408 5081
rect 14364 5045 14408 5061
rect 14483 5077 14532 5087
rect 14483 5057 14494 5077
rect 14514 5057 14532 5077
rect 14483 5045 14532 5057
rect 14582 5081 14626 5087
rect 14582 5061 14597 5081
rect 14617 5061 14626 5081
rect 14582 5045 14626 5061
rect 14696 5081 14740 5087
rect 14696 5061 14705 5081
rect 14725 5061 14740 5081
rect 14696 5045 14740 5061
rect 14790 5077 14839 5087
rect 14790 5057 14808 5077
rect 14828 5057 14839 5077
rect 15419 5069 15430 5089
rect 15450 5069 15468 5089
rect 15419 5059 15468 5069
rect 15518 5085 15562 5101
rect 15518 5065 15533 5085
rect 15553 5065 15562 5085
rect 15518 5059 15562 5065
rect 15632 5085 15676 5101
rect 15632 5065 15641 5085
rect 15661 5065 15676 5085
rect 15632 5059 15676 5065
rect 15726 5089 15775 5101
rect 15726 5069 15744 5089
rect 15764 5069 15775 5089
rect 15726 5059 15775 5069
rect 15850 5085 15894 5101
rect 15850 5065 15859 5085
rect 15879 5065 15894 5085
rect 15850 5059 15894 5065
rect 15944 5089 15993 5101
rect 15944 5069 15962 5089
rect 15982 5069 15993 5089
rect 15944 5059 15993 5069
rect 14790 5045 14839 5057
rect 888 4779 937 4791
rect 4727 4824 4776 4834
rect 4727 4804 4738 4824
rect 4758 4804 4776 4824
rect 4727 4792 4776 4804
rect 4826 4828 4870 4834
rect 4826 4808 4841 4828
rect 4861 4808 4870 4828
rect 4826 4792 4870 4808
rect 4945 4824 4994 4834
rect 4945 4804 4956 4824
rect 4976 4804 4994 4824
rect 4945 4792 4994 4804
rect 5044 4828 5088 4834
rect 5044 4808 5059 4828
rect 5079 4808 5088 4828
rect 5044 4792 5088 4808
rect 5158 4828 5202 4834
rect 5158 4808 5167 4828
rect 5187 4808 5202 4828
rect 5158 4792 5202 4808
rect 5252 4824 5301 4834
rect 5252 4804 5270 4824
rect 5290 4804 5301 4824
rect 5252 4792 5301 4804
rect 9104 4836 9153 4846
rect 9104 4816 9115 4836
rect 9135 4816 9153 4836
rect 9104 4804 9153 4816
rect 9203 4840 9247 4846
rect 9203 4820 9218 4840
rect 9238 4820 9247 4840
rect 9203 4804 9247 4820
rect 9322 4836 9371 4846
rect 9322 4816 9333 4836
rect 9353 4816 9371 4836
rect 9322 4804 9371 4816
rect 9421 4840 9465 4846
rect 9421 4820 9436 4840
rect 9456 4820 9465 4840
rect 9421 4804 9465 4820
rect 9535 4840 9579 4846
rect 9535 4820 9544 4840
rect 9564 4820 9579 4840
rect 9535 4804 9579 4820
rect 9629 4836 9678 4846
rect 9629 4816 9647 4836
rect 9667 4816 9678 4836
rect 9629 4804 9678 4816
rect 13468 4849 13517 4859
rect 13468 4829 13479 4849
rect 13499 4829 13517 4849
rect 13468 4817 13517 4829
rect 13567 4853 13611 4859
rect 13567 4833 13582 4853
rect 13602 4833 13611 4853
rect 13567 4817 13611 4833
rect 13686 4849 13735 4859
rect 13686 4829 13697 4849
rect 13717 4829 13735 4849
rect 13686 4817 13735 4829
rect 13785 4853 13829 4859
rect 13785 4833 13800 4853
rect 13820 4833 13829 4853
rect 13785 4817 13829 4833
rect 13899 4853 13943 4859
rect 13899 4833 13908 4853
rect 13928 4833 13943 4853
rect 13899 4817 13943 4833
rect 13993 4849 14042 4859
rect 13993 4829 14011 4849
rect 14031 4829 14042 4849
rect 13993 4817 14042 4829
rect 3396 4667 3445 4679
rect 3396 4647 3407 4667
rect 3427 4647 3445 4667
rect 3396 4637 3445 4647
rect 3495 4663 3539 4679
rect 3495 4643 3510 4663
rect 3530 4643 3539 4663
rect 3495 4637 3539 4643
rect 3609 4663 3653 4679
rect 3609 4643 3618 4663
rect 3638 4643 3653 4663
rect 3609 4637 3653 4643
rect 3703 4667 3752 4679
rect 3703 4647 3721 4667
rect 3741 4647 3752 4667
rect 3703 4637 3752 4647
rect 3827 4663 3871 4679
rect 3827 4643 3836 4663
rect 3856 4643 3871 4663
rect 3827 4637 3871 4643
rect 3921 4667 3970 4679
rect 3921 4647 3939 4667
rect 3959 4647 3970 4667
rect 3921 4637 3970 4647
rect 7760 4680 7809 4692
rect 7760 4660 7771 4680
rect 7791 4660 7809 4680
rect 7760 4650 7809 4660
rect 7859 4676 7903 4692
rect 7859 4656 7874 4676
rect 7894 4656 7903 4676
rect 7859 4650 7903 4656
rect 7973 4676 8017 4692
rect 7973 4656 7982 4676
rect 8002 4656 8017 4676
rect 7973 4650 8017 4656
rect 8067 4680 8116 4692
rect 8067 4660 8085 4680
rect 8105 4660 8116 4680
rect 8067 4650 8116 4660
rect 8191 4676 8235 4692
rect 8191 4656 8200 4676
rect 8220 4656 8235 4676
rect 8191 4650 8235 4656
rect 8285 4680 8334 4692
rect 8285 4660 8303 4680
rect 8323 4660 8334 4680
rect 8285 4650 8334 4660
rect 12137 4692 12186 4704
rect 12137 4672 12148 4692
rect 12168 4672 12186 4692
rect 12137 4662 12186 4672
rect 12236 4688 12280 4704
rect 12236 4668 12251 4688
rect 12271 4668 12280 4688
rect 12236 4662 12280 4668
rect 12350 4688 12394 4704
rect 12350 4668 12359 4688
rect 12379 4668 12394 4688
rect 12350 4662 12394 4668
rect 12444 4692 12493 4704
rect 12444 4672 12462 4692
rect 12482 4672 12493 4692
rect 12444 4662 12493 4672
rect 12568 4688 12612 4704
rect 12568 4668 12577 4688
rect 12597 4668 12612 4688
rect 12568 4662 12612 4668
rect 12662 4692 12711 4704
rect 12662 4672 12680 4692
rect 12700 4672 12711 4692
rect 12662 4662 12711 4672
rect 16501 4705 16550 4717
rect 2599 4439 2648 4451
rect 1445 4427 1494 4437
rect 1445 4407 1456 4427
rect 1476 4407 1494 4427
rect 1445 4395 1494 4407
rect 1544 4431 1588 4437
rect 1544 4411 1559 4431
rect 1579 4411 1588 4431
rect 1544 4395 1588 4411
rect 1663 4427 1712 4437
rect 1663 4407 1674 4427
rect 1694 4407 1712 4427
rect 1663 4395 1712 4407
rect 1762 4431 1806 4437
rect 1762 4411 1777 4431
rect 1797 4411 1806 4431
rect 1762 4395 1806 4411
rect 1876 4431 1920 4437
rect 1876 4411 1885 4431
rect 1905 4411 1920 4431
rect 1876 4395 1920 4411
rect 1970 4427 2019 4437
rect 1970 4407 1988 4427
rect 2008 4407 2019 4427
rect 2599 4419 2610 4439
rect 2630 4419 2648 4439
rect 2599 4409 2648 4419
rect 2698 4435 2742 4451
rect 2698 4415 2713 4435
rect 2733 4415 2742 4435
rect 2698 4409 2742 4415
rect 2812 4435 2856 4451
rect 2812 4415 2821 4435
rect 2841 4415 2856 4435
rect 2812 4409 2856 4415
rect 2906 4439 2955 4451
rect 2906 4419 2924 4439
rect 2944 4419 2955 4439
rect 2906 4409 2955 4419
rect 3030 4435 3074 4451
rect 3030 4415 3039 4435
rect 3059 4415 3074 4435
rect 3030 4409 3074 4415
rect 3124 4439 3173 4451
rect 3124 4419 3142 4439
rect 3162 4419 3173 4439
rect 3124 4409 3173 4419
rect 16501 4685 16512 4705
rect 16532 4685 16550 4705
rect 16501 4675 16550 4685
rect 16600 4701 16644 4717
rect 16600 4681 16615 4701
rect 16635 4681 16644 4701
rect 16600 4675 16644 4681
rect 16714 4701 16758 4717
rect 16714 4681 16723 4701
rect 16743 4681 16758 4701
rect 16714 4675 16758 4681
rect 16808 4705 16857 4717
rect 16808 4685 16826 4705
rect 16846 4685 16857 4705
rect 16808 4675 16857 4685
rect 16932 4701 16976 4717
rect 16932 4681 16941 4701
rect 16961 4681 16976 4701
rect 16932 4675 16976 4681
rect 17026 4705 17075 4717
rect 17026 4685 17044 4705
rect 17064 4685 17075 4705
rect 17026 4675 17075 4685
rect 6963 4452 7012 4464
rect 5809 4440 5858 4450
rect 5809 4420 5820 4440
rect 5840 4420 5858 4440
rect 1970 4395 2019 4407
rect 5809 4408 5858 4420
rect 5908 4444 5952 4450
rect 5908 4424 5923 4444
rect 5943 4424 5952 4444
rect 5908 4408 5952 4424
rect 6027 4440 6076 4450
rect 6027 4420 6038 4440
rect 6058 4420 6076 4440
rect 6027 4408 6076 4420
rect 6126 4444 6170 4450
rect 6126 4424 6141 4444
rect 6161 4424 6170 4444
rect 6126 4408 6170 4424
rect 6240 4444 6284 4450
rect 6240 4424 6249 4444
rect 6269 4424 6284 4444
rect 6240 4408 6284 4424
rect 6334 4440 6383 4450
rect 6334 4420 6352 4440
rect 6372 4420 6383 4440
rect 6963 4432 6974 4452
rect 6994 4432 7012 4452
rect 6963 4422 7012 4432
rect 7062 4448 7106 4464
rect 7062 4428 7077 4448
rect 7097 4428 7106 4448
rect 7062 4422 7106 4428
rect 7176 4448 7220 4464
rect 7176 4428 7185 4448
rect 7205 4428 7220 4448
rect 7176 4422 7220 4428
rect 7270 4452 7319 4464
rect 7270 4432 7288 4452
rect 7308 4432 7319 4452
rect 7270 4422 7319 4432
rect 7394 4448 7438 4464
rect 7394 4428 7403 4448
rect 7423 4428 7438 4448
rect 7394 4422 7438 4428
rect 7488 4452 7537 4464
rect 7488 4432 7506 4452
rect 7526 4432 7537 4452
rect 7488 4422 7537 4432
rect 11340 4464 11389 4476
rect 10186 4452 10235 4462
rect 10186 4432 10197 4452
rect 10217 4432 10235 4452
rect 6334 4408 6383 4420
rect 10186 4420 10235 4432
rect 10285 4456 10329 4462
rect 10285 4436 10300 4456
rect 10320 4436 10329 4456
rect 10285 4420 10329 4436
rect 10404 4452 10453 4462
rect 10404 4432 10415 4452
rect 10435 4432 10453 4452
rect 10404 4420 10453 4432
rect 10503 4456 10547 4462
rect 10503 4436 10518 4456
rect 10538 4436 10547 4456
rect 10503 4420 10547 4436
rect 10617 4456 10661 4462
rect 10617 4436 10626 4456
rect 10646 4436 10661 4456
rect 10617 4420 10661 4436
rect 10711 4452 10760 4462
rect 10711 4432 10729 4452
rect 10749 4432 10760 4452
rect 11340 4444 11351 4464
rect 11371 4444 11389 4464
rect 11340 4434 11389 4444
rect 11439 4460 11483 4476
rect 11439 4440 11454 4460
rect 11474 4440 11483 4460
rect 11439 4434 11483 4440
rect 11553 4460 11597 4476
rect 11553 4440 11562 4460
rect 11582 4440 11597 4460
rect 11553 4434 11597 4440
rect 11647 4464 11696 4476
rect 11647 4444 11665 4464
rect 11685 4444 11696 4464
rect 11647 4434 11696 4444
rect 11771 4460 11815 4476
rect 11771 4440 11780 4460
rect 11800 4440 11815 4460
rect 11771 4434 11815 4440
rect 11865 4464 11914 4476
rect 11865 4444 11883 4464
rect 11903 4444 11914 4464
rect 11865 4434 11914 4444
rect 15704 4477 15753 4489
rect 14550 4465 14599 4475
rect 14550 4445 14561 4465
rect 14581 4445 14599 4465
rect 10711 4420 10760 4432
rect 3397 4255 3446 4267
rect 3397 4235 3408 4255
rect 3428 4235 3446 4255
rect 343 4205 392 4215
rect 343 4185 354 4205
rect 374 4185 392 4205
rect 343 4173 392 4185
rect 442 4209 486 4215
rect 442 4189 457 4209
rect 477 4189 486 4209
rect 442 4173 486 4189
rect 561 4205 610 4215
rect 561 4185 572 4205
rect 592 4185 610 4205
rect 561 4173 610 4185
rect 660 4209 704 4215
rect 660 4189 675 4209
rect 695 4189 704 4209
rect 660 4173 704 4189
rect 774 4209 818 4215
rect 774 4189 783 4209
rect 803 4189 818 4209
rect 774 4173 818 4189
rect 868 4205 917 4215
rect 3397 4225 3446 4235
rect 3496 4251 3540 4267
rect 3496 4231 3511 4251
rect 3531 4231 3540 4251
rect 3496 4225 3540 4231
rect 3610 4251 3654 4267
rect 3610 4231 3619 4251
rect 3639 4231 3654 4251
rect 3610 4225 3654 4231
rect 3704 4255 3753 4267
rect 3704 4235 3722 4255
rect 3742 4235 3753 4255
rect 3704 4225 3753 4235
rect 3828 4251 3872 4267
rect 3828 4231 3837 4251
rect 3857 4231 3872 4251
rect 3828 4225 3872 4231
rect 3922 4255 3971 4267
rect 3922 4235 3940 4255
rect 3960 4235 3971 4255
rect 3922 4225 3971 4235
rect 868 4185 886 4205
rect 906 4185 917 4205
rect 868 4173 917 4185
rect 14550 4433 14599 4445
rect 14649 4469 14693 4475
rect 14649 4449 14664 4469
rect 14684 4449 14693 4469
rect 14649 4433 14693 4449
rect 14768 4465 14817 4475
rect 14768 4445 14779 4465
rect 14799 4445 14817 4465
rect 14768 4433 14817 4445
rect 14867 4469 14911 4475
rect 14867 4449 14882 4469
rect 14902 4449 14911 4469
rect 14867 4433 14911 4449
rect 14981 4469 15025 4475
rect 14981 4449 14990 4469
rect 15010 4449 15025 4469
rect 14981 4433 15025 4449
rect 15075 4465 15124 4475
rect 15075 4445 15093 4465
rect 15113 4445 15124 4465
rect 15704 4457 15715 4477
rect 15735 4457 15753 4477
rect 15704 4447 15753 4457
rect 15803 4473 15847 4489
rect 15803 4453 15818 4473
rect 15838 4453 15847 4473
rect 15803 4447 15847 4453
rect 15917 4473 15961 4489
rect 15917 4453 15926 4473
rect 15946 4453 15961 4473
rect 15917 4447 15961 4453
rect 16011 4477 16060 4489
rect 16011 4457 16029 4477
rect 16049 4457 16060 4477
rect 16011 4447 16060 4457
rect 16135 4473 16179 4489
rect 16135 4453 16144 4473
rect 16164 4453 16179 4473
rect 16135 4447 16179 4453
rect 16229 4477 16278 4489
rect 16229 4457 16247 4477
rect 16267 4457 16278 4477
rect 16229 4447 16278 4457
rect 15075 4433 15124 4445
rect 7761 4268 7810 4280
rect 7761 4248 7772 4268
rect 7792 4248 7810 4268
rect 4707 4218 4756 4228
rect 4707 4198 4718 4218
rect 4738 4198 4756 4218
rect 4707 4186 4756 4198
rect 4806 4222 4850 4228
rect 4806 4202 4821 4222
rect 4841 4202 4850 4222
rect 4806 4186 4850 4202
rect 4925 4218 4974 4228
rect 4925 4198 4936 4218
rect 4956 4198 4974 4218
rect 4925 4186 4974 4198
rect 5024 4222 5068 4228
rect 5024 4202 5039 4222
rect 5059 4202 5068 4222
rect 5024 4186 5068 4202
rect 5138 4222 5182 4228
rect 5138 4202 5147 4222
rect 5167 4202 5182 4222
rect 5138 4186 5182 4202
rect 5232 4218 5281 4228
rect 7761 4238 7810 4248
rect 7860 4264 7904 4280
rect 7860 4244 7875 4264
rect 7895 4244 7904 4264
rect 7860 4238 7904 4244
rect 7974 4264 8018 4280
rect 7974 4244 7983 4264
rect 8003 4244 8018 4264
rect 7974 4238 8018 4244
rect 8068 4268 8117 4280
rect 8068 4248 8086 4268
rect 8106 4248 8117 4268
rect 8068 4238 8117 4248
rect 8192 4264 8236 4280
rect 8192 4244 8201 4264
rect 8221 4244 8236 4264
rect 8192 4238 8236 4244
rect 8286 4268 8335 4280
rect 8286 4248 8304 4268
rect 8324 4248 8335 4268
rect 8286 4238 8335 4248
rect 5232 4198 5250 4218
rect 5270 4198 5281 4218
rect 5232 4186 5281 4198
rect 12138 4280 12187 4292
rect 12138 4260 12149 4280
rect 12169 4260 12187 4280
rect 9084 4230 9133 4240
rect 9084 4210 9095 4230
rect 9115 4210 9133 4230
rect 9084 4198 9133 4210
rect 9183 4234 9227 4240
rect 9183 4214 9198 4234
rect 9218 4214 9227 4234
rect 9183 4198 9227 4214
rect 9302 4230 9351 4240
rect 9302 4210 9313 4230
rect 9333 4210 9351 4230
rect 9302 4198 9351 4210
rect 9401 4234 9445 4240
rect 9401 4214 9416 4234
rect 9436 4214 9445 4234
rect 9401 4198 9445 4214
rect 9515 4234 9559 4240
rect 9515 4214 9524 4234
rect 9544 4214 9559 4234
rect 9515 4198 9559 4214
rect 9609 4230 9658 4240
rect 12138 4250 12187 4260
rect 12237 4276 12281 4292
rect 12237 4256 12252 4276
rect 12272 4256 12281 4276
rect 12237 4250 12281 4256
rect 12351 4276 12395 4292
rect 12351 4256 12360 4276
rect 12380 4256 12395 4276
rect 12351 4250 12395 4256
rect 12445 4280 12494 4292
rect 12445 4260 12463 4280
rect 12483 4260 12494 4280
rect 12445 4250 12494 4260
rect 12569 4276 12613 4292
rect 12569 4256 12578 4276
rect 12598 4256 12613 4276
rect 12569 4250 12613 4256
rect 12663 4280 12712 4292
rect 12663 4260 12681 4280
rect 12701 4260 12712 4280
rect 12663 4250 12712 4260
rect 9609 4210 9627 4230
rect 9647 4210 9658 4230
rect 9609 4198 9658 4210
rect 1141 4021 1190 4031
rect 1141 4001 1152 4021
rect 1172 4001 1190 4021
rect 1141 3989 1190 4001
rect 1240 4025 1284 4031
rect 1240 4005 1255 4025
rect 1275 4005 1284 4025
rect 1240 3989 1284 4005
rect 1359 4021 1408 4031
rect 1359 4001 1370 4021
rect 1390 4001 1408 4021
rect 1359 3989 1408 4001
rect 1458 4025 1502 4031
rect 1458 4005 1473 4025
rect 1493 4005 1502 4025
rect 1458 3989 1502 4005
rect 1572 4025 1616 4031
rect 1572 4005 1581 4025
rect 1601 4005 1616 4025
rect 1572 3989 1616 4005
rect 1666 4021 1715 4031
rect 1666 4001 1684 4021
rect 1704 4001 1715 4021
rect 1666 3989 1715 4001
rect 2500 4029 2549 4041
rect 2500 4009 2511 4029
rect 2531 4009 2549 4029
rect 2500 3999 2549 4009
rect 2599 4025 2643 4041
rect 2599 4005 2614 4025
rect 2634 4005 2643 4025
rect 2599 3999 2643 4005
rect 2713 4025 2757 4041
rect 2713 4005 2722 4025
rect 2742 4005 2757 4025
rect 2713 3999 2757 4005
rect 2807 4029 2856 4041
rect 2807 4009 2825 4029
rect 2845 4009 2856 4029
rect 2807 3999 2856 4009
rect 2931 4025 2975 4041
rect 2931 4005 2940 4025
rect 2960 4005 2975 4025
rect 2931 3999 2975 4005
rect 3025 4029 3074 4041
rect 16502 4293 16551 4305
rect 16502 4273 16513 4293
rect 16533 4273 16551 4293
rect 13448 4243 13497 4253
rect 13448 4223 13459 4243
rect 13479 4223 13497 4243
rect 13448 4211 13497 4223
rect 13547 4247 13591 4253
rect 13547 4227 13562 4247
rect 13582 4227 13591 4247
rect 13547 4211 13591 4227
rect 13666 4243 13715 4253
rect 13666 4223 13677 4243
rect 13697 4223 13715 4243
rect 13666 4211 13715 4223
rect 13765 4247 13809 4253
rect 13765 4227 13780 4247
rect 13800 4227 13809 4247
rect 13765 4211 13809 4227
rect 13879 4247 13923 4253
rect 13879 4227 13888 4247
rect 13908 4227 13923 4247
rect 13879 4211 13923 4227
rect 13973 4243 14022 4253
rect 16502 4263 16551 4273
rect 16601 4289 16645 4305
rect 16601 4269 16616 4289
rect 16636 4269 16645 4289
rect 16601 4263 16645 4269
rect 16715 4289 16759 4305
rect 16715 4269 16724 4289
rect 16744 4269 16759 4289
rect 16715 4263 16759 4269
rect 16809 4293 16858 4305
rect 16809 4273 16827 4293
rect 16847 4273 16858 4293
rect 16809 4263 16858 4273
rect 16933 4289 16977 4305
rect 16933 4269 16942 4289
rect 16962 4269 16977 4289
rect 16933 4263 16977 4269
rect 17027 4293 17076 4305
rect 17027 4273 17045 4293
rect 17065 4273 17076 4293
rect 17027 4263 17076 4273
rect 13973 4223 13991 4243
rect 14011 4223 14022 4243
rect 13973 4211 14022 4223
rect 3025 4009 3043 4029
rect 3063 4009 3074 4029
rect 3025 3999 3074 4009
rect 5505 4034 5554 4044
rect 5505 4014 5516 4034
rect 5536 4014 5554 4034
rect 5505 4002 5554 4014
rect 5604 4038 5648 4044
rect 5604 4018 5619 4038
rect 5639 4018 5648 4038
rect 5604 4002 5648 4018
rect 5723 4034 5772 4044
rect 5723 4014 5734 4034
rect 5754 4014 5772 4034
rect 5723 4002 5772 4014
rect 5822 4038 5866 4044
rect 5822 4018 5837 4038
rect 5857 4018 5866 4038
rect 5822 4002 5866 4018
rect 5936 4038 5980 4044
rect 5936 4018 5945 4038
rect 5965 4018 5980 4038
rect 5936 4002 5980 4018
rect 6030 4034 6079 4044
rect 6030 4014 6048 4034
rect 6068 4014 6079 4034
rect 6030 4002 6079 4014
rect 6864 4042 6913 4054
rect 6864 4022 6875 4042
rect 6895 4022 6913 4042
rect 6864 4012 6913 4022
rect 6963 4038 7007 4054
rect 6963 4018 6978 4038
rect 6998 4018 7007 4038
rect 6963 4012 7007 4018
rect 7077 4038 7121 4054
rect 7077 4018 7086 4038
rect 7106 4018 7121 4038
rect 7077 4012 7121 4018
rect 7171 4042 7220 4054
rect 7171 4022 7189 4042
rect 7209 4022 7220 4042
rect 7171 4012 7220 4022
rect 7295 4038 7339 4054
rect 7295 4018 7304 4038
rect 7324 4018 7339 4038
rect 7295 4012 7339 4018
rect 7389 4042 7438 4054
rect 7389 4022 7407 4042
rect 7427 4022 7438 4042
rect 7389 4012 7438 4022
rect 9882 4046 9931 4056
rect 9882 4026 9893 4046
rect 9913 4026 9931 4046
rect 9882 4014 9931 4026
rect 9981 4050 10025 4056
rect 9981 4030 9996 4050
rect 10016 4030 10025 4050
rect 9981 4014 10025 4030
rect 10100 4046 10149 4056
rect 10100 4026 10111 4046
rect 10131 4026 10149 4046
rect 10100 4014 10149 4026
rect 10199 4050 10243 4056
rect 10199 4030 10214 4050
rect 10234 4030 10243 4050
rect 10199 4014 10243 4030
rect 10313 4050 10357 4056
rect 10313 4030 10322 4050
rect 10342 4030 10357 4050
rect 10313 4014 10357 4030
rect 10407 4046 10456 4056
rect 10407 4026 10425 4046
rect 10445 4026 10456 4046
rect 10407 4014 10456 4026
rect 11241 4054 11290 4066
rect 11241 4034 11252 4054
rect 11272 4034 11290 4054
rect 11241 4024 11290 4034
rect 11340 4050 11384 4066
rect 11340 4030 11355 4050
rect 11375 4030 11384 4050
rect 11340 4024 11384 4030
rect 11454 4050 11498 4066
rect 11454 4030 11463 4050
rect 11483 4030 11498 4050
rect 11454 4024 11498 4030
rect 11548 4054 11597 4066
rect 11548 4034 11566 4054
rect 11586 4034 11597 4054
rect 11548 4024 11597 4034
rect 11672 4050 11716 4066
rect 11672 4030 11681 4050
rect 11701 4030 11716 4050
rect 11672 4024 11716 4030
rect 11766 4054 11815 4066
rect 11766 4034 11784 4054
rect 11804 4034 11815 4054
rect 11766 4024 11815 4034
rect 14246 4059 14295 4069
rect 14246 4039 14257 4059
rect 14277 4039 14295 4059
rect 344 3793 393 3803
rect 344 3773 355 3793
rect 375 3773 393 3793
rect 344 3761 393 3773
rect 443 3797 487 3803
rect 443 3777 458 3797
rect 478 3777 487 3797
rect 443 3761 487 3777
rect 562 3793 611 3803
rect 562 3773 573 3793
rect 593 3773 611 3793
rect 562 3761 611 3773
rect 661 3797 705 3803
rect 661 3777 676 3797
rect 696 3777 705 3797
rect 661 3761 705 3777
rect 775 3797 819 3803
rect 775 3777 784 3797
rect 804 3777 819 3797
rect 775 3761 819 3777
rect 869 3793 918 3803
rect 869 3773 887 3793
rect 907 3773 918 3793
rect 14246 4027 14295 4039
rect 14345 4063 14389 4069
rect 14345 4043 14360 4063
rect 14380 4043 14389 4063
rect 14345 4027 14389 4043
rect 14464 4059 14513 4069
rect 14464 4039 14475 4059
rect 14495 4039 14513 4059
rect 14464 4027 14513 4039
rect 14563 4063 14607 4069
rect 14563 4043 14578 4063
rect 14598 4043 14607 4063
rect 14563 4027 14607 4043
rect 14677 4063 14721 4069
rect 14677 4043 14686 4063
rect 14706 4043 14721 4063
rect 14677 4027 14721 4043
rect 14771 4059 14820 4069
rect 14771 4039 14789 4059
rect 14809 4039 14820 4059
rect 14771 4027 14820 4039
rect 15605 4067 15654 4079
rect 15605 4047 15616 4067
rect 15636 4047 15654 4067
rect 15605 4037 15654 4047
rect 15704 4063 15748 4079
rect 15704 4043 15719 4063
rect 15739 4043 15748 4063
rect 15704 4037 15748 4043
rect 15818 4063 15862 4079
rect 15818 4043 15827 4063
rect 15847 4043 15862 4063
rect 15818 4037 15862 4043
rect 15912 4067 15961 4079
rect 15912 4047 15930 4067
rect 15950 4047 15961 4067
rect 15912 4037 15961 4047
rect 16036 4063 16080 4079
rect 16036 4043 16045 4063
rect 16065 4043 16080 4063
rect 16036 4037 16080 4043
rect 16130 4067 16179 4079
rect 16130 4047 16148 4067
rect 16168 4047 16179 4067
rect 16130 4037 16179 4047
rect 869 3761 918 3773
rect 4708 3806 4757 3816
rect 4708 3786 4719 3806
rect 4739 3786 4757 3806
rect 4708 3774 4757 3786
rect 4807 3810 4851 3816
rect 4807 3790 4822 3810
rect 4842 3790 4851 3810
rect 4807 3774 4851 3790
rect 4926 3806 4975 3816
rect 4926 3786 4937 3806
rect 4957 3786 4975 3806
rect 4926 3774 4975 3786
rect 5025 3810 5069 3816
rect 5025 3790 5040 3810
rect 5060 3790 5069 3810
rect 5025 3774 5069 3790
rect 5139 3810 5183 3816
rect 5139 3790 5148 3810
rect 5168 3790 5183 3810
rect 5139 3774 5183 3790
rect 5233 3806 5282 3816
rect 5233 3786 5251 3806
rect 5271 3786 5282 3806
rect 5233 3774 5282 3786
rect 9085 3818 9134 3828
rect 9085 3798 9096 3818
rect 9116 3798 9134 3818
rect 9085 3786 9134 3798
rect 9184 3822 9228 3828
rect 9184 3802 9199 3822
rect 9219 3802 9228 3822
rect 9184 3786 9228 3802
rect 9303 3818 9352 3828
rect 9303 3798 9314 3818
rect 9334 3798 9352 3818
rect 9303 3786 9352 3798
rect 9402 3822 9446 3828
rect 9402 3802 9417 3822
rect 9437 3802 9446 3822
rect 9402 3786 9446 3802
rect 9516 3822 9560 3828
rect 9516 3802 9525 3822
rect 9545 3802 9560 3822
rect 9516 3786 9560 3802
rect 9610 3818 9659 3828
rect 9610 3798 9628 3818
rect 9648 3798 9659 3818
rect 9610 3786 9659 3798
rect 13449 3831 13498 3841
rect 13449 3811 13460 3831
rect 13480 3811 13498 3831
rect 13449 3799 13498 3811
rect 13548 3835 13592 3841
rect 13548 3815 13563 3835
rect 13583 3815 13592 3835
rect 13548 3799 13592 3815
rect 13667 3831 13716 3841
rect 13667 3811 13678 3831
rect 13698 3811 13716 3831
rect 13667 3799 13716 3811
rect 13766 3835 13810 3841
rect 13766 3815 13781 3835
rect 13801 3815 13810 3835
rect 13766 3799 13810 3815
rect 13880 3835 13924 3841
rect 13880 3815 13889 3835
rect 13909 3815 13924 3835
rect 13880 3799 13924 3815
rect 13974 3831 14023 3841
rect 13974 3811 13992 3831
rect 14012 3811 14023 3831
rect 13974 3799 14023 3811
rect 3379 3649 3428 3661
rect 3379 3629 3390 3649
rect 3410 3629 3428 3649
rect 3379 3619 3428 3629
rect 3478 3645 3522 3661
rect 3478 3625 3493 3645
rect 3513 3625 3522 3645
rect 3478 3619 3522 3625
rect 3592 3645 3636 3661
rect 3592 3625 3601 3645
rect 3621 3625 3636 3645
rect 3592 3619 3636 3625
rect 3686 3649 3735 3661
rect 3686 3629 3704 3649
rect 3724 3629 3735 3649
rect 3686 3619 3735 3629
rect 3810 3645 3854 3661
rect 3810 3625 3819 3645
rect 3839 3625 3854 3645
rect 3810 3619 3854 3625
rect 3904 3649 3953 3661
rect 3904 3629 3922 3649
rect 3942 3629 3953 3649
rect 3904 3619 3953 3629
rect 7743 3662 7792 3674
rect 7743 3642 7754 3662
rect 7774 3642 7792 3662
rect 7743 3632 7792 3642
rect 7842 3658 7886 3674
rect 7842 3638 7857 3658
rect 7877 3638 7886 3658
rect 7842 3632 7886 3638
rect 7956 3658 8000 3674
rect 7956 3638 7965 3658
rect 7985 3638 8000 3658
rect 7956 3632 8000 3638
rect 8050 3662 8099 3674
rect 8050 3642 8068 3662
rect 8088 3642 8099 3662
rect 8050 3632 8099 3642
rect 8174 3658 8218 3674
rect 8174 3638 8183 3658
rect 8203 3638 8218 3658
rect 8174 3632 8218 3638
rect 8268 3662 8317 3674
rect 8268 3642 8286 3662
rect 8306 3642 8317 3662
rect 8268 3632 8317 3642
rect 12120 3674 12169 3686
rect 12120 3654 12131 3674
rect 12151 3654 12169 3674
rect 12120 3644 12169 3654
rect 12219 3670 12263 3686
rect 12219 3650 12234 3670
rect 12254 3650 12263 3670
rect 12219 3644 12263 3650
rect 12333 3670 12377 3686
rect 12333 3650 12342 3670
rect 12362 3650 12377 3670
rect 12333 3644 12377 3650
rect 12427 3674 12476 3686
rect 12427 3654 12445 3674
rect 12465 3654 12476 3674
rect 12427 3644 12476 3654
rect 12551 3670 12595 3686
rect 12551 3650 12560 3670
rect 12580 3650 12595 3670
rect 12551 3644 12595 3650
rect 12645 3674 12694 3686
rect 12645 3654 12663 3674
rect 12683 3654 12694 3674
rect 12645 3644 12694 3654
rect 16484 3687 16533 3699
rect 1223 3413 1272 3423
rect 1223 3393 1234 3413
rect 1254 3393 1272 3413
rect 1223 3381 1272 3393
rect 1322 3417 1366 3423
rect 1322 3397 1337 3417
rect 1357 3397 1366 3417
rect 1322 3381 1366 3397
rect 1441 3413 1490 3423
rect 1441 3393 1452 3413
rect 1472 3393 1490 3413
rect 1441 3381 1490 3393
rect 1540 3417 1584 3423
rect 1540 3397 1555 3417
rect 1575 3397 1584 3417
rect 1540 3381 1584 3397
rect 1654 3417 1698 3423
rect 1654 3397 1663 3417
rect 1683 3397 1698 3417
rect 1654 3381 1698 3397
rect 1748 3413 1797 3423
rect 1748 3393 1766 3413
rect 1786 3393 1797 3413
rect 1748 3381 1797 3393
rect 2582 3421 2631 3433
rect 2582 3401 2593 3421
rect 2613 3401 2631 3421
rect 2582 3391 2631 3401
rect 2681 3417 2725 3433
rect 2681 3397 2696 3417
rect 2716 3397 2725 3417
rect 2681 3391 2725 3397
rect 2795 3417 2839 3433
rect 2795 3397 2804 3417
rect 2824 3397 2839 3417
rect 2795 3391 2839 3397
rect 2889 3421 2938 3433
rect 2889 3401 2907 3421
rect 2927 3401 2938 3421
rect 2889 3391 2938 3401
rect 3013 3417 3057 3433
rect 3013 3397 3022 3417
rect 3042 3397 3057 3417
rect 3013 3391 3057 3397
rect 3107 3421 3156 3433
rect 16484 3667 16495 3687
rect 16515 3667 16533 3687
rect 16484 3657 16533 3667
rect 16583 3683 16627 3699
rect 16583 3663 16598 3683
rect 16618 3663 16627 3683
rect 16583 3657 16627 3663
rect 16697 3683 16741 3699
rect 16697 3663 16706 3683
rect 16726 3663 16741 3683
rect 16697 3657 16741 3663
rect 16791 3687 16840 3699
rect 16791 3667 16809 3687
rect 16829 3667 16840 3687
rect 16791 3657 16840 3667
rect 16915 3683 16959 3699
rect 16915 3663 16924 3683
rect 16944 3663 16959 3683
rect 16915 3657 16959 3663
rect 17009 3687 17058 3699
rect 17009 3667 17027 3687
rect 17047 3667 17058 3687
rect 17009 3657 17058 3667
rect 3107 3401 3125 3421
rect 3145 3401 3156 3421
rect 3107 3391 3156 3401
rect 5587 3426 5636 3436
rect 5587 3406 5598 3426
rect 5618 3406 5636 3426
rect 5587 3394 5636 3406
rect 5686 3430 5730 3436
rect 5686 3410 5701 3430
rect 5721 3410 5730 3430
rect 5686 3394 5730 3410
rect 5805 3426 5854 3436
rect 5805 3406 5816 3426
rect 5836 3406 5854 3426
rect 5805 3394 5854 3406
rect 5904 3430 5948 3436
rect 5904 3410 5919 3430
rect 5939 3410 5948 3430
rect 5904 3394 5948 3410
rect 6018 3430 6062 3436
rect 6018 3410 6027 3430
rect 6047 3410 6062 3430
rect 6018 3394 6062 3410
rect 6112 3426 6161 3436
rect 6112 3406 6130 3426
rect 6150 3406 6161 3426
rect 6112 3394 6161 3406
rect 6946 3434 6995 3446
rect 6946 3414 6957 3434
rect 6977 3414 6995 3434
rect 6946 3404 6995 3414
rect 7045 3430 7089 3446
rect 7045 3410 7060 3430
rect 7080 3410 7089 3430
rect 7045 3404 7089 3410
rect 7159 3430 7203 3446
rect 7159 3410 7168 3430
rect 7188 3410 7203 3430
rect 7159 3404 7203 3410
rect 7253 3434 7302 3446
rect 7253 3414 7271 3434
rect 7291 3414 7302 3434
rect 7253 3404 7302 3414
rect 7377 3430 7421 3446
rect 7377 3410 7386 3430
rect 7406 3410 7421 3430
rect 7377 3404 7421 3410
rect 7471 3434 7520 3446
rect 7471 3414 7489 3434
rect 7509 3414 7520 3434
rect 7471 3404 7520 3414
rect 9964 3438 10013 3448
rect 9964 3418 9975 3438
rect 9995 3418 10013 3438
rect 9964 3406 10013 3418
rect 10063 3442 10107 3448
rect 10063 3422 10078 3442
rect 10098 3422 10107 3442
rect 10063 3406 10107 3422
rect 10182 3438 10231 3448
rect 10182 3418 10193 3438
rect 10213 3418 10231 3438
rect 10182 3406 10231 3418
rect 10281 3442 10325 3448
rect 10281 3422 10296 3442
rect 10316 3422 10325 3442
rect 10281 3406 10325 3422
rect 10395 3442 10439 3448
rect 10395 3422 10404 3442
rect 10424 3422 10439 3442
rect 10395 3406 10439 3422
rect 10489 3438 10538 3448
rect 10489 3418 10507 3438
rect 10527 3418 10538 3438
rect 10489 3406 10538 3418
rect 11323 3446 11372 3458
rect 11323 3426 11334 3446
rect 11354 3426 11372 3446
rect 11323 3416 11372 3426
rect 11422 3442 11466 3458
rect 11422 3422 11437 3442
rect 11457 3422 11466 3442
rect 11422 3416 11466 3422
rect 11536 3442 11580 3458
rect 11536 3422 11545 3442
rect 11565 3422 11580 3442
rect 11536 3416 11580 3422
rect 11630 3446 11679 3458
rect 11630 3426 11648 3446
rect 11668 3426 11679 3446
rect 11630 3416 11679 3426
rect 11754 3442 11798 3458
rect 11754 3422 11763 3442
rect 11783 3422 11798 3442
rect 11754 3416 11798 3422
rect 11848 3446 11897 3458
rect 11848 3426 11866 3446
rect 11886 3426 11897 3446
rect 11848 3416 11897 3426
rect 14328 3451 14377 3461
rect 14328 3431 14339 3451
rect 14359 3431 14377 3451
rect 3380 3237 3429 3249
rect 3380 3217 3391 3237
rect 3411 3217 3429 3237
rect 326 3187 375 3197
rect 326 3167 337 3187
rect 357 3167 375 3187
rect 326 3155 375 3167
rect 425 3191 469 3197
rect 425 3171 440 3191
rect 460 3171 469 3191
rect 425 3155 469 3171
rect 544 3187 593 3197
rect 544 3167 555 3187
rect 575 3167 593 3187
rect 544 3155 593 3167
rect 643 3191 687 3197
rect 643 3171 658 3191
rect 678 3171 687 3191
rect 643 3155 687 3171
rect 757 3191 801 3197
rect 757 3171 766 3191
rect 786 3171 801 3191
rect 757 3155 801 3171
rect 851 3187 900 3197
rect 3380 3207 3429 3217
rect 3479 3233 3523 3249
rect 3479 3213 3494 3233
rect 3514 3213 3523 3233
rect 3479 3207 3523 3213
rect 3593 3233 3637 3249
rect 3593 3213 3602 3233
rect 3622 3213 3637 3233
rect 3593 3207 3637 3213
rect 3687 3237 3736 3249
rect 3687 3217 3705 3237
rect 3725 3217 3736 3237
rect 3687 3207 3736 3217
rect 3811 3233 3855 3249
rect 3811 3213 3820 3233
rect 3840 3213 3855 3233
rect 3811 3207 3855 3213
rect 3905 3237 3954 3249
rect 3905 3217 3923 3237
rect 3943 3217 3954 3237
rect 3905 3207 3954 3217
rect 851 3167 869 3187
rect 889 3167 900 3187
rect 851 3155 900 3167
rect 14328 3419 14377 3431
rect 14427 3455 14471 3461
rect 14427 3435 14442 3455
rect 14462 3435 14471 3455
rect 14427 3419 14471 3435
rect 14546 3451 14595 3461
rect 14546 3431 14557 3451
rect 14577 3431 14595 3451
rect 14546 3419 14595 3431
rect 14645 3455 14689 3461
rect 14645 3435 14660 3455
rect 14680 3435 14689 3455
rect 14645 3419 14689 3435
rect 14759 3455 14803 3461
rect 14759 3435 14768 3455
rect 14788 3435 14803 3455
rect 14759 3419 14803 3435
rect 14853 3451 14902 3461
rect 14853 3431 14871 3451
rect 14891 3431 14902 3451
rect 14853 3419 14902 3431
rect 15687 3459 15736 3471
rect 15687 3439 15698 3459
rect 15718 3439 15736 3459
rect 15687 3429 15736 3439
rect 15786 3455 15830 3471
rect 15786 3435 15801 3455
rect 15821 3435 15830 3455
rect 15786 3429 15830 3435
rect 15900 3455 15944 3471
rect 15900 3435 15909 3455
rect 15929 3435 15944 3455
rect 15900 3429 15944 3435
rect 15994 3459 16043 3471
rect 15994 3439 16012 3459
rect 16032 3439 16043 3459
rect 15994 3429 16043 3439
rect 16118 3455 16162 3471
rect 16118 3435 16127 3455
rect 16147 3435 16162 3455
rect 16118 3429 16162 3435
rect 16212 3459 16261 3471
rect 16212 3439 16230 3459
rect 16250 3439 16261 3459
rect 16212 3429 16261 3439
rect 7744 3250 7793 3262
rect 7744 3230 7755 3250
rect 7775 3230 7793 3250
rect 4690 3200 4739 3210
rect 4690 3180 4701 3200
rect 4721 3180 4739 3200
rect 4690 3168 4739 3180
rect 4789 3204 4833 3210
rect 4789 3184 4804 3204
rect 4824 3184 4833 3204
rect 4789 3168 4833 3184
rect 4908 3200 4957 3210
rect 4908 3180 4919 3200
rect 4939 3180 4957 3200
rect 4908 3168 4957 3180
rect 5007 3204 5051 3210
rect 5007 3184 5022 3204
rect 5042 3184 5051 3204
rect 5007 3168 5051 3184
rect 5121 3204 5165 3210
rect 5121 3184 5130 3204
rect 5150 3184 5165 3204
rect 5121 3168 5165 3184
rect 5215 3200 5264 3210
rect 7744 3220 7793 3230
rect 7843 3246 7887 3262
rect 7843 3226 7858 3246
rect 7878 3226 7887 3246
rect 7843 3220 7887 3226
rect 7957 3246 8001 3262
rect 7957 3226 7966 3246
rect 7986 3226 8001 3246
rect 7957 3220 8001 3226
rect 8051 3250 8100 3262
rect 8051 3230 8069 3250
rect 8089 3230 8100 3250
rect 8051 3220 8100 3230
rect 8175 3246 8219 3262
rect 8175 3226 8184 3246
rect 8204 3226 8219 3246
rect 8175 3220 8219 3226
rect 8269 3250 8318 3262
rect 8269 3230 8287 3250
rect 8307 3230 8318 3250
rect 8269 3220 8318 3230
rect 5215 3180 5233 3200
rect 5253 3180 5264 3200
rect 5215 3168 5264 3180
rect 12121 3262 12170 3274
rect 12121 3242 12132 3262
rect 12152 3242 12170 3262
rect 9067 3212 9116 3222
rect 9067 3192 9078 3212
rect 9098 3192 9116 3212
rect 9067 3180 9116 3192
rect 9166 3216 9210 3222
rect 9166 3196 9181 3216
rect 9201 3196 9210 3216
rect 9166 3180 9210 3196
rect 9285 3212 9334 3222
rect 9285 3192 9296 3212
rect 9316 3192 9334 3212
rect 9285 3180 9334 3192
rect 9384 3216 9428 3222
rect 9384 3196 9399 3216
rect 9419 3196 9428 3216
rect 9384 3180 9428 3196
rect 9498 3216 9542 3222
rect 9498 3196 9507 3216
rect 9527 3196 9542 3216
rect 9498 3180 9542 3196
rect 9592 3212 9641 3222
rect 12121 3232 12170 3242
rect 12220 3258 12264 3274
rect 12220 3238 12235 3258
rect 12255 3238 12264 3258
rect 12220 3232 12264 3238
rect 12334 3258 12378 3274
rect 12334 3238 12343 3258
rect 12363 3238 12378 3258
rect 12334 3232 12378 3238
rect 12428 3262 12477 3274
rect 12428 3242 12446 3262
rect 12466 3242 12477 3262
rect 12428 3232 12477 3242
rect 12552 3258 12596 3274
rect 12552 3238 12561 3258
rect 12581 3238 12596 3258
rect 12552 3232 12596 3238
rect 12646 3262 12695 3274
rect 12646 3242 12664 3262
rect 12684 3242 12695 3262
rect 12646 3232 12695 3242
rect 9592 3192 9610 3212
rect 9630 3192 9641 3212
rect 9592 3180 9641 3192
rect 2417 3013 2466 3025
rect 1124 3003 1173 3013
rect 1124 2983 1135 3003
rect 1155 2983 1173 3003
rect 1124 2971 1173 2983
rect 1223 3007 1267 3013
rect 1223 2987 1238 3007
rect 1258 2987 1267 3007
rect 1223 2971 1267 2987
rect 1342 3003 1391 3013
rect 1342 2983 1353 3003
rect 1373 2983 1391 3003
rect 1342 2971 1391 2983
rect 1441 3007 1485 3013
rect 1441 2987 1456 3007
rect 1476 2987 1485 3007
rect 1441 2971 1485 2987
rect 1555 3007 1599 3013
rect 1555 2987 1564 3007
rect 1584 2987 1599 3007
rect 1555 2971 1599 2987
rect 1649 3003 1698 3013
rect 1649 2983 1667 3003
rect 1687 2983 1698 3003
rect 2417 2993 2428 3013
rect 2448 2993 2466 3013
rect 2417 2983 2466 2993
rect 2516 3009 2560 3025
rect 2516 2989 2531 3009
rect 2551 2989 2560 3009
rect 2516 2983 2560 2989
rect 2630 3009 2674 3025
rect 2630 2989 2639 3009
rect 2659 2989 2674 3009
rect 2630 2983 2674 2989
rect 2724 3013 2773 3025
rect 2724 2993 2742 3013
rect 2762 2993 2773 3013
rect 2724 2983 2773 2993
rect 2848 3009 2892 3025
rect 2848 2989 2857 3009
rect 2877 2989 2892 3009
rect 2848 2983 2892 2989
rect 2942 3013 2991 3025
rect 16485 3275 16534 3287
rect 16485 3255 16496 3275
rect 16516 3255 16534 3275
rect 13431 3225 13480 3235
rect 13431 3205 13442 3225
rect 13462 3205 13480 3225
rect 13431 3193 13480 3205
rect 13530 3229 13574 3235
rect 13530 3209 13545 3229
rect 13565 3209 13574 3229
rect 13530 3193 13574 3209
rect 13649 3225 13698 3235
rect 13649 3205 13660 3225
rect 13680 3205 13698 3225
rect 13649 3193 13698 3205
rect 13748 3229 13792 3235
rect 13748 3209 13763 3229
rect 13783 3209 13792 3229
rect 13748 3193 13792 3209
rect 13862 3229 13906 3235
rect 13862 3209 13871 3229
rect 13891 3209 13906 3229
rect 13862 3193 13906 3209
rect 13956 3225 14005 3235
rect 16485 3245 16534 3255
rect 16584 3271 16628 3287
rect 16584 3251 16599 3271
rect 16619 3251 16628 3271
rect 16584 3245 16628 3251
rect 16698 3271 16742 3287
rect 16698 3251 16707 3271
rect 16727 3251 16742 3271
rect 16698 3245 16742 3251
rect 16792 3275 16841 3287
rect 16792 3255 16810 3275
rect 16830 3255 16841 3275
rect 16792 3245 16841 3255
rect 16916 3271 16960 3287
rect 16916 3251 16925 3271
rect 16945 3251 16960 3271
rect 16916 3245 16960 3251
rect 17010 3275 17059 3287
rect 17010 3255 17028 3275
rect 17048 3255 17059 3275
rect 17010 3245 17059 3255
rect 13956 3205 13974 3225
rect 13994 3205 14005 3225
rect 13956 3193 14005 3205
rect 6781 3026 6830 3038
rect 2942 2993 2960 3013
rect 2980 2993 2991 3013
rect 2942 2983 2991 2993
rect 1649 2971 1698 2983
rect 5488 3016 5537 3026
rect 5488 2996 5499 3016
rect 5519 2996 5537 3016
rect 5488 2984 5537 2996
rect 5587 3020 5631 3026
rect 5587 3000 5602 3020
rect 5622 3000 5631 3020
rect 5587 2984 5631 3000
rect 5706 3016 5755 3026
rect 5706 2996 5717 3016
rect 5737 2996 5755 3016
rect 5706 2984 5755 2996
rect 5805 3020 5849 3026
rect 5805 3000 5820 3020
rect 5840 3000 5849 3020
rect 5805 2984 5849 3000
rect 5919 3020 5963 3026
rect 5919 3000 5928 3020
rect 5948 3000 5963 3020
rect 5919 2984 5963 3000
rect 6013 3016 6062 3026
rect 6013 2996 6031 3016
rect 6051 2996 6062 3016
rect 6781 3006 6792 3026
rect 6812 3006 6830 3026
rect 6781 2996 6830 3006
rect 6880 3022 6924 3038
rect 6880 3002 6895 3022
rect 6915 3002 6924 3022
rect 6880 2996 6924 3002
rect 6994 3022 7038 3038
rect 6994 3002 7003 3022
rect 7023 3002 7038 3022
rect 6994 2996 7038 3002
rect 7088 3026 7137 3038
rect 7088 3006 7106 3026
rect 7126 3006 7137 3026
rect 7088 2996 7137 3006
rect 7212 3022 7256 3038
rect 7212 3002 7221 3022
rect 7241 3002 7256 3022
rect 7212 2996 7256 3002
rect 7306 3026 7355 3038
rect 11158 3038 11207 3050
rect 7306 3006 7324 3026
rect 7344 3006 7355 3026
rect 7306 2996 7355 3006
rect 6013 2984 6062 2996
rect 9865 3028 9914 3038
rect 9865 3008 9876 3028
rect 9896 3008 9914 3028
rect 9865 2996 9914 3008
rect 9964 3032 10008 3038
rect 9964 3012 9979 3032
rect 9999 3012 10008 3032
rect 9964 2996 10008 3012
rect 10083 3028 10132 3038
rect 10083 3008 10094 3028
rect 10114 3008 10132 3028
rect 10083 2996 10132 3008
rect 10182 3032 10226 3038
rect 10182 3012 10197 3032
rect 10217 3012 10226 3032
rect 10182 2996 10226 3012
rect 10296 3032 10340 3038
rect 10296 3012 10305 3032
rect 10325 3012 10340 3032
rect 10296 2996 10340 3012
rect 10390 3028 10439 3038
rect 10390 3008 10408 3028
rect 10428 3008 10439 3028
rect 11158 3018 11169 3038
rect 11189 3018 11207 3038
rect 11158 3008 11207 3018
rect 11257 3034 11301 3050
rect 11257 3014 11272 3034
rect 11292 3014 11301 3034
rect 11257 3008 11301 3014
rect 11371 3034 11415 3050
rect 11371 3014 11380 3034
rect 11400 3014 11415 3034
rect 11371 3008 11415 3014
rect 11465 3038 11514 3050
rect 11465 3018 11483 3038
rect 11503 3018 11514 3038
rect 11465 3008 11514 3018
rect 11589 3034 11633 3050
rect 11589 3014 11598 3034
rect 11618 3014 11633 3034
rect 11589 3008 11633 3014
rect 11683 3038 11732 3050
rect 15522 3051 15571 3063
rect 11683 3018 11701 3038
rect 11721 3018 11732 3038
rect 11683 3008 11732 3018
rect 10390 2996 10439 3008
rect 327 2775 376 2785
rect 327 2755 338 2775
rect 358 2755 376 2775
rect 327 2743 376 2755
rect 426 2779 470 2785
rect 426 2759 441 2779
rect 461 2759 470 2779
rect 426 2743 470 2759
rect 545 2775 594 2785
rect 545 2755 556 2775
rect 576 2755 594 2775
rect 545 2743 594 2755
rect 644 2779 688 2785
rect 644 2759 659 2779
rect 679 2759 688 2779
rect 644 2743 688 2759
rect 758 2779 802 2785
rect 758 2759 767 2779
rect 787 2759 802 2779
rect 758 2743 802 2759
rect 852 2775 901 2785
rect 852 2755 870 2775
rect 890 2755 901 2775
rect 14229 3041 14278 3051
rect 14229 3021 14240 3041
rect 14260 3021 14278 3041
rect 14229 3009 14278 3021
rect 14328 3045 14372 3051
rect 14328 3025 14343 3045
rect 14363 3025 14372 3045
rect 14328 3009 14372 3025
rect 14447 3041 14496 3051
rect 14447 3021 14458 3041
rect 14478 3021 14496 3041
rect 14447 3009 14496 3021
rect 14546 3045 14590 3051
rect 14546 3025 14561 3045
rect 14581 3025 14590 3045
rect 14546 3009 14590 3025
rect 14660 3045 14704 3051
rect 14660 3025 14669 3045
rect 14689 3025 14704 3045
rect 14660 3009 14704 3025
rect 14754 3041 14803 3051
rect 14754 3021 14772 3041
rect 14792 3021 14803 3041
rect 15522 3031 15533 3051
rect 15553 3031 15571 3051
rect 15522 3021 15571 3031
rect 15621 3047 15665 3063
rect 15621 3027 15636 3047
rect 15656 3027 15665 3047
rect 15621 3021 15665 3027
rect 15735 3047 15779 3063
rect 15735 3027 15744 3047
rect 15764 3027 15779 3047
rect 15735 3021 15779 3027
rect 15829 3051 15878 3063
rect 15829 3031 15847 3051
rect 15867 3031 15878 3051
rect 15829 3021 15878 3031
rect 15953 3047 15997 3063
rect 15953 3027 15962 3047
rect 15982 3027 15997 3047
rect 15953 3021 15997 3027
rect 16047 3051 16096 3063
rect 16047 3031 16065 3051
rect 16085 3031 16096 3051
rect 16047 3021 16096 3031
rect 14754 3009 14803 3021
rect 852 2743 901 2755
rect 4691 2788 4740 2798
rect 4691 2768 4702 2788
rect 4722 2768 4740 2788
rect 4691 2756 4740 2768
rect 4790 2792 4834 2798
rect 4790 2772 4805 2792
rect 4825 2772 4834 2792
rect 4790 2756 4834 2772
rect 4909 2788 4958 2798
rect 4909 2768 4920 2788
rect 4940 2768 4958 2788
rect 4909 2756 4958 2768
rect 5008 2792 5052 2798
rect 5008 2772 5023 2792
rect 5043 2772 5052 2792
rect 5008 2756 5052 2772
rect 5122 2792 5166 2798
rect 5122 2772 5131 2792
rect 5151 2772 5166 2792
rect 5122 2756 5166 2772
rect 5216 2788 5265 2798
rect 5216 2768 5234 2788
rect 5254 2768 5265 2788
rect 5216 2756 5265 2768
rect 9068 2800 9117 2810
rect 9068 2780 9079 2800
rect 9099 2780 9117 2800
rect 9068 2768 9117 2780
rect 9167 2804 9211 2810
rect 9167 2784 9182 2804
rect 9202 2784 9211 2804
rect 9167 2768 9211 2784
rect 9286 2800 9335 2810
rect 9286 2780 9297 2800
rect 9317 2780 9335 2800
rect 9286 2768 9335 2780
rect 9385 2804 9429 2810
rect 9385 2784 9400 2804
rect 9420 2784 9429 2804
rect 9385 2768 9429 2784
rect 9499 2804 9543 2810
rect 9499 2784 9508 2804
rect 9528 2784 9543 2804
rect 9499 2768 9543 2784
rect 9593 2800 9642 2810
rect 9593 2780 9611 2800
rect 9631 2780 9642 2800
rect 9593 2768 9642 2780
rect 13432 2813 13481 2823
rect 13432 2793 13443 2813
rect 13463 2793 13481 2813
rect 13432 2781 13481 2793
rect 13531 2817 13575 2823
rect 13531 2797 13546 2817
rect 13566 2797 13575 2817
rect 13531 2781 13575 2797
rect 13650 2813 13699 2823
rect 13650 2793 13661 2813
rect 13681 2793 13699 2813
rect 13650 2781 13699 2793
rect 13749 2817 13793 2823
rect 13749 2797 13764 2817
rect 13784 2797 13793 2817
rect 13749 2781 13793 2797
rect 13863 2817 13907 2823
rect 13863 2797 13872 2817
rect 13892 2797 13907 2817
rect 13863 2781 13907 2797
rect 13957 2813 14006 2823
rect 13957 2793 13975 2813
rect 13995 2793 14006 2813
rect 13957 2781 14006 2793
rect 3359 2631 3408 2643
rect 3359 2611 3370 2631
rect 3390 2611 3408 2631
rect 3359 2601 3408 2611
rect 3458 2627 3502 2643
rect 3458 2607 3473 2627
rect 3493 2607 3502 2627
rect 3458 2601 3502 2607
rect 3572 2627 3616 2643
rect 3572 2607 3581 2627
rect 3601 2607 3616 2627
rect 3572 2601 3616 2607
rect 3666 2631 3715 2643
rect 3666 2611 3684 2631
rect 3704 2611 3715 2631
rect 3666 2601 3715 2611
rect 3790 2627 3834 2643
rect 3790 2607 3799 2627
rect 3819 2607 3834 2627
rect 3790 2601 3834 2607
rect 3884 2631 3933 2643
rect 3884 2611 3902 2631
rect 3922 2611 3933 2631
rect 3884 2601 3933 2611
rect 7723 2644 7772 2656
rect 7723 2624 7734 2644
rect 7754 2624 7772 2644
rect 7723 2614 7772 2624
rect 7822 2640 7866 2656
rect 7822 2620 7837 2640
rect 7857 2620 7866 2640
rect 7822 2614 7866 2620
rect 7936 2640 7980 2656
rect 7936 2620 7945 2640
rect 7965 2620 7980 2640
rect 7936 2614 7980 2620
rect 8030 2644 8079 2656
rect 8030 2624 8048 2644
rect 8068 2624 8079 2644
rect 8030 2614 8079 2624
rect 8154 2640 8198 2656
rect 8154 2620 8163 2640
rect 8183 2620 8198 2640
rect 8154 2614 8198 2620
rect 8248 2644 8297 2656
rect 8248 2624 8266 2644
rect 8286 2624 8297 2644
rect 8248 2614 8297 2624
rect 12100 2656 12149 2668
rect 12100 2636 12111 2656
rect 12131 2636 12149 2656
rect 12100 2626 12149 2636
rect 12199 2652 12243 2668
rect 12199 2632 12214 2652
rect 12234 2632 12243 2652
rect 12199 2626 12243 2632
rect 12313 2652 12357 2668
rect 12313 2632 12322 2652
rect 12342 2632 12357 2652
rect 12313 2626 12357 2632
rect 12407 2656 12456 2668
rect 12407 2636 12425 2656
rect 12445 2636 12456 2656
rect 12407 2626 12456 2636
rect 12531 2652 12575 2668
rect 12531 2632 12540 2652
rect 12560 2632 12575 2652
rect 12531 2626 12575 2632
rect 12625 2656 12674 2668
rect 12625 2636 12643 2656
rect 12663 2636 12674 2656
rect 12625 2626 12674 2636
rect 16464 2669 16513 2681
rect 2562 2403 2611 2415
rect 1269 2393 1318 2403
rect 1269 2373 1280 2393
rect 1300 2373 1318 2393
rect 1269 2361 1318 2373
rect 1368 2397 1412 2403
rect 1368 2377 1383 2397
rect 1403 2377 1412 2397
rect 1368 2361 1412 2377
rect 1487 2393 1536 2403
rect 1487 2373 1498 2393
rect 1518 2373 1536 2393
rect 1487 2361 1536 2373
rect 1586 2397 1630 2403
rect 1586 2377 1601 2397
rect 1621 2377 1630 2397
rect 1586 2361 1630 2377
rect 1700 2397 1744 2403
rect 1700 2377 1709 2397
rect 1729 2377 1744 2397
rect 1700 2361 1744 2377
rect 1794 2393 1843 2403
rect 1794 2373 1812 2393
rect 1832 2373 1843 2393
rect 2562 2383 2573 2403
rect 2593 2383 2611 2403
rect 2562 2373 2611 2383
rect 2661 2399 2705 2415
rect 2661 2379 2676 2399
rect 2696 2379 2705 2399
rect 2661 2373 2705 2379
rect 2775 2399 2819 2415
rect 2775 2379 2784 2399
rect 2804 2379 2819 2399
rect 2775 2373 2819 2379
rect 2869 2403 2918 2415
rect 2869 2383 2887 2403
rect 2907 2383 2918 2403
rect 2869 2373 2918 2383
rect 2993 2399 3037 2415
rect 2993 2379 3002 2399
rect 3022 2379 3037 2399
rect 2993 2373 3037 2379
rect 3087 2403 3136 2415
rect 3087 2383 3105 2403
rect 3125 2383 3136 2403
rect 3087 2373 3136 2383
rect 16464 2649 16475 2669
rect 16495 2649 16513 2669
rect 16464 2639 16513 2649
rect 16563 2665 16607 2681
rect 16563 2645 16578 2665
rect 16598 2645 16607 2665
rect 16563 2639 16607 2645
rect 16677 2665 16721 2681
rect 16677 2645 16686 2665
rect 16706 2645 16721 2665
rect 16677 2639 16721 2645
rect 16771 2669 16820 2681
rect 16771 2649 16789 2669
rect 16809 2649 16820 2669
rect 16771 2639 16820 2649
rect 16895 2665 16939 2681
rect 16895 2645 16904 2665
rect 16924 2645 16939 2665
rect 16895 2639 16939 2645
rect 16989 2669 17038 2681
rect 16989 2649 17007 2669
rect 17027 2649 17038 2669
rect 16989 2639 17038 2649
rect 6926 2416 6975 2428
rect 5633 2406 5682 2416
rect 5633 2386 5644 2406
rect 5664 2386 5682 2406
rect 1794 2361 1843 2373
rect 5633 2374 5682 2386
rect 5732 2410 5776 2416
rect 5732 2390 5747 2410
rect 5767 2390 5776 2410
rect 5732 2374 5776 2390
rect 5851 2406 5900 2416
rect 5851 2386 5862 2406
rect 5882 2386 5900 2406
rect 5851 2374 5900 2386
rect 5950 2410 5994 2416
rect 5950 2390 5965 2410
rect 5985 2390 5994 2410
rect 5950 2374 5994 2390
rect 6064 2410 6108 2416
rect 6064 2390 6073 2410
rect 6093 2390 6108 2410
rect 6064 2374 6108 2390
rect 6158 2406 6207 2416
rect 6158 2386 6176 2406
rect 6196 2386 6207 2406
rect 6926 2396 6937 2416
rect 6957 2396 6975 2416
rect 6926 2386 6975 2396
rect 7025 2412 7069 2428
rect 7025 2392 7040 2412
rect 7060 2392 7069 2412
rect 7025 2386 7069 2392
rect 7139 2412 7183 2428
rect 7139 2392 7148 2412
rect 7168 2392 7183 2412
rect 7139 2386 7183 2392
rect 7233 2416 7282 2428
rect 7233 2396 7251 2416
rect 7271 2396 7282 2416
rect 7233 2386 7282 2396
rect 7357 2412 7401 2428
rect 7357 2392 7366 2412
rect 7386 2392 7401 2412
rect 7357 2386 7401 2392
rect 7451 2416 7500 2428
rect 7451 2396 7469 2416
rect 7489 2396 7500 2416
rect 7451 2386 7500 2396
rect 11303 2428 11352 2440
rect 10010 2418 10059 2428
rect 10010 2398 10021 2418
rect 10041 2398 10059 2418
rect 6158 2374 6207 2386
rect 10010 2386 10059 2398
rect 10109 2422 10153 2428
rect 10109 2402 10124 2422
rect 10144 2402 10153 2422
rect 10109 2386 10153 2402
rect 10228 2418 10277 2428
rect 10228 2398 10239 2418
rect 10259 2398 10277 2418
rect 10228 2386 10277 2398
rect 10327 2422 10371 2428
rect 10327 2402 10342 2422
rect 10362 2402 10371 2422
rect 10327 2386 10371 2402
rect 10441 2422 10485 2428
rect 10441 2402 10450 2422
rect 10470 2402 10485 2422
rect 10441 2386 10485 2402
rect 10535 2418 10584 2428
rect 10535 2398 10553 2418
rect 10573 2398 10584 2418
rect 11303 2408 11314 2428
rect 11334 2408 11352 2428
rect 11303 2398 11352 2408
rect 11402 2424 11446 2440
rect 11402 2404 11417 2424
rect 11437 2404 11446 2424
rect 11402 2398 11446 2404
rect 11516 2424 11560 2440
rect 11516 2404 11525 2424
rect 11545 2404 11560 2424
rect 11516 2398 11560 2404
rect 11610 2428 11659 2440
rect 11610 2408 11628 2428
rect 11648 2408 11659 2428
rect 11610 2398 11659 2408
rect 11734 2424 11778 2440
rect 11734 2404 11743 2424
rect 11763 2404 11778 2424
rect 11734 2398 11778 2404
rect 11828 2428 11877 2440
rect 11828 2408 11846 2428
rect 11866 2408 11877 2428
rect 11828 2398 11877 2408
rect 15667 2441 15716 2453
rect 14374 2431 14423 2441
rect 14374 2411 14385 2431
rect 14405 2411 14423 2431
rect 10535 2386 10584 2398
rect 3360 2219 3409 2231
rect 3360 2199 3371 2219
rect 3391 2199 3409 2219
rect 306 2169 355 2179
rect 306 2149 317 2169
rect 337 2149 355 2169
rect 306 2137 355 2149
rect 405 2173 449 2179
rect 405 2153 420 2173
rect 440 2153 449 2173
rect 405 2137 449 2153
rect 524 2169 573 2179
rect 524 2149 535 2169
rect 555 2149 573 2169
rect 524 2137 573 2149
rect 623 2173 667 2179
rect 623 2153 638 2173
rect 658 2153 667 2173
rect 623 2137 667 2153
rect 737 2173 781 2179
rect 737 2153 746 2173
rect 766 2153 781 2173
rect 737 2137 781 2153
rect 831 2169 880 2179
rect 3360 2189 3409 2199
rect 3459 2215 3503 2231
rect 3459 2195 3474 2215
rect 3494 2195 3503 2215
rect 3459 2189 3503 2195
rect 3573 2215 3617 2231
rect 3573 2195 3582 2215
rect 3602 2195 3617 2215
rect 3573 2189 3617 2195
rect 3667 2219 3716 2231
rect 3667 2199 3685 2219
rect 3705 2199 3716 2219
rect 3667 2189 3716 2199
rect 3791 2215 3835 2231
rect 3791 2195 3800 2215
rect 3820 2195 3835 2215
rect 3791 2189 3835 2195
rect 3885 2219 3934 2231
rect 3885 2199 3903 2219
rect 3923 2199 3934 2219
rect 3885 2189 3934 2199
rect 831 2149 849 2169
rect 869 2149 880 2169
rect 831 2137 880 2149
rect 14374 2399 14423 2411
rect 14473 2435 14517 2441
rect 14473 2415 14488 2435
rect 14508 2415 14517 2435
rect 14473 2399 14517 2415
rect 14592 2431 14641 2441
rect 14592 2411 14603 2431
rect 14623 2411 14641 2431
rect 14592 2399 14641 2411
rect 14691 2435 14735 2441
rect 14691 2415 14706 2435
rect 14726 2415 14735 2435
rect 14691 2399 14735 2415
rect 14805 2435 14849 2441
rect 14805 2415 14814 2435
rect 14834 2415 14849 2435
rect 14805 2399 14849 2415
rect 14899 2431 14948 2441
rect 14899 2411 14917 2431
rect 14937 2411 14948 2431
rect 15667 2421 15678 2441
rect 15698 2421 15716 2441
rect 15667 2411 15716 2421
rect 15766 2437 15810 2453
rect 15766 2417 15781 2437
rect 15801 2417 15810 2437
rect 15766 2411 15810 2417
rect 15880 2437 15924 2453
rect 15880 2417 15889 2437
rect 15909 2417 15924 2437
rect 15880 2411 15924 2417
rect 15974 2441 16023 2453
rect 15974 2421 15992 2441
rect 16012 2421 16023 2441
rect 15974 2411 16023 2421
rect 16098 2437 16142 2453
rect 16098 2417 16107 2437
rect 16127 2417 16142 2437
rect 16098 2411 16142 2417
rect 16192 2441 16241 2453
rect 16192 2421 16210 2441
rect 16230 2421 16241 2441
rect 16192 2411 16241 2421
rect 14899 2399 14948 2411
rect 7724 2232 7773 2244
rect 7724 2212 7735 2232
rect 7755 2212 7773 2232
rect 4670 2182 4719 2192
rect 4670 2162 4681 2182
rect 4701 2162 4719 2182
rect 4670 2150 4719 2162
rect 4769 2186 4813 2192
rect 4769 2166 4784 2186
rect 4804 2166 4813 2186
rect 4769 2150 4813 2166
rect 4888 2182 4937 2192
rect 4888 2162 4899 2182
rect 4919 2162 4937 2182
rect 4888 2150 4937 2162
rect 4987 2186 5031 2192
rect 4987 2166 5002 2186
rect 5022 2166 5031 2186
rect 4987 2150 5031 2166
rect 5101 2186 5145 2192
rect 5101 2166 5110 2186
rect 5130 2166 5145 2186
rect 5101 2150 5145 2166
rect 5195 2182 5244 2192
rect 7724 2202 7773 2212
rect 7823 2228 7867 2244
rect 7823 2208 7838 2228
rect 7858 2208 7867 2228
rect 7823 2202 7867 2208
rect 7937 2228 7981 2244
rect 7937 2208 7946 2228
rect 7966 2208 7981 2228
rect 7937 2202 7981 2208
rect 8031 2232 8080 2244
rect 8031 2212 8049 2232
rect 8069 2212 8080 2232
rect 8031 2202 8080 2212
rect 8155 2228 8199 2244
rect 8155 2208 8164 2228
rect 8184 2208 8199 2228
rect 8155 2202 8199 2208
rect 8249 2232 8298 2244
rect 8249 2212 8267 2232
rect 8287 2212 8298 2232
rect 8249 2202 8298 2212
rect 5195 2162 5213 2182
rect 5233 2162 5244 2182
rect 5195 2150 5244 2162
rect 12101 2244 12150 2256
rect 12101 2224 12112 2244
rect 12132 2224 12150 2244
rect 9047 2194 9096 2204
rect 9047 2174 9058 2194
rect 9078 2174 9096 2194
rect 9047 2162 9096 2174
rect 9146 2198 9190 2204
rect 9146 2178 9161 2198
rect 9181 2178 9190 2198
rect 9146 2162 9190 2178
rect 9265 2194 9314 2204
rect 9265 2174 9276 2194
rect 9296 2174 9314 2194
rect 9265 2162 9314 2174
rect 9364 2198 9408 2204
rect 9364 2178 9379 2198
rect 9399 2178 9408 2198
rect 9364 2162 9408 2178
rect 9478 2198 9522 2204
rect 9478 2178 9487 2198
rect 9507 2178 9522 2198
rect 9478 2162 9522 2178
rect 9572 2194 9621 2204
rect 12101 2214 12150 2224
rect 12200 2240 12244 2256
rect 12200 2220 12215 2240
rect 12235 2220 12244 2240
rect 12200 2214 12244 2220
rect 12314 2240 12358 2256
rect 12314 2220 12323 2240
rect 12343 2220 12358 2240
rect 12314 2214 12358 2220
rect 12408 2244 12457 2256
rect 12408 2224 12426 2244
rect 12446 2224 12457 2244
rect 12408 2214 12457 2224
rect 12532 2240 12576 2256
rect 12532 2220 12541 2240
rect 12561 2220 12576 2240
rect 12532 2214 12576 2220
rect 12626 2244 12675 2256
rect 12626 2224 12644 2244
rect 12664 2224 12675 2244
rect 12626 2214 12675 2224
rect 9572 2174 9590 2194
rect 9610 2174 9621 2194
rect 9572 2162 9621 2174
rect 1104 1985 1153 1995
rect 1104 1965 1115 1985
rect 1135 1965 1153 1985
rect 1104 1953 1153 1965
rect 1203 1989 1247 1995
rect 1203 1969 1218 1989
rect 1238 1969 1247 1989
rect 1203 1953 1247 1969
rect 1322 1985 1371 1995
rect 1322 1965 1333 1985
rect 1353 1965 1371 1985
rect 1322 1953 1371 1965
rect 1421 1989 1465 1995
rect 1421 1969 1436 1989
rect 1456 1969 1465 1989
rect 1421 1953 1465 1969
rect 1535 1989 1579 1995
rect 1535 1969 1544 1989
rect 1564 1969 1579 1989
rect 1535 1953 1579 1969
rect 1629 1985 1678 1995
rect 1629 1965 1647 1985
rect 1667 1965 1678 1985
rect 1629 1953 1678 1965
rect 2463 1993 2512 2005
rect 2463 1973 2474 1993
rect 2494 1973 2512 1993
rect 2463 1963 2512 1973
rect 2562 1989 2606 2005
rect 2562 1969 2577 1989
rect 2597 1969 2606 1989
rect 2562 1963 2606 1969
rect 2676 1989 2720 2005
rect 2676 1969 2685 1989
rect 2705 1969 2720 1989
rect 2676 1963 2720 1969
rect 2770 1993 2819 2005
rect 2770 1973 2788 1993
rect 2808 1973 2819 1993
rect 2770 1963 2819 1973
rect 2894 1989 2938 2005
rect 2894 1969 2903 1989
rect 2923 1969 2938 1989
rect 2894 1963 2938 1969
rect 2988 1993 3037 2005
rect 16465 2257 16514 2269
rect 16465 2237 16476 2257
rect 16496 2237 16514 2257
rect 13411 2207 13460 2217
rect 13411 2187 13422 2207
rect 13442 2187 13460 2207
rect 13411 2175 13460 2187
rect 13510 2211 13554 2217
rect 13510 2191 13525 2211
rect 13545 2191 13554 2211
rect 13510 2175 13554 2191
rect 13629 2207 13678 2217
rect 13629 2187 13640 2207
rect 13660 2187 13678 2207
rect 13629 2175 13678 2187
rect 13728 2211 13772 2217
rect 13728 2191 13743 2211
rect 13763 2191 13772 2211
rect 13728 2175 13772 2191
rect 13842 2211 13886 2217
rect 13842 2191 13851 2211
rect 13871 2191 13886 2211
rect 13842 2175 13886 2191
rect 13936 2207 13985 2217
rect 16465 2227 16514 2237
rect 16564 2253 16608 2269
rect 16564 2233 16579 2253
rect 16599 2233 16608 2253
rect 16564 2227 16608 2233
rect 16678 2253 16722 2269
rect 16678 2233 16687 2253
rect 16707 2233 16722 2253
rect 16678 2227 16722 2233
rect 16772 2257 16821 2269
rect 16772 2237 16790 2257
rect 16810 2237 16821 2257
rect 16772 2227 16821 2237
rect 16896 2253 16940 2269
rect 16896 2233 16905 2253
rect 16925 2233 16940 2253
rect 16896 2227 16940 2233
rect 16990 2257 17039 2269
rect 16990 2237 17008 2257
rect 17028 2237 17039 2257
rect 16990 2227 17039 2237
rect 13936 2187 13954 2207
rect 13974 2187 13985 2207
rect 13936 2175 13985 2187
rect 2988 1973 3006 1993
rect 3026 1973 3037 1993
rect 2988 1963 3037 1973
rect 5468 1998 5517 2008
rect 5468 1978 5479 1998
rect 5499 1978 5517 1998
rect 5468 1966 5517 1978
rect 5567 2002 5611 2008
rect 5567 1982 5582 2002
rect 5602 1982 5611 2002
rect 5567 1966 5611 1982
rect 5686 1998 5735 2008
rect 5686 1978 5697 1998
rect 5717 1978 5735 1998
rect 5686 1966 5735 1978
rect 5785 2002 5829 2008
rect 5785 1982 5800 2002
rect 5820 1982 5829 2002
rect 5785 1966 5829 1982
rect 5899 2002 5943 2008
rect 5899 1982 5908 2002
rect 5928 1982 5943 2002
rect 5899 1966 5943 1982
rect 5993 1998 6042 2008
rect 5993 1978 6011 1998
rect 6031 1978 6042 1998
rect 5993 1966 6042 1978
rect 6827 2006 6876 2018
rect 6827 1986 6838 2006
rect 6858 1986 6876 2006
rect 6827 1976 6876 1986
rect 6926 2002 6970 2018
rect 6926 1982 6941 2002
rect 6961 1982 6970 2002
rect 6926 1976 6970 1982
rect 7040 2002 7084 2018
rect 7040 1982 7049 2002
rect 7069 1982 7084 2002
rect 7040 1976 7084 1982
rect 7134 2006 7183 2018
rect 7134 1986 7152 2006
rect 7172 1986 7183 2006
rect 7134 1976 7183 1986
rect 7258 2002 7302 2018
rect 7258 1982 7267 2002
rect 7287 1982 7302 2002
rect 7258 1976 7302 1982
rect 7352 2006 7401 2018
rect 7352 1986 7370 2006
rect 7390 1986 7401 2006
rect 7352 1976 7401 1986
rect 9845 2010 9894 2020
rect 9845 1990 9856 2010
rect 9876 1990 9894 2010
rect 9845 1978 9894 1990
rect 9944 2014 9988 2020
rect 9944 1994 9959 2014
rect 9979 1994 9988 2014
rect 9944 1978 9988 1994
rect 10063 2010 10112 2020
rect 10063 1990 10074 2010
rect 10094 1990 10112 2010
rect 10063 1978 10112 1990
rect 10162 2014 10206 2020
rect 10162 1994 10177 2014
rect 10197 1994 10206 2014
rect 10162 1978 10206 1994
rect 10276 2014 10320 2020
rect 10276 1994 10285 2014
rect 10305 1994 10320 2014
rect 10276 1978 10320 1994
rect 10370 2010 10419 2020
rect 10370 1990 10388 2010
rect 10408 1990 10419 2010
rect 10370 1978 10419 1990
rect 11204 2018 11253 2030
rect 11204 1998 11215 2018
rect 11235 1998 11253 2018
rect 11204 1988 11253 1998
rect 11303 2014 11347 2030
rect 11303 1994 11318 2014
rect 11338 1994 11347 2014
rect 11303 1988 11347 1994
rect 11417 2014 11461 2030
rect 11417 1994 11426 2014
rect 11446 1994 11461 2014
rect 11417 1988 11461 1994
rect 11511 2018 11560 2030
rect 11511 1998 11529 2018
rect 11549 1998 11560 2018
rect 11511 1988 11560 1998
rect 11635 2014 11679 2030
rect 11635 1994 11644 2014
rect 11664 1994 11679 2014
rect 11635 1988 11679 1994
rect 11729 2018 11778 2030
rect 11729 1998 11747 2018
rect 11767 1998 11778 2018
rect 11729 1988 11778 1998
rect 14209 2023 14258 2033
rect 14209 2003 14220 2023
rect 14240 2003 14258 2023
rect 307 1757 356 1767
rect 307 1737 318 1757
rect 338 1737 356 1757
rect 307 1725 356 1737
rect 406 1761 450 1767
rect 406 1741 421 1761
rect 441 1741 450 1761
rect 406 1725 450 1741
rect 525 1757 574 1767
rect 525 1737 536 1757
rect 556 1737 574 1757
rect 525 1725 574 1737
rect 624 1761 668 1767
rect 624 1741 639 1761
rect 659 1741 668 1761
rect 624 1725 668 1741
rect 738 1761 782 1767
rect 738 1741 747 1761
rect 767 1741 782 1761
rect 738 1725 782 1741
rect 832 1757 881 1767
rect 832 1737 850 1757
rect 870 1737 881 1757
rect 14209 1991 14258 2003
rect 14308 2027 14352 2033
rect 14308 2007 14323 2027
rect 14343 2007 14352 2027
rect 14308 1991 14352 2007
rect 14427 2023 14476 2033
rect 14427 2003 14438 2023
rect 14458 2003 14476 2023
rect 14427 1991 14476 2003
rect 14526 2027 14570 2033
rect 14526 2007 14541 2027
rect 14561 2007 14570 2027
rect 14526 1991 14570 2007
rect 14640 2027 14684 2033
rect 14640 2007 14649 2027
rect 14669 2007 14684 2027
rect 14640 1991 14684 2007
rect 14734 2023 14783 2033
rect 14734 2003 14752 2023
rect 14772 2003 14783 2023
rect 14734 1991 14783 2003
rect 15568 2031 15617 2043
rect 15568 2011 15579 2031
rect 15599 2011 15617 2031
rect 15568 2001 15617 2011
rect 15667 2027 15711 2043
rect 15667 2007 15682 2027
rect 15702 2007 15711 2027
rect 15667 2001 15711 2007
rect 15781 2027 15825 2043
rect 15781 2007 15790 2027
rect 15810 2007 15825 2027
rect 15781 2001 15825 2007
rect 15875 2031 15924 2043
rect 15875 2011 15893 2031
rect 15913 2011 15924 2031
rect 15875 2001 15924 2011
rect 15999 2027 16043 2043
rect 15999 2007 16008 2027
rect 16028 2007 16043 2027
rect 15999 2001 16043 2007
rect 16093 2031 16142 2043
rect 16093 2011 16111 2031
rect 16131 2011 16142 2031
rect 16093 2001 16142 2011
rect 832 1725 881 1737
rect 4671 1770 4720 1780
rect 4671 1750 4682 1770
rect 4702 1750 4720 1770
rect 4671 1738 4720 1750
rect 4770 1774 4814 1780
rect 4770 1754 4785 1774
rect 4805 1754 4814 1774
rect 4770 1738 4814 1754
rect 4889 1770 4938 1780
rect 4889 1750 4900 1770
rect 4920 1750 4938 1770
rect 4889 1738 4938 1750
rect 4988 1774 5032 1780
rect 4988 1754 5003 1774
rect 5023 1754 5032 1774
rect 4988 1738 5032 1754
rect 5102 1774 5146 1780
rect 5102 1754 5111 1774
rect 5131 1754 5146 1774
rect 5102 1738 5146 1754
rect 5196 1770 5245 1780
rect 5196 1750 5214 1770
rect 5234 1750 5245 1770
rect 5196 1738 5245 1750
rect 9048 1782 9097 1792
rect 9048 1762 9059 1782
rect 9079 1762 9097 1782
rect 9048 1750 9097 1762
rect 9147 1786 9191 1792
rect 9147 1766 9162 1786
rect 9182 1766 9191 1786
rect 9147 1750 9191 1766
rect 9266 1782 9315 1792
rect 9266 1762 9277 1782
rect 9297 1762 9315 1782
rect 9266 1750 9315 1762
rect 9365 1786 9409 1792
rect 9365 1766 9380 1786
rect 9400 1766 9409 1786
rect 9365 1750 9409 1766
rect 9479 1786 9523 1792
rect 9479 1766 9488 1786
rect 9508 1766 9523 1786
rect 9479 1750 9523 1766
rect 9573 1782 9622 1792
rect 9573 1762 9591 1782
rect 9611 1762 9622 1782
rect 9573 1750 9622 1762
rect 13412 1795 13461 1805
rect 13412 1775 13423 1795
rect 13443 1775 13461 1795
rect 13412 1763 13461 1775
rect 13511 1799 13555 1805
rect 13511 1779 13526 1799
rect 13546 1779 13555 1799
rect 13511 1763 13555 1779
rect 13630 1795 13679 1805
rect 13630 1775 13641 1795
rect 13661 1775 13679 1795
rect 13630 1763 13679 1775
rect 13729 1799 13773 1805
rect 13729 1779 13744 1799
rect 13764 1779 13773 1799
rect 13729 1763 13773 1779
rect 13843 1799 13887 1805
rect 13843 1779 13852 1799
rect 13872 1779 13887 1799
rect 13843 1763 13887 1779
rect 13937 1795 13986 1805
rect 13937 1775 13955 1795
rect 13975 1775 13986 1795
rect 13937 1763 13986 1775
rect 3342 1613 3391 1625
rect 3342 1593 3353 1613
rect 3373 1593 3391 1613
rect 3342 1583 3391 1593
rect 3441 1609 3485 1625
rect 3441 1589 3456 1609
rect 3476 1589 3485 1609
rect 3441 1583 3485 1589
rect 3555 1609 3599 1625
rect 3555 1589 3564 1609
rect 3584 1589 3599 1609
rect 3555 1583 3599 1589
rect 3649 1613 3698 1625
rect 3649 1593 3667 1613
rect 3687 1593 3698 1613
rect 3649 1583 3698 1593
rect 3773 1609 3817 1625
rect 3773 1589 3782 1609
rect 3802 1589 3817 1609
rect 3773 1583 3817 1589
rect 3867 1613 3916 1625
rect 3867 1593 3885 1613
rect 3905 1593 3916 1613
rect 3867 1583 3916 1593
rect 7706 1626 7755 1638
rect 7706 1606 7717 1626
rect 7737 1606 7755 1626
rect 7706 1596 7755 1606
rect 7805 1622 7849 1638
rect 7805 1602 7820 1622
rect 7840 1602 7849 1622
rect 7805 1596 7849 1602
rect 7919 1622 7963 1638
rect 7919 1602 7928 1622
rect 7948 1602 7963 1622
rect 7919 1596 7963 1602
rect 8013 1626 8062 1638
rect 8013 1606 8031 1626
rect 8051 1606 8062 1626
rect 8013 1596 8062 1606
rect 8137 1622 8181 1638
rect 8137 1602 8146 1622
rect 8166 1602 8181 1622
rect 8137 1596 8181 1602
rect 8231 1626 8280 1638
rect 8231 1606 8249 1626
rect 8269 1606 8280 1626
rect 8231 1596 8280 1606
rect 12083 1638 12132 1650
rect 12083 1618 12094 1638
rect 12114 1618 12132 1638
rect 12083 1608 12132 1618
rect 12182 1634 12226 1650
rect 12182 1614 12197 1634
rect 12217 1614 12226 1634
rect 12182 1608 12226 1614
rect 12296 1634 12340 1650
rect 12296 1614 12305 1634
rect 12325 1614 12340 1634
rect 12296 1608 12340 1614
rect 12390 1638 12439 1650
rect 12390 1618 12408 1638
rect 12428 1618 12439 1638
rect 12390 1608 12439 1618
rect 12514 1634 12558 1650
rect 12514 1614 12523 1634
rect 12543 1614 12558 1634
rect 12514 1608 12558 1614
rect 12608 1638 12657 1650
rect 12608 1618 12626 1638
rect 12646 1618 12657 1638
rect 12608 1608 12657 1618
rect 16447 1651 16496 1663
rect 1186 1377 1235 1387
rect 1186 1357 1197 1377
rect 1217 1357 1235 1377
rect 1186 1345 1235 1357
rect 1285 1381 1329 1387
rect 1285 1361 1300 1381
rect 1320 1361 1329 1381
rect 1285 1345 1329 1361
rect 1404 1377 1453 1387
rect 1404 1357 1415 1377
rect 1435 1357 1453 1377
rect 1404 1345 1453 1357
rect 1503 1381 1547 1387
rect 1503 1361 1518 1381
rect 1538 1361 1547 1381
rect 1503 1345 1547 1361
rect 1617 1381 1661 1387
rect 1617 1361 1626 1381
rect 1646 1361 1661 1381
rect 1617 1345 1661 1361
rect 1711 1377 1760 1387
rect 1711 1357 1729 1377
rect 1749 1357 1760 1377
rect 1711 1345 1760 1357
rect 2545 1385 2594 1397
rect 2545 1365 2556 1385
rect 2576 1365 2594 1385
rect 2545 1355 2594 1365
rect 2644 1381 2688 1397
rect 2644 1361 2659 1381
rect 2679 1361 2688 1381
rect 2644 1355 2688 1361
rect 2758 1381 2802 1397
rect 2758 1361 2767 1381
rect 2787 1361 2802 1381
rect 2758 1355 2802 1361
rect 2852 1385 2901 1397
rect 2852 1365 2870 1385
rect 2890 1365 2901 1385
rect 2852 1355 2901 1365
rect 2976 1381 3020 1397
rect 2976 1361 2985 1381
rect 3005 1361 3020 1381
rect 2976 1355 3020 1361
rect 3070 1385 3119 1397
rect 16447 1631 16458 1651
rect 16478 1631 16496 1651
rect 16447 1621 16496 1631
rect 16546 1647 16590 1663
rect 16546 1627 16561 1647
rect 16581 1627 16590 1647
rect 16546 1621 16590 1627
rect 16660 1647 16704 1663
rect 16660 1627 16669 1647
rect 16689 1627 16704 1647
rect 16660 1621 16704 1627
rect 16754 1651 16803 1663
rect 16754 1631 16772 1651
rect 16792 1631 16803 1651
rect 16754 1621 16803 1631
rect 16878 1647 16922 1663
rect 16878 1627 16887 1647
rect 16907 1627 16922 1647
rect 16878 1621 16922 1627
rect 16972 1651 17021 1663
rect 16972 1631 16990 1651
rect 17010 1631 17021 1651
rect 16972 1621 17021 1631
rect 3070 1365 3088 1385
rect 3108 1365 3119 1385
rect 3070 1355 3119 1365
rect 5550 1390 5599 1400
rect 5550 1370 5561 1390
rect 5581 1370 5599 1390
rect 5550 1358 5599 1370
rect 5649 1394 5693 1400
rect 5649 1374 5664 1394
rect 5684 1374 5693 1394
rect 5649 1358 5693 1374
rect 5768 1390 5817 1400
rect 5768 1370 5779 1390
rect 5799 1370 5817 1390
rect 5768 1358 5817 1370
rect 5867 1394 5911 1400
rect 5867 1374 5882 1394
rect 5902 1374 5911 1394
rect 5867 1358 5911 1374
rect 5981 1394 6025 1400
rect 5981 1374 5990 1394
rect 6010 1374 6025 1394
rect 5981 1358 6025 1374
rect 6075 1390 6124 1400
rect 6075 1370 6093 1390
rect 6113 1370 6124 1390
rect 6075 1358 6124 1370
rect 6909 1398 6958 1410
rect 6909 1378 6920 1398
rect 6940 1378 6958 1398
rect 6909 1368 6958 1378
rect 7008 1394 7052 1410
rect 7008 1374 7023 1394
rect 7043 1374 7052 1394
rect 7008 1368 7052 1374
rect 7122 1394 7166 1410
rect 7122 1374 7131 1394
rect 7151 1374 7166 1394
rect 7122 1368 7166 1374
rect 7216 1398 7265 1410
rect 7216 1378 7234 1398
rect 7254 1378 7265 1398
rect 7216 1368 7265 1378
rect 7340 1394 7384 1410
rect 7340 1374 7349 1394
rect 7369 1374 7384 1394
rect 7340 1368 7384 1374
rect 7434 1398 7483 1410
rect 7434 1378 7452 1398
rect 7472 1378 7483 1398
rect 7434 1368 7483 1378
rect 9927 1402 9976 1412
rect 9927 1382 9938 1402
rect 9958 1382 9976 1402
rect 9927 1370 9976 1382
rect 10026 1406 10070 1412
rect 10026 1386 10041 1406
rect 10061 1386 10070 1406
rect 10026 1370 10070 1386
rect 10145 1402 10194 1412
rect 10145 1382 10156 1402
rect 10176 1382 10194 1402
rect 10145 1370 10194 1382
rect 10244 1406 10288 1412
rect 10244 1386 10259 1406
rect 10279 1386 10288 1406
rect 10244 1370 10288 1386
rect 10358 1406 10402 1412
rect 10358 1386 10367 1406
rect 10387 1386 10402 1406
rect 10358 1370 10402 1386
rect 10452 1402 10501 1412
rect 10452 1382 10470 1402
rect 10490 1382 10501 1402
rect 10452 1370 10501 1382
rect 11286 1410 11335 1422
rect 11286 1390 11297 1410
rect 11317 1390 11335 1410
rect 11286 1380 11335 1390
rect 11385 1406 11429 1422
rect 11385 1386 11400 1406
rect 11420 1386 11429 1406
rect 11385 1380 11429 1386
rect 11499 1406 11543 1422
rect 11499 1386 11508 1406
rect 11528 1386 11543 1406
rect 11499 1380 11543 1386
rect 11593 1410 11642 1422
rect 11593 1390 11611 1410
rect 11631 1390 11642 1410
rect 11593 1380 11642 1390
rect 11717 1406 11761 1422
rect 11717 1386 11726 1406
rect 11746 1386 11761 1406
rect 11717 1380 11761 1386
rect 11811 1410 11860 1422
rect 11811 1390 11829 1410
rect 11849 1390 11860 1410
rect 11811 1380 11860 1390
rect 14291 1415 14340 1425
rect 14291 1395 14302 1415
rect 14322 1395 14340 1415
rect 3343 1201 3392 1213
rect 3343 1181 3354 1201
rect 3374 1181 3392 1201
rect 289 1151 338 1161
rect 289 1131 300 1151
rect 320 1131 338 1151
rect 289 1119 338 1131
rect 388 1155 432 1161
rect 388 1135 403 1155
rect 423 1135 432 1155
rect 388 1119 432 1135
rect 507 1151 556 1161
rect 507 1131 518 1151
rect 538 1131 556 1151
rect 507 1119 556 1131
rect 606 1155 650 1161
rect 606 1135 621 1155
rect 641 1135 650 1155
rect 606 1119 650 1135
rect 720 1155 764 1161
rect 720 1135 729 1155
rect 749 1135 764 1155
rect 720 1119 764 1135
rect 814 1151 863 1161
rect 3343 1171 3392 1181
rect 3442 1197 3486 1213
rect 3442 1177 3457 1197
rect 3477 1177 3486 1197
rect 3442 1171 3486 1177
rect 3556 1197 3600 1213
rect 3556 1177 3565 1197
rect 3585 1177 3600 1197
rect 3556 1171 3600 1177
rect 3650 1201 3699 1213
rect 3650 1181 3668 1201
rect 3688 1181 3699 1201
rect 3650 1171 3699 1181
rect 3774 1197 3818 1213
rect 3774 1177 3783 1197
rect 3803 1177 3818 1197
rect 3774 1171 3818 1177
rect 3868 1201 3917 1213
rect 3868 1181 3886 1201
rect 3906 1181 3917 1201
rect 3868 1171 3917 1181
rect 814 1131 832 1151
rect 852 1131 863 1151
rect 814 1119 863 1131
rect 14291 1383 14340 1395
rect 14390 1419 14434 1425
rect 14390 1399 14405 1419
rect 14425 1399 14434 1419
rect 14390 1383 14434 1399
rect 14509 1415 14558 1425
rect 14509 1395 14520 1415
rect 14540 1395 14558 1415
rect 14509 1383 14558 1395
rect 14608 1419 14652 1425
rect 14608 1399 14623 1419
rect 14643 1399 14652 1419
rect 14608 1383 14652 1399
rect 14722 1419 14766 1425
rect 14722 1399 14731 1419
rect 14751 1399 14766 1419
rect 14722 1383 14766 1399
rect 14816 1415 14865 1425
rect 14816 1395 14834 1415
rect 14854 1395 14865 1415
rect 14816 1383 14865 1395
rect 15650 1423 15699 1435
rect 15650 1403 15661 1423
rect 15681 1403 15699 1423
rect 15650 1393 15699 1403
rect 15749 1419 15793 1435
rect 15749 1399 15764 1419
rect 15784 1399 15793 1419
rect 15749 1393 15793 1399
rect 15863 1419 15907 1435
rect 15863 1399 15872 1419
rect 15892 1399 15907 1419
rect 15863 1393 15907 1399
rect 15957 1423 16006 1435
rect 15957 1403 15975 1423
rect 15995 1403 16006 1423
rect 15957 1393 16006 1403
rect 16081 1419 16125 1435
rect 16081 1399 16090 1419
rect 16110 1399 16125 1419
rect 16081 1393 16125 1399
rect 16175 1423 16224 1435
rect 16175 1403 16193 1423
rect 16213 1403 16224 1423
rect 16175 1393 16224 1403
rect 7707 1214 7756 1226
rect 7707 1194 7718 1214
rect 7738 1194 7756 1214
rect 4653 1164 4702 1174
rect 4653 1144 4664 1164
rect 4684 1144 4702 1164
rect 4653 1132 4702 1144
rect 4752 1168 4796 1174
rect 4752 1148 4767 1168
rect 4787 1148 4796 1168
rect 4752 1132 4796 1148
rect 4871 1164 4920 1174
rect 4871 1144 4882 1164
rect 4902 1144 4920 1164
rect 4871 1132 4920 1144
rect 4970 1168 5014 1174
rect 4970 1148 4985 1168
rect 5005 1148 5014 1168
rect 4970 1132 5014 1148
rect 5084 1168 5128 1174
rect 5084 1148 5093 1168
rect 5113 1148 5128 1168
rect 5084 1132 5128 1148
rect 5178 1164 5227 1174
rect 7707 1184 7756 1194
rect 7806 1210 7850 1226
rect 7806 1190 7821 1210
rect 7841 1190 7850 1210
rect 7806 1184 7850 1190
rect 7920 1210 7964 1226
rect 7920 1190 7929 1210
rect 7949 1190 7964 1210
rect 7920 1184 7964 1190
rect 8014 1214 8063 1226
rect 8014 1194 8032 1214
rect 8052 1194 8063 1214
rect 8014 1184 8063 1194
rect 8138 1210 8182 1226
rect 8138 1190 8147 1210
rect 8167 1190 8182 1210
rect 8138 1184 8182 1190
rect 8232 1214 8281 1226
rect 8232 1194 8250 1214
rect 8270 1194 8281 1214
rect 8232 1184 8281 1194
rect 5178 1144 5196 1164
rect 5216 1144 5227 1164
rect 5178 1132 5227 1144
rect 12084 1226 12133 1238
rect 12084 1206 12095 1226
rect 12115 1206 12133 1226
rect 9030 1176 9079 1186
rect 9030 1156 9041 1176
rect 9061 1156 9079 1176
rect 9030 1144 9079 1156
rect 9129 1180 9173 1186
rect 9129 1160 9144 1180
rect 9164 1160 9173 1180
rect 9129 1144 9173 1160
rect 9248 1176 9297 1186
rect 9248 1156 9259 1176
rect 9279 1156 9297 1176
rect 9248 1144 9297 1156
rect 9347 1180 9391 1186
rect 9347 1160 9362 1180
rect 9382 1160 9391 1180
rect 9347 1144 9391 1160
rect 9461 1180 9505 1186
rect 9461 1160 9470 1180
rect 9490 1160 9505 1180
rect 9461 1144 9505 1160
rect 9555 1176 9604 1186
rect 12084 1196 12133 1206
rect 12183 1222 12227 1238
rect 12183 1202 12198 1222
rect 12218 1202 12227 1222
rect 12183 1196 12227 1202
rect 12297 1222 12341 1238
rect 12297 1202 12306 1222
rect 12326 1202 12341 1222
rect 12297 1196 12341 1202
rect 12391 1226 12440 1238
rect 12391 1206 12409 1226
rect 12429 1206 12440 1226
rect 12391 1196 12440 1206
rect 12515 1222 12559 1238
rect 12515 1202 12524 1222
rect 12544 1202 12559 1222
rect 12515 1196 12559 1202
rect 12609 1226 12658 1238
rect 12609 1206 12627 1226
rect 12647 1206 12658 1226
rect 12609 1196 12658 1206
rect 9555 1156 9573 1176
rect 9593 1156 9604 1176
rect 9555 1144 9604 1156
rect 16448 1239 16497 1251
rect 16448 1219 16459 1239
rect 16479 1219 16497 1239
rect 13394 1189 13443 1199
rect 13394 1169 13405 1189
rect 13425 1169 13443 1189
rect 13394 1157 13443 1169
rect 13493 1193 13537 1199
rect 13493 1173 13508 1193
rect 13528 1173 13537 1193
rect 13493 1157 13537 1173
rect 13612 1189 13661 1199
rect 13612 1169 13623 1189
rect 13643 1169 13661 1189
rect 13612 1157 13661 1169
rect 13711 1193 13755 1199
rect 13711 1173 13726 1193
rect 13746 1173 13755 1193
rect 13711 1157 13755 1173
rect 13825 1193 13869 1199
rect 13825 1173 13834 1193
rect 13854 1173 13869 1193
rect 13825 1157 13869 1173
rect 13919 1189 13968 1199
rect 16448 1209 16497 1219
rect 16547 1235 16591 1251
rect 16547 1215 16562 1235
rect 16582 1215 16591 1235
rect 16547 1209 16591 1215
rect 16661 1235 16705 1251
rect 16661 1215 16670 1235
rect 16690 1215 16705 1235
rect 16661 1209 16705 1215
rect 16755 1239 16804 1251
rect 16755 1219 16773 1239
rect 16793 1219 16804 1239
rect 16755 1209 16804 1219
rect 16879 1235 16923 1251
rect 16879 1215 16888 1235
rect 16908 1215 16923 1235
rect 16879 1209 16923 1215
rect 16973 1239 17022 1251
rect 16973 1219 16991 1239
rect 17011 1219 17022 1239
rect 16973 1209 17022 1219
rect 13919 1169 13937 1189
rect 13957 1169 13968 1189
rect 13919 1157 13968 1169
rect 1087 967 1136 977
rect 1087 947 1098 967
rect 1118 947 1136 967
rect 1087 935 1136 947
rect 1186 971 1230 977
rect 1186 951 1201 971
rect 1221 951 1230 971
rect 1186 935 1230 951
rect 1305 967 1354 977
rect 1305 947 1316 967
rect 1336 947 1354 967
rect 1305 935 1354 947
rect 1404 971 1448 977
rect 1404 951 1419 971
rect 1439 951 1448 971
rect 1404 935 1448 951
rect 1518 971 1562 977
rect 1518 951 1527 971
rect 1547 951 1562 971
rect 1518 935 1562 951
rect 1612 967 1661 977
rect 1612 947 1630 967
rect 1650 947 1661 967
rect 1612 935 1661 947
rect 5451 980 5500 990
rect 5451 960 5462 980
rect 5482 960 5500 980
rect 5451 948 5500 960
rect 5550 984 5594 990
rect 5550 964 5565 984
rect 5585 964 5594 984
rect 5550 948 5594 964
rect 5669 980 5718 990
rect 5669 960 5680 980
rect 5700 960 5718 980
rect 5669 948 5718 960
rect 5768 984 5812 990
rect 5768 964 5783 984
rect 5803 964 5812 984
rect 5768 948 5812 964
rect 5882 984 5926 990
rect 5882 964 5891 984
rect 5911 964 5926 984
rect 5882 948 5926 964
rect 5976 980 6025 990
rect 5976 960 5994 980
rect 6014 960 6025 980
rect 5976 948 6025 960
rect 9828 992 9877 1002
rect 9828 972 9839 992
rect 9859 972 9877 992
rect 9828 960 9877 972
rect 9927 996 9971 1002
rect 9927 976 9942 996
rect 9962 976 9971 996
rect 9927 960 9971 976
rect 10046 992 10095 1002
rect 10046 972 10057 992
rect 10077 972 10095 992
rect 10046 960 10095 972
rect 10145 996 10189 1002
rect 10145 976 10160 996
rect 10180 976 10189 996
rect 10145 960 10189 976
rect 10259 996 10303 1002
rect 10259 976 10268 996
rect 10288 976 10303 996
rect 10259 960 10303 976
rect 10353 992 10402 1002
rect 10353 972 10371 992
rect 10391 972 10402 992
rect 10353 960 10402 972
rect 14192 1005 14241 1015
rect 14192 985 14203 1005
rect 14223 985 14241 1005
rect 290 739 339 749
rect 290 719 301 739
rect 321 719 339 739
rect 290 707 339 719
rect 389 743 433 749
rect 389 723 404 743
rect 424 723 433 743
rect 389 707 433 723
rect 508 739 557 749
rect 508 719 519 739
rect 539 719 557 739
rect 508 707 557 719
rect 607 743 651 749
rect 607 723 622 743
rect 642 723 651 743
rect 607 707 651 723
rect 721 743 765 749
rect 721 723 730 743
rect 750 723 765 743
rect 721 707 765 723
rect 815 739 864 749
rect 815 719 833 739
rect 853 719 864 739
rect 14192 973 14241 985
rect 14291 1009 14335 1015
rect 14291 989 14306 1009
rect 14326 989 14335 1009
rect 14291 973 14335 989
rect 14410 1005 14459 1015
rect 14410 985 14421 1005
rect 14441 985 14459 1005
rect 14410 973 14459 985
rect 14509 1009 14553 1015
rect 14509 989 14524 1009
rect 14544 989 14553 1009
rect 14509 973 14553 989
rect 14623 1009 14667 1015
rect 14623 989 14632 1009
rect 14652 989 14667 1009
rect 14623 973 14667 989
rect 14717 1005 14766 1015
rect 14717 985 14735 1005
rect 14755 985 14766 1005
rect 14717 973 14766 985
rect 815 707 864 719
rect 4654 752 4703 762
rect 4654 732 4665 752
rect 4685 732 4703 752
rect 4654 720 4703 732
rect 4753 756 4797 762
rect 4753 736 4768 756
rect 4788 736 4797 756
rect 4753 720 4797 736
rect 4872 752 4921 762
rect 4872 732 4883 752
rect 4903 732 4921 752
rect 4872 720 4921 732
rect 4971 756 5015 762
rect 4971 736 4986 756
rect 5006 736 5015 756
rect 4971 720 5015 736
rect 5085 756 5129 762
rect 5085 736 5094 756
rect 5114 736 5129 756
rect 5085 720 5129 736
rect 5179 752 5228 762
rect 5179 732 5197 752
rect 5217 732 5228 752
rect 5179 720 5228 732
rect 9031 764 9080 774
rect 9031 744 9042 764
rect 9062 744 9080 764
rect 9031 732 9080 744
rect 9130 768 9174 774
rect 9130 748 9145 768
rect 9165 748 9174 768
rect 9130 732 9174 748
rect 9249 764 9298 774
rect 9249 744 9260 764
rect 9280 744 9298 764
rect 9249 732 9298 744
rect 9348 768 9392 774
rect 9348 748 9363 768
rect 9383 748 9392 768
rect 9348 732 9392 748
rect 9462 768 9506 774
rect 9462 748 9471 768
rect 9491 748 9506 768
rect 9462 732 9506 748
rect 9556 764 9605 774
rect 9556 744 9574 764
rect 9594 744 9605 764
rect 9556 732 9605 744
rect 13395 777 13444 787
rect 13395 757 13406 777
rect 13426 757 13444 777
rect 13395 745 13444 757
rect 13494 781 13538 787
rect 13494 761 13509 781
rect 13529 761 13538 781
rect 13494 745 13538 761
rect 13613 777 13662 787
rect 13613 757 13624 777
rect 13644 757 13662 777
rect 13613 745 13662 757
rect 13712 781 13756 787
rect 13712 761 13727 781
rect 13747 761 13756 781
rect 13712 745 13756 761
rect 13826 781 13870 787
rect 13826 761 13835 781
rect 13855 761 13870 781
rect 13826 745 13870 761
rect 13920 777 13969 787
rect 13920 757 13938 777
rect 13958 757 13969 777
rect 13920 745 13969 757
rect 5867 176 5916 186
rect 1503 163 1552 173
rect 1503 143 1514 163
rect 1534 143 1552 163
rect 1503 131 1552 143
rect 1602 167 1646 173
rect 1602 147 1617 167
rect 1637 147 1646 167
rect 1602 131 1646 147
rect 1721 163 1770 173
rect 1721 143 1732 163
rect 1752 143 1770 163
rect 1721 131 1770 143
rect 1820 167 1864 173
rect 1820 147 1835 167
rect 1855 147 1864 167
rect 1820 131 1864 147
rect 1934 167 1978 173
rect 1934 147 1943 167
rect 1963 147 1978 167
rect 1934 131 1978 147
rect 2028 163 2077 173
rect 2028 143 2046 163
rect 2066 143 2077 163
rect 2028 131 2077 143
rect 5867 156 5878 176
rect 5898 156 5916 176
rect 5867 144 5916 156
rect 5966 180 6010 186
rect 5966 160 5981 180
rect 6001 160 6010 180
rect 5966 144 6010 160
rect 6085 176 6134 186
rect 6085 156 6096 176
rect 6116 156 6134 176
rect 6085 144 6134 156
rect 6184 180 6228 186
rect 6184 160 6199 180
rect 6219 160 6228 180
rect 6184 144 6228 160
rect 6298 180 6342 186
rect 6298 160 6307 180
rect 6327 160 6342 180
rect 6298 144 6342 160
rect 6392 176 6441 186
rect 6392 156 6410 176
rect 6430 156 6441 176
rect 6392 144 6441 156
rect 14608 201 14657 211
rect 10244 188 10293 198
rect 10244 168 10255 188
rect 10275 168 10293 188
rect 10244 156 10293 168
rect 10343 192 10387 198
rect 10343 172 10358 192
rect 10378 172 10387 192
rect 10343 156 10387 172
rect 10462 188 10511 198
rect 10462 168 10473 188
rect 10493 168 10511 188
rect 10462 156 10511 168
rect 10561 192 10605 198
rect 10561 172 10576 192
rect 10596 172 10605 192
rect 10561 156 10605 172
rect 10675 192 10719 198
rect 10675 172 10684 192
rect 10704 172 10719 192
rect 10675 156 10719 172
rect 10769 188 10818 198
rect 10769 168 10787 188
rect 10807 168 10818 188
rect 10769 156 10818 168
rect 14608 181 14619 201
rect 14639 181 14657 201
rect 14608 169 14657 181
rect 14707 205 14751 211
rect 14707 185 14722 205
rect 14742 185 14751 205
rect 14707 169 14751 185
rect 14826 201 14875 211
rect 14826 181 14837 201
rect 14857 181 14875 201
rect 14826 169 14875 181
rect 14925 205 14969 211
rect 14925 185 14940 205
rect 14960 185 14969 205
rect 14925 169 14969 185
rect 15039 205 15083 211
rect 15039 185 15048 205
rect 15068 185 15083 205
rect 15039 169 15083 185
rect 15133 201 15182 211
rect 15133 181 15151 201
rect 15171 181 15182 201
rect 15133 169 15182 181
rect 8440 113 8489 123
rect 3992 89 4041 99
rect 3992 69 4003 89
rect 4023 69 4041 89
rect 3992 57 4041 69
rect 4091 93 4135 99
rect 4091 73 4106 93
rect 4126 73 4135 93
rect 4091 57 4135 73
rect 4210 89 4259 99
rect 4210 69 4221 89
rect 4241 69 4259 89
rect 4210 57 4259 69
rect 4309 93 4353 99
rect 4309 73 4324 93
rect 4344 73 4353 93
rect 4309 57 4353 73
rect 4423 93 4467 99
rect 4423 73 4432 93
rect 4452 73 4467 93
rect 4423 57 4467 73
rect 4517 89 4566 99
rect 4517 69 4535 89
rect 4555 69 4566 89
rect 8440 93 8451 113
rect 8471 93 8489 113
rect 8440 81 8489 93
rect 8539 117 8583 123
rect 8539 97 8554 117
rect 8574 97 8583 117
rect 8539 81 8583 97
rect 8658 113 8707 123
rect 8658 93 8669 113
rect 8689 93 8707 113
rect 8658 81 8707 93
rect 8757 117 8801 123
rect 8757 97 8772 117
rect 8792 97 8801 117
rect 8757 81 8801 97
rect 8871 117 8915 123
rect 8871 97 8880 117
rect 8900 97 8915 117
rect 8871 81 8915 97
rect 8965 113 9014 123
rect 8965 93 8983 113
rect 9003 93 9014 113
rect 8965 81 9014 93
rect 12733 114 12782 124
rect 12733 94 12744 114
rect 12764 94 12782 114
rect 12733 82 12782 94
rect 12832 118 12876 124
rect 12832 98 12847 118
rect 12867 98 12876 118
rect 12832 82 12876 98
rect 12951 114 13000 124
rect 12951 94 12962 114
rect 12982 94 13000 114
rect 12951 82 13000 94
rect 13050 118 13094 124
rect 13050 98 13065 118
rect 13085 98 13094 118
rect 13050 82 13094 98
rect 13164 118 13208 124
rect 13164 98 13173 118
rect 13193 98 13208 118
rect 13164 82 13208 98
rect 13258 114 13307 124
rect 13258 94 13276 114
rect 13296 94 13307 114
rect 13258 82 13307 94
rect 4517 57 4566 69
<< pdiff >>
rect 3474 8590 3518 8632
rect 3474 8570 3486 8590
rect 3506 8570 3518 8590
rect 3474 8563 3518 8570
rect 3473 8532 3518 8563
rect 3568 8590 3610 8632
rect 3568 8570 3582 8590
rect 3602 8570 3610 8590
rect 3568 8532 3610 8570
rect 3684 8590 3726 8632
rect 3684 8570 3692 8590
rect 3712 8570 3726 8590
rect 3684 8532 3726 8570
rect 3776 8590 3820 8632
rect 3776 8570 3788 8590
rect 3808 8570 3820 8590
rect 3776 8532 3820 8570
rect 3902 8590 3944 8632
rect 3902 8570 3910 8590
rect 3930 8570 3944 8590
rect 3902 8532 3944 8570
rect 3994 8590 4038 8632
rect 3994 8570 4006 8590
rect 4026 8570 4038 8590
rect 3994 8532 4038 8570
rect 7838 8603 7882 8645
rect 7838 8583 7850 8603
rect 7870 8583 7882 8603
rect 7838 8576 7882 8583
rect 7837 8545 7882 8576
rect 7932 8603 7974 8645
rect 7932 8583 7946 8603
rect 7966 8583 7974 8603
rect 7932 8545 7974 8583
rect 8048 8603 8090 8645
rect 8048 8583 8056 8603
rect 8076 8583 8090 8603
rect 8048 8545 8090 8583
rect 8140 8603 8184 8645
rect 8140 8583 8152 8603
rect 8172 8583 8184 8603
rect 8140 8545 8184 8583
rect 8266 8603 8308 8645
rect 8266 8583 8274 8603
rect 8294 8583 8308 8603
rect 8266 8545 8308 8583
rect 8358 8603 8402 8645
rect 8358 8583 8370 8603
rect 8390 8583 8402 8603
rect 8358 8545 8402 8583
rect 12215 8615 12259 8657
rect 12215 8595 12227 8615
rect 12247 8595 12259 8615
rect 12215 8588 12259 8595
rect 12214 8557 12259 8588
rect 12309 8615 12351 8657
rect 12309 8595 12323 8615
rect 12343 8595 12351 8615
rect 12309 8557 12351 8595
rect 12425 8615 12467 8657
rect 12425 8595 12433 8615
rect 12453 8595 12467 8615
rect 12425 8557 12467 8595
rect 12517 8615 12561 8657
rect 12517 8595 12529 8615
rect 12549 8595 12561 8615
rect 12517 8557 12561 8595
rect 12643 8615 12685 8657
rect 12643 8595 12651 8615
rect 12671 8595 12685 8615
rect 12643 8557 12685 8595
rect 12735 8615 12779 8657
rect 12735 8595 12747 8615
rect 12767 8595 12779 8615
rect 12735 8557 12779 8595
rect 16579 8628 16623 8670
rect 16579 8608 16591 8628
rect 16611 8608 16623 8628
rect 16579 8601 16623 8608
rect 16578 8570 16623 8601
rect 16673 8628 16715 8670
rect 16673 8608 16687 8628
rect 16707 8608 16715 8628
rect 16673 8570 16715 8608
rect 16789 8628 16831 8670
rect 16789 8608 16797 8628
rect 16817 8608 16831 8628
rect 16789 8570 16831 8608
rect 16881 8628 16925 8670
rect 16881 8608 16893 8628
rect 16913 8608 16925 8628
rect 16881 8570 16925 8608
rect 17007 8628 17049 8670
rect 17007 8608 17015 8628
rect 17035 8608 17049 8628
rect 17007 8570 17049 8608
rect 17099 8628 17143 8670
rect 17099 8608 17111 8628
rect 17131 8608 17143 8628
rect 17099 8570 17143 8608
rect 421 8426 465 8464
rect 421 8406 433 8426
rect 453 8406 465 8426
rect 421 8364 465 8406
rect 515 8426 557 8464
rect 515 8406 529 8426
rect 549 8406 557 8426
rect 515 8364 557 8406
rect 639 8426 683 8464
rect 639 8406 651 8426
rect 671 8406 683 8426
rect 639 8364 683 8406
rect 733 8426 775 8464
rect 733 8406 747 8426
rect 767 8406 775 8426
rect 733 8364 775 8406
rect 849 8426 891 8464
rect 849 8406 857 8426
rect 877 8406 891 8426
rect 849 8364 891 8406
rect 941 8433 986 8464
rect 941 8426 985 8433
rect 941 8406 953 8426
rect 973 8406 985 8426
rect 941 8364 985 8406
rect 4785 8439 4829 8477
rect 4785 8419 4797 8439
rect 4817 8419 4829 8439
rect 2677 8362 2721 8404
rect 2677 8342 2689 8362
rect 2709 8342 2721 8362
rect 2677 8335 2721 8342
rect 2676 8304 2721 8335
rect 2771 8362 2813 8404
rect 2771 8342 2785 8362
rect 2805 8342 2813 8362
rect 2771 8304 2813 8342
rect 2887 8362 2929 8404
rect 2887 8342 2895 8362
rect 2915 8342 2929 8362
rect 2887 8304 2929 8342
rect 2979 8362 3023 8404
rect 2979 8342 2991 8362
rect 3011 8342 3023 8362
rect 2979 8304 3023 8342
rect 3105 8362 3147 8404
rect 3105 8342 3113 8362
rect 3133 8342 3147 8362
rect 3105 8304 3147 8342
rect 3197 8362 3241 8404
rect 4785 8377 4829 8419
rect 4879 8439 4921 8477
rect 4879 8419 4893 8439
rect 4913 8419 4921 8439
rect 4879 8377 4921 8419
rect 5003 8439 5047 8477
rect 5003 8419 5015 8439
rect 5035 8419 5047 8439
rect 5003 8377 5047 8419
rect 5097 8439 5139 8477
rect 5097 8419 5111 8439
rect 5131 8419 5139 8439
rect 5097 8377 5139 8419
rect 5213 8439 5255 8477
rect 5213 8419 5221 8439
rect 5241 8419 5255 8439
rect 5213 8377 5255 8419
rect 5305 8446 5350 8477
rect 5305 8439 5349 8446
rect 5305 8419 5317 8439
rect 5337 8419 5349 8439
rect 5305 8377 5349 8419
rect 9162 8451 9206 8489
rect 9162 8431 9174 8451
rect 9194 8431 9206 8451
rect 3197 8342 3209 8362
rect 3229 8342 3241 8362
rect 3197 8304 3241 8342
rect 1219 8242 1263 8280
rect 1219 8222 1231 8242
rect 1251 8222 1263 8242
rect 1219 8180 1263 8222
rect 1313 8242 1355 8280
rect 1313 8222 1327 8242
rect 1347 8222 1355 8242
rect 1313 8180 1355 8222
rect 1437 8242 1481 8280
rect 1437 8222 1449 8242
rect 1469 8222 1481 8242
rect 1437 8180 1481 8222
rect 1531 8242 1573 8280
rect 1531 8222 1545 8242
rect 1565 8222 1573 8242
rect 1531 8180 1573 8222
rect 1647 8242 1689 8280
rect 1647 8222 1655 8242
rect 1675 8222 1689 8242
rect 1647 8180 1689 8222
rect 1739 8249 1784 8280
rect 1739 8242 1783 8249
rect 1739 8222 1751 8242
rect 1771 8222 1783 8242
rect 1739 8180 1783 8222
rect 7041 8375 7085 8417
rect 7041 8355 7053 8375
rect 7073 8355 7085 8375
rect 7041 8348 7085 8355
rect 7040 8317 7085 8348
rect 7135 8375 7177 8417
rect 7135 8355 7149 8375
rect 7169 8355 7177 8375
rect 7135 8317 7177 8355
rect 7251 8375 7293 8417
rect 7251 8355 7259 8375
rect 7279 8355 7293 8375
rect 7251 8317 7293 8355
rect 7343 8375 7387 8417
rect 7343 8355 7355 8375
rect 7375 8355 7387 8375
rect 7343 8317 7387 8355
rect 7469 8375 7511 8417
rect 7469 8355 7477 8375
rect 7497 8355 7511 8375
rect 7469 8317 7511 8355
rect 7561 8375 7605 8417
rect 9162 8389 9206 8431
rect 9256 8451 9298 8489
rect 9256 8431 9270 8451
rect 9290 8431 9298 8451
rect 9256 8389 9298 8431
rect 9380 8451 9424 8489
rect 9380 8431 9392 8451
rect 9412 8431 9424 8451
rect 9380 8389 9424 8431
rect 9474 8451 9516 8489
rect 9474 8431 9488 8451
rect 9508 8431 9516 8451
rect 9474 8389 9516 8431
rect 9590 8451 9632 8489
rect 9590 8431 9598 8451
rect 9618 8431 9632 8451
rect 9590 8389 9632 8431
rect 9682 8458 9727 8489
rect 9682 8451 9726 8458
rect 9682 8431 9694 8451
rect 9714 8431 9726 8451
rect 9682 8389 9726 8431
rect 13526 8464 13570 8502
rect 13526 8444 13538 8464
rect 13558 8444 13570 8464
rect 7561 8355 7573 8375
rect 7593 8355 7605 8375
rect 7561 8317 7605 8355
rect 5583 8255 5627 8293
rect 5583 8235 5595 8255
rect 5615 8235 5627 8255
rect 3475 8178 3519 8220
rect 3475 8158 3487 8178
rect 3507 8158 3519 8178
rect 3475 8151 3519 8158
rect 3474 8120 3519 8151
rect 3569 8178 3611 8220
rect 3569 8158 3583 8178
rect 3603 8158 3611 8178
rect 3569 8120 3611 8158
rect 3685 8178 3727 8220
rect 3685 8158 3693 8178
rect 3713 8158 3727 8178
rect 3685 8120 3727 8158
rect 3777 8178 3821 8220
rect 3777 8158 3789 8178
rect 3809 8158 3821 8178
rect 3777 8120 3821 8158
rect 3903 8178 3945 8220
rect 3903 8158 3911 8178
rect 3931 8158 3945 8178
rect 3903 8120 3945 8158
rect 3995 8178 4039 8220
rect 5583 8193 5627 8235
rect 5677 8255 5719 8293
rect 5677 8235 5691 8255
rect 5711 8235 5719 8255
rect 5677 8193 5719 8235
rect 5801 8255 5845 8293
rect 5801 8235 5813 8255
rect 5833 8235 5845 8255
rect 5801 8193 5845 8235
rect 5895 8255 5937 8293
rect 5895 8235 5909 8255
rect 5929 8235 5937 8255
rect 5895 8193 5937 8235
rect 6011 8255 6053 8293
rect 6011 8235 6019 8255
rect 6039 8235 6053 8255
rect 6011 8193 6053 8235
rect 6103 8262 6148 8293
rect 6103 8255 6147 8262
rect 6103 8235 6115 8255
rect 6135 8235 6147 8255
rect 6103 8193 6147 8235
rect 11418 8387 11462 8429
rect 11418 8367 11430 8387
rect 11450 8367 11462 8387
rect 11418 8360 11462 8367
rect 11417 8329 11462 8360
rect 11512 8387 11554 8429
rect 11512 8367 11526 8387
rect 11546 8367 11554 8387
rect 11512 8329 11554 8367
rect 11628 8387 11670 8429
rect 11628 8367 11636 8387
rect 11656 8367 11670 8387
rect 11628 8329 11670 8367
rect 11720 8387 11764 8429
rect 11720 8367 11732 8387
rect 11752 8367 11764 8387
rect 11720 8329 11764 8367
rect 11846 8387 11888 8429
rect 11846 8367 11854 8387
rect 11874 8367 11888 8387
rect 11846 8329 11888 8367
rect 11938 8387 11982 8429
rect 13526 8402 13570 8444
rect 13620 8464 13662 8502
rect 13620 8444 13634 8464
rect 13654 8444 13662 8464
rect 13620 8402 13662 8444
rect 13744 8464 13788 8502
rect 13744 8444 13756 8464
rect 13776 8444 13788 8464
rect 13744 8402 13788 8444
rect 13838 8464 13880 8502
rect 13838 8444 13852 8464
rect 13872 8444 13880 8464
rect 13838 8402 13880 8444
rect 13954 8464 13996 8502
rect 13954 8444 13962 8464
rect 13982 8444 13996 8464
rect 13954 8402 13996 8444
rect 14046 8471 14091 8502
rect 14046 8464 14090 8471
rect 14046 8444 14058 8464
rect 14078 8444 14090 8464
rect 14046 8402 14090 8444
rect 11938 8367 11950 8387
rect 11970 8367 11982 8387
rect 11938 8329 11982 8367
rect 9960 8267 10004 8305
rect 9960 8247 9972 8267
rect 9992 8247 10004 8267
rect 3995 8158 4007 8178
rect 4027 8158 4039 8178
rect 3995 8120 4039 8158
rect 7839 8191 7883 8233
rect 7839 8171 7851 8191
rect 7871 8171 7883 8191
rect 7839 8164 7883 8171
rect 7838 8133 7883 8164
rect 7933 8191 7975 8233
rect 7933 8171 7947 8191
rect 7967 8171 7975 8191
rect 7933 8133 7975 8171
rect 8049 8191 8091 8233
rect 8049 8171 8057 8191
rect 8077 8171 8091 8191
rect 8049 8133 8091 8171
rect 8141 8191 8185 8233
rect 8141 8171 8153 8191
rect 8173 8171 8185 8191
rect 8141 8133 8185 8171
rect 8267 8191 8309 8233
rect 8267 8171 8275 8191
rect 8295 8171 8309 8191
rect 8267 8133 8309 8171
rect 8359 8191 8403 8233
rect 9960 8205 10004 8247
rect 10054 8267 10096 8305
rect 10054 8247 10068 8267
rect 10088 8247 10096 8267
rect 10054 8205 10096 8247
rect 10178 8267 10222 8305
rect 10178 8247 10190 8267
rect 10210 8247 10222 8267
rect 10178 8205 10222 8247
rect 10272 8267 10314 8305
rect 10272 8247 10286 8267
rect 10306 8247 10314 8267
rect 10272 8205 10314 8247
rect 10388 8267 10430 8305
rect 10388 8247 10396 8267
rect 10416 8247 10430 8267
rect 10388 8205 10430 8247
rect 10480 8274 10525 8305
rect 10480 8267 10524 8274
rect 10480 8247 10492 8267
rect 10512 8247 10524 8267
rect 10480 8205 10524 8247
rect 15782 8400 15826 8442
rect 15782 8380 15794 8400
rect 15814 8380 15826 8400
rect 15782 8373 15826 8380
rect 15781 8342 15826 8373
rect 15876 8400 15918 8442
rect 15876 8380 15890 8400
rect 15910 8380 15918 8400
rect 15876 8342 15918 8380
rect 15992 8400 16034 8442
rect 15992 8380 16000 8400
rect 16020 8380 16034 8400
rect 15992 8342 16034 8380
rect 16084 8400 16128 8442
rect 16084 8380 16096 8400
rect 16116 8380 16128 8400
rect 16084 8342 16128 8380
rect 16210 8400 16252 8442
rect 16210 8380 16218 8400
rect 16238 8380 16252 8400
rect 16210 8342 16252 8380
rect 16302 8400 16346 8442
rect 16302 8380 16314 8400
rect 16334 8380 16346 8400
rect 16302 8342 16346 8380
rect 14324 8280 14368 8318
rect 14324 8260 14336 8280
rect 14356 8260 14368 8280
rect 8359 8171 8371 8191
rect 8391 8171 8403 8191
rect 8359 8133 8403 8171
rect 422 8014 466 8052
rect 422 7994 434 8014
rect 454 7994 466 8014
rect 422 7952 466 7994
rect 516 8014 558 8052
rect 516 7994 530 8014
rect 550 7994 558 8014
rect 516 7952 558 7994
rect 640 8014 684 8052
rect 640 7994 652 8014
rect 672 7994 684 8014
rect 640 7952 684 7994
rect 734 8014 776 8052
rect 734 7994 748 8014
rect 768 7994 776 8014
rect 734 7952 776 7994
rect 850 8014 892 8052
rect 850 7994 858 8014
rect 878 7994 892 8014
rect 850 7952 892 7994
rect 942 8021 987 8052
rect 942 8014 986 8021
rect 942 7994 954 8014
rect 974 7994 986 8014
rect 12216 8203 12260 8245
rect 12216 8183 12228 8203
rect 12248 8183 12260 8203
rect 12216 8176 12260 8183
rect 12215 8145 12260 8176
rect 12310 8203 12352 8245
rect 12310 8183 12324 8203
rect 12344 8183 12352 8203
rect 12310 8145 12352 8183
rect 12426 8203 12468 8245
rect 12426 8183 12434 8203
rect 12454 8183 12468 8203
rect 12426 8145 12468 8183
rect 12518 8203 12562 8245
rect 12518 8183 12530 8203
rect 12550 8183 12562 8203
rect 12518 8145 12562 8183
rect 12644 8203 12686 8245
rect 12644 8183 12652 8203
rect 12672 8183 12686 8203
rect 12644 8145 12686 8183
rect 12736 8203 12780 8245
rect 14324 8218 14368 8260
rect 14418 8280 14460 8318
rect 14418 8260 14432 8280
rect 14452 8260 14460 8280
rect 14418 8218 14460 8260
rect 14542 8280 14586 8318
rect 14542 8260 14554 8280
rect 14574 8260 14586 8280
rect 14542 8218 14586 8260
rect 14636 8280 14678 8318
rect 14636 8260 14650 8280
rect 14670 8260 14678 8280
rect 14636 8218 14678 8260
rect 14752 8280 14794 8318
rect 14752 8260 14760 8280
rect 14780 8260 14794 8280
rect 14752 8218 14794 8260
rect 14844 8287 14889 8318
rect 14844 8280 14888 8287
rect 14844 8260 14856 8280
rect 14876 8260 14888 8280
rect 14844 8218 14888 8260
rect 12736 8183 12748 8203
rect 12768 8183 12780 8203
rect 12736 8145 12780 8183
rect 4786 8027 4830 8065
rect 942 7952 986 7994
rect 2578 7952 2622 7994
rect 2578 7932 2590 7952
rect 2610 7932 2622 7952
rect 2578 7925 2622 7932
rect 2577 7894 2622 7925
rect 2672 7952 2714 7994
rect 2672 7932 2686 7952
rect 2706 7932 2714 7952
rect 2672 7894 2714 7932
rect 2788 7952 2830 7994
rect 2788 7932 2796 7952
rect 2816 7932 2830 7952
rect 2788 7894 2830 7932
rect 2880 7952 2924 7994
rect 2880 7932 2892 7952
rect 2912 7932 2924 7952
rect 2880 7894 2924 7932
rect 3006 7952 3048 7994
rect 3006 7932 3014 7952
rect 3034 7932 3048 7952
rect 3006 7894 3048 7932
rect 3098 7952 3142 7994
rect 4786 8007 4798 8027
rect 4818 8007 4830 8027
rect 3098 7932 3110 7952
rect 3130 7932 3142 7952
rect 4786 7965 4830 8007
rect 4880 8027 4922 8065
rect 4880 8007 4894 8027
rect 4914 8007 4922 8027
rect 4880 7965 4922 8007
rect 5004 8027 5048 8065
rect 5004 8007 5016 8027
rect 5036 8007 5048 8027
rect 5004 7965 5048 8007
rect 5098 8027 5140 8065
rect 5098 8007 5112 8027
rect 5132 8007 5140 8027
rect 5098 7965 5140 8007
rect 5214 8027 5256 8065
rect 5214 8007 5222 8027
rect 5242 8007 5256 8027
rect 5214 7965 5256 8007
rect 5306 8034 5351 8065
rect 5306 8027 5350 8034
rect 5306 8007 5318 8027
rect 5338 8007 5350 8027
rect 16580 8216 16624 8258
rect 16580 8196 16592 8216
rect 16612 8196 16624 8216
rect 16580 8189 16624 8196
rect 16579 8158 16624 8189
rect 16674 8216 16716 8258
rect 16674 8196 16688 8216
rect 16708 8196 16716 8216
rect 16674 8158 16716 8196
rect 16790 8216 16832 8258
rect 16790 8196 16798 8216
rect 16818 8196 16832 8216
rect 16790 8158 16832 8196
rect 16882 8216 16926 8258
rect 16882 8196 16894 8216
rect 16914 8196 16926 8216
rect 16882 8158 16926 8196
rect 17008 8216 17050 8258
rect 17008 8196 17016 8216
rect 17036 8196 17050 8216
rect 17008 8158 17050 8196
rect 17100 8216 17144 8258
rect 17100 8196 17112 8216
rect 17132 8196 17144 8216
rect 17100 8158 17144 8196
rect 9163 8039 9207 8077
rect 5306 7965 5350 8007
rect 6942 7965 6986 8007
rect 3098 7894 3142 7932
rect 6942 7945 6954 7965
rect 6974 7945 6986 7965
rect 6942 7938 6986 7945
rect 6941 7907 6986 7938
rect 7036 7965 7078 8007
rect 7036 7945 7050 7965
rect 7070 7945 7078 7965
rect 7036 7907 7078 7945
rect 7152 7965 7194 8007
rect 7152 7945 7160 7965
rect 7180 7945 7194 7965
rect 7152 7907 7194 7945
rect 7244 7965 7288 8007
rect 7244 7945 7256 7965
rect 7276 7945 7288 7965
rect 7244 7907 7288 7945
rect 7370 7965 7412 8007
rect 7370 7945 7378 7965
rect 7398 7945 7412 7965
rect 7370 7907 7412 7945
rect 7462 7965 7506 8007
rect 9163 8019 9175 8039
rect 9195 8019 9207 8039
rect 7462 7945 7474 7965
rect 7494 7945 7506 7965
rect 9163 7977 9207 8019
rect 9257 8039 9299 8077
rect 9257 8019 9271 8039
rect 9291 8019 9299 8039
rect 9257 7977 9299 8019
rect 9381 8039 9425 8077
rect 9381 8019 9393 8039
rect 9413 8019 9425 8039
rect 9381 7977 9425 8019
rect 9475 8039 9517 8077
rect 9475 8019 9489 8039
rect 9509 8019 9517 8039
rect 9475 7977 9517 8019
rect 9591 8039 9633 8077
rect 9591 8019 9599 8039
rect 9619 8019 9633 8039
rect 9591 7977 9633 8019
rect 9683 8046 9728 8077
rect 9683 8039 9727 8046
rect 9683 8019 9695 8039
rect 9715 8019 9727 8039
rect 13527 8052 13571 8090
rect 9683 7977 9727 8019
rect 11319 7977 11363 8019
rect 7462 7907 7506 7945
rect 11319 7957 11331 7977
rect 11351 7957 11363 7977
rect 11319 7950 11363 7957
rect 11318 7919 11363 7950
rect 11413 7977 11455 8019
rect 11413 7957 11427 7977
rect 11447 7957 11455 7977
rect 11413 7919 11455 7957
rect 11529 7977 11571 8019
rect 11529 7957 11537 7977
rect 11557 7957 11571 7977
rect 11529 7919 11571 7957
rect 11621 7977 11665 8019
rect 11621 7957 11633 7977
rect 11653 7957 11665 7977
rect 11621 7919 11665 7957
rect 11747 7977 11789 8019
rect 11747 7957 11755 7977
rect 11775 7957 11789 7977
rect 11747 7919 11789 7957
rect 11839 7977 11883 8019
rect 13527 8032 13539 8052
rect 13559 8032 13571 8052
rect 11839 7957 11851 7977
rect 11871 7957 11883 7977
rect 13527 7990 13571 8032
rect 13621 8052 13663 8090
rect 13621 8032 13635 8052
rect 13655 8032 13663 8052
rect 13621 7990 13663 8032
rect 13745 8052 13789 8090
rect 13745 8032 13757 8052
rect 13777 8032 13789 8052
rect 13745 7990 13789 8032
rect 13839 8052 13881 8090
rect 13839 8032 13853 8052
rect 13873 8032 13881 8052
rect 13839 7990 13881 8032
rect 13955 8052 13997 8090
rect 13955 8032 13963 8052
rect 13983 8032 13997 8052
rect 13955 7990 13997 8032
rect 14047 8059 14092 8090
rect 14047 8052 14091 8059
rect 14047 8032 14059 8052
rect 14079 8032 14091 8052
rect 14047 7990 14091 8032
rect 15683 7990 15727 8032
rect 11839 7919 11883 7957
rect 15683 7970 15695 7990
rect 15715 7970 15727 7990
rect 15683 7963 15727 7970
rect 15682 7932 15727 7963
rect 15777 7990 15819 8032
rect 15777 7970 15791 7990
rect 15811 7970 15819 7990
rect 15777 7932 15819 7970
rect 15893 7990 15935 8032
rect 15893 7970 15901 7990
rect 15921 7970 15935 7990
rect 15893 7932 15935 7970
rect 15985 7990 16029 8032
rect 15985 7970 15997 7990
rect 16017 7970 16029 7990
rect 15985 7932 16029 7970
rect 16111 7990 16153 8032
rect 16111 7970 16119 7990
rect 16139 7970 16153 7990
rect 16111 7932 16153 7970
rect 16203 7990 16247 8032
rect 16203 7970 16215 7990
rect 16235 7970 16247 7990
rect 16203 7932 16247 7970
rect 1301 7634 1345 7672
rect 1301 7614 1313 7634
rect 1333 7614 1345 7634
rect 1301 7572 1345 7614
rect 1395 7634 1437 7672
rect 1395 7614 1409 7634
rect 1429 7614 1437 7634
rect 1395 7572 1437 7614
rect 1519 7634 1563 7672
rect 1519 7614 1531 7634
rect 1551 7614 1563 7634
rect 1519 7572 1563 7614
rect 1613 7634 1655 7672
rect 1613 7614 1627 7634
rect 1647 7614 1655 7634
rect 1613 7572 1655 7614
rect 1729 7634 1771 7672
rect 1729 7614 1737 7634
rect 1757 7614 1771 7634
rect 1729 7572 1771 7614
rect 1821 7641 1866 7672
rect 1821 7634 1865 7641
rect 1821 7614 1833 7634
rect 1853 7614 1865 7634
rect 5665 7647 5709 7685
rect 1821 7572 1865 7614
rect 3457 7572 3501 7614
rect 3457 7552 3469 7572
rect 3489 7552 3501 7572
rect 3457 7545 3501 7552
rect 3456 7514 3501 7545
rect 3551 7572 3593 7614
rect 3551 7552 3565 7572
rect 3585 7552 3593 7572
rect 3551 7514 3593 7552
rect 3667 7572 3709 7614
rect 3667 7552 3675 7572
rect 3695 7552 3709 7572
rect 3667 7514 3709 7552
rect 3759 7572 3803 7614
rect 3759 7552 3771 7572
rect 3791 7552 3803 7572
rect 3759 7514 3803 7552
rect 3885 7572 3927 7614
rect 3885 7552 3893 7572
rect 3913 7552 3927 7572
rect 3885 7514 3927 7552
rect 3977 7572 4021 7614
rect 5665 7627 5677 7647
rect 5697 7627 5709 7647
rect 3977 7552 3989 7572
rect 4009 7552 4021 7572
rect 5665 7585 5709 7627
rect 5759 7647 5801 7685
rect 5759 7627 5773 7647
rect 5793 7627 5801 7647
rect 5759 7585 5801 7627
rect 5883 7647 5927 7685
rect 5883 7627 5895 7647
rect 5915 7627 5927 7647
rect 5883 7585 5927 7627
rect 5977 7647 6019 7685
rect 5977 7627 5991 7647
rect 6011 7627 6019 7647
rect 5977 7585 6019 7627
rect 6093 7647 6135 7685
rect 6093 7627 6101 7647
rect 6121 7627 6135 7647
rect 6093 7585 6135 7627
rect 6185 7654 6230 7685
rect 6185 7647 6229 7654
rect 6185 7627 6197 7647
rect 6217 7627 6229 7647
rect 10042 7659 10086 7697
rect 6185 7585 6229 7627
rect 7821 7585 7865 7627
rect 3977 7514 4021 7552
rect 7821 7565 7833 7585
rect 7853 7565 7865 7585
rect 7821 7558 7865 7565
rect 7820 7527 7865 7558
rect 7915 7585 7957 7627
rect 7915 7565 7929 7585
rect 7949 7565 7957 7585
rect 7915 7527 7957 7565
rect 8031 7585 8073 7627
rect 8031 7565 8039 7585
rect 8059 7565 8073 7585
rect 8031 7527 8073 7565
rect 8123 7585 8167 7627
rect 8123 7565 8135 7585
rect 8155 7565 8167 7585
rect 8123 7527 8167 7565
rect 8249 7585 8291 7627
rect 8249 7565 8257 7585
rect 8277 7565 8291 7585
rect 8249 7527 8291 7565
rect 8341 7585 8385 7627
rect 10042 7639 10054 7659
rect 10074 7639 10086 7659
rect 8341 7565 8353 7585
rect 8373 7565 8385 7585
rect 10042 7597 10086 7639
rect 10136 7659 10178 7697
rect 10136 7639 10150 7659
rect 10170 7639 10178 7659
rect 10136 7597 10178 7639
rect 10260 7659 10304 7697
rect 10260 7639 10272 7659
rect 10292 7639 10304 7659
rect 10260 7597 10304 7639
rect 10354 7659 10396 7697
rect 10354 7639 10368 7659
rect 10388 7639 10396 7659
rect 10354 7597 10396 7639
rect 10470 7659 10512 7697
rect 10470 7639 10478 7659
rect 10498 7639 10512 7659
rect 10470 7597 10512 7639
rect 10562 7666 10607 7697
rect 10562 7659 10606 7666
rect 10562 7639 10574 7659
rect 10594 7639 10606 7659
rect 14406 7672 14450 7710
rect 10562 7597 10606 7639
rect 12198 7597 12242 7639
rect 8341 7527 8385 7565
rect 404 7408 448 7446
rect 404 7388 416 7408
rect 436 7388 448 7408
rect 404 7346 448 7388
rect 498 7408 540 7446
rect 498 7388 512 7408
rect 532 7388 540 7408
rect 498 7346 540 7388
rect 622 7408 666 7446
rect 622 7388 634 7408
rect 654 7388 666 7408
rect 622 7346 666 7388
rect 716 7408 758 7446
rect 716 7388 730 7408
rect 750 7388 758 7408
rect 716 7346 758 7388
rect 832 7408 874 7446
rect 832 7388 840 7408
rect 860 7388 874 7408
rect 832 7346 874 7388
rect 924 7415 969 7446
rect 924 7408 968 7415
rect 924 7388 936 7408
rect 956 7388 968 7408
rect 924 7346 968 7388
rect 12198 7577 12210 7597
rect 12230 7577 12242 7597
rect 12198 7570 12242 7577
rect 12197 7539 12242 7570
rect 12292 7597 12334 7639
rect 12292 7577 12306 7597
rect 12326 7577 12334 7597
rect 12292 7539 12334 7577
rect 12408 7597 12450 7639
rect 12408 7577 12416 7597
rect 12436 7577 12450 7597
rect 12408 7539 12450 7577
rect 12500 7597 12544 7639
rect 12500 7577 12512 7597
rect 12532 7577 12544 7597
rect 12500 7539 12544 7577
rect 12626 7597 12668 7639
rect 12626 7577 12634 7597
rect 12654 7577 12668 7597
rect 12626 7539 12668 7577
rect 12718 7597 12762 7639
rect 14406 7652 14418 7672
rect 14438 7652 14450 7672
rect 12718 7577 12730 7597
rect 12750 7577 12762 7597
rect 14406 7610 14450 7652
rect 14500 7672 14542 7710
rect 14500 7652 14514 7672
rect 14534 7652 14542 7672
rect 14500 7610 14542 7652
rect 14624 7672 14668 7710
rect 14624 7652 14636 7672
rect 14656 7652 14668 7672
rect 14624 7610 14668 7652
rect 14718 7672 14760 7710
rect 14718 7652 14732 7672
rect 14752 7652 14760 7672
rect 14718 7610 14760 7652
rect 14834 7672 14876 7710
rect 14834 7652 14842 7672
rect 14862 7652 14876 7672
rect 14834 7610 14876 7652
rect 14926 7679 14971 7710
rect 14926 7672 14970 7679
rect 14926 7652 14938 7672
rect 14958 7652 14970 7672
rect 14926 7610 14970 7652
rect 16562 7610 16606 7652
rect 12718 7539 12762 7577
rect 4768 7421 4812 7459
rect 4768 7401 4780 7421
rect 4800 7401 4812 7421
rect 2660 7344 2704 7386
rect 2660 7324 2672 7344
rect 2692 7324 2704 7344
rect 2660 7317 2704 7324
rect 2659 7286 2704 7317
rect 2754 7344 2796 7386
rect 2754 7324 2768 7344
rect 2788 7324 2796 7344
rect 2754 7286 2796 7324
rect 2870 7344 2912 7386
rect 2870 7324 2878 7344
rect 2898 7324 2912 7344
rect 2870 7286 2912 7324
rect 2962 7344 3006 7386
rect 2962 7324 2974 7344
rect 2994 7324 3006 7344
rect 2962 7286 3006 7324
rect 3088 7344 3130 7386
rect 3088 7324 3096 7344
rect 3116 7324 3130 7344
rect 3088 7286 3130 7324
rect 3180 7344 3224 7386
rect 4768 7359 4812 7401
rect 4862 7421 4904 7459
rect 4862 7401 4876 7421
rect 4896 7401 4904 7421
rect 4862 7359 4904 7401
rect 4986 7421 5030 7459
rect 4986 7401 4998 7421
rect 5018 7401 5030 7421
rect 4986 7359 5030 7401
rect 5080 7421 5122 7459
rect 5080 7401 5094 7421
rect 5114 7401 5122 7421
rect 5080 7359 5122 7401
rect 5196 7421 5238 7459
rect 5196 7401 5204 7421
rect 5224 7401 5238 7421
rect 5196 7359 5238 7401
rect 5288 7428 5333 7459
rect 5288 7421 5332 7428
rect 5288 7401 5300 7421
rect 5320 7401 5332 7421
rect 5288 7359 5332 7401
rect 16562 7590 16574 7610
rect 16594 7590 16606 7610
rect 16562 7583 16606 7590
rect 16561 7552 16606 7583
rect 16656 7610 16698 7652
rect 16656 7590 16670 7610
rect 16690 7590 16698 7610
rect 16656 7552 16698 7590
rect 16772 7610 16814 7652
rect 16772 7590 16780 7610
rect 16800 7590 16814 7610
rect 16772 7552 16814 7590
rect 16864 7610 16908 7652
rect 16864 7590 16876 7610
rect 16896 7590 16908 7610
rect 16864 7552 16908 7590
rect 16990 7610 17032 7652
rect 16990 7590 16998 7610
rect 17018 7590 17032 7610
rect 16990 7552 17032 7590
rect 17082 7610 17126 7652
rect 17082 7590 17094 7610
rect 17114 7590 17126 7610
rect 17082 7552 17126 7590
rect 9145 7433 9189 7471
rect 9145 7413 9157 7433
rect 9177 7413 9189 7433
rect 3180 7324 3192 7344
rect 3212 7324 3224 7344
rect 3180 7286 3224 7324
rect 1202 7224 1246 7262
rect 1202 7204 1214 7224
rect 1234 7204 1246 7224
rect 1202 7162 1246 7204
rect 1296 7224 1338 7262
rect 1296 7204 1310 7224
rect 1330 7204 1338 7224
rect 1296 7162 1338 7204
rect 1420 7224 1464 7262
rect 1420 7204 1432 7224
rect 1452 7204 1464 7224
rect 1420 7162 1464 7204
rect 1514 7224 1556 7262
rect 1514 7204 1528 7224
rect 1548 7204 1556 7224
rect 1514 7162 1556 7204
rect 1630 7224 1672 7262
rect 1630 7204 1638 7224
rect 1658 7204 1672 7224
rect 1630 7162 1672 7204
rect 1722 7231 1767 7262
rect 1722 7224 1766 7231
rect 1722 7204 1734 7224
rect 1754 7204 1766 7224
rect 1722 7162 1766 7204
rect 7024 7357 7068 7399
rect 7024 7337 7036 7357
rect 7056 7337 7068 7357
rect 7024 7330 7068 7337
rect 7023 7299 7068 7330
rect 7118 7357 7160 7399
rect 7118 7337 7132 7357
rect 7152 7337 7160 7357
rect 7118 7299 7160 7337
rect 7234 7357 7276 7399
rect 7234 7337 7242 7357
rect 7262 7337 7276 7357
rect 7234 7299 7276 7337
rect 7326 7357 7370 7399
rect 7326 7337 7338 7357
rect 7358 7337 7370 7357
rect 7326 7299 7370 7337
rect 7452 7357 7494 7399
rect 7452 7337 7460 7357
rect 7480 7337 7494 7357
rect 7452 7299 7494 7337
rect 7544 7357 7588 7399
rect 9145 7371 9189 7413
rect 9239 7433 9281 7471
rect 9239 7413 9253 7433
rect 9273 7413 9281 7433
rect 9239 7371 9281 7413
rect 9363 7433 9407 7471
rect 9363 7413 9375 7433
rect 9395 7413 9407 7433
rect 9363 7371 9407 7413
rect 9457 7433 9499 7471
rect 9457 7413 9471 7433
rect 9491 7413 9499 7433
rect 9457 7371 9499 7413
rect 9573 7433 9615 7471
rect 9573 7413 9581 7433
rect 9601 7413 9615 7433
rect 9573 7371 9615 7413
rect 9665 7440 9710 7471
rect 9665 7433 9709 7440
rect 9665 7413 9677 7433
rect 9697 7413 9709 7433
rect 9665 7371 9709 7413
rect 13509 7446 13553 7484
rect 13509 7426 13521 7446
rect 13541 7426 13553 7446
rect 7544 7337 7556 7357
rect 7576 7337 7588 7357
rect 7544 7299 7588 7337
rect 5566 7237 5610 7275
rect 5566 7217 5578 7237
rect 5598 7217 5610 7237
rect 3458 7160 3502 7202
rect 3458 7140 3470 7160
rect 3490 7140 3502 7160
rect 3458 7133 3502 7140
rect 3457 7102 3502 7133
rect 3552 7160 3594 7202
rect 3552 7140 3566 7160
rect 3586 7140 3594 7160
rect 3552 7102 3594 7140
rect 3668 7160 3710 7202
rect 3668 7140 3676 7160
rect 3696 7140 3710 7160
rect 3668 7102 3710 7140
rect 3760 7160 3804 7202
rect 3760 7140 3772 7160
rect 3792 7140 3804 7160
rect 3760 7102 3804 7140
rect 3886 7160 3928 7202
rect 3886 7140 3894 7160
rect 3914 7140 3928 7160
rect 3886 7102 3928 7140
rect 3978 7160 4022 7202
rect 5566 7175 5610 7217
rect 5660 7237 5702 7275
rect 5660 7217 5674 7237
rect 5694 7217 5702 7237
rect 5660 7175 5702 7217
rect 5784 7237 5828 7275
rect 5784 7217 5796 7237
rect 5816 7217 5828 7237
rect 5784 7175 5828 7217
rect 5878 7237 5920 7275
rect 5878 7217 5892 7237
rect 5912 7217 5920 7237
rect 5878 7175 5920 7217
rect 5994 7237 6036 7275
rect 5994 7217 6002 7237
rect 6022 7217 6036 7237
rect 5994 7175 6036 7217
rect 6086 7244 6131 7275
rect 6086 7237 6130 7244
rect 6086 7217 6098 7237
rect 6118 7217 6130 7237
rect 6086 7175 6130 7217
rect 11401 7369 11445 7411
rect 11401 7349 11413 7369
rect 11433 7349 11445 7369
rect 11401 7342 11445 7349
rect 11400 7311 11445 7342
rect 11495 7369 11537 7411
rect 11495 7349 11509 7369
rect 11529 7349 11537 7369
rect 11495 7311 11537 7349
rect 11611 7369 11653 7411
rect 11611 7349 11619 7369
rect 11639 7349 11653 7369
rect 11611 7311 11653 7349
rect 11703 7369 11747 7411
rect 11703 7349 11715 7369
rect 11735 7349 11747 7369
rect 11703 7311 11747 7349
rect 11829 7369 11871 7411
rect 11829 7349 11837 7369
rect 11857 7349 11871 7369
rect 11829 7311 11871 7349
rect 11921 7369 11965 7411
rect 13509 7384 13553 7426
rect 13603 7446 13645 7484
rect 13603 7426 13617 7446
rect 13637 7426 13645 7446
rect 13603 7384 13645 7426
rect 13727 7446 13771 7484
rect 13727 7426 13739 7446
rect 13759 7426 13771 7446
rect 13727 7384 13771 7426
rect 13821 7446 13863 7484
rect 13821 7426 13835 7446
rect 13855 7426 13863 7446
rect 13821 7384 13863 7426
rect 13937 7446 13979 7484
rect 13937 7426 13945 7446
rect 13965 7426 13979 7446
rect 13937 7384 13979 7426
rect 14029 7453 14074 7484
rect 14029 7446 14073 7453
rect 14029 7426 14041 7446
rect 14061 7426 14073 7446
rect 14029 7384 14073 7426
rect 11921 7349 11933 7369
rect 11953 7349 11965 7369
rect 11921 7311 11965 7349
rect 9943 7249 9987 7287
rect 9943 7229 9955 7249
rect 9975 7229 9987 7249
rect 3978 7140 3990 7160
rect 4010 7140 4022 7160
rect 3978 7102 4022 7140
rect 7822 7173 7866 7215
rect 7822 7153 7834 7173
rect 7854 7153 7866 7173
rect 7822 7146 7866 7153
rect 7821 7115 7866 7146
rect 7916 7173 7958 7215
rect 7916 7153 7930 7173
rect 7950 7153 7958 7173
rect 7916 7115 7958 7153
rect 8032 7173 8074 7215
rect 8032 7153 8040 7173
rect 8060 7153 8074 7173
rect 8032 7115 8074 7153
rect 8124 7173 8168 7215
rect 8124 7153 8136 7173
rect 8156 7153 8168 7173
rect 8124 7115 8168 7153
rect 8250 7173 8292 7215
rect 8250 7153 8258 7173
rect 8278 7153 8292 7173
rect 8250 7115 8292 7153
rect 8342 7173 8386 7215
rect 9943 7187 9987 7229
rect 10037 7249 10079 7287
rect 10037 7229 10051 7249
rect 10071 7229 10079 7249
rect 10037 7187 10079 7229
rect 10161 7249 10205 7287
rect 10161 7229 10173 7249
rect 10193 7229 10205 7249
rect 10161 7187 10205 7229
rect 10255 7249 10297 7287
rect 10255 7229 10269 7249
rect 10289 7229 10297 7249
rect 10255 7187 10297 7229
rect 10371 7249 10413 7287
rect 10371 7229 10379 7249
rect 10399 7229 10413 7249
rect 10371 7187 10413 7229
rect 10463 7256 10508 7287
rect 10463 7249 10507 7256
rect 10463 7229 10475 7249
rect 10495 7229 10507 7249
rect 10463 7187 10507 7229
rect 15765 7382 15809 7424
rect 15765 7362 15777 7382
rect 15797 7362 15809 7382
rect 15765 7355 15809 7362
rect 15764 7324 15809 7355
rect 15859 7382 15901 7424
rect 15859 7362 15873 7382
rect 15893 7362 15901 7382
rect 15859 7324 15901 7362
rect 15975 7382 16017 7424
rect 15975 7362 15983 7382
rect 16003 7362 16017 7382
rect 15975 7324 16017 7362
rect 16067 7382 16111 7424
rect 16067 7362 16079 7382
rect 16099 7362 16111 7382
rect 16067 7324 16111 7362
rect 16193 7382 16235 7424
rect 16193 7362 16201 7382
rect 16221 7362 16235 7382
rect 16193 7324 16235 7362
rect 16285 7382 16329 7424
rect 16285 7362 16297 7382
rect 16317 7362 16329 7382
rect 16285 7324 16329 7362
rect 14307 7262 14351 7300
rect 14307 7242 14319 7262
rect 14339 7242 14351 7262
rect 8342 7153 8354 7173
rect 8374 7153 8386 7173
rect 8342 7115 8386 7153
rect 405 6996 449 7034
rect 405 6976 417 6996
rect 437 6976 449 6996
rect 405 6934 449 6976
rect 499 6996 541 7034
rect 499 6976 513 6996
rect 533 6976 541 6996
rect 499 6934 541 6976
rect 623 6996 667 7034
rect 623 6976 635 6996
rect 655 6976 667 6996
rect 623 6934 667 6976
rect 717 6996 759 7034
rect 717 6976 731 6996
rect 751 6976 759 6996
rect 717 6934 759 6976
rect 833 6996 875 7034
rect 833 6976 841 6996
rect 861 6976 875 6996
rect 833 6934 875 6976
rect 925 7003 970 7034
rect 925 6996 969 7003
rect 925 6976 937 6996
rect 957 6976 969 6996
rect 12199 7185 12243 7227
rect 12199 7165 12211 7185
rect 12231 7165 12243 7185
rect 12199 7158 12243 7165
rect 12198 7127 12243 7158
rect 12293 7185 12335 7227
rect 12293 7165 12307 7185
rect 12327 7165 12335 7185
rect 12293 7127 12335 7165
rect 12409 7185 12451 7227
rect 12409 7165 12417 7185
rect 12437 7165 12451 7185
rect 12409 7127 12451 7165
rect 12501 7185 12545 7227
rect 12501 7165 12513 7185
rect 12533 7165 12545 7185
rect 12501 7127 12545 7165
rect 12627 7185 12669 7227
rect 12627 7165 12635 7185
rect 12655 7165 12669 7185
rect 12627 7127 12669 7165
rect 12719 7185 12763 7227
rect 14307 7200 14351 7242
rect 14401 7262 14443 7300
rect 14401 7242 14415 7262
rect 14435 7242 14443 7262
rect 14401 7200 14443 7242
rect 14525 7262 14569 7300
rect 14525 7242 14537 7262
rect 14557 7242 14569 7262
rect 14525 7200 14569 7242
rect 14619 7262 14661 7300
rect 14619 7242 14633 7262
rect 14653 7242 14661 7262
rect 14619 7200 14661 7242
rect 14735 7262 14777 7300
rect 14735 7242 14743 7262
rect 14763 7242 14777 7262
rect 14735 7200 14777 7242
rect 14827 7269 14872 7300
rect 14827 7262 14871 7269
rect 14827 7242 14839 7262
rect 14859 7242 14871 7262
rect 14827 7200 14871 7242
rect 12719 7165 12731 7185
rect 12751 7165 12763 7185
rect 12719 7127 12763 7165
rect 4769 7009 4813 7047
rect 925 6934 969 6976
rect 2495 6936 2539 6978
rect 2495 6916 2507 6936
rect 2527 6916 2539 6936
rect 2495 6909 2539 6916
rect 2494 6878 2539 6909
rect 2589 6936 2631 6978
rect 2589 6916 2603 6936
rect 2623 6916 2631 6936
rect 2589 6878 2631 6916
rect 2705 6936 2747 6978
rect 2705 6916 2713 6936
rect 2733 6916 2747 6936
rect 2705 6878 2747 6916
rect 2797 6936 2841 6978
rect 2797 6916 2809 6936
rect 2829 6916 2841 6936
rect 2797 6878 2841 6916
rect 2923 6936 2965 6978
rect 2923 6916 2931 6936
rect 2951 6916 2965 6936
rect 2923 6878 2965 6916
rect 3015 6936 3059 6978
rect 4769 6989 4781 7009
rect 4801 6989 4813 7009
rect 3015 6916 3027 6936
rect 3047 6916 3059 6936
rect 4769 6947 4813 6989
rect 4863 7009 4905 7047
rect 4863 6989 4877 7009
rect 4897 6989 4905 7009
rect 4863 6947 4905 6989
rect 4987 7009 5031 7047
rect 4987 6989 4999 7009
rect 5019 6989 5031 7009
rect 4987 6947 5031 6989
rect 5081 7009 5123 7047
rect 5081 6989 5095 7009
rect 5115 6989 5123 7009
rect 5081 6947 5123 6989
rect 5197 7009 5239 7047
rect 5197 6989 5205 7009
rect 5225 6989 5239 7009
rect 5197 6947 5239 6989
rect 5289 7016 5334 7047
rect 5289 7009 5333 7016
rect 5289 6989 5301 7009
rect 5321 6989 5333 7009
rect 16563 7198 16607 7240
rect 16563 7178 16575 7198
rect 16595 7178 16607 7198
rect 16563 7171 16607 7178
rect 16562 7140 16607 7171
rect 16657 7198 16699 7240
rect 16657 7178 16671 7198
rect 16691 7178 16699 7198
rect 16657 7140 16699 7178
rect 16773 7198 16815 7240
rect 16773 7178 16781 7198
rect 16801 7178 16815 7198
rect 16773 7140 16815 7178
rect 16865 7198 16909 7240
rect 16865 7178 16877 7198
rect 16897 7178 16909 7198
rect 16865 7140 16909 7178
rect 16991 7198 17033 7240
rect 16991 7178 16999 7198
rect 17019 7178 17033 7198
rect 16991 7140 17033 7178
rect 17083 7198 17127 7240
rect 17083 7178 17095 7198
rect 17115 7178 17127 7198
rect 17083 7140 17127 7178
rect 9146 7021 9190 7059
rect 5289 6947 5333 6989
rect 6859 6949 6903 6991
rect 3015 6878 3059 6916
rect 6859 6929 6871 6949
rect 6891 6929 6903 6949
rect 6859 6922 6903 6929
rect 6858 6891 6903 6922
rect 6953 6949 6995 6991
rect 6953 6929 6967 6949
rect 6987 6929 6995 6949
rect 6953 6891 6995 6929
rect 7069 6949 7111 6991
rect 7069 6929 7077 6949
rect 7097 6929 7111 6949
rect 7069 6891 7111 6929
rect 7161 6949 7205 6991
rect 7161 6929 7173 6949
rect 7193 6929 7205 6949
rect 7161 6891 7205 6929
rect 7287 6949 7329 6991
rect 7287 6929 7295 6949
rect 7315 6929 7329 6949
rect 7287 6891 7329 6929
rect 7379 6949 7423 6991
rect 9146 7001 9158 7021
rect 9178 7001 9190 7021
rect 7379 6929 7391 6949
rect 7411 6929 7423 6949
rect 9146 6959 9190 7001
rect 9240 7021 9282 7059
rect 9240 7001 9254 7021
rect 9274 7001 9282 7021
rect 9240 6959 9282 7001
rect 9364 7021 9408 7059
rect 9364 7001 9376 7021
rect 9396 7001 9408 7021
rect 9364 6959 9408 7001
rect 9458 7021 9500 7059
rect 9458 7001 9472 7021
rect 9492 7001 9500 7021
rect 9458 6959 9500 7001
rect 9574 7021 9616 7059
rect 9574 7001 9582 7021
rect 9602 7001 9616 7021
rect 9574 6959 9616 7001
rect 9666 7028 9711 7059
rect 9666 7021 9710 7028
rect 9666 7001 9678 7021
rect 9698 7001 9710 7021
rect 13510 7034 13554 7072
rect 9666 6959 9710 7001
rect 11236 6961 11280 7003
rect 7379 6891 7423 6929
rect 11236 6941 11248 6961
rect 11268 6941 11280 6961
rect 11236 6934 11280 6941
rect 11235 6903 11280 6934
rect 11330 6961 11372 7003
rect 11330 6941 11344 6961
rect 11364 6941 11372 6961
rect 11330 6903 11372 6941
rect 11446 6961 11488 7003
rect 11446 6941 11454 6961
rect 11474 6941 11488 6961
rect 11446 6903 11488 6941
rect 11538 6961 11582 7003
rect 11538 6941 11550 6961
rect 11570 6941 11582 6961
rect 11538 6903 11582 6941
rect 11664 6961 11706 7003
rect 11664 6941 11672 6961
rect 11692 6941 11706 6961
rect 11664 6903 11706 6941
rect 11756 6961 11800 7003
rect 13510 7014 13522 7034
rect 13542 7014 13554 7034
rect 11756 6941 11768 6961
rect 11788 6941 11800 6961
rect 13510 6972 13554 7014
rect 13604 7034 13646 7072
rect 13604 7014 13618 7034
rect 13638 7014 13646 7034
rect 13604 6972 13646 7014
rect 13728 7034 13772 7072
rect 13728 7014 13740 7034
rect 13760 7014 13772 7034
rect 13728 6972 13772 7014
rect 13822 7034 13864 7072
rect 13822 7014 13836 7034
rect 13856 7014 13864 7034
rect 13822 6972 13864 7014
rect 13938 7034 13980 7072
rect 13938 7014 13946 7034
rect 13966 7014 13980 7034
rect 13938 6972 13980 7014
rect 14030 7041 14075 7072
rect 14030 7034 14074 7041
rect 14030 7014 14042 7034
rect 14062 7014 14074 7034
rect 14030 6972 14074 7014
rect 15600 6974 15644 7016
rect 11756 6903 11800 6941
rect 15600 6954 15612 6974
rect 15632 6954 15644 6974
rect 15600 6947 15644 6954
rect 15599 6916 15644 6947
rect 15694 6974 15736 7016
rect 15694 6954 15708 6974
rect 15728 6954 15736 6974
rect 15694 6916 15736 6954
rect 15810 6974 15852 7016
rect 15810 6954 15818 6974
rect 15838 6954 15852 6974
rect 15810 6916 15852 6954
rect 15902 6974 15946 7016
rect 15902 6954 15914 6974
rect 15934 6954 15946 6974
rect 15902 6916 15946 6954
rect 16028 6974 16070 7016
rect 16028 6954 16036 6974
rect 16056 6954 16070 6974
rect 16028 6916 16070 6954
rect 16120 6974 16164 7016
rect 16120 6954 16132 6974
rect 16152 6954 16164 6974
rect 16120 6916 16164 6954
rect 1347 6614 1391 6652
rect 1347 6594 1359 6614
rect 1379 6594 1391 6614
rect 1347 6552 1391 6594
rect 1441 6614 1483 6652
rect 1441 6594 1455 6614
rect 1475 6594 1483 6614
rect 1441 6552 1483 6594
rect 1565 6614 1609 6652
rect 1565 6594 1577 6614
rect 1597 6594 1609 6614
rect 1565 6552 1609 6594
rect 1659 6614 1701 6652
rect 1659 6594 1673 6614
rect 1693 6594 1701 6614
rect 1659 6552 1701 6594
rect 1775 6614 1817 6652
rect 1775 6594 1783 6614
rect 1803 6594 1817 6614
rect 1775 6552 1817 6594
rect 1867 6621 1912 6652
rect 1867 6614 1911 6621
rect 1867 6594 1879 6614
rect 1899 6594 1911 6614
rect 5711 6627 5755 6665
rect 1867 6552 1911 6594
rect 3437 6554 3481 6596
rect 3437 6534 3449 6554
rect 3469 6534 3481 6554
rect 3437 6527 3481 6534
rect 3436 6496 3481 6527
rect 3531 6554 3573 6596
rect 3531 6534 3545 6554
rect 3565 6534 3573 6554
rect 3531 6496 3573 6534
rect 3647 6554 3689 6596
rect 3647 6534 3655 6554
rect 3675 6534 3689 6554
rect 3647 6496 3689 6534
rect 3739 6554 3783 6596
rect 3739 6534 3751 6554
rect 3771 6534 3783 6554
rect 3739 6496 3783 6534
rect 3865 6554 3907 6596
rect 3865 6534 3873 6554
rect 3893 6534 3907 6554
rect 3865 6496 3907 6534
rect 3957 6554 4001 6596
rect 5711 6607 5723 6627
rect 5743 6607 5755 6627
rect 3957 6534 3969 6554
rect 3989 6534 4001 6554
rect 5711 6565 5755 6607
rect 5805 6627 5847 6665
rect 5805 6607 5819 6627
rect 5839 6607 5847 6627
rect 5805 6565 5847 6607
rect 5929 6627 5973 6665
rect 5929 6607 5941 6627
rect 5961 6607 5973 6627
rect 5929 6565 5973 6607
rect 6023 6627 6065 6665
rect 6023 6607 6037 6627
rect 6057 6607 6065 6627
rect 6023 6565 6065 6607
rect 6139 6627 6181 6665
rect 6139 6607 6147 6627
rect 6167 6607 6181 6627
rect 6139 6565 6181 6607
rect 6231 6634 6276 6665
rect 6231 6627 6275 6634
rect 6231 6607 6243 6627
rect 6263 6607 6275 6627
rect 10088 6639 10132 6677
rect 6231 6565 6275 6607
rect 7801 6567 7845 6609
rect 3957 6496 4001 6534
rect 7801 6547 7813 6567
rect 7833 6547 7845 6567
rect 7801 6540 7845 6547
rect 7800 6509 7845 6540
rect 7895 6567 7937 6609
rect 7895 6547 7909 6567
rect 7929 6547 7937 6567
rect 7895 6509 7937 6547
rect 8011 6567 8053 6609
rect 8011 6547 8019 6567
rect 8039 6547 8053 6567
rect 8011 6509 8053 6547
rect 8103 6567 8147 6609
rect 8103 6547 8115 6567
rect 8135 6547 8147 6567
rect 8103 6509 8147 6547
rect 8229 6567 8271 6609
rect 8229 6547 8237 6567
rect 8257 6547 8271 6567
rect 8229 6509 8271 6547
rect 8321 6567 8365 6609
rect 10088 6619 10100 6639
rect 10120 6619 10132 6639
rect 8321 6547 8333 6567
rect 8353 6547 8365 6567
rect 10088 6577 10132 6619
rect 10182 6639 10224 6677
rect 10182 6619 10196 6639
rect 10216 6619 10224 6639
rect 10182 6577 10224 6619
rect 10306 6639 10350 6677
rect 10306 6619 10318 6639
rect 10338 6619 10350 6639
rect 10306 6577 10350 6619
rect 10400 6639 10442 6677
rect 10400 6619 10414 6639
rect 10434 6619 10442 6639
rect 10400 6577 10442 6619
rect 10516 6639 10558 6677
rect 10516 6619 10524 6639
rect 10544 6619 10558 6639
rect 10516 6577 10558 6619
rect 10608 6646 10653 6677
rect 10608 6639 10652 6646
rect 10608 6619 10620 6639
rect 10640 6619 10652 6639
rect 14452 6652 14496 6690
rect 10608 6577 10652 6619
rect 12178 6579 12222 6621
rect 8321 6509 8365 6547
rect 384 6390 428 6428
rect 384 6370 396 6390
rect 416 6370 428 6390
rect 384 6328 428 6370
rect 478 6390 520 6428
rect 478 6370 492 6390
rect 512 6370 520 6390
rect 478 6328 520 6370
rect 602 6390 646 6428
rect 602 6370 614 6390
rect 634 6370 646 6390
rect 602 6328 646 6370
rect 696 6390 738 6428
rect 696 6370 710 6390
rect 730 6370 738 6390
rect 696 6328 738 6370
rect 812 6390 854 6428
rect 812 6370 820 6390
rect 840 6370 854 6390
rect 812 6328 854 6370
rect 904 6397 949 6428
rect 904 6390 948 6397
rect 904 6370 916 6390
rect 936 6370 948 6390
rect 904 6328 948 6370
rect 12178 6559 12190 6579
rect 12210 6559 12222 6579
rect 12178 6552 12222 6559
rect 12177 6521 12222 6552
rect 12272 6579 12314 6621
rect 12272 6559 12286 6579
rect 12306 6559 12314 6579
rect 12272 6521 12314 6559
rect 12388 6579 12430 6621
rect 12388 6559 12396 6579
rect 12416 6559 12430 6579
rect 12388 6521 12430 6559
rect 12480 6579 12524 6621
rect 12480 6559 12492 6579
rect 12512 6559 12524 6579
rect 12480 6521 12524 6559
rect 12606 6579 12648 6621
rect 12606 6559 12614 6579
rect 12634 6559 12648 6579
rect 12606 6521 12648 6559
rect 12698 6579 12742 6621
rect 14452 6632 14464 6652
rect 14484 6632 14496 6652
rect 12698 6559 12710 6579
rect 12730 6559 12742 6579
rect 14452 6590 14496 6632
rect 14546 6652 14588 6690
rect 14546 6632 14560 6652
rect 14580 6632 14588 6652
rect 14546 6590 14588 6632
rect 14670 6652 14714 6690
rect 14670 6632 14682 6652
rect 14702 6632 14714 6652
rect 14670 6590 14714 6632
rect 14764 6652 14806 6690
rect 14764 6632 14778 6652
rect 14798 6632 14806 6652
rect 14764 6590 14806 6632
rect 14880 6652 14922 6690
rect 14880 6632 14888 6652
rect 14908 6632 14922 6652
rect 14880 6590 14922 6632
rect 14972 6659 15017 6690
rect 14972 6652 15016 6659
rect 14972 6632 14984 6652
rect 15004 6632 15016 6652
rect 14972 6590 15016 6632
rect 16542 6592 16586 6634
rect 12698 6521 12742 6559
rect 4748 6403 4792 6441
rect 4748 6383 4760 6403
rect 4780 6383 4792 6403
rect 2640 6326 2684 6368
rect 2640 6306 2652 6326
rect 2672 6306 2684 6326
rect 2640 6299 2684 6306
rect 2639 6268 2684 6299
rect 2734 6326 2776 6368
rect 2734 6306 2748 6326
rect 2768 6306 2776 6326
rect 2734 6268 2776 6306
rect 2850 6326 2892 6368
rect 2850 6306 2858 6326
rect 2878 6306 2892 6326
rect 2850 6268 2892 6306
rect 2942 6326 2986 6368
rect 2942 6306 2954 6326
rect 2974 6306 2986 6326
rect 2942 6268 2986 6306
rect 3068 6326 3110 6368
rect 3068 6306 3076 6326
rect 3096 6306 3110 6326
rect 3068 6268 3110 6306
rect 3160 6326 3204 6368
rect 4748 6341 4792 6383
rect 4842 6403 4884 6441
rect 4842 6383 4856 6403
rect 4876 6383 4884 6403
rect 4842 6341 4884 6383
rect 4966 6403 5010 6441
rect 4966 6383 4978 6403
rect 4998 6383 5010 6403
rect 4966 6341 5010 6383
rect 5060 6403 5102 6441
rect 5060 6383 5074 6403
rect 5094 6383 5102 6403
rect 5060 6341 5102 6383
rect 5176 6403 5218 6441
rect 5176 6383 5184 6403
rect 5204 6383 5218 6403
rect 5176 6341 5218 6383
rect 5268 6410 5313 6441
rect 5268 6403 5312 6410
rect 5268 6383 5280 6403
rect 5300 6383 5312 6403
rect 5268 6341 5312 6383
rect 16542 6572 16554 6592
rect 16574 6572 16586 6592
rect 16542 6565 16586 6572
rect 16541 6534 16586 6565
rect 16636 6592 16678 6634
rect 16636 6572 16650 6592
rect 16670 6572 16678 6592
rect 16636 6534 16678 6572
rect 16752 6592 16794 6634
rect 16752 6572 16760 6592
rect 16780 6572 16794 6592
rect 16752 6534 16794 6572
rect 16844 6592 16888 6634
rect 16844 6572 16856 6592
rect 16876 6572 16888 6592
rect 16844 6534 16888 6572
rect 16970 6592 17012 6634
rect 16970 6572 16978 6592
rect 16998 6572 17012 6592
rect 16970 6534 17012 6572
rect 17062 6592 17106 6634
rect 17062 6572 17074 6592
rect 17094 6572 17106 6592
rect 17062 6534 17106 6572
rect 9125 6415 9169 6453
rect 9125 6395 9137 6415
rect 9157 6395 9169 6415
rect 3160 6306 3172 6326
rect 3192 6306 3204 6326
rect 3160 6268 3204 6306
rect 1182 6206 1226 6244
rect 1182 6186 1194 6206
rect 1214 6186 1226 6206
rect 1182 6144 1226 6186
rect 1276 6206 1318 6244
rect 1276 6186 1290 6206
rect 1310 6186 1318 6206
rect 1276 6144 1318 6186
rect 1400 6206 1444 6244
rect 1400 6186 1412 6206
rect 1432 6186 1444 6206
rect 1400 6144 1444 6186
rect 1494 6206 1536 6244
rect 1494 6186 1508 6206
rect 1528 6186 1536 6206
rect 1494 6144 1536 6186
rect 1610 6206 1652 6244
rect 1610 6186 1618 6206
rect 1638 6186 1652 6206
rect 1610 6144 1652 6186
rect 1702 6213 1747 6244
rect 1702 6206 1746 6213
rect 1702 6186 1714 6206
rect 1734 6186 1746 6206
rect 1702 6144 1746 6186
rect 7004 6339 7048 6381
rect 7004 6319 7016 6339
rect 7036 6319 7048 6339
rect 7004 6312 7048 6319
rect 7003 6281 7048 6312
rect 7098 6339 7140 6381
rect 7098 6319 7112 6339
rect 7132 6319 7140 6339
rect 7098 6281 7140 6319
rect 7214 6339 7256 6381
rect 7214 6319 7222 6339
rect 7242 6319 7256 6339
rect 7214 6281 7256 6319
rect 7306 6339 7350 6381
rect 7306 6319 7318 6339
rect 7338 6319 7350 6339
rect 7306 6281 7350 6319
rect 7432 6339 7474 6381
rect 7432 6319 7440 6339
rect 7460 6319 7474 6339
rect 7432 6281 7474 6319
rect 7524 6339 7568 6381
rect 9125 6353 9169 6395
rect 9219 6415 9261 6453
rect 9219 6395 9233 6415
rect 9253 6395 9261 6415
rect 9219 6353 9261 6395
rect 9343 6415 9387 6453
rect 9343 6395 9355 6415
rect 9375 6395 9387 6415
rect 9343 6353 9387 6395
rect 9437 6415 9479 6453
rect 9437 6395 9451 6415
rect 9471 6395 9479 6415
rect 9437 6353 9479 6395
rect 9553 6415 9595 6453
rect 9553 6395 9561 6415
rect 9581 6395 9595 6415
rect 9553 6353 9595 6395
rect 9645 6422 9690 6453
rect 9645 6415 9689 6422
rect 9645 6395 9657 6415
rect 9677 6395 9689 6415
rect 9645 6353 9689 6395
rect 13489 6428 13533 6466
rect 13489 6408 13501 6428
rect 13521 6408 13533 6428
rect 7524 6319 7536 6339
rect 7556 6319 7568 6339
rect 7524 6281 7568 6319
rect 5546 6219 5590 6257
rect 5546 6199 5558 6219
rect 5578 6199 5590 6219
rect 3438 6142 3482 6184
rect 3438 6122 3450 6142
rect 3470 6122 3482 6142
rect 3438 6115 3482 6122
rect 3437 6084 3482 6115
rect 3532 6142 3574 6184
rect 3532 6122 3546 6142
rect 3566 6122 3574 6142
rect 3532 6084 3574 6122
rect 3648 6142 3690 6184
rect 3648 6122 3656 6142
rect 3676 6122 3690 6142
rect 3648 6084 3690 6122
rect 3740 6142 3784 6184
rect 3740 6122 3752 6142
rect 3772 6122 3784 6142
rect 3740 6084 3784 6122
rect 3866 6142 3908 6184
rect 3866 6122 3874 6142
rect 3894 6122 3908 6142
rect 3866 6084 3908 6122
rect 3958 6142 4002 6184
rect 5546 6157 5590 6199
rect 5640 6219 5682 6257
rect 5640 6199 5654 6219
rect 5674 6199 5682 6219
rect 5640 6157 5682 6199
rect 5764 6219 5808 6257
rect 5764 6199 5776 6219
rect 5796 6199 5808 6219
rect 5764 6157 5808 6199
rect 5858 6219 5900 6257
rect 5858 6199 5872 6219
rect 5892 6199 5900 6219
rect 5858 6157 5900 6199
rect 5974 6219 6016 6257
rect 5974 6199 5982 6219
rect 6002 6199 6016 6219
rect 5974 6157 6016 6199
rect 6066 6226 6111 6257
rect 6066 6219 6110 6226
rect 6066 6199 6078 6219
rect 6098 6199 6110 6219
rect 6066 6157 6110 6199
rect 11381 6351 11425 6393
rect 11381 6331 11393 6351
rect 11413 6331 11425 6351
rect 11381 6324 11425 6331
rect 11380 6293 11425 6324
rect 11475 6351 11517 6393
rect 11475 6331 11489 6351
rect 11509 6331 11517 6351
rect 11475 6293 11517 6331
rect 11591 6351 11633 6393
rect 11591 6331 11599 6351
rect 11619 6331 11633 6351
rect 11591 6293 11633 6331
rect 11683 6351 11727 6393
rect 11683 6331 11695 6351
rect 11715 6331 11727 6351
rect 11683 6293 11727 6331
rect 11809 6351 11851 6393
rect 11809 6331 11817 6351
rect 11837 6331 11851 6351
rect 11809 6293 11851 6331
rect 11901 6351 11945 6393
rect 13489 6366 13533 6408
rect 13583 6428 13625 6466
rect 13583 6408 13597 6428
rect 13617 6408 13625 6428
rect 13583 6366 13625 6408
rect 13707 6428 13751 6466
rect 13707 6408 13719 6428
rect 13739 6408 13751 6428
rect 13707 6366 13751 6408
rect 13801 6428 13843 6466
rect 13801 6408 13815 6428
rect 13835 6408 13843 6428
rect 13801 6366 13843 6408
rect 13917 6428 13959 6466
rect 13917 6408 13925 6428
rect 13945 6408 13959 6428
rect 13917 6366 13959 6408
rect 14009 6435 14054 6466
rect 14009 6428 14053 6435
rect 14009 6408 14021 6428
rect 14041 6408 14053 6428
rect 14009 6366 14053 6408
rect 11901 6331 11913 6351
rect 11933 6331 11945 6351
rect 11901 6293 11945 6331
rect 9923 6231 9967 6269
rect 9923 6211 9935 6231
rect 9955 6211 9967 6231
rect 3958 6122 3970 6142
rect 3990 6122 4002 6142
rect 3958 6084 4002 6122
rect 7802 6155 7846 6197
rect 7802 6135 7814 6155
rect 7834 6135 7846 6155
rect 7802 6128 7846 6135
rect 7801 6097 7846 6128
rect 7896 6155 7938 6197
rect 7896 6135 7910 6155
rect 7930 6135 7938 6155
rect 7896 6097 7938 6135
rect 8012 6155 8054 6197
rect 8012 6135 8020 6155
rect 8040 6135 8054 6155
rect 8012 6097 8054 6135
rect 8104 6155 8148 6197
rect 8104 6135 8116 6155
rect 8136 6135 8148 6155
rect 8104 6097 8148 6135
rect 8230 6155 8272 6197
rect 8230 6135 8238 6155
rect 8258 6135 8272 6155
rect 8230 6097 8272 6135
rect 8322 6155 8366 6197
rect 9923 6169 9967 6211
rect 10017 6231 10059 6269
rect 10017 6211 10031 6231
rect 10051 6211 10059 6231
rect 10017 6169 10059 6211
rect 10141 6231 10185 6269
rect 10141 6211 10153 6231
rect 10173 6211 10185 6231
rect 10141 6169 10185 6211
rect 10235 6231 10277 6269
rect 10235 6211 10249 6231
rect 10269 6211 10277 6231
rect 10235 6169 10277 6211
rect 10351 6231 10393 6269
rect 10351 6211 10359 6231
rect 10379 6211 10393 6231
rect 10351 6169 10393 6211
rect 10443 6238 10488 6269
rect 10443 6231 10487 6238
rect 10443 6211 10455 6231
rect 10475 6211 10487 6231
rect 10443 6169 10487 6211
rect 15745 6364 15789 6406
rect 15745 6344 15757 6364
rect 15777 6344 15789 6364
rect 15745 6337 15789 6344
rect 15744 6306 15789 6337
rect 15839 6364 15881 6406
rect 15839 6344 15853 6364
rect 15873 6344 15881 6364
rect 15839 6306 15881 6344
rect 15955 6364 15997 6406
rect 15955 6344 15963 6364
rect 15983 6344 15997 6364
rect 15955 6306 15997 6344
rect 16047 6364 16091 6406
rect 16047 6344 16059 6364
rect 16079 6344 16091 6364
rect 16047 6306 16091 6344
rect 16173 6364 16215 6406
rect 16173 6344 16181 6364
rect 16201 6344 16215 6364
rect 16173 6306 16215 6344
rect 16265 6364 16309 6406
rect 16265 6344 16277 6364
rect 16297 6344 16309 6364
rect 16265 6306 16309 6344
rect 14287 6244 14331 6282
rect 14287 6224 14299 6244
rect 14319 6224 14331 6244
rect 8322 6135 8334 6155
rect 8354 6135 8366 6155
rect 8322 6097 8366 6135
rect 385 5978 429 6016
rect 385 5958 397 5978
rect 417 5958 429 5978
rect 385 5916 429 5958
rect 479 5978 521 6016
rect 479 5958 493 5978
rect 513 5958 521 5978
rect 479 5916 521 5958
rect 603 5978 647 6016
rect 603 5958 615 5978
rect 635 5958 647 5978
rect 603 5916 647 5958
rect 697 5978 739 6016
rect 697 5958 711 5978
rect 731 5958 739 5978
rect 697 5916 739 5958
rect 813 5978 855 6016
rect 813 5958 821 5978
rect 841 5958 855 5978
rect 813 5916 855 5958
rect 905 5985 950 6016
rect 905 5978 949 5985
rect 905 5958 917 5978
rect 937 5958 949 5978
rect 12179 6167 12223 6209
rect 12179 6147 12191 6167
rect 12211 6147 12223 6167
rect 12179 6140 12223 6147
rect 12178 6109 12223 6140
rect 12273 6167 12315 6209
rect 12273 6147 12287 6167
rect 12307 6147 12315 6167
rect 12273 6109 12315 6147
rect 12389 6167 12431 6209
rect 12389 6147 12397 6167
rect 12417 6147 12431 6167
rect 12389 6109 12431 6147
rect 12481 6167 12525 6209
rect 12481 6147 12493 6167
rect 12513 6147 12525 6167
rect 12481 6109 12525 6147
rect 12607 6167 12649 6209
rect 12607 6147 12615 6167
rect 12635 6147 12649 6167
rect 12607 6109 12649 6147
rect 12699 6167 12743 6209
rect 14287 6182 14331 6224
rect 14381 6244 14423 6282
rect 14381 6224 14395 6244
rect 14415 6224 14423 6244
rect 14381 6182 14423 6224
rect 14505 6244 14549 6282
rect 14505 6224 14517 6244
rect 14537 6224 14549 6244
rect 14505 6182 14549 6224
rect 14599 6244 14641 6282
rect 14599 6224 14613 6244
rect 14633 6224 14641 6244
rect 14599 6182 14641 6224
rect 14715 6244 14757 6282
rect 14715 6224 14723 6244
rect 14743 6224 14757 6244
rect 14715 6182 14757 6224
rect 14807 6251 14852 6282
rect 14807 6244 14851 6251
rect 14807 6224 14819 6244
rect 14839 6224 14851 6244
rect 14807 6182 14851 6224
rect 12699 6147 12711 6167
rect 12731 6147 12743 6167
rect 12699 6109 12743 6147
rect 4749 5991 4793 6029
rect 905 5916 949 5958
rect 2541 5916 2585 5958
rect 2541 5896 2553 5916
rect 2573 5896 2585 5916
rect 2541 5889 2585 5896
rect 2540 5858 2585 5889
rect 2635 5916 2677 5958
rect 2635 5896 2649 5916
rect 2669 5896 2677 5916
rect 2635 5858 2677 5896
rect 2751 5916 2793 5958
rect 2751 5896 2759 5916
rect 2779 5896 2793 5916
rect 2751 5858 2793 5896
rect 2843 5916 2887 5958
rect 2843 5896 2855 5916
rect 2875 5896 2887 5916
rect 2843 5858 2887 5896
rect 2969 5916 3011 5958
rect 2969 5896 2977 5916
rect 2997 5896 3011 5916
rect 2969 5858 3011 5896
rect 3061 5916 3105 5958
rect 4749 5971 4761 5991
rect 4781 5971 4793 5991
rect 3061 5896 3073 5916
rect 3093 5896 3105 5916
rect 4749 5929 4793 5971
rect 4843 5991 4885 6029
rect 4843 5971 4857 5991
rect 4877 5971 4885 5991
rect 4843 5929 4885 5971
rect 4967 5991 5011 6029
rect 4967 5971 4979 5991
rect 4999 5971 5011 5991
rect 4967 5929 5011 5971
rect 5061 5991 5103 6029
rect 5061 5971 5075 5991
rect 5095 5971 5103 5991
rect 5061 5929 5103 5971
rect 5177 5991 5219 6029
rect 5177 5971 5185 5991
rect 5205 5971 5219 5991
rect 5177 5929 5219 5971
rect 5269 5998 5314 6029
rect 5269 5991 5313 5998
rect 5269 5971 5281 5991
rect 5301 5971 5313 5991
rect 16543 6180 16587 6222
rect 16543 6160 16555 6180
rect 16575 6160 16587 6180
rect 16543 6153 16587 6160
rect 16542 6122 16587 6153
rect 16637 6180 16679 6222
rect 16637 6160 16651 6180
rect 16671 6160 16679 6180
rect 16637 6122 16679 6160
rect 16753 6180 16795 6222
rect 16753 6160 16761 6180
rect 16781 6160 16795 6180
rect 16753 6122 16795 6160
rect 16845 6180 16889 6222
rect 16845 6160 16857 6180
rect 16877 6160 16889 6180
rect 16845 6122 16889 6160
rect 16971 6180 17013 6222
rect 16971 6160 16979 6180
rect 16999 6160 17013 6180
rect 16971 6122 17013 6160
rect 17063 6180 17107 6222
rect 17063 6160 17075 6180
rect 17095 6160 17107 6180
rect 17063 6122 17107 6160
rect 9126 6003 9170 6041
rect 5269 5929 5313 5971
rect 6905 5929 6949 5971
rect 3061 5858 3105 5896
rect 6905 5909 6917 5929
rect 6937 5909 6949 5929
rect 6905 5902 6949 5909
rect 6904 5871 6949 5902
rect 6999 5929 7041 5971
rect 6999 5909 7013 5929
rect 7033 5909 7041 5929
rect 6999 5871 7041 5909
rect 7115 5929 7157 5971
rect 7115 5909 7123 5929
rect 7143 5909 7157 5929
rect 7115 5871 7157 5909
rect 7207 5929 7251 5971
rect 7207 5909 7219 5929
rect 7239 5909 7251 5929
rect 7207 5871 7251 5909
rect 7333 5929 7375 5971
rect 7333 5909 7341 5929
rect 7361 5909 7375 5929
rect 7333 5871 7375 5909
rect 7425 5929 7469 5971
rect 9126 5983 9138 6003
rect 9158 5983 9170 6003
rect 7425 5909 7437 5929
rect 7457 5909 7469 5929
rect 9126 5941 9170 5983
rect 9220 6003 9262 6041
rect 9220 5983 9234 6003
rect 9254 5983 9262 6003
rect 9220 5941 9262 5983
rect 9344 6003 9388 6041
rect 9344 5983 9356 6003
rect 9376 5983 9388 6003
rect 9344 5941 9388 5983
rect 9438 6003 9480 6041
rect 9438 5983 9452 6003
rect 9472 5983 9480 6003
rect 9438 5941 9480 5983
rect 9554 6003 9596 6041
rect 9554 5983 9562 6003
rect 9582 5983 9596 6003
rect 9554 5941 9596 5983
rect 9646 6010 9691 6041
rect 9646 6003 9690 6010
rect 9646 5983 9658 6003
rect 9678 5983 9690 6003
rect 13490 6016 13534 6054
rect 9646 5941 9690 5983
rect 11282 5941 11326 5983
rect 7425 5871 7469 5909
rect 11282 5921 11294 5941
rect 11314 5921 11326 5941
rect 11282 5914 11326 5921
rect 11281 5883 11326 5914
rect 11376 5941 11418 5983
rect 11376 5921 11390 5941
rect 11410 5921 11418 5941
rect 11376 5883 11418 5921
rect 11492 5941 11534 5983
rect 11492 5921 11500 5941
rect 11520 5921 11534 5941
rect 11492 5883 11534 5921
rect 11584 5941 11628 5983
rect 11584 5921 11596 5941
rect 11616 5921 11628 5941
rect 11584 5883 11628 5921
rect 11710 5941 11752 5983
rect 11710 5921 11718 5941
rect 11738 5921 11752 5941
rect 11710 5883 11752 5921
rect 11802 5941 11846 5983
rect 13490 5996 13502 6016
rect 13522 5996 13534 6016
rect 11802 5921 11814 5941
rect 11834 5921 11846 5941
rect 13490 5954 13534 5996
rect 13584 6016 13626 6054
rect 13584 5996 13598 6016
rect 13618 5996 13626 6016
rect 13584 5954 13626 5996
rect 13708 6016 13752 6054
rect 13708 5996 13720 6016
rect 13740 5996 13752 6016
rect 13708 5954 13752 5996
rect 13802 6016 13844 6054
rect 13802 5996 13816 6016
rect 13836 5996 13844 6016
rect 13802 5954 13844 5996
rect 13918 6016 13960 6054
rect 13918 5996 13926 6016
rect 13946 5996 13960 6016
rect 13918 5954 13960 5996
rect 14010 6023 14055 6054
rect 14010 6016 14054 6023
rect 14010 5996 14022 6016
rect 14042 5996 14054 6016
rect 14010 5954 14054 5996
rect 15646 5954 15690 5996
rect 11802 5883 11846 5921
rect 15646 5934 15658 5954
rect 15678 5934 15690 5954
rect 15646 5927 15690 5934
rect 15645 5896 15690 5927
rect 15740 5954 15782 5996
rect 15740 5934 15754 5954
rect 15774 5934 15782 5954
rect 15740 5896 15782 5934
rect 15856 5954 15898 5996
rect 15856 5934 15864 5954
rect 15884 5934 15898 5954
rect 15856 5896 15898 5934
rect 15948 5954 15992 5996
rect 15948 5934 15960 5954
rect 15980 5934 15992 5954
rect 15948 5896 15992 5934
rect 16074 5954 16116 5996
rect 16074 5934 16082 5954
rect 16102 5934 16116 5954
rect 16074 5896 16116 5934
rect 16166 5954 16210 5996
rect 16166 5934 16178 5954
rect 16198 5934 16210 5954
rect 16166 5896 16210 5934
rect 1264 5598 1308 5636
rect 1264 5578 1276 5598
rect 1296 5578 1308 5598
rect 1264 5536 1308 5578
rect 1358 5598 1400 5636
rect 1358 5578 1372 5598
rect 1392 5578 1400 5598
rect 1358 5536 1400 5578
rect 1482 5598 1526 5636
rect 1482 5578 1494 5598
rect 1514 5578 1526 5598
rect 1482 5536 1526 5578
rect 1576 5598 1618 5636
rect 1576 5578 1590 5598
rect 1610 5578 1618 5598
rect 1576 5536 1618 5578
rect 1692 5598 1734 5636
rect 1692 5578 1700 5598
rect 1720 5578 1734 5598
rect 1692 5536 1734 5578
rect 1784 5605 1829 5636
rect 1784 5598 1828 5605
rect 1784 5578 1796 5598
rect 1816 5578 1828 5598
rect 5628 5611 5672 5649
rect 1784 5536 1828 5578
rect 3420 5536 3464 5578
rect 3420 5516 3432 5536
rect 3452 5516 3464 5536
rect 3420 5509 3464 5516
rect 3419 5478 3464 5509
rect 3514 5536 3556 5578
rect 3514 5516 3528 5536
rect 3548 5516 3556 5536
rect 3514 5478 3556 5516
rect 3630 5536 3672 5578
rect 3630 5516 3638 5536
rect 3658 5516 3672 5536
rect 3630 5478 3672 5516
rect 3722 5536 3766 5578
rect 3722 5516 3734 5536
rect 3754 5516 3766 5536
rect 3722 5478 3766 5516
rect 3848 5536 3890 5578
rect 3848 5516 3856 5536
rect 3876 5516 3890 5536
rect 3848 5478 3890 5516
rect 3940 5536 3984 5578
rect 5628 5591 5640 5611
rect 5660 5591 5672 5611
rect 3940 5516 3952 5536
rect 3972 5516 3984 5536
rect 5628 5549 5672 5591
rect 5722 5611 5764 5649
rect 5722 5591 5736 5611
rect 5756 5591 5764 5611
rect 5722 5549 5764 5591
rect 5846 5611 5890 5649
rect 5846 5591 5858 5611
rect 5878 5591 5890 5611
rect 5846 5549 5890 5591
rect 5940 5611 5982 5649
rect 5940 5591 5954 5611
rect 5974 5591 5982 5611
rect 5940 5549 5982 5591
rect 6056 5611 6098 5649
rect 6056 5591 6064 5611
rect 6084 5591 6098 5611
rect 6056 5549 6098 5591
rect 6148 5618 6193 5649
rect 6148 5611 6192 5618
rect 6148 5591 6160 5611
rect 6180 5591 6192 5611
rect 10005 5623 10049 5661
rect 6148 5549 6192 5591
rect 7784 5549 7828 5591
rect 3940 5478 3984 5516
rect 7784 5529 7796 5549
rect 7816 5529 7828 5549
rect 7784 5522 7828 5529
rect 7783 5491 7828 5522
rect 7878 5549 7920 5591
rect 7878 5529 7892 5549
rect 7912 5529 7920 5549
rect 7878 5491 7920 5529
rect 7994 5549 8036 5591
rect 7994 5529 8002 5549
rect 8022 5529 8036 5549
rect 7994 5491 8036 5529
rect 8086 5549 8130 5591
rect 8086 5529 8098 5549
rect 8118 5529 8130 5549
rect 8086 5491 8130 5529
rect 8212 5549 8254 5591
rect 8212 5529 8220 5549
rect 8240 5529 8254 5549
rect 8212 5491 8254 5529
rect 8304 5549 8348 5591
rect 10005 5603 10017 5623
rect 10037 5603 10049 5623
rect 8304 5529 8316 5549
rect 8336 5529 8348 5549
rect 10005 5561 10049 5603
rect 10099 5623 10141 5661
rect 10099 5603 10113 5623
rect 10133 5603 10141 5623
rect 10099 5561 10141 5603
rect 10223 5623 10267 5661
rect 10223 5603 10235 5623
rect 10255 5603 10267 5623
rect 10223 5561 10267 5603
rect 10317 5623 10359 5661
rect 10317 5603 10331 5623
rect 10351 5603 10359 5623
rect 10317 5561 10359 5603
rect 10433 5623 10475 5661
rect 10433 5603 10441 5623
rect 10461 5603 10475 5623
rect 10433 5561 10475 5603
rect 10525 5630 10570 5661
rect 10525 5623 10569 5630
rect 10525 5603 10537 5623
rect 10557 5603 10569 5623
rect 14369 5636 14413 5674
rect 10525 5561 10569 5603
rect 12161 5561 12205 5603
rect 8304 5491 8348 5529
rect 367 5372 411 5410
rect 367 5352 379 5372
rect 399 5352 411 5372
rect 367 5310 411 5352
rect 461 5372 503 5410
rect 461 5352 475 5372
rect 495 5352 503 5372
rect 461 5310 503 5352
rect 585 5372 629 5410
rect 585 5352 597 5372
rect 617 5352 629 5372
rect 585 5310 629 5352
rect 679 5372 721 5410
rect 679 5352 693 5372
rect 713 5352 721 5372
rect 679 5310 721 5352
rect 795 5372 837 5410
rect 795 5352 803 5372
rect 823 5352 837 5372
rect 795 5310 837 5352
rect 887 5379 932 5410
rect 887 5372 931 5379
rect 887 5352 899 5372
rect 919 5352 931 5372
rect 887 5310 931 5352
rect 12161 5541 12173 5561
rect 12193 5541 12205 5561
rect 12161 5534 12205 5541
rect 12160 5503 12205 5534
rect 12255 5561 12297 5603
rect 12255 5541 12269 5561
rect 12289 5541 12297 5561
rect 12255 5503 12297 5541
rect 12371 5561 12413 5603
rect 12371 5541 12379 5561
rect 12399 5541 12413 5561
rect 12371 5503 12413 5541
rect 12463 5561 12507 5603
rect 12463 5541 12475 5561
rect 12495 5541 12507 5561
rect 12463 5503 12507 5541
rect 12589 5561 12631 5603
rect 12589 5541 12597 5561
rect 12617 5541 12631 5561
rect 12589 5503 12631 5541
rect 12681 5561 12725 5603
rect 14369 5616 14381 5636
rect 14401 5616 14413 5636
rect 12681 5541 12693 5561
rect 12713 5541 12725 5561
rect 14369 5574 14413 5616
rect 14463 5636 14505 5674
rect 14463 5616 14477 5636
rect 14497 5616 14505 5636
rect 14463 5574 14505 5616
rect 14587 5636 14631 5674
rect 14587 5616 14599 5636
rect 14619 5616 14631 5636
rect 14587 5574 14631 5616
rect 14681 5636 14723 5674
rect 14681 5616 14695 5636
rect 14715 5616 14723 5636
rect 14681 5574 14723 5616
rect 14797 5636 14839 5674
rect 14797 5616 14805 5636
rect 14825 5616 14839 5636
rect 14797 5574 14839 5616
rect 14889 5643 14934 5674
rect 14889 5636 14933 5643
rect 14889 5616 14901 5636
rect 14921 5616 14933 5636
rect 14889 5574 14933 5616
rect 16525 5574 16569 5616
rect 12681 5503 12725 5541
rect 4731 5385 4775 5423
rect 4731 5365 4743 5385
rect 4763 5365 4775 5385
rect 2623 5308 2667 5350
rect 2623 5288 2635 5308
rect 2655 5288 2667 5308
rect 2623 5281 2667 5288
rect 2622 5250 2667 5281
rect 2717 5308 2759 5350
rect 2717 5288 2731 5308
rect 2751 5288 2759 5308
rect 2717 5250 2759 5288
rect 2833 5308 2875 5350
rect 2833 5288 2841 5308
rect 2861 5288 2875 5308
rect 2833 5250 2875 5288
rect 2925 5308 2969 5350
rect 2925 5288 2937 5308
rect 2957 5288 2969 5308
rect 2925 5250 2969 5288
rect 3051 5308 3093 5350
rect 3051 5288 3059 5308
rect 3079 5288 3093 5308
rect 3051 5250 3093 5288
rect 3143 5308 3187 5350
rect 4731 5323 4775 5365
rect 4825 5385 4867 5423
rect 4825 5365 4839 5385
rect 4859 5365 4867 5385
rect 4825 5323 4867 5365
rect 4949 5385 4993 5423
rect 4949 5365 4961 5385
rect 4981 5365 4993 5385
rect 4949 5323 4993 5365
rect 5043 5385 5085 5423
rect 5043 5365 5057 5385
rect 5077 5365 5085 5385
rect 5043 5323 5085 5365
rect 5159 5385 5201 5423
rect 5159 5365 5167 5385
rect 5187 5365 5201 5385
rect 5159 5323 5201 5365
rect 5251 5392 5296 5423
rect 5251 5385 5295 5392
rect 5251 5365 5263 5385
rect 5283 5365 5295 5385
rect 5251 5323 5295 5365
rect 16525 5554 16537 5574
rect 16557 5554 16569 5574
rect 16525 5547 16569 5554
rect 16524 5516 16569 5547
rect 16619 5574 16661 5616
rect 16619 5554 16633 5574
rect 16653 5554 16661 5574
rect 16619 5516 16661 5554
rect 16735 5574 16777 5616
rect 16735 5554 16743 5574
rect 16763 5554 16777 5574
rect 16735 5516 16777 5554
rect 16827 5574 16871 5616
rect 16827 5554 16839 5574
rect 16859 5554 16871 5574
rect 16827 5516 16871 5554
rect 16953 5574 16995 5616
rect 16953 5554 16961 5574
rect 16981 5554 16995 5574
rect 16953 5516 16995 5554
rect 17045 5574 17089 5616
rect 17045 5554 17057 5574
rect 17077 5554 17089 5574
rect 17045 5516 17089 5554
rect 9108 5397 9152 5435
rect 9108 5377 9120 5397
rect 9140 5377 9152 5397
rect 3143 5288 3155 5308
rect 3175 5288 3187 5308
rect 3143 5250 3187 5288
rect 1165 5188 1209 5226
rect 1165 5168 1177 5188
rect 1197 5168 1209 5188
rect 1165 5126 1209 5168
rect 1259 5188 1301 5226
rect 1259 5168 1273 5188
rect 1293 5168 1301 5188
rect 1259 5126 1301 5168
rect 1383 5188 1427 5226
rect 1383 5168 1395 5188
rect 1415 5168 1427 5188
rect 1383 5126 1427 5168
rect 1477 5188 1519 5226
rect 1477 5168 1491 5188
rect 1511 5168 1519 5188
rect 1477 5126 1519 5168
rect 1593 5188 1635 5226
rect 1593 5168 1601 5188
rect 1621 5168 1635 5188
rect 1593 5126 1635 5168
rect 1685 5195 1730 5226
rect 1685 5188 1729 5195
rect 1685 5168 1697 5188
rect 1717 5168 1729 5188
rect 1685 5126 1729 5168
rect 6987 5321 7031 5363
rect 6987 5301 6999 5321
rect 7019 5301 7031 5321
rect 6987 5294 7031 5301
rect 6986 5263 7031 5294
rect 7081 5321 7123 5363
rect 7081 5301 7095 5321
rect 7115 5301 7123 5321
rect 7081 5263 7123 5301
rect 7197 5321 7239 5363
rect 7197 5301 7205 5321
rect 7225 5301 7239 5321
rect 7197 5263 7239 5301
rect 7289 5321 7333 5363
rect 7289 5301 7301 5321
rect 7321 5301 7333 5321
rect 7289 5263 7333 5301
rect 7415 5321 7457 5363
rect 7415 5301 7423 5321
rect 7443 5301 7457 5321
rect 7415 5263 7457 5301
rect 7507 5321 7551 5363
rect 9108 5335 9152 5377
rect 9202 5397 9244 5435
rect 9202 5377 9216 5397
rect 9236 5377 9244 5397
rect 9202 5335 9244 5377
rect 9326 5397 9370 5435
rect 9326 5377 9338 5397
rect 9358 5377 9370 5397
rect 9326 5335 9370 5377
rect 9420 5397 9462 5435
rect 9420 5377 9434 5397
rect 9454 5377 9462 5397
rect 9420 5335 9462 5377
rect 9536 5397 9578 5435
rect 9536 5377 9544 5397
rect 9564 5377 9578 5397
rect 9536 5335 9578 5377
rect 9628 5404 9673 5435
rect 9628 5397 9672 5404
rect 9628 5377 9640 5397
rect 9660 5377 9672 5397
rect 9628 5335 9672 5377
rect 13472 5410 13516 5448
rect 13472 5390 13484 5410
rect 13504 5390 13516 5410
rect 7507 5301 7519 5321
rect 7539 5301 7551 5321
rect 7507 5263 7551 5301
rect 5529 5201 5573 5239
rect 5529 5181 5541 5201
rect 5561 5181 5573 5201
rect 3421 5124 3465 5166
rect 3421 5104 3433 5124
rect 3453 5104 3465 5124
rect 3421 5097 3465 5104
rect 3420 5066 3465 5097
rect 3515 5124 3557 5166
rect 3515 5104 3529 5124
rect 3549 5104 3557 5124
rect 3515 5066 3557 5104
rect 3631 5124 3673 5166
rect 3631 5104 3639 5124
rect 3659 5104 3673 5124
rect 3631 5066 3673 5104
rect 3723 5124 3767 5166
rect 3723 5104 3735 5124
rect 3755 5104 3767 5124
rect 3723 5066 3767 5104
rect 3849 5124 3891 5166
rect 3849 5104 3857 5124
rect 3877 5104 3891 5124
rect 3849 5066 3891 5104
rect 3941 5124 3985 5166
rect 5529 5139 5573 5181
rect 5623 5201 5665 5239
rect 5623 5181 5637 5201
rect 5657 5181 5665 5201
rect 5623 5139 5665 5181
rect 5747 5201 5791 5239
rect 5747 5181 5759 5201
rect 5779 5181 5791 5201
rect 5747 5139 5791 5181
rect 5841 5201 5883 5239
rect 5841 5181 5855 5201
rect 5875 5181 5883 5201
rect 5841 5139 5883 5181
rect 5957 5201 5999 5239
rect 5957 5181 5965 5201
rect 5985 5181 5999 5201
rect 5957 5139 5999 5181
rect 6049 5208 6094 5239
rect 6049 5201 6093 5208
rect 6049 5181 6061 5201
rect 6081 5181 6093 5201
rect 6049 5139 6093 5181
rect 11364 5333 11408 5375
rect 11364 5313 11376 5333
rect 11396 5313 11408 5333
rect 11364 5306 11408 5313
rect 11363 5275 11408 5306
rect 11458 5333 11500 5375
rect 11458 5313 11472 5333
rect 11492 5313 11500 5333
rect 11458 5275 11500 5313
rect 11574 5333 11616 5375
rect 11574 5313 11582 5333
rect 11602 5313 11616 5333
rect 11574 5275 11616 5313
rect 11666 5333 11710 5375
rect 11666 5313 11678 5333
rect 11698 5313 11710 5333
rect 11666 5275 11710 5313
rect 11792 5333 11834 5375
rect 11792 5313 11800 5333
rect 11820 5313 11834 5333
rect 11792 5275 11834 5313
rect 11884 5333 11928 5375
rect 13472 5348 13516 5390
rect 13566 5410 13608 5448
rect 13566 5390 13580 5410
rect 13600 5390 13608 5410
rect 13566 5348 13608 5390
rect 13690 5410 13734 5448
rect 13690 5390 13702 5410
rect 13722 5390 13734 5410
rect 13690 5348 13734 5390
rect 13784 5410 13826 5448
rect 13784 5390 13798 5410
rect 13818 5390 13826 5410
rect 13784 5348 13826 5390
rect 13900 5410 13942 5448
rect 13900 5390 13908 5410
rect 13928 5390 13942 5410
rect 13900 5348 13942 5390
rect 13992 5417 14037 5448
rect 13992 5410 14036 5417
rect 13992 5390 14004 5410
rect 14024 5390 14036 5410
rect 13992 5348 14036 5390
rect 11884 5313 11896 5333
rect 11916 5313 11928 5333
rect 11884 5275 11928 5313
rect 9906 5213 9950 5251
rect 9906 5193 9918 5213
rect 9938 5193 9950 5213
rect 3941 5104 3953 5124
rect 3973 5104 3985 5124
rect 3941 5066 3985 5104
rect 7785 5137 7829 5179
rect 7785 5117 7797 5137
rect 7817 5117 7829 5137
rect 7785 5110 7829 5117
rect 7784 5079 7829 5110
rect 7879 5137 7921 5179
rect 7879 5117 7893 5137
rect 7913 5117 7921 5137
rect 7879 5079 7921 5117
rect 7995 5137 8037 5179
rect 7995 5117 8003 5137
rect 8023 5117 8037 5137
rect 7995 5079 8037 5117
rect 8087 5137 8131 5179
rect 8087 5117 8099 5137
rect 8119 5117 8131 5137
rect 8087 5079 8131 5117
rect 8213 5137 8255 5179
rect 8213 5117 8221 5137
rect 8241 5117 8255 5137
rect 8213 5079 8255 5117
rect 8305 5137 8349 5179
rect 9906 5151 9950 5193
rect 10000 5213 10042 5251
rect 10000 5193 10014 5213
rect 10034 5193 10042 5213
rect 10000 5151 10042 5193
rect 10124 5213 10168 5251
rect 10124 5193 10136 5213
rect 10156 5193 10168 5213
rect 10124 5151 10168 5193
rect 10218 5213 10260 5251
rect 10218 5193 10232 5213
rect 10252 5193 10260 5213
rect 10218 5151 10260 5193
rect 10334 5213 10376 5251
rect 10334 5193 10342 5213
rect 10362 5193 10376 5213
rect 10334 5151 10376 5193
rect 10426 5220 10471 5251
rect 10426 5213 10470 5220
rect 10426 5193 10438 5213
rect 10458 5193 10470 5213
rect 10426 5151 10470 5193
rect 15728 5346 15772 5388
rect 15728 5326 15740 5346
rect 15760 5326 15772 5346
rect 15728 5319 15772 5326
rect 15727 5288 15772 5319
rect 15822 5346 15864 5388
rect 15822 5326 15836 5346
rect 15856 5326 15864 5346
rect 15822 5288 15864 5326
rect 15938 5346 15980 5388
rect 15938 5326 15946 5346
rect 15966 5326 15980 5346
rect 15938 5288 15980 5326
rect 16030 5346 16074 5388
rect 16030 5326 16042 5346
rect 16062 5326 16074 5346
rect 16030 5288 16074 5326
rect 16156 5346 16198 5388
rect 16156 5326 16164 5346
rect 16184 5326 16198 5346
rect 16156 5288 16198 5326
rect 16248 5346 16292 5388
rect 16248 5326 16260 5346
rect 16280 5326 16292 5346
rect 16248 5288 16292 5326
rect 14270 5226 14314 5264
rect 14270 5206 14282 5226
rect 14302 5206 14314 5226
rect 8305 5117 8317 5137
rect 8337 5117 8349 5137
rect 8305 5079 8349 5117
rect 368 4960 412 4998
rect 368 4940 380 4960
rect 400 4940 412 4960
rect 368 4898 412 4940
rect 462 4960 504 4998
rect 462 4940 476 4960
rect 496 4940 504 4960
rect 462 4898 504 4940
rect 586 4960 630 4998
rect 586 4940 598 4960
rect 618 4940 630 4960
rect 586 4898 630 4940
rect 680 4960 722 4998
rect 680 4940 694 4960
rect 714 4940 722 4960
rect 680 4898 722 4940
rect 796 4960 838 4998
rect 796 4940 804 4960
rect 824 4940 838 4960
rect 796 4898 838 4940
rect 888 4967 933 4998
rect 888 4960 932 4967
rect 888 4940 900 4960
rect 920 4940 932 4960
rect 12162 5149 12206 5191
rect 12162 5129 12174 5149
rect 12194 5129 12206 5149
rect 12162 5122 12206 5129
rect 12161 5091 12206 5122
rect 12256 5149 12298 5191
rect 12256 5129 12270 5149
rect 12290 5129 12298 5149
rect 12256 5091 12298 5129
rect 12372 5149 12414 5191
rect 12372 5129 12380 5149
rect 12400 5129 12414 5149
rect 12372 5091 12414 5129
rect 12464 5149 12508 5191
rect 12464 5129 12476 5149
rect 12496 5129 12508 5149
rect 12464 5091 12508 5129
rect 12590 5149 12632 5191
rect 12590 5129 12598 5149
rect 12618 5129 12632 5149
rect 12590 5091 12632 5129
rect 12682 5149 12726 5191
rect 14270 5164 14314 5206
rect 14364 5226 14406 5264
rect 14364 5206 14378 5226
rect 14398 5206 14406 5226
rect 14364 5164 14406 5206
rect 14488 5226 14532 5264
rect 14488 5206 14500 5226
rect 14520 5206 14532 5226
rect 14488 5164 14532 5206
rect 14582 5226 14624 5264
rect 14582 5206 14596 5226
rect 14616 5206 14624 5226
rect 14582 5164 14624 5206
rect 14698 5226 14740 5264
rect 14698 5206 14706 5226
rect 14726 5206 14740 5226
rect 14698 5164 14740 5206
rect 14790 5233 14835 5264
rect 14790 5226 14834 5233
rect 14790 5206 14802 5226
rect 14822 5206 14834 5226
rect 14790 5164 14834 5206
rect 12682 5129 12694 5149
rect 12714 5129 12726 5149
rect 12682 5091 12726 5129
rect 4732 4973 4776 5011
rect 888 4898 932 4940
rect 2319 4902 2363 4944
rect 2319 4882 2331 4902
rect 2351 4882 2363 4902
rect 2319 4875 2363 4882
rect 2318 4844 2363 4875
rect 2413 4902 2455 4944
rect 2413 4882 2427 4902
rect 2447 4882 2455 4902
rect 2413 4844 2455 4882
rect 2529 4902 2571 4944
rect 2529 4882 2537 4902
rect 2557 4882 2571 4902
rect 2529 4844 2571 4882
rect 2621 4902 2665 4944
rect 2621 4882 2633 4902
rect 2653 4882 2665 4902
rect 2621 4844 2665 4882
rect 2747 4902 2789 4944
rect 2747 4882 2755 4902
rect 2775 4882 2789 4902
rect 2747 4844 2789 4882
rect 2839 4902 2883 4944
rect 4732 4953 4744 4973
rect 4764 4953 4776 4973
rect 2839 4882 2851 4902
rect 2871 4882 2883 4902
rect 4732 4911 4776 4953
rect 4826 4973 4868 5011
rect 4826 4953 4840 4973
rect 4860 4953 4868 4973
rect 4826 4911 4868 4953
rect 4950 4973 4994 5011
rect 4950 4953 4962 4973
rect 4982 4953 4994 4973
rect 4950 4911 4994 4953
rect 5044 4973 5086 5011
rect 5044 4953 5058 4973
rect 5078 4953 5086 4973
rect 5044 4911 5086 4953
rect 5160 4973 5202 5011
rect 5160 4953 5168 4973
rect 5188 4953 5202 4973
rect 5160 4911 5202 4953
rect 5252 4980 5297 5011
rect 5252 4973 5296 4980
rect 5252 4953 5264 4973
rect 5284 4953 5296 4973
rect 16526 5162 16570 5204
rect 16526 5142 16538 5162
rect 16558 5142 16570 5162
rect 16526 5135 16570 5142
rect 16525 5104 16570 5135
rect 16620 5162 16662 5204
rect 16620 5142 16634 5162
rect 16654 5142 16662 5162
rect 16620 5104 16662 5142
rect 16736 5162 16778 5204
rect 16736 5142 16744 5162
rect 16764 5142 16778 5162
rect 16736 5104 16778 5142
rect 16828 5162 16872 5204
rect 16828 5142 16840 5162
rect 16860 5142 16872 5162
rect 16828 5104 16872 5142
rect 16954 5162 16996 5204
rect 16954 5142 16962 5162
rect 16982 5142 16996 5162
rect 16954 5104 16996 5142
rect 17046 5162 17090 5204
rect 17046 5142 17058 5162
rect 17078 5142 17090 5162
rect 17046 5104 17090 5142
rect 9109 4985 9153 5023
rect 5252 4911 5296 4953
rect 6683 4915 6727 4957
rect 2839 4844 2883 4882
rect 6683 4895 6695 4915
rect 6715 4895 6727 4915
rect 6683 4888 6727 4895
rect 6682 4857 6727 4888
rect 6777 4915 6819 4957
rect 6777 4895 6791 4915
rect 6811 4895 6819 4915
rect 6777 4857 6819 4895
rect 6893 4915 6935 4957
rect 6893 4895 6901 4915
rect 6921 4895 6935 4915
rect 6893 4857 6935 4895
rect 6985 4915 7029 4957
rect 6985 4895 6997 4915
rect 7017 4895 7029 4915
rect 6985 4857 7029 4895
rect 7111 4915 7153 4957
rect 7111 4895 7119 4915
rect 7139 4895 7153 4915
rect 7111 4857 7153 4895
rect 7203 4915 7247 4957
rect 9109 4965 9121 4985
rect 9141 4965 9153 4985
rect 7203 4895 7215 4915
rect 7235 4895 7247 4915
rect 9109 4923 9153 4965
rect 9203 4985 9245 5023
rect 9203 4965 9217 4985
rect 9237 4965 9245 4985
rect 9203 4923 9245 4965
rect 9327 4985 9371 5023
rect 9327 4965 9339 4985
rect 9359 4965 9371 4985
rect 9327 4923 9371 4965
rect 9421 4985 9463 5023
rect 9421 4965 9435 4985
rect 9455 4965 9463 4985
rect 9421 4923 9463 4965
rect 9537 4985 9579 5023
rect 9537 4965 9545 4985
rect 9565 4965 9579 4985
rect 9537 4923 9579 4965
rect 9629 4992 9674 5023
rect 9629 4985 9673 4992
rect 9629 4965 9641 4985
rect 9661 4965 9673 4985
rect 13473 4998 13517 5036
rect 9629 4923 9673 4965
rect 11060 4927 11104 4969
rect 7203 4857 7247 4895
rect 11060 4907 11072 4927
rect 11092 4907 11104 4927
rect 11060 4900 11104 4907
rect 11059 4869 11104 4900
rect 11154 4927 11196 4969
rect 11154 4907 11168 4927
rect 11188 4907 11196 4927
rect 11154 4869 11196 4907
rect 11270 4927 11312 4969
rect 11270 4907 11278 4927
rect 11298 4907 11312 4927
rect 11270 4869 11312 4907
rect 11362 4927 11406 4969
rect 11362 4907 11374 4927
rect 11394 4907 11406 4927
rect 11362 4869 11406 4907
rect 11488 4927 11530 4969
rect 11488 4907 11496 4927
rect 11516 4907 11530 4927
rect 11488 4869 11530 4907
rect 11580 4927 11624 4969
rect 13473 4978 13485 4998
rect 13505 4978 13517 4998
rect 11580 4907 11592 4927
rect 11612 4907 11624 4927
rect 13473 4936 13517 4978
rect 13567 4998 13609 5036
rect 13567 4978 13581 4998
rect 13601 4978 13609 4998
rect 13567 4936 13609 4978
rect 13691 4998 13735 5036
rect 13691 4978 13703 4998
rect 13723 4978 13735 4998
rect 13691 4936 13735 4978
rect 13785 4998 13827 5036
rect 13785 4978 13799 4998
rect 13819 4978 13827 4998
rect 13785 4936 13827 4978
rect 13901 4998 13943 5036
rect 13901 4978 13909 4998
rect 13929 4978 13943 4998
rect 13901 4936 13943 4978
rect 13993 5005 14038 5036
rect 13993 4998 14037 5005
rect 13993 4978 14005 4998
rect 14025 4978 14037 4998
rect 13993 4936 14037 4978
rect 15424 4940 15468 4982
rect 11580 4869 11624 4907
rect 15424 4920 15436 4940
rect 15456 4920 15468 4940
rect 15424 4913 15468 4920
rect 15423 4882 15468 4913
rect 15518 4940 15560 4982
rect 15518 4920 15532 4940
rect 15552 4920 15560 4940
rect 15518 4882 15560 4920
rect 15634 4940 15676 4982
rect 15634 4920 15642 4940
rect 15662 4920 15676 4940
rect 15634 4882 15676 4920
rect 15726 4940 15770 4982
rect 15726 4920 15738 4940
rect 15758 4920 15770 4940
rect 15726 4882 15770 4920
rect 15852 4940 15894 4982
rect 15852 4920 15860 4940
rect 15880 4920 15894 4940
rect 15852 4882 15894 4920
rect 15944 4940 15988 4982
rect 15944 4920 15956 4940
rect 15976 4920 15988 4940
rect 15944 4882 15988 4920
rect 1450 4576 1494 4614
rect 1450 4556 1462 4576
rect 1482 4556 1494 4576
rect 1450 4514 1494 4556
rect 1544 4576 1586 4614
rect 1544 4556 1558 4576
rect 1578 4556 1586 4576
rect 1544 4514 1586 4556
rect 1668 4576 1712 4614
rect 1668 4556 1680 4576
rect 1700 4556 1712 4576
rect 1668 4514 1712 4556
rect 1762 4576 1804 4614
rect 1762 4556 1776 4576
rect 1796 4556 1804 4576
rect 1762 4514 1804 4556
rect 1878 4576 1920 4614
rect 1878 4556 1886 4576
rect 1906 4556 1920 4576
rect 1878 4514 1920 4556
rect 1970 4583 2015 4614
rect 1970 4576 2014 4583
rect 1970 4556 1982 4576
rect 2002 4556 2014 4576
rect 5814 4589 5858 4627
rect 1970 4514 2014 4556
rect 3401 4518 3445 4560
rect 3401 4498 3413 4518
rect 3433 4498 3445 4518
rect 3401 4491 3445 4498
rect 3400 4460 3445 4491
rect 3495 4518 3537 4560
rect 3495 4498 3509 4518
rect 3529 4498 3537 4518
rect 3495 4460 3537 4498
rect 3611 4518 3653 4560
rect 3611 4498 3619 4518
rect 3639 4498 3653 4518
rect 3611 4460 3653 4498
rect 3703 4518 3747 4560
rect 3703 4498 3715 4518
rect 3735 4498 3747 4518
rect 3703 4460 3747 4498
rect 3829 4518 3871 4560
rect 3829 4498 3837 4518
rect 3857 4498 3871 4518
rect 3829 4460 3871 4498
rect 3921 4518 3965 4560
rect 5814 4569 5826 4589
rect 5846 4569 5858 4589
rect 3921 4498 3933 4518
rect 3953 4498 3965 4518
rect 5814 4527 5858 4569
rect 5908 4589 5950 4627
rect 5908 4569 5922 4589
rect 5942 4569 5950 4589
rect 5908 4527 5950 4569
rect 6032 4589 6076 4627
rect 6032 4569 6044 4589
rect 6064 4569 6076 4589
rect 6032 4527 6076 4569
rect 6126 4589 6168 4627
rect 6126 4569 6140 4589
rect 6160 4569 6168 4589
rect 6126 4527 6168 4569
rect 6242 4589 6284 4627
rect 6242 4569 6250 4589
rect 6270 4569 6284 4589
rect 6242 4527 6284 4569
rect 6334 4596 6379 4627
rect 6334 4589 6378 4596
rect 6334 4569 6346 4589
rect 6366 4569 6378 4589
rect 10191 4601 10235 4639
rect 6334 4527 6378 4569
rect 7765 4531 7809 4573
rect 3921 4460 3965 4498
rect 7765 4511 7777 4531
rect 7797 4511 7809 4531
rect 7765 4504 7809 4511
rect 7764 4473 7809 4504
rect 7859 4531 7901 4573
rect 7859 4511 7873 4531
rect 7893 4511 7901 4531
rect 7859 4473 7901 4511
rect 7975 4531 8017 4573
rect 7975 4511 7983 4531
rect 8003 4511 8017 4531
rect 7975 4473 8017 4511
rect 8067 4531 8111 4573
rect 8067 4511 8079 4531
rect 8099 4511 8111 4531
rect 8067 4473 8111 4511
rect 8193 4531 8235 4573
rect 8193 4511 8201 4531
rect 8221 4511 8235 4531
rect 8193 4473 8235 4511
rect 8285 4531 8329 4573
rect 10191 4581 10203 4601
rect 10223 4581 10235 4601
rect 8285 4511 8297 4531
rect 8317 4511 8329 4531
rect 10191 4539 10235 4581
rect 10285 4601 10327 4639
rect 10285 4581 10299 4601
rect 10319 4581 10327 4601
rect 10285 4539 10327 4581
rect 10409 4601 10453 4639
rect 10409 4581 10421 4601
rect 10441 4581 10453 4601
rect 10409 4539 10453 4581
rect 10503 4601 10545 4639
rect 10503 4581 10517 4601
rect 10537 4581 10545 4601
rect 10503 4539 10545 4581
rect 10619 4601 10661 4639
rect 10619 4581 10627 4601
rect 10647 4581 10661 4601
rect 10619 4539 10661 4581
rect 10711 4608 10756 4639
rect 10711 4601 10755 4608
rect 10711 4581 10723 4601
rect 10743 4581 10755 4601
rect 14555 4614 14599 4652
rect 10711 4539 10755 4581
rect 12142 4543 12186 4585
rect 8285 4473 8329 4511
rect 348 4354 392 4392
rect 348 4334 360 4354
rect 380 4334 392 4354
rect 348 4292 392 4334
rect 442 4354 484 4392
rect 442 4334 456 4354
rect 476 4334 484 4354
rect 442 4292 484 4334
rect 566 4354 610 4392
rect 566 4334 578 4354
rect 598 4334 610 4354
rect 566 4292 610 4334
rect 660 4354 702 4392
rect 660 4334 674 4354
rect 694 4334 702 4354
rect 660 4292 702 4334
rect 776 4354 818 4392
rect 776 4334 784 4354
rect 804 4334 818 4354
rect 776 4292 818 4334
rect 868 4361 913 4392
rect 868 4354 912 4361
rect 868 4334 880 4354
rect 900 4334 912 4354
rect 868 4292 912 4334
rect 12142 4523 12154 4543
rect 12174 4523 12186 4543
rect 12142 4516 12186 4523
rect 12141 4485 12186 4516
rect 12236 4543 12278 4585
rect 12236 4523 12250 4543
rect 12270 4523 12278 4543
rect 12236 4485 12278 4523
rect 12352 4543 12394 4585
rect 12352 4523 12360 4543
rect 12380 4523 12394 4543
rect 12352 4485 12394 4523
rect 12444 4543 12488 4585
rect 12444 4523 12456 4543
rect 12476 4523 12488 4543
rect 12444 4485 12488 4523
rect 12570 4543 12612 4585
rect 12570 4523 12578 4543
rect 12598 4523 12612 4543
rect 12570 4485 12612 4523
rect 12662 4543 12706 4585
rect 14555 4594 14567 4614
rect 14587 4594 14599 4614
rect 12662 4523 12674 4543
rect 12694 4523 12706 4543
rect 14555 4552 14599 4594
rect 14649 4614 14691 4652
rect 14649 4594 14663 4614
rect 14683 4594 14691 4614
rect 14649 4552 14691 4594
rect 14773 4614 14817 4652
rect 14773 4594 14785 4614
rect 14805 4594 14817 4614
rect 14773 4552 14817 4594
rect 14867 4614 14909 4652
rect 14867 4594 14881 4614
rect 14901 4594 14909 4614
rect 14867 4552 14909 4594
rect 14983 4614 15025 4652
rect 14983 4594 14991 4614
rect 15011 4594 15025 4614
rect 14983 4552 15025 4594
rect 15075 4621 15120 4652
rect 15075 4614 15119 4621
rect 15075 4594 15087 4614
rect 15107 4594 15119 4614
rect 15075 4552 15119 4594
rect 16506 4556 16550 4598
rect 12662 4485 12706 4523
rect 4712 4367 4756 4405
rect 4712 4347 4724 4367
rect 4744 4347 4756 4367
rect 2604 4290 2648 4332
rect 2604 4270 2616 4290
rect 2636 4270 2648 4290
rect 2604 4263 2648 4270
rect 2603 4232 2648 4263
rect 2698 4290 2740 4332
rect 2698 4270 2712 4290
rect 2732 4270 2740 4290
rect 2698 4232 2740 4270
rect 2814 4290 2856 4332
rect 2814 4270 2822 4290
rect 2842 4270 2856 4290
rect 2814 4232 2856 4270
rect 2906 4290 2950 4332
rect 2906 4270 2918 4290
rect 2938 4270 2950 4290
rect 2906 4232 2950 4270
rect 3032 4290 3074 4332
rect 3032 4270 3040 4290
rect 3060 4270 3074 4290
rect 3032 4232 3074 4270
rect 3124 4290 3168 4332
rect 4712 4305 4756 4347
rect 4806 4367 4848 4405
rect 4806 4347 4820 4367
rect 4840 4347 4848 4367
rect 4806 4305 4848 4347
rect 4930 4367 4974 4405
rect 4930 4347 4942 4367
rect 4962 4347 4974 4367
rect 4930 4305 4974 4347
rect 5024 4367 5066 4405
rect 5024 4347 5038 4367
rect 5058 4347 5066 4367
rect 5024 4305 5066 4347
rect 5140 4367 5182 4405
rect 5140 4347 5148 4367
rect 5168 4347 5182 4367
rect 5140 4305 5182 4347
rect 5232 4374 5277 4405
rect 5232 4367 5276 4374
rect 5232 4347 5244 4367
rect 5264 4347 5276 4367
rect 5232 4305 5276 4347
rect 16506 4536 16518 4556
rect 16538 4536 16550 4556
rect 16506 4529 16550 4536
rect 16505 4498 16550 4529
rect 16600 4556 16642 4598
rect 16600 4536 16614 4556
rect 16634 4536 16642 4556
rect 16600 4498 16642 4536
rect 16716 4556 16758 4598
rect 16716 4536 16724 4556
rect 16744 4536 16758 4556
rect 16716 4498 16758 4536
rect 16808 4556 16852 4598
rect 16808 4536 16820 4556
rect 16840 4536 16852 4556
rect 16808 4498 16852 4536
rect 16934 4556 16976 4598
rect 16934 4536 16942 4556
rect 16962 4536 16976 4556
rect 16934 4498 16976 4536
rect 17026 4556 17070 4598
rect 17026 4536 17038 4556
rect 17058 4536 17070 4556
rect 17026 4498 17070 4536
rect 9089 4379 9133 4417
rect 9089 4359 9101 4379
rect 9121 4359 9133 4379
rect 3124 4270 3136 4290
rect 3156 4270 3168 4290
rect 3124 4232 3168 4270
rect 1146 4170 1190 4208
rect 1146 4150 1158 4170
rect 1178 4150 1190 4170
rect 1146 4108 1190 4150
rect 1240 4170 1282 4208
rect 1240 4150 1254 4170
rect 1274 4150 1282 4170
rect 1240 4108 1282 4150
rect 1364 4170 1408 4208
rect 1364 4150 1376 4170
rect 1396 4150 1408 4170
rect 1364 4108 1408 4150
rect 1458 4170 1500 4208
rect 1458 4150 1472 4170
rect 1492 4150 1500 4170
rect 1458 4108 1500 4150
rect 1574 4170 1616 4208
rect 1574 4150 1582 4170
rect 1602 4150 1616 4170
rect 1574 4108 1616 4150
rect 1666 4177 1711 4208
rect 1666 4170 1710 4177
rect 1666 4150 1678 4170
rect 1698 4150 1710 4170
rect 1666 4108 1710 4150
rect 6968 4303 7012 4345
rect 6968 4283 6980 4303
rect 7000 4283 7012 4303
rect 6968 4276 7012 4283
rect 6967 4245 7012 4276
rect 7062 4303 7104 4345
rect 7062 4283 7076 4303
rect 7096 4283 7104 4303
rect 7062 4245 7104 4283
rect 7178 4303 7220 4345
rect 7178 4283 7186 4303
rect 7206 4283 7220 4303
rect 7178 4245 7220 4283
rect 7270 4303 7314 4345
rect 7270 4283 7282 4303
rect 7302 4283 7314 4303
rect 7270 4245 7314 4283
rect 7396 4303 7438 4345
rect 7396 4283 7404 4303
rect 7424 4283 7438 4303
rect 7396 4245 7438 4283
rect 7488 4303 7532 4345
rect 9089 4317 9133 4359
rect 9183 4379 9225 4417
rect 9183 4359 9197 4379
rect 9217 4359 9225 4379
rect 9183 4317 9225 4359
rect 9307 4379 9351 4417
rect 9307 4359 9319 4379
rect 9339 4359 9351 4379
rect 9307 4317 9351 4359
rect 9401 4379 9443 4417
rect 9401 4359 9415 4379
rect 9435 4359 9443 4379
rect 9401 4317 9443 4359
rect 9517 4379 9559 4417
rect 9517 4359 9525 4379
rect 9545 4359 9559 4379
rect 9517 4317 9559 4359
rect 9609 4386 9654 4417
rect 9609 4379 9653 4386
rect 9609 4359 9621 4379
rect 9641 4359 9653 4379
rect 9609 4317 9653 4359
rect 13453 4392 13497 4430
rect 13453 4372 13465 4392
rect 13485 4372 13497 4392
rect 7488 4283 7500 4303
rect 7520 4283 7532 4303
rect 7488 4245 7532 4283
rect 5510 4183 5554 4221
rect 5510 4163 5522 4183
rect 5542 4163 5554 4183
rect 3402 4106 3446 4148
rect 3402 4086 3414 4106
rect 3434 4086 3446 4106
rect 3402 4079 3446 4086
rect 3401 4048 3446 4079
rect 3496 4106 3538 4148
rect 3496 4086 3510 4106
rect 3530 4086 3538 4106
rect 3496 4048 3538 4086
rect 3612 4106 3654 4148
rect 3612 4086 3620 4106
rect 3640 4086 3654 4106
rect 3612 4048 3654 4086
rect 3704 4106 3748 4148
rect 3704 4086 3716 4106
rect 3736 4086 3748 4106
rect 3704 4048 3748 4086
rect 3830 4106 3872 4148
rect 3830 4086 3838 4106
rect 3858 4086 3872 4106
rect 3830 4048 3872 4086
rect 3922 4106 3966 4148
rect 5510 4121 5554 4163
rect 5604 4183 5646 4221
rect 5604 4163 5618 4183
rect 5638 4163 5646 4183
rect 5604 4121 5646 4163
rect 5728 4183 5772 4221
rect 5728 4163 5740 4183
rect 5760 4163 5772 4183
rect 5728 4121 5772 4163
rect 5822 4183 5864 4221
rect 5822 4163 5836 4183
rect 5856 4163 5864 4183
rect 5822 4121 5864 4163
rect 5938 4183 5980 4221
rect 5938 4163 5946 4183
rect 5966 4163 5980 4183
rect 5938 4121 5980 4163
rect 6030 4190 6075 4221
rect 6030 4183 6074 4190
rect 6030 4163 6042 4183
rect 6062 4163 6074 4183
rect 6030 4121 6074 4163
rect 11345 4315 11389 4357
rect 11345 4295 11357 4315
rect 11377 4295 11389 4315
rect 11345 4288 11389 4295
rect 11344 4257 11389 4288
rect 11439 4315 11481 4357
rect 11439 4295 11453 4315
rect 11473 4295 11481 4315
rect 11439 4257 11481 4295
rect 11555 4315 11597 4357
rect 11555 4295 11563 4315
rect 11583 4295 11597 4315
rect 11555 4257 11597 4295
rect 11647 4315 11691 4357
rect 11647 4295 11659 4315
rect 11679 4295 11691 4315
rect 11647 4257 11691 4295
rect 11773 4315 11815 4357
rect 11773 4295 11781 4315
rect 11801 4295 11815 4315
rect 11773 4257 11815 4295
rect 11865 4315 11909 4357
rect 13453 4330 13497 4372
rect 13547 4392 13589 4430
rect 13547 4372 13561 4392
rect 13581 4372 13589 4392
rect 13547 4330 13589 4372
rect 13671 4392 13715 4430
rect 13671 4372 13683 4392
rect 13703 4372 13715 4392
rect 13671 4330 13715 4372
rect 13765 4392 13807 4430
rect 13765 4372 13779 4392
rect 13799 4372 13807 4392
rect 13765 4330 13807 4372
rect 13881 4392 13923 4430
rect 13881 4372 13889 4392
rect 13909 4372 13923 4392
rect 13881 4330 13923 4372
rect 13973 4399 14018 4430
rect 13973 4392 14017 4399
rect 13973 4372 13985 4392
rect 14005 4372 14017 4392
rect 13973 4330 14017 4372
rect 11865 4295 11877 4315
rect 11897 4295 11909 4315
rect 11865 4257 11909 4295
rect 9887 4195 9931 4233
rect 9887 4175 9899 4195
rect 9919 4175 9931 4195
rect 3922 4086 3934 4106
rect 3954 4086 3966 4106
rect 3922 4048 3966 4086
rect 7766 4119 7810 4161
rect 7766 4099 7778 4119
rect 7798 4099 7810 4119
rect 7766 4092 7810 4099
rect 7765 4061 7810 4092
rect 7860 4119 7902 4161
rect 7860 4099 7874 4119
rect 7894 4099 7902 4119
rect 7860 4061 7902 4099
rect 7976 4119 8018 4161
rect 7976 4099 7984 4119
rect 8004 4099 8018 4119
rect 7976 4061 8018 4099
rect 8068 4119 8112 4161
rect 8068 4099 8080 4119
rect 8100 4099 8112 4119
rect 8068 4061 8112 4099
rect 8194 4119 8236 4161
rect 8194 4099 8202 4119
rect 8222 4099 8236 4119
rect 8194 4061 8236 4099
rect 8286 4119 8330 4161
rect 9887 4133 9931 4175
rect 9981 4195 10023 4233
rect 9981 4175 9995 4195
rect 10015 4175 10023 4195
rect 9981 4133 10023 4175
rect 10105 4195 10149 4233
rect 10105 4175 10117 4195
rect 10137 4175 10149 4195
rect 10105 4133 10149 4175
rect 10199 4195 10241 4233
rect 10199 4175 10213 4195
rect 10233 4175 10241 4195
rect 10199 4133 10241 4175
rect 10315 4195 10357 4233
rect 10315 4175 10323 4195
rect 10343 4175 10357 4195
rect 10315 4133 10357 4175
rect 10407 4202 10452 4233
rect 10407 4195 10451 4202
rect 10407 4175 10419 4195
rect 10439 4175 10451 4195
rect 10407 4133 10451 4175
rect 15709 4328 15753 4370
rect 15709 4308 15721 4328
rect 15741 4308 15753 4328
rect 15709 4301 15753 4308
rect 15708 4270 15753 4301
rect 15803 4328 15845 4370
rect 15803 4308 15817 4328
rect 15837 4308 15845 4328
rect 15803 4270 15845 4308
rect 15919 4328 15961 4370
rect 15919 4308 15927 4328
rect 15947 4308 15961 4328
rect 15919 4270 15961 4308
rect 16011 4328 16055 4370
rect 16011 4308 16023 4328
rect 16043 4308 16055 4328
rect 16011 4270 16055 4308
rect 16137 4328 16179 4370
rect 16137 4308 16145 4328
rect 16165 4308 16179 4328
rect 16137 4270 16179 4308
rect 16229 4328 16273 4370
rect 16229 4308 16241 4328
rect 16261 4308 16273 4328
rect 16229 4270 16273 4308
rect 14251 4208 14295 4246
rect 14251 4188 14263 4208
rect 14283 4188 14295 4208
rect 8286 4099 8298 4119
rect 8318 4099 8330 4119
rect 8286 4061 8330 4099
rect 349 3942 393 3980
rect 349 3922 361 3942
rect 381 3922 393 3942
rect 349 3880 393 3922
rect 443 3942 485 3980
rect 443 3922 457 3942
rect 477 3922 485 3942
rect 443 3880 485 3922
rect 567 3942 611 3980
rect 567 3922 579 3942
rect 599 3922 611 3942
rect 567 3880 611 3922
rect 661 3942 703 3980
rect 661 3922 675 3942
rect 695 3922 703 3942
rect 661 3880 703 3922
rect 777 3942 819 3980
rect 777 3922 785 3942
rect 805 3922 819 3942
rect 777 3880 819 3922
rect 869 3949 914 3980
rect 869 3942 913 3949
rect 869 3922 881 3942
rect 901 3922 913 3942
rect 12143 4131 12187 4173
rect 12143 4111 12155 4131
rect 12175 4111 12187 4131
rect 12143 4104 12187 4111
rect 12142 4073 12187 4104
rect 12237 4131 12279 4173
rect 12237 4111 12251 4131
rect 12271 4111 12279 4131
rect 12237 4073 12279 4111
rect 12353 4131 12395 4173
rect 12353 4111 12361 4131
rect 12381 4111 12395 4131
rect 12353 4073 12395 4111
rect 12445 4131 12489 4173
rect 12445 4111 12457 4131
rect 12477 4111 12489 4131
rect 12445 4073 12489 4111
rect 12571 4131 12613 4173
rect 12571 4111 12579 4131
rect 12599 4111 12613 4131
rect 12571 4073 12613 4111
rect 12663 4131 12707 4173
rect 14251 4146 14295 4188
rect 14345 4208 14387 4246
rect 14345 4188 14359 4208
rect 14379 4188 14387 4208
rect 14345 4146 14387 4188
rect 14469 4208 14513 4246
rect 14469 4188 14481 4208
rect 14501 4188 14513 4208
rect 14469 4146 14513 4188
rect 14563 4208 14605 4246
rect 14563 4188 14577 4208
rect 14597 4188 14605 4208
rect 14563 4146 14605 4188
rect 14679 4208 14721 4246
rect 14679 4188 14687 4208
rect 14707 4188 14721 4208
rect 14679 4146 14721 4188
rect 14771 4215 14816 4246
rect 14771 4208 14815 4215
rect 14771 4188 14783 4208
rect 14803 4188 14815 4208
rect 14771 4146 14815 4188
rect 12663 4111 12675 4131
rect 12695 4111 12707 4131
rect 12663 4073 12707 4111
rect 4713 3955 4757 3993
rect 869 3880 913 3922
rect 2505 3880 2549 3922
rect 2505 3860 2517 3880
rect 2537 3860 2549 3880
rect 2505 3853 2549 3860
rect 2504 3822 2549 3853
rect 2599 3880 2641 3922
rect 2599 3860 2613 3880
rect 2633 3860 2641 3880
rect 2599 3822 2641 3860
rect 2715 3880 2757 3922
rect 2715 3860 2723 3880
rect 2743 3860 2757 3880
rect 2715 3822 2757 3860
rect 2807 3880 2851 3922
rect 2807 3860 2819 3880
rect 2839 3860 2851 3880
rect 2807 3822 2851 3860
rect 2933 3880 2975 3922
rect 2933 3860 2941 3880
rect 2961 3860 2975 3880
rect 2933 3822 2975 3860
rect 3025 3880 3069 3922
rect 4713 3935 4725 3955
rect 4745 3935 4757 3955
rect 3025 3860 3037 3880
rect 3057 3860 3069 3880
rect 4713 3893 4757 3935
rect 4807 3955 4849 3993
rect 4807 3935 4821 3955
rect 4841 3935 4849 3955
rect 4807 3893 4849 3935
rect 4931 3955 4975 3993
rect 4931 3935 4943 3955
rect 4963 3935 4975 3955
rect 4931 3893 4975 3935
rect 5025 3955 5067 3993
rect 5025 3935 5039 3955
rect 5059 3935 5067 3955
rect 5025 3893 5067 3935
rect 5141 3955 5183 3993
rect 5141 3935 5149 3955
rect 5169 3935 5183 3955
rect 5141 3893 5183 3935
rect 5233 3962 5278 3993
rect 5233 3955 5277 3962
rect 5233 3935 5245 3955
rect 5265 3935 5277 3955
rect 16507 4144 16551 4186
rect 16507 4124 16519 4144
rect 16539 4124 16551 4144
rect 16507 4117 16551 4124
rect 16506 4086 16551 4117
rect 16601 4144 16643 4186
rect 16601 4124 16615 4144
rect 16635 4124 16643 4144
rect 16601 4086 16643 4124
rect 16717 4144 16759 4186
rect 16717 4124 16725 4144
rect 16745 4124 16759 4144
rect 16717 4086 16759 4124
rect 16809 4144 16853 4186
rect 16809 4124 16821 4144
rect 16841 4124 16853 4144
rect 16809 4086 16853 4124
rect 16935 4144 16977 4186
rect 16935 4124 16943 4144
rect 16963 4124 16977 4144
rect 16935 4086 16977 4124
rect 17027 4144 17071 4186
rect 17027 4124 17039 4144
rect 17059 4124 17071 4144
rect 17027 4086 17071 4124
rect 9090 3967 9134 4005
rect 5233 3893 5277 3935
rect 6869 3893 6913 3935
rect 3025 3822 3069 3860
rect 6869 3873 6881 3893
rect 6901 3873 6913 3893
rect 6869 3866 6913 3873
rect 6868 3835 6913 3866
rect 6963 3893 7005 3935
rect 6963 3873 6977 3893
rect 6997 3873 7005 3893
rect 6963 3835 7005 3873
rect 7079 3893 7121 3935
rect 7079 3873 7087 3893
rect 7107 3873 7121 3893
rect 7079 3835 7121 3873
rect 7171 3893 7215 3935
rect 7171 3873 7183 3893
rect 7203 3873 7215 3893
rect 7171 3835 7215 3873
rect 7297 3893 7339 3935
rect 7297 3873 7305 3893
rect 7325 3873 7339 3893
rect 7297 3835 7339 3873
rect 7389 3893 7433 3935
rect 9090 3947 9102 3967
rect 9122 3947 9134 3967
rect 7389 3873 7401 3893
rect 7421 3873 7433 3893
rect 9090 3905 9134 3947
rect 9184 3967 9226 4005
rect 9184 3947 9198 3967
rect 9218 3947 9226 3967
rect 9184 3905 9226 3947
rect 9308 3967 9352 4005
rect 9308 3947 9320 3967
rect 9340 3947 9352 3967
rect 9308 3905 9352 3947
rect 9402 3967 9444 4005
rect 9402 3947 9416 3967
rect 9436 3947 9444 3967
rect 9402 3905 9444 3947
rect 9518 3967 9560 4005
rect 9518 3947 9526 3967
rect 9546 3947 9560 3967
rect 9518 3905 9560 3947
rect 9610 3974 9655 4005
rect 9610 3967 9654 3974
rect 9610 3947 9622 3967
rect 9642 3947 9654 3967
rect 13454 3980 13498 4018
rect 9610 3905 9654 3947
rect 11246 3905 11290 3947
rect 7389 3835 7433 3873
rect 11246 3885 11258 3905
rect 11278 3885 11290 3905
rect 11246 3878 11290 3885
rect 11245 3847 11290 3878
rect 11340 3905 11382 3947
rect 11340 3885 11354 3905
rect 11374 3885 11382 3905
rect 11340 3847 11382 3885
rect 11456 3905 11498 3947
rect 11456 3885 11464 3905
rect 11484 3885 11498 3905
rect 11456 3847 11498 3885
rect 11548 3905 11592 3947
rect 11548 3885 11560 3905
rect 11580 3885 11592 3905
rect 11548 3847 11592 3885
rect 11674 3905 11716 3947
rect 11674 3885 11682 3905
rect 11702 3885 11716 3905
rect 11674 3847 11716 3885
rect 11766 3905 11810 3947
rect 13454 3960 13466 3980
rect 13486 3960 13498 3980
rect 11766 3885 11778 3905
rect 11798 3885 11810 3905
rect 13454 3918 13498 3960
rect 13548 3980 13590 4018
rect 13548 3960 13562 3980
rect 13582 3960 13590 3980
rect 13548 3918 13590 3960
rect 13672 3980 13716 4018
rect 13672 3960 13684 3980
rect 13704 3960 13716 3980
rect 13672 3918 13716 3960
rect 13766 3980 13808 4018
rect 13766 3960 13780 3980
rect 13800 3960 13808 3980
rect 13766 3918 13808 3960
rect 13882 3980 13924 4018
rect 13882 3960 13890 3980
rect 13910 3960 13924 3980
rect 13882 3918 13924 3960
rect 13974 3987 14019 4018
rect 13974 3980 14018 3987
rect 13974 3960 13986 3980
rect 14006 3960 14018 3980
rect 13974 3918 14018 3960
rect 15610 3918 15654 3960
rect 11766 3847 11810 3885
rect 15610 3898 15622 3918
rect 15642 3898 15654 3918
rect 15610 3891 15654 3898
rect 15609 3860 15654 3891
rect 15704 3918 15746 3960
rect 15704 3898 15718 3918
rect 15738 3898 15746 3918
rect 15704 3860 15746 3898
rect 15820 3918 15862 3960
rect 15820 3898 15828 3918
rect 15848 3898 15862 3918
rect 15820 3860 15862 3898
rect 15912 3918 15956 3960
rect 15912 3898 15924 3918
rect 15944 3898 15956 3918
rect 15912 3860 15956 3898
rect 16038 3918 16080 3960
rect 16038 3898 16046 3918
rect 16066 3898 16080 3918
rect 16038 3860 16080 3898
rect 16130 3918 16174 3960
rect 16130 3898 16142 3918
rect 16162 3898 16174 3918
rect 16130 3860 16174 3898
rect 1228 3562 1272 3600
rect 1228 3542 1240 3562
rect 1260 3542 1272 3562
rect 1228 3500 1272 3542
rect 1322 3562 1364 3600
rect 1322 3542 1336 3562
rect 1356 3542 1364 3562
rect 1322 3500 1364 3542
rect 1446 3562 1490 3600
rect 1446 3542 1458 3562
rect 1478 3542 1490 3562
rect 1446 3500 1490 3542
rect 1540 3562 1582 3600
rect 1540 3542 1554 3562
rect 1574 3542 1582 3562
rect 1540 3500 1582 3542
rect 1656 3562 1698 3600
rect 1656 3542 1664 3562
rect 1684 3542 1698 3562
rect 1656 3500 1698 3542
rect 1748 3569 1793 3600
rect 1748 3562 1792 3569
rect 1748 3542 1760 3562
rect 1780 3542 1792 3562
rect 5592 3575 5636 3613
rect 1748 3500 1792 3542
rect 3384 3500 3428 3542
rect 3384 3480 3396 3500
rect 3416 3480 3428 3500
rect 3384 3473 3428 3480
rect 3383 3442 3428 3473
rect 3478 3500 3520 3542
rect 3478 3480 3492 3500
rect 3512 3480 3520 3500
rect 3478 3442 3520 3480
rect 3594 3500 3636 3542
rect 3594 3480 3602 3500
rect 3622 3480 3636 3500
rect 3594 3442 3636 3480
rect 3686 3500 3730 3542
rect 3686 3480 3698 3500
rect 3718 3480 3730 3500
rect 3686 3442 3730 3480
rect 3812 3500 3854 3542
rect 3812 3480 3820 3500
rect 3840 3480 3854 3500
rect 3812 3442 3854 3480
rect 3904 3500 3948 3542
rect 5592 3555 5604 3575
rect 5624 3555 5636 3575
rect 3904 3480 3916 3500
rect 3936 3480 3948 3500
rect 5592 3513 5636 3555
rect 5686 3575 5728 3613
rect 5686 3555 5700 3575
rect 5720 3555 5728 3575
rect 5686 3513 5728 3555
rect 5810 3575 5854 3613
rect 5810 3555 5822 3575
rect 5842 3555 5854 3575
rect 5810 3513 5854 3555
rect 5904 3575 5946 3613
rect 5904 3555 5918 3575
rect 5938 3555 5946 3575
rect 5904 3513 5946 3555
rect 6020 3575 6062 3613
rect 6020 3555 6028 3575
rect 6048 3555 6062 3575
rect 6020 3513 6062 3555
rect 6112 3582 6157 3613
rect 6112 3575 6156 3582
rect 6112 3555 6124 3575
rect 6144 3555 6156 3575
rect 9969 3587 10013 3625
rect 6112 3513 6156 3555
rect 7748 3513 7792 3555
rect 3904 3442 3948 3480
rect 7748 3493 7760 3513
rect 7780 3493 7792 3513
rect 7748 3486 7792 3493
rect 7747 3455 7792 3486
rect 7842 3513 7884 3555
rect 7842 3493 7856 3513
rect 7876 3493 7884 3513
rect 7842 3455 7884 3493
rect 7958 3513 8000 3555
rect 7958 3493 7966 3513
rect 7986 3493 8000 3513
rect 7958 3455 8000 3493
rect 8050 3513 8094 3555
rect 8050 3493 8062 3513
rect 8082 3493 8094 3513
rect 8050 3455 8094 3493
rect 8176 3513 8218 3555
rect 8176 3493 8184 3513
rect 8204 3493 8218 3513
rect 8176 3455 8218 3493
rect 8268 3513 8312 3555
rect 9969 3567 9981 3587
rect 10001 3567 10013 3587
rect 8268 3493 8280 3513
rect 8300 3493 8312 3513
rect 9969 3525 10013 3567
rect 10063 3587 10105 3625
rect 10063 3567 10077 3587
rect 10097 3567 10105 3587
rect 10063 3525 10105 3567
rect 10187 3587 10231 3625
rect 10187 3567 10199 3587
rect 10219 3567 10231 3587
rect 10187 3525 10231 3567
rect 10281 3587 10323 3625
rect 10281 3567 10295 3587
rect 10315 3567 10323 3587
rect 10281 3525 10323 3567
rect 10397 3587 10439 3625
rect 10397 3567 10405 3587
rect 10425 3567 10439 3587
rect 10397 3525 10439 3567
rect 10489 3594 10534 3625
rect 10489 3587 10533 3594
rect 10489 3567 10501 3587
rect 10521 3567 10533 3587
rect 14333 3600 14377 3638
rect 10489 3525 10533 3567
rect 12125 3525 12169 3567
rect 8268 3455 8312 3493
rect 331 3336 375 3374
rect 331 3316 343 3336
rect 363 3316 375 3336
rect 331 3274 375 3316
rect 425 3336 467 3374
rect 425 3316 439 3336
rect 459 3316 467 3336
rect 425 3274 467 3316
rect 549 3336 593 3374
rect 549 3316 561 3336
rect 581 3316 593 3336
rect 549 3274 593 3316
rect 643 3336 685 3374
rect 643 3316 657 3336
rect 677 3316 685 3336
rect 643 3274 685 3316
rect 759 3336 801 3374
rect 759 3316 767 3336
rect 787 3316 801 3336
rect 759 3274 801 3316
rect 851 3343 896 3374
rect 851 3336 895 3343
rect 851 3316 863 3336
rect 883 3316 895 3336
rect 851 3274 895 3316
rect 12125 3505 12137 3525
rect 12157 3505 12169 3525
rect 12125 3498 12169 3505
rect 12124 3467 12169 3498
rect 12219 3525 12261 3567
rect 12219 3505 12233 3525
rect 12253 3505 12261 3525
rect 12219 3467 12261 3505
rect 12335 3525 12377 3567
rect 12335 3505 12343 3525
rect 12363 3505 12377 3525
rect 12335 3467 12377 3505
rect 12427 3525 12471 3567
rect 12427 3505 12439 3525
rect 12459 3505 12471 3525
rect 12427 3467 12471 3505
rect 12553 3525 12595 3567
rect 12553 3505 12561 3525
rect 12581 3505 12595 3525
rect 12553 3467 12595 3505
rect 12645 3525 12689 3567
rect 14333 3580 14345 3600
rect 14365 3580 14377 3600
rect 12645 3505 12657 3525
rect 12677 3505 12689 3525
rect 14333 3538 14377 3580
rect 14427 3600 14469 3638
rect 14427 3580 14441 3600
rect 14461 3580 14469 3600
rect 14427 3538 14469 3580
rect 14551 3600 14595 3638
rect 14551 3580 14563 3600
rect 14583 3580 14595 3600
rect 14551 3538 14595 3580
rect 14645 3600 14687 3638
rect 14645 3580 14659 3600
rect 14679 3580 14687 3600
rect 14645 3538 14687 3580
rect 14761 3600 14803 3638
rect 14761 3580 14769 3600
rect 14789 3580 14803 3600
rect 14761 3538 14803 3580
rect 14853 3607 14898 3638
rect 14853 3600 14897 3607
rect 14853 3580 14865 3600
rect 14885 3580 14897 3600
rect 14853 3538 14897 3580
rect 16489 3538 16533 3580
rect 12645 3467 12689 3505
rect 4695 3349 4739 3387
rect 4695 3329 4707 3349
rect 4727 3329 4739 3349
rect 2587 3272 2631 3314
rect 2587 3252 2599 3272
rect 2619 3252 2631 3272
rect 2587 3245 2631 3252
rect 2586 3214 2631 3245
rect 2681 3272 2723 3314
rect 2681 3252 2695 3272
rect 2715 3252 2723 3272
rect 2681 3214 2723 3252
rect 2797 3272 2839 3314
rect 2797 3252 2805 3272
rect 2825 3252 2839 3272
rect 2797 3214 2839 3252
rect 2889 3272 2933 3314
rect 2889 3252 2901 3272
rect 2921 3252 2933 3272
rect 2889 3214 2933 3252
rect 3015 3272 3057 3314
rect 3015 3252 3023 3272
rect 3043 3252 3057 3272
rect 3015 3214 3057 3252
rect 3107 3272 3151 3314
rect 4695 3287 4739 3329
rect 4789 3349 4831 3387
rect 4789 3329 4803 3349
rect 4823 3329 4831 3349
rect 4789 3287 4831 3329
rect 4913 3349 4957 3387
rect 4913 3329 4925 3349
rect 4945 3329 4957 3349
rect 4913 3287 4957 3329
rect 5007 3349 5049 3387
rect 5007 3329 5021 3349
rect 5041 3329 5049 3349
rect 5007 3287 5049 3329
rect 5123 3349 5165 3387
rect 5123 3329 5131 3349
rect 5151 3329 5165 3349
rect 5123 3287 5165 3329
rect 5215 3356 5260 3387
rect 5215 3349 5259 3356
rect 5215 3329 5227 3349
rect 5247 3329 5259 3349
rect 5215 3287 5259 3329
rect 16489 3518 16501 3538
rect 16521 3518 16533 3538
rect 16489 3511 16533 3518
rect 16488 3480 16533 3511
rect 16583 3538 16625 3580
rect 16583 3518 16597 3538
rect 16617 3518 16625 3538
rect 16583 3480 16625 3518
rect 16699 3538 16741 3580
rect 16699 3518 16707 3538
rect 16727 3518 16741 3538
rect 16699 3480 16741 3518
rect 16791 3538 16835 3580
rect 16791 3518 16803 3538
rect 16823 3518 16835 3538
rect 16791 3480 16835 3518
rect 16917 3538 16959 3580
rect 16917 3518 16925 3538
rect 16945 3518 16959 3538
rect 16917 3480 16959 3518
rect 17009 3538 17053 3580
rect 17009 3518 17021 3538
rect 17041 3518 17053 3538
rect 17009 3480 17053 3518
rect 9072 3361 9116 3399
rect 9072 3341 9084 3361
rect 9104 3341 9116 3361
rect 3107 3252 3119 3272
rect 3139 3252 3151 3272
rect 3107 3214 3151 3252
rect 1129 3152 1173 3190
rect 1129 3132 1141 3152
rect 1161 3132 1173 3152
rect 1129 3090 1173 3132
rect 1223 3152 1265 3190
rect 1223 3132 1237 3152
rect 1257 3132 1265 3152
rect 1223 3090 1265 3132
rect 1347 3152 1391 3190
rect 1347 3132 1359 3152
rect 1379 3132 1391 3152
rect 1347 3090 1391 3132
rect 1441 3152 1483 3190
rect 1441 3132 1455 3152
rect 1475 3132 1483 3152
rect 1441 3090 1483 3132
rect 1557 3152 1599 3190
rect 1557 3132 1565 3152
rect 1585 3132 1599 3152
rect 1557 3090 1599 3132
rect 1649 3159 1694 3190
rect 1649 3152 1693 3159
rect 1649 3132 1661 3152
rect 1681 3132 1693 3152
rect 1649 3090 1693 3132
rect 6951 3285 6995 3327
rect 6951 3265 6963 3285
rect 6983 3265 6995 3285
rect 6951 3258 6995 3265
rect 6950 3227 6995 3258
rect 7045 3285 7087 3327
rect 7045 3265 7059 3285
rect 7079 3265 7087 3285
rect 7045 3227 7087 3265
rect 7161 3285 7203 3327
rect 7161 3265 7169 3285
rect 7189 3265 7203 3285
rect 7161 3227 7203 3265
rect 7253 3285 7297 3327
rect 7253 3265 7265 3285
rect 7285 3265 7297 3285
rect 7253 3227 7297 3265
rect 7379 3285 7421 3327
rect 7379 3265 7387 3285
rect 7407 3265 7421 3285
rect 7379 3227 7421 3265
rect 7471 3285 7515 3327
rect 9072 3299 9116 3341
rect 9166 3361 9208 3399
rect 9166 3341 9180 3361
rect 9200 3341 9208 3361
rect 9166 3299 9208 3341
rect 9290 3361 9334 3399
rect 9290 3341 9302 3361
rect 9322 3341 9334 3361
rect 9290 3299 9334 3341
rect 9384 3361 9426 3399
rect 9384 3341 9398 3361
rect 9418 3341 9426 3361
rect 9384 3299 9426 3341
rect 9500 3361 9542 3399
rect 9500 3341 9508 3361
rect 9528 3341 9542 3361
rect 9500 3299 9542 3341
rect 9592 3368 9637 3399
rect 9592 3361 9636 3368
rect 9592 3341 9604 3361
rect 9624 3341 9636 3361
rect 9592 3299 9636 3341
rect 13436 3374 13480 3412
rect 13436 3354 13448 3374
rect 13468 3354 13480 3374
rect 7471 3265 7483 3285
rect 7503 3265 7515 3285
rect 7471 3227 7515 3265
rect 5493 3165 5537 3203
rect 5493 3145 5505 3165
rect 5525 3145 5537 3165
rect 3385 3088 3429 3130
rect 3385 3068 3397 3088
rect 3417 3068 3429 3088
rect 3385 3061 3429 3068
rect 3384 3030 3429 3061
rect 3479 3088 3521 3130
rect 3479 3068 3493 3088
rect 3513 3068 3521 3088
rect 3479 3030 3521 3068
rect 3595 3088 3637 3130
rect 3595 3068 3603 3088
rect 3623 3068 3637 3088
rect 3595 3030 3637 3068
rect 3687 3088 3731 3130
rect 3687 3068 3699 3088
rect 3719 3068 3731 3088
rect 3687 3030 3731 3068
rect 3813 3088 3855 3130
rect 3813 3068 3821 3088
rect 3841 3068 3855 3088
rect 3813 3030 3855 3068
rect 3905 3088 3949 3130
rect 5493 3103 5537 3145
rect 5587 3165 5629 3203
rect 5587 3145 5601 3165
rect 5621 3145 5629 3165
rect 5587 3103 5629 3145
rect 5711 3165 5755 3203
rect 5711 3145 5723 3165
rect 5743 3145 5755 3165
rect 5711 3103 5755 3145
rect 5805 3165 5847 3203
rect 5805 3145 5819 3165
rect 5839 3145 5847 3165
rect 5805 3103 5847 3145
rect 5921 3165 5963 3203
rect 5921 3145 5929 3165
rect 5949 3145 5963 3165
rect 5921 3103 5963 3145
rect 6013 3172 6058 3203
rect 6013 3165 6057 3172
rect 6013 3145 6025 3165
rect 6045 3145 6057 3165
rect 6013 3103 6057 3145
rect 11328 3297 11372 3339
rect 11328 3277 11340 3297
rect 11360 3277 11372 3297
rect 11328 3270 11372 3277
rect 11327 3239 11372 3270
rect 11422 3297 11464 3339
rect 11422 3277 11436 3297
rect 11456 3277 11464 3297
rect 11422 3239 11464 3277
rect 11538 3297 11580 3339
rect 11538 3277 11546 3297
rect 11566 3277 11580 3297
rect 11538 3239 11580 3277
rect 11630 3297 11674 3339
rect 11630 3277 11642 3297
rect 11662 3277 11674 3297
rect 11630 3239 11674 3277
rect 11756 3297 11798 3339
rect 11756 3277 11764 3297
rect 11784 3277 11798 3297
rect 11756 3239 11798 3277
rect 11848 3297 11892 3339
rect 13436 3312 13480 3354
rect 13530 3374 13572 3412
rect 13530 3354 13544 3374
rect 13564 3354 13572 3374
rect 13530 3312 13572 3354
rect 13654 3374 13698 3412
rect 13654 3354 13666 3374
rect 13686 3354 13698 3374
rect 13654 3312 13698 3354
rect 13748 3374 13790 3412
rect 13748 3354 13762 3374
rect 13782 3354 13790 3374
rect 13748 3312 13790 3354
rect 13864 3374 13906 3412
rect 13864 3354 13872 3374
rect 13892 3354 13906 3374
rect 13864 3312 13906 3354
rect 13956 3381 14001 3412
rect 13956 3374 14000 3381
rect 13956 3354 13968 3374
rect 13988 3354 14000 3374
rect 13956 3312 14000 3354
rect 11848 3277 11860 3297
rect 11880 3277 11892 3297
rect 11848 3239 11892 3277
rect 9870 3177 9914 3215
rect 9870 3157 9882 3177
rect 9902 3157 9914 3177
rect 3905 3068 3917 3088
rect 3937 3068 3949 3088
rect 3905 3030 3949 3068
rect 7749 3101 7793 3143
rect 7749 3081 7761 3101
rect 7781 3081 7793 3101
rect 7749 3074 7793 3081
rect 7748 3043 7793 3074
rect 7843 3101 7885 3143
rect 7843 3081 7857 3101
rect 7877 3081 7885 3101
rect 7843 3043 7885 3081
rect 7959 3101 8001 3143
rect 7959 3081 7967 3101
rect 7987 3081 8001 3101
rect 7959 3043 8001 3081
rect 8051 3101 8095 3143
rect 8051 3081 8063 3101
rect 8083 3081 8095 3101
rect 8051 3043 8095 3081
rect 8177 3101 8219 3143
rect 8177 3081 8185 3101
rect 8205 3081 8219 3101
rect 8177 3043 8219 3081
rect 8269 3101 8313 3143
rect 9870 3115 9914 3157
rect 9964 3177 10006 3215
rect 9964 3157 9978 3177
rect 9998 3157 10006 3177
rect 9964 3115 10006 3157
rect 10088 3177 10132 3215
rect 10088 3157 10100 3177
rect 10120 3157 10132 3177
rect 10088 3115 10132 3157
rect 10182 3177 10224 3215
rect 10182 3157 10196 3177
rect 10216 3157 10224 3177
rect 10182 3115 10224 3157
rect 10298 3177 10340 3215
rect 10298 3157 10306 3177
rect 10326 3157 10340 3177
rect 10298 3115 10340 3157
rect 10390 3184 10435 3215
rect 10390 3177 10434 3184
rect 10390 3157 10402 3177
rect 10422 3157 10434 3177
rect 10390 3115 10434 3157
rect 15692 3310 15736 3352
rect 15692 3290 15704 3310
rect 15724 3290 15736 3310
rect 15692 3283 15736 3290
rect 15691 3252 15736 3283
rect 15786 3310 15828 3352
rect 15786 3290 15800 3310
rect 15820 3290 15828 3310
rect 15786 3252 15828 3290
rect 15902 3310 15944 3352
rect 15902 3290 15910 3310
rect 15930 3290 15944 3310
rect 15902 3252 15944 3290
rect 15994 3310 16038 3352
rect 15994 3290 16006 3310
rect 16026 3290 16038 3310
rect 15994 3252 16038 3290
rect 16120 3310 16162 3352
rect 16120 3290 16128 3310
rect 16148 3290 16162 3310
rect 16120 3252 16162 3290
rect 16212 3310 16256 3352
rect 16212 3290 16224 3310
rect 16244 3290 16256 3310
rect 16212 3252 16256 3290
rect 14234 3190 14278 3228
rect 14234 3170 14246 3190
rect 14266 3170 14278 3190
rect 8269 3081 8281 3101
rect 8301 3081 8313 3101
rect 8269 3043 8313 3081
rect 332 2924 376 2962
rect 332 2904 344 2924
rect 364 2904 376 2924
rect 332 2862 376 2904
rect 426 2924 468 2962
rect 426 2904 440 2924
rect 460 2904 468 2924
rect 426 2862 468 2904
rect 550 2924 594 2962
rect 550 2904 562 2924
rect 582 2904 594 2924
rect 550 2862 594 2904
rect 644 2924 686 2962
rect 644 2904 658 2924
rect 678 2904 686 2924
rect 644 2862 686 2904
rect 760 2924 802 2962
rect 760 2904 768 2924
rect 788 2904 802 2924
rect 760 2862 802 2904
rect 852 2931 897 2962
rect 852 2924 896 2931
rect 852 2904 864 2924
rect 884 2904 896 2924
rect 12126 3113 12170 3155
rect 12126 3093 12138 3113
rect 12158 3093 12170 3113
rect 12126 3086 12170 3093
rect 12125 3055 12170 3086
rect 12220 3113 12262 3155
rect 12220 3093 12234 3113
rect 12254 3093 12262 3113
rect 12220 3055 12262 3093
rect 12336 3113 12378 3155
rect 12336 3093 12344 3113
rect 12364 3093 12378 3113
rect 12336 3055 12378 3093
rect 12428 3113 12472 3155
rect 12428 3093 12440 3113
rect 12460 3093 12472 3113
rect 12428 3055 12472 3093
rect 12554 3113 12596 3155
rect 12554 3093 12562 3113
rect 12582 3093 12596 3113
rect 12554 3055 12596 3093
rect 12646 3113 12690 3155
rect 14234 3128 14278 3170
rect 14328 3190 14370 3228
rect 14328 3170 14342 3190
rect 14362 3170 14370 3190
rect 14328 3128 14370 3170
rect 14452 3190 14496 3228
rect 14452 3170 14464 3190
rect 14484 3170 14496 3190
rect 14452 3128 14496 3170
rect 14546 3190 14588 3228
rect 14546 3170 14560 3190
rect 14580 3170 14588 3190
rect 14546 3128 14588 3170
rect 14662 3190 14704 3228
rect 14662 3170 14670 3190
rect 14690 3170 14704 3190
rect 14662 3128 14704 3170
rect 14754 3197 14799 3228
rect 14754 3190 14798 3197
rect 14754 3170 14766 3190
rect 14786 3170 14798 3190
rect 14754 3128 14798 3170
rect 12646 3093 12658 3113
rect 12678 3093 12690 3113
rect 12646 3055 12690 3093
rect 4696 2937 4740 2975
rect 852 2862 896 2904
rect 2422 2864 2466 2906
rect 2422 2844 2434 2864
rect 2454 2844 2466 2864
rect 2422 2837 2466 2844
rect 2421 2806 2466 2837
rect 2516 2864 2558 2906
rect 2516 2844 2530 2864
rect 2550 2844 2558 2864
rect 2516 2806 2558 2844
rect 2632 2864 2674 2906
rect 2632 2844 2640 2864
rect 2660 2844 2674 2864
rect 2632 2806 2674 2844
rect 2724 2864 2768 2906
rect 2724 2844 2736 2864
rect 2756 2844 2768 2864
rect 2724 2806 2768 2844
rect 2850 2864 2892 2906
rect 2850 2844 2858 2864
rect 2878 2844 2892 2864
rect 2850 2806 2892 2844
rect 2942 2864 2986 2906
rect 4696 2917 4708 2937
rect 4728 2917 4740 2937
rect 2942 2844 2954 2864
rect 2974 2844 2986 2864
rect 4696 2875 4740 2917
rect 4790 2937 4832 2975
rect 4790 2917 4804 2937
rect 4824 2917 4832 2937
rect 4790 2875 4832 2917
rect 4914 2937 4958 2975
rect 4914 2917 4926 2937
rect 4946 2917 4958 2937
rect 4914 2875 4958 2917
rect 5008 2937 5050 2975
rect 5008 2917 5022 2937
rect 5042 2917 5050 2937
rect 5008 2875 5050 2917
rect 5124 2937 5166 2975
rect 5124 2917 5132 2937
rect 5152 2917 5166 2937
rect 5124 2875 5166 2917
rect 5216 2944 5261 2975
rect 5216 2937 5260 2944
rect 5216 2917 5228 2937
rect 5248 2917 5260 2937
rect 16490 3126 16534 3168
rect 16490 3106 16502 3126
rect 16522 3106 16534 3126
rect 16490 3099 16534 3106
rect 16489 3068 16534 3099
rect 16584 3126 16626 3168
rect 16584 3106 16598 3126
rect 16618 3106 16626 3126
rect 16584 3068 16626 3106
rect 16700 3126 16742 3168
rect 16700 3106 16708 3126
rect 16728 3106 16742 3126
rect 16700 3068 16742 3106
rect 16792 3126 16836 3168
rect 16792 3106 16804 3126
rect 16824 3106 16836 3126
rect 16792 3068 16836 3106
rect 16918 3126 16960 3168
rect 16918 3106 16926 3126
rect 16946 3106 16960 3126
rect 16918 3068 16960 3106
rect 17010 3126 17054 3168
rect 17010 3106 17022 3126
rect 17042 3106 17054 3126
rect 17010 3068 17054 3106
rect 9073 2949 9117 2987
rect 5216 2875 5260 2917
rect 6786 2877 6830 2919
rect 2942 2806 2986 2844
rect 6786 2857 6798 2877
rect 6818 2857 6830 2877
rect 6786 2850 6830 2857
rect 6785 2819 6830 2850
rect 6880 2877 6922 2919
rect 6880 2857 6894 2877
rect 6914 2857 6922 2877
rect 6880 2819 6922 2857
rect 6996 2877 7038 2919
rect 6996 2857 7004 2877
rect 7024 2857 7038 2877
rect 6996 2819 7038 2857
rect 7088 2877 7132 2919
rect 7088 2857 7100 2877
rect 7120 2857 7132 2877
rect 7088 2819 7132 2857
rect 7214 2877 7256 2919
rect 7214 2857 7222 2877
rect 7242 2857 7256 2877
rect 7214 2819 7256 2857
rect 7306 2877 7350 2919
rect 9073 2929 9085 2949
rect 9105 2929 9117 2949
rect 7306 2857 7318 2877
rect 7338 2857 7350 2877
rect 9073 2887 9117 2929
rect 9167 2949 9209 2987
rect 9167 2929 9181 2949
rect 9201 2929 9209 2949
rect 9167 2887 9209 2929
rect 9291 2949 9335 2987
rect 9291 2929 9303 2949
rect 9323 2929 9335 2949
rect 9291 2887 9335 2929
rect 9385 2949 9427 2987
rect 9385 2929 9399 2949
rect 9419 2929 9427 2949
rect 9385 2887 9427 2929
rect 9501 2949 9543 2987
rect 9501 2929 9509 2949
rect 9529 2929 9543 2949
rect 9501 2887 9543 2929
rect 9593 2956 9638 2987
rect 9593 2949 9637 2956
rect 9593 2929 9605 2949
rect 9625 2929 9637 2949
rect 13437 2962 13481 3000
rect 9593 2887 9637 2929
rect 11163 2889 11207 2931
rect 7306 2819 7350 2857
rect 11163 2869 11175 2889
rect 11195 2869 11207 2889
rect 11163 2862 11207 2869
rect 11162 2831 11207 2862
rect 11257 2889 11299 2931
rect 11257 2869 11271 2889
rect 11291 2869 11299 2889
rect 11257 2831 11299 2869
rect 11373 2889 11415 2931
rect 11373 2869 11381 2889
rect 11401 2869 11415 2889
rect 11373 2831 11415 2869
rect 11465 2889 11509 2931
rect 11465 2869 11477 2889
rect 11497 2869 11509 2889
rect 11465 2831 11509 2869
rect 11591 2889 11633 2931
rect 11591 2869 11599 2889
rect 11619 2869 11633 2889
rect 11591 2831 11633 2869
rect 11683 2889 11727 2931
rect 13437 2942 13449 2962
rect 13469 2942 13481 2962
rect 11683 2869 11695 2889
rect 11715 2869 11727 2889
rect 13437 2900 13481 2942
rect 13531 2962 13573 3000
rect 13531 2942 13545 2962
rect 13565 2942 13573 2962
rect 13531 2900 13573 2942
rect 13655 2962 13699 3000
rect 13655 2942 13667 2962
rect 13687 2942 13699 2962
rect 13655 2900 13699 2942
rect 13749 2962 13791 3000
rect 13749 2942 13763 2962
rect 13783 2942 13791 2962
rect 13749 2900 13791 2942
rect 13865 2962 13907 3000
rect 13865 2942 13873 2962
rect 13893 2942 13907 2962
rect 13865 2900 13907 2942
rect 13957 2969 14002 3000
rect 13957 2962 14001 2969
rect 13957 2942 13969 2962
rect 13989 2942 14001 2962
rect 13957 2900 14001 2942
rect 15527 2902 15571 2944
rect 11683 2831 11727 2869
rect 15527 2882 15539 2902
rect 15559 2882 15571 2902
rect 15527 2875 15571 2882
rect 15526 2844 15571 2875
rect 15621 2902 15663 2944
rect 15621 2882 15635 2902
rect 15655 2882 15663 2902
rect 15621 2844 15663 2882
rect 15737 2902 15779 2944
rect 15737 2882 15745 2902
rect 15765 2882 15779 2902
rect 15737 2844 15779 2882
rect 15829 2902 15873 2944
rect 15829 2882 15841 2902
rect 15861 2882 15873 2902
rect 15829 2844 15873 2882
rect 15955 2902 15997 2944
rect 15955 2882 15963 2902
rect 15983 2882 15997 2902
rect 15955 2844 15997 2882
rect 16047 2902 16091 2944
rect 16047 2882 16059 2902
rect 16079 2882 16091 2902
rect 16047 2844 16091 2882
rect 1274 2542 1318 2580
rect 1274 2522 1286 2542
rect 1306 2522 1318 2542
rect 1274 2480 1318 2522
rect 1368 2542 1410 2580
rect 1368 2522 1382 2542
rect 1402 2522 1410 2542
rect 1368 2480 1410 2522
rect 1492 2542 1536 2580
rect 1492 2522 1504 2542
rect 1524 2522 1536 2542
rect 1492 2480 1536 2522
rect 1586 2542 1628 2580
rect 1586 2522 1600 2542
rect 1620 2522 1628 2542
rect 1586 2480 1628 2522
rect 1702 2542 1744 2580
rect 1702 2522 1710 2542
rect 1730 2522 1744 2542
rect 1702 2480 1744 2522
rect 1794 2549 1839 2580
rect 1794 2542 1838 2549
rect 1794 2522 1806 2542
rect 1826 2522 1838 2542
rect 5638 2555 5682 2593
rect 1794 2480 1838 2522
rect 3364 2482 3408 2524
rect 3364 2462 3376 2482
rect 3396 2462 3408 2482
rect 3364 2455 3408 2462
rect 3363 2424 3408 2455
rect 3458 2482 3500 2524
rect 3458 2462 3472 2482
rect 3492 2462 3500 2482
rect 3458 2424 3500 2462
rect 3574 2482 3616 2524
rect 3574 2462 3582 2482
rect 3602 2462 3616 2482
rect 3574 2424 3616 2462
rect 3666 2482 3710 2524
rect 3666 2462 3678 2482
rect 3698 2462 3710 2482
rect 3666 2424 3710 2462
rect 3792 2482 3834 2524
rect 3792 2462 3800 2482
rect 3820 2462 3834 2482
rect 3792 2424 3834 2462
rect 3884 2482 3928 2524
rect 5638 2535 5650 2555
rect 5670 2535 5682 2555
rect 3884 2462 3896 2482
rect 3916 2462 3928 2482
rect 5638 2493 5682 2535
rect 5732 2555 5774 2593
rect 5732 2535 5746 2555
rect 5766 2535 5774 2555
rect 5732 2493 5774 2535
rect 5856 2555 5900 2593
rect 5856 2535 5868 2555
rect 5888 2535 5900 2555
rect 5856 2493 5900 2535
rect 5950 2555 5992 2593
rect 5950 2535 5964 2555
rect 5984 2535 5992 2555
rect 5950 2493 5992 2535
rect 6066 2555 6108 2593
rect 6066 2535 6074 2555
rect 6094 2535 6108 2555
rect 6066 2493 6108 2535
rect 6158 2562 6203 2593
rect 6158 2555 6202 2562
rect 6158 2535 6170 2555
rect 6190 2535 6202 2555
rect 10015 2567 10059 2605
rect 6158 2493 6202 2535
rect 7728 2495 7772 2537
rect 3884 2424 3928 2462
rect 7728 2475 7740 2495
rect 7760 2475 7772 2495
rect 7728 2468 7772 2475
rect 7727 2437 7772 2468
rect 7822 2495 7864 2537
rect 7822 2475 7836 2495
rect 7856 2475 7864 2495
rect 7822 2437 7864 2475
rect 7938 2495 7980 2537
rect 7938 2475 7946 2495
rect 7966 2475 7980 2495
rect 7938 2437 7980 2475
rect 8030 2495 8074 2537
rect 8030 2475 8042 2495
rect 8062 2475 8074 2495
rect 8030 2437 8074 2475
rect 8156 2495 8198 2537
rect 8156 2475 8164 2495
rect 8184 2475 8198 2495
rect 8156 2437 8198 2475
rect 8248 2495 8292 2537
rect 10015 2547 10027 2567
rect 10047 2547 10059 2567
rect 8248 2475 8260 2495
rect 8280 2475 8292 2495
rect 10015 2505 10059 2547
rect 10109 2567 10151 2605
rect 10109 2547 10123 2567
rect 10143 2547 10151 2567
rect 10109 2505 10151 2547
rect 10233 2567 10277 2605
rect 10233 2547 10245 2567
rect 10265 2547 10277 2567
rect 10233 2505 10277 2547
rect 10327 2567 10369 2605
rect 10327 2547 10341 2567
rect 10361 2547 10369 2567
rect 10327 2505 10369 2547
rect 10443 2567 10485 2605
rect 10443 2547 10451 2567
rect 10471 2547 10485 2567
rect 10443 2505 10485 2547
rect 10535 2574 10580 2605
rect 10535 2567 10579 2574
rect 10535 2547 10547 2567
rect 10567 2547 10579 2567
rect 14379 2580 14423 2618
rect 10535 2505 10579 2547
rect 12105 2507 12149 2549
rect 8248 2437 8292 2475
rect 311 2318 355 2356
rect 311 2298 323 2318
rect 343 2298 355 2318
rect 311 2256 355 2298
rect 405 2318 447 2356
rect 405 2298 419 2318
rect 439 2298 447 2318
rect 405 2256 447 2298
rect 529 2318 573 2356
rect 529 2298 541 2318
rect 561 2298 573 2318
rect 529 2256 573 2298
rect 623 2318 665 2356
rect 623 2298 637 2318
rect 657 2298 665 2318
rect 623 2256 665 2298
rect 739 2318 781 2356
rect 739 2298 747 2318
rect 767 2298 781 2318
rect 739 2256 781 2298
rect 831 2325 876 2356
rect 831 2318 875 2325
rect 831 2298 843 2318
rect 863 2298 875 2318
rect 831 2256 875 2298
rect 12105 2487 12117 2507
rect 12137 2487 12149 2507
rect 12105 2480 12149 2487
rect 12104 2449 12149 2480
rect 12199 2507 12241 2549
rect 12199 2487 12213 2507
rect 12233 2487 12241 2507
rect 12199 2449 12241 2487
rect 12315 2507 12357 2549
rect 12315 2487 12323 2507
rect 12343 2487 12357 2507
rect 12315 2449 12357 2487
rect 12407 2507 12451 2549
rect 12407 2487 12419 2507
rect 12439 2487 12451 2507
rect 12407 2449 12451 2487
rect 12533 2507 12575 2549
rect 12533 2487 12541 2507
rect 12561 2487 12575 2507
rect 12533 2449 12575 2487
rect 12625 2507 12669 2549
rect 14379 2560 14391 2580
rect 14411 2560 14423 2580
rect 12625 2487 12637 2507
rect 12657 2487 12669 2507
rect 14379 2518 14423 2560
rect 14473 2580 14515 2618
rect 14473 2560 14487 2580
rect 14507 2560 14515 2580
rect 14473 2518 14515 2560
rect 14597 2580 14641 2618
rect 14597 2560 14609 2580
rect 14629 2560 14641 2580
rect 14597 2518 14641 2560
rect 14691 2580 14733 2618
rect 14691 2560 14705 2580
rect 14725 2560 14733 2580
rect 14691 2518 14733 2560
rect 14807 2580 14849 2618
rect 14807 2560 14815 2580
rect 14835 2560 14849 2580
rect 14807 2518 14849 2560
rect 14899 2587 14944 2618
rect 14899 2580 14943 2587
rect 14899 2560 14911 2580
rect 14931 2560 14943 2580
rect 14899 2518 14943 2560
rect 16469 2520 16513 2562
rect 12625 2449 12669 2487
rect 4675 2331 4719 2369
rect 4675 2311 4687 2331
rect 4707 2311 4719 2331
rect 2567 2254 2611 2296
rect 2567 2234 2579 2254
rect 2599 2234 2611 2254
rect 2567 2227 2611 2234
rect 2566 2196 2611 2227
rect 2661 2254 2703 2296
rect 2661 2234 2675 2254
rect 2695 2234 2703 2254
rect 2661 2196 2703 2234
rect 2777 2254 2819 2296
rect 2777 2234 2785 2254
rect 2805 2234 2819 2254
rect 2777 2196 2819 2234
rect 2869 2254 2913 2296
rect 2869 2234 2881 2254
rect 2901 2234 2913 2254
rect 2869 2196 2913 2234
rect 2995 2254 3037 2296
rect 2995 2234 3003 2254
rect 3023 2234 3037 2254
rect 2995 2196 3037 2234
rect 3087 2254 3131 2296
rect 4675 2269 4719 2311
rect 4769 2331 4811 2369
rect 4769 2311 4783 2331
rect 4803 2311 4811 2331
rect 4769 2269 4811 2311
rect 4893 2331 4937 2369
rect 4893 2311 4905 2331
rect 4925 2311 4937 2331
rect 4893 2269 4937 2311
rect 4987 2331 5029 2369
rect 4987 2311 5001 2331
rect 5021 2311 5029 2331
rect 4987 2269 5029 2311
rect 5103 2331 5145 2369
rect 5103 2311 5111 2331
rect 5131 2311 5145 2331
rect 5103 2269 5145 2311
rect 5195 2338 5240 2369
rect 5195 2331 5239 2338
rect 5195 2311 5207 2331
rect 5227 2311 5239 2331
rect 5195 2269 5239 2311
rect 16469 2500 16481 2520
rect 16501 2500 16513 2520
rect 16469 2493 16513 2500
rect 16468 2462 16513 2493
rect 16563 2520 16605 2562
rect 16563 2500 16577 2520
rect 16597 2500 16605 2520
rect 16563 2462 16605 2500
rect 16679 2520 16721 2562
rect 16679 2500 16687 2520
rect 16707 2500 16721 2520
rect 16679 2462 16721 2500
rect 16771 2520 16815 2562
rect 16771 2500 16783 2520
rect 16803 2500 16815 2520
rect 16771 2462 16815 2500
rect 16897 2520 16939 2562
rect 16897 2500 16905 2520
rect 16925 2500 16939 2520
rect 16897 2462 16939 2500
rect 16989 2520 17033 2562
rect 16989 2500 17001 2520
rect 17021 2500 17033 2520
rect 16989 2462 17033 2500
rect 9052 2343 9096 2381
rect 9052 2323 9064 2343
rect 9084 2323 9096 2343
rect 3087 2234 3099 2254
rect 3119 2234 3131 2254
rect 3087 2196 3131 2234
rect 1109 2134 1153 2172
rect 1109 2114 1121 2134
rect 1141 2114 1153 2134
rect 1109 2072 1153 2114
rect 1203 2134 1245 2172
rect 1203 2114 1217 2134
rect 1237 2114 1245 2134
rect 1203 2072 1245 2114
rect 1327 2134 1371 2172
rect 1327 2114 1339 2134
rect 1359 2114 1371 2134
rect 1327 2072 1371 2114
rect 1421 2134 1463 2172
rect 1421 2114 1435 2134
rect 1455 2114 1463 2134
rect 1421 2072 1463 2114
rect 1537 2134 1579 2172
rect 1537 2114 1545 2134
rect 1565 2114 1579 2134
rect 1537 2072 1579 2114
rect 1629 2141 1674 2172
rect 1629 2134 1673 2141
rect 1629 2114 1641 2134
rect 1661 2114 1673 2134
rect 1629 2072 1673 2114
rect 6931 2267 6975 2309
rect 6931 2247 6943 2267
rect 6963 2247 6975 2267
rect 6931 2240 6975 2247
rect 6930 2209 6975 2240
rect 7025 2267 7067 2309
rect 7025 2247 7039 2267
rect 7059 2247 7067 2267
rect 7025 2209 7067 2247
rect 7141 2267 7183 2309
rect 7141 2247 7149 2267
rect 7169 2247 7183 2267
rect 7141 2209 7183 2247
rect 7233 2267 7277 2309
rect 7233 2247 7245 2267
rect 7265 2247 7277 2267
rect 7233 2209 7277 2247
rect 7359 2267 7401 2309
rect 7359 2247 7367 2267
rect 7387 2247 7401 2267
rect 7359 2209 7401 2247
rect 7451 2267 7495 2309
rect 9052 2281 9096 2323
rect 9146 2343 9188 2381
rect 9146 2323 9160 2343
rect 9180 2323 9188 2343
rect 9146 2281 9188 2323
rect 9270 2343 9314 2381
rect 9270 2323 9282 2343
rect 9302 2323 9314 2343
rect 9270 2281 9314 2323
rect 9364 2343 9406 2381
rect 9364 2323 9378 2343
rect 9398 2323 9406 2343
rect 9364 2281 9406 2323
rect 9480 2343 9522 2381
rect 9480 2323 9488 2343
rect 9508 2323 9522 2343
rect 9480 2281 9522 2323
rect 9572 2350 9617 2381
rect 9572 2343 9616 2350
rect 9572 2323 9584 2343
rect 9604 2323 9616 2343
rect 9572 2281 9616 2323
rect 13416 2356 13460 2394
rect 13416 2336 13428 2356
rect 13448 2336 13460 2356
rect 7451 2247 7463 2267
rect 7483 2247 7495 2267
rect 7451 2209 7495 2247
rect 5473 2147 5517 2185
rect 5473 2127 5485 2147
rect 5505 2127 5517 2147
rect 3365 2070 3409 2112
rect 3365 2050 3377 2070
rect 3397 2050 3409 2070
rect 3365 2043 3409 2050
rect 3364 2012 3409 2043
rect 3459 2070 3501 2112
rect 3459 2050 3473 2070
rect 3493 2050 3501 2070
rect 3459 2012 3501 2050
rect 3575 2070 3617 2112
rect 3575 2050 3583 2070
rect 3603 2050 3617 2070
rect 3575 2012 3617 2050
rect 3667 2070 3711 2112
rect 3667 2050 3679 2070
rect 3699 2050 3711 2070
rect 3667 2012 3711 2050
rect 3793 2070 3835 2112
rect 3793 2050 3801 2070
rect 3821 2050 3835 2070
rect 3793 2012 3835 2050
rect 3885 2070 3929 2112
rect 5473 2085 5517 2127
rect 5567 2147 5609 2185
rect 5567 2127 5581 2147
rect 5601 2127 5609 2147
rect 5567 2085 5609 2127
rect 5691 2147 5735 2185
rect 5691 2127 5703 2147
rect 5723 2127 5735 2147
rect 5691 2085 5735 2127
rect 5785 2147 5827 2185
rect 5785 2127 5799 2147
rect 5819 2127 5827 2147
rect 5785 2085 5827 2127
rect 5901 2147 5943 2185
rect 5901 2127 5909 2147
rect 5929 2127 5943 2147
rect 5901 2085 5943 2127
rect 5993 2154 6038 2185
rect 5993 2147 6037 2154
rect 5993 2127 6005 2147
rect 6025 2127 6037 2147
rect 5993 2085 6037 2127
rect 11308 2279 11352 2321
rect 11308 2259 11320 2279
rect 11340 2259 11352 2279
rect 11308 2252 11352 2259
rect 11307 2221 11352 2252
rect 11402 2279 11444 2321
rect 11402 2259 11416 2279
rect 11436 2259 11444 2279
rect 11402 2221 11444 2259
rect 11518 2279 11560 2321
rect 11518 2259 11526 2279
rect 11546 2259 11560 2279
rect 11518 2221 11560 2259
rect 11610 2279 11654 2321
rect 11610 2259 11622 2279
rect 11642 2259 11654 2279
rect 11610 2221 11654 2259
rect 11736 2279 11778 2321
rect 11736 2259 11744 2279
rect 11764 2259 11778 2279
rect 11736 2221 11778 2259
rect 11828 2279 11872 2321
rect 13416 2294 13460 2336
rect 13510 2356 13552 2394
rect 13510 2336 13524 2356
rect 13544 2336 13552 2356
rect 13510 2294 13552 2336
rect 13634 2356 13678 2394
rect 13634 2336 13646 2356
rect 13666 2336 13678 2356
rect 13634 2294 13678 2336
rect 13728 2356 13770 2394
rect 13728 2336 13742 2356
rect 13762 2336 13770 2356
rect 13728 2294 13770 2336
rect 13844 2356 13886 2394
rect 13844 2336 13852 2356
rect 13872 2336 13886 2356
rect 13844 2294 13886 2336
rect 13936 2363 13981 2394
rect 13936 2356 13980 2363
rect 13936 2336 13948 2356
rect 13968 2336 13980 2356
rect 13936 2294 13980 2336
rect 11828 2259 11840 2279
rect 11860 2259 11872 2279
rect 11828 2221 11872 2259
rect 9850 2159 9894 2197
rect 9850 2139 9862 2159
rect 9882 2139 9894 2159
rect 3885 2050 3897 2070
rect 3917 2050 3929 2070
rect 3885 2012 3929 2050
rect 7729 2083 7773 2125
rect 7729 2063 7741 2083
rect 7761 2063 7773 2083
rect 7729 2056 7773 2063
rect 7728 2025 7773 2056
rect 7823 2083 7865 2125
rect 7823 2063 7837 2083
rect 7857 2063 7865 2083
rect 7823 2025 7865 2063
rect 7939 2083 7981 2125
rect 7939 2063 7947 2083
rect 7967 2063 7981 2083
rect 7939 2025 7981 2063
rect 8031 2083 8075 2125
rect 8031 2063 8043 2083
rect 8063 2063 8075 2083
rect 8031 2025 8075 2063
rect 8157 2083 8199 2125
rect 8157 2063 8165 2083
rect 8185 2063 8199 2083
rect 8157 2025 8199 2063
rect 8249 2083 8293 2125
rect 9850 2097 9894 2139
rect 9944 2159 9986 2197
rect 9944 2139 9958 2159
rect 9978 2139 9986 2159
rect 9944 2097 9986 2139
rect 10068 2159 10112 2197
rect 10068 2139 10080 2159
rect 10100 2139 10112 2159
rect 10068 2097 10112 2139
rect 10162 2159 10204 2197
rect 10162 2139 10176 2159
rect 10196 2139 10204 2159
rect 10162 2097 10204 2139
rect 10278 2159 10320 2197
rect 10278 2139 10286 2159
rect 10306 2139 10320 2159
rect 10278 2097 10320 2139
rect 10370 2166 10415 2197
rect 10370 2159 10414 2166
rect 10370 2139 10382 2159
rect 10402 2139 10414 2159
rect 10370 2097 10414 2139
rect 15672 2292 15716 2334
rect 15672 2272 15684 2292
rect 15704 2272 15716 2292
rect 15672 2265 15716 2272
rect 15671 2234 15716 2265
rect 15766 2292 15808 2334
rect 15766 2272 15780 2292
rect 15800 2272 15808 2292
rect 15766 2234 15808 2272
rect 15882 2292 15924 2334
rect 15882 2272 15890 2292
rect 15910 2272 15924 2292
rect 15882 2234 15924 2272
rect 15974 2292 16018 2334
rect 15974 2272 15986 2292
rect 16006 2272 16018 2292
rect 15974 2234 16018 2272
rect 16100 2292 16142 2334
rect 16100 2272 16108 2292
rect 16128 2272 16142 2292
rect 16100 2234 16142 2272
rect 16192 2292 16236 2334
rect 16192 2272 16204 2292
rect 16224 2272 16236 2292
rect 16192 2234 16236 2272
rect 14214 2172 14258 2210
rect 14214 2152 14226 2172
rect 14246 2152 14258 2172
rect 8249 2063 8261 2083
rect 8281 2063 8293 2083
rect 8249 2025 8293 2063
rect 312 1906 356 1944
rect 312 1886 324 1906
rect 344 1886 356 1906
rect 312 1844 356 1886
rect 406 1906 448 1944
rect 406 1886 420 1906
rect 440 1886 448 1906
rect 406 1844 448 1886
rect 530 1906 574 1944
rect 530 1886 542 1906
rect 562 1886 574 1906
rect 530 1844 574 1886
rect 624 1906 666 1944
rect 624 1886 638 1906
rect 658 1886 666 1906
rect 624 1844 666 1886
rect 740 1906 782 1944
rect 740 1886 748 1906
rect 768 1886 782 1906
rect 740 1844 782 1886
rect 832 1913 877 1944
rect 832 1906 876 1913
rect 832 1886 844 1906
rect 864 1886 876 1906
rect 12106 2095 12150 2137
rect 12106 2075 12118 2095
rect 12138 2075 12150 2095
rect 12106 2068 12150 2075
rect 12105 2037 12150 2068
rect 12200 2095 12242 2137
rect 12200 2075 12214 2095
rect 12234 2075 12242 2095
rect 12200 2037 12242 2075
rect 12316 2095 12358 2137
rect 12316 2075 12324 2095
rect 12344 2075 12358 2095
rect 12316 2037 12358 2075
rect 12408 2095 12452 2137
rect 12408 2075 12420 2095
rect 12440 2075 12452 2095
rect 12408 2037 12452 2075
rect 12534 2095 12576 2137
rect 12534 2075 12542 2095
rect 12562 2075 12576 2095
rect 12534 2037 12576 2075
rect 12626 2095 12670 2137
rect 14214 2110 14258 2152
rect 14308 2172 14350 2210
rect 14308 2152 14322 2172
rect 14342 2152 14350 2172
rect 14308 2110 14350 2152
rect 14432 2172 14476 2210
rect 14432 2152 14444 2172
rect 14464 2152 14476 2172
rect 14432 2110 14476 2152
rect 14526 2172 14568 2210
rect 14526 2152 14540 2172
rect 14560 2152 14568 2172
rect 14526 2110 14568 2152
rect 14642 2172 14684 2210
rect 14642 2152 14650 2172
rect 14670 2152 14684 2172
rect 14642 2110 14684 2152
rect 14734 2179 14779 2210
rect 14734 2172 14778 2179
rect 14734 2152 14746 2172
rect 14766 2152 14778 2172
rect 14734 2110 14778 2152
rect 12626 2075 12638 2095
rect 12658 2075 12670 2095
rect 12626 2037 12670 2075
rect 4676 1919 4720 1957
rect 832 1844 876 1886
rect 2468 1844 2512 1886
rect 2468 1824 2480 1844
rect 2500 1824 2512 1844
rect 2468 1817 2512 1824
rect 2467 1786 2512 1817
rect 2562 1844 2604 1886
rect 2562 1824 2576 1844
rect 2596 1824 2604 1844
rect 2562 1786 2604 1824
rect 2678 1844 2720 1886
rect 2678 1824 2686 1844
rect 2706 1824 2720 1844
rect 2678 1786 2720 1824
rect 2770 1844 2814 1886
rect 2770 1824 2782 1844
rect 2802 1824 2814 1844
rect 2770 1786 2814 1824
rect 2896 1844 2938 1886
rect 2896 1824 2904 1844
rect 2924 1824 2938 1844
rect 2896 1786 2938 1824
rect 2988 1844 3032 1886
rect 4676 1899 4688 1919
rect 4708 1899 4720 1919
rect 2988 1824 3000 1844
rect 3020 1824 3032 1844
rect 4676 1857 4720 1899
rect 4770 1919 4812 1957
rect 4770 1899 4784 1919
rect 4804 1899 4812 1919
rect 4770 1857 4812 1899
rect 4894 1919 4938 1957
rect 4894 1899 4906 1919
rect 4926 1899 4938 1919
rect 4894 1857 4938 1899
rect 4988 1919 5030 1957
rect 4988 1899 5002 1919
rect 5022 1899 5030 1919
rect 4988 1857 5030 1899
rect 5104 1919 5146 1957
rect 5104 1899 5112 1919
rect 5132 1899 5146 1919
rect 5104 1857 5146 1899
rect 5196 1926 5241 1957
rect 5196 1919 5240 1926
rect 5196 1899 5208 1919
rect 5228 1899 5240 1919
rect 16470 2108 16514 2150
rect 16470 2088 16482 2108
rect 16502 2088 16514 2108
rect 16470 2081 16514 2088
rect 16469 2050 16514 2081
rect 16564 2108 16606 2150
rect 16564 2088 16578 2108
rect 16598 2088 16606 2108
rect 16564 2050 16606 2088
rect 16680 2108 16722 2150
rect 16680 2088 16688 2108
rect 16708 2088 16722 2108
rect 16680 2050 16722 2088
rect 16772 2108 16816 2150
rect 16772 2088 16784 2108
rect 16804 2088 16816 2108
rect 16772 2050 16816 2088
rect 16898 2108 16940 2150
rect 16898 2088 16906 2108
rect 16926 2088 16940 2108
rect 16898 2050 16940 2088
rect 16990 2108 17034 2150
rect 16990 2088 17002 2108
rect 17022 2088 17034 2108
rect 16990 2050 17034 2088
rect 9053 1931 9097 1969
rect 5196 1857 5240 1899
rect 6832 1857 6876 1899
rect 2988 1786 3032 1824
rect 6832 1837 6844 1857
rect 6864 1837 6876 1857
rect 6832 1830 6876 1837
rect 6831 1799 6876 1830
rect 6926 1857 6968 1899
rect 6926 1837 6940 1857
rect 6960 1837 6968 1857
rect 6926 1799 6968 1837
rect 7042 1857 7084 1899
rect 7042 1837 7050 1857
rect 7070 1837 7084 1857
rect 7042 1799 7084 1837
rect 7134 1857 7178 1899
rect 7134 1837 7146 1857
rect 7166 1837 7178 1857
rect 7134 1799 7178 1837
rect 7260 1857 7302 1899
rect 7260 1837 7268 1857
rect 7288 1837 7302 1857
rect 7260 1799 7302 1837
rect 7352 1857 7396 1899
rect 9053 1911 9065 1931
rect 9085 1911 9097 1931
rect 7352 1837 7364 1857
rect 7384 1837 7396 1857
rect 9053 1869 9097 1911
rect 9147 1931 9189 1969
rect 9147 1911 9161 1931
rect 9181 1911 9189 1931
rect 9147 1869 9189 1911
rect 9271 1931 9315 1969
rect 9271 1911 9283 1931
rect 9303 1911 9315 1931
rect 9271 1869 9315 1911
rect 9365 1931 9407 1969
rect 9365 1911 9379 1931
rect 9399 1911 9407 1931
rect 9365 1869 9407 1911
rect 9481 1931 9523 1969
rect 9481 1911 9489 1931
rect 9509 1911 9523 1931
rect 9481 1869 9523 1911
rect 9573 1938 9618 1969
rect 9573 1931 9617 1938
rect 9573 1911 9585 1931
rect 9605 1911 9617 1931
rect 13417 1944 13461 1982
rect 9573 1869 9617 1911
rect 11209 1869 11253 1911
rect 7352 1799 7396 1837
rect 11209 1849 11221 1869
rect 11241 1849 11253 1869
rect 11209 1842 11253 1849
rect 11208 1811 11253 1842
rect 11303 1869 11345 1911
rect 11303 1849 11317 1869
rect 11337 1849 11345 1869
rect 11303 1811 11345 1849
rect 11419 1869 11461 1911
rect 11419 1849 11427 1869
rect 11447 1849 11461 1869
rect 11419 1811 11461 1849
rect 11511 1869 11555 1911
rect 11511 1849 11523 1869
rect 11543 1849 11555 1869
rect 11511 1811 11555 1849
rect 11637 1869 11679 1911
rect 11637 1849 11645 1869
rect 11665 1849 11679 1869
rect 11637 1811 11679 1849
rect 11729 1869 11773 1911
rect 13417 1924 13429 1944
rect 13449 1924 13461 1944
rect 11729 1849 11741 1869
rect 11761 1849 11773 1869
rect 13417 1882 13461 1924
rect 13511 1944 13553 1982
rect 13511 1924 13525 1944
rect 13545 1924 13553 1944
rect 13511 1882 13553 1924
rect 13635 1944 13679 1982
rect 13635 1924 13647 1944
rect 13667 1924 13679 1944
rect 13635 1882 13679 1924
rect 13729 1944 13771 1982
rect 13729 1924 13743 1944
rect 13763 1924 13771 1944
rect 13729 1882 13771 1924
rect 13845 1944 13887 1982
rect 13845 1924 13853 1944
rect 13873 1924 13887 1944
rect 13845 1882 13887 1924
rect 13937 1951 13982 1982
rect 13937 1944 13981 1951
rect 13937 1924 13949 1944
rect 13969 1924 13981 1944
rect 13937 1882 13981 1924
rect 15573 1882 15617 1924
rect 11729 1811 11773 1849
rect 15573 1862 15585 1882
rect 15605 1862 15617 1882
rect 15573 1855 15617 1862
rect 15572 1824 15617 1855
rect 15667 1882 15709 1924
rect 15667 1862 15681 1882
rect 15701 1862 15709 1882
rect 15667 1824 15709 1862
rect 15783 1882 15825 1924
rect 15783 1862 15791 1882
rect 15811 1862 15825 1882
rect 15783 1824 15825 1862
rect 15875 1882 15919 1924
rect 15875 1862 15887 1882
rect 15907 1862 15919 1882
rect 15875 1824 15919 1862
rect 16001 1882 16043 1924
rect 16001 1862 16009 1882
rect 16029 1862 16043 1882
rect 16001 1824 16043 1862
rect 16093 1882 16137 1924
rect 16093 1862 16105 1882
rect 16125 1862 16137 1882
rect 16093 1824 16137 1862
rect 1191 1526 1235 1564
rect 1191 1506 1203 1526
rect 1223 1506 1235 1526
rect 1191 1464 1235 1506
rect 1285 1526 1327 1564
rect 1285 1506 1299 1526
rect 1319 1506 1327 1526
rect 1285 1464 1327 1506
rect 1409 1526 1453 1564
rect 1409 1506 1421 1526
rect 1441 1506 1453 1526
rect 1409 1464 1453 1506
rect 1503 1526 1545 1564
rect 1503 1506 1517 1526
rect 1537 1506 1545 1526
rect 1503 1464 1545 1506
rect 1619 1526 1661 1564
rect 1619 1506 1627 1526
rect 1647 1506 1661 1526
rect 1619 1464 1661 1506
rect 1711 1533 1756 1564
rect 1711 1526 1755 1533
rect 1711 1506 1723 1526
rect 1743 1506 1755 1526
rect 5555 1539 5599 1577
rect 1711 1464 1755 1506
rect 3347 1464 3391 1506
rect 3347 1444 3359 1464
rect 3379 1444 3391 1464
rect 3347 1437 3391 1444
rect 3346 1406 3391 1437
rect 3441 1464 3483 1506
rect 3441 1444 3455 1464
rect 3475 1444 3483 1464
rect 3441 1406 3483 1444
rect 3557 1464 3599 1506
rect 3557 1444 3565 1464
rect 3585 1444 3599 1464
rect 3557 1406 3599 1444
rect 3649 1464 3693 1506
rect 3649 1444 3661 1464
rect 3681 1444 3693 1464
rect 3649 1406 3693 1444
rect 3775 1464 3817 1506
rect 3775 1444 3783 1464
rect 3803 1444 3817 1464
rect 3775 1406 3817 1444
rect 3867 1464 3911 1506
rect 5555 1519 5567 1539
rect 5587 1519 5599 1539
rect 3867 1444 3879 1464
rect 3899 1444 3911 1464
rect 5555 1477 5599 1519
rect 5649 1539 5691 1577
rect 5649 1519 5663 1539
rect 5683 1519 5691 1539
rect 5649 1477 5691 1519
rect 5773 1539 5817 1577
rect 5773 1519 5785 1539
rect 5805 1519 5817 1539
rect 5773 1477 5817 1519
rect 5867 1539 5909 1577
rect 5867 1519 5881 1539
rect 5901 1519 5909 1539
rect 5867 1477 5909 1519
rect 5983 1539 6025 1577
rect 5983 1519 5991 1539
rect 6011 1519 6025 1539
rect 5983 1477 6025 1519
rect 6075 1546 6120 1577
rect 6075 1539 6119 1546
rect 6075 1519 6087 1539
rect 6107 1519 6119 1539
rect 9932 1551 9976 1589
rect 6075 1477 6119 1519
rect 7711 1477 7755 1519
rect 3867 1406 3911 1444
rect 7711 1457 7723 1477
rect 7743 1457 7755 1477
rect 7711 1450 7755 1457
rect 7710 1419 7755 1450
rect 7805 1477 7847 1519
rect 7805 1457 7819 1477
rect 7839 1457 7847 1477
rect 7805 1419 7847 1457
rect 7921 1477 7963 1519
rect 7921 1457 7929 1477
rect 7949 1457 7963 1477
rect 7921 1419 7963 1457
rect 8013 1477 8057 1519
rect 8013 1457 8025 1477
rect 8045 1457 8057 1477
rect 8013 1419 8057 1457
rect 8139 1477 8181 1519
rect 8139 1457 8147 1477
rect 8167 1457 8181 1477
rect 8139 1419 8181 1457
rect 8231 1477 8275 1519
rect 9932 1531 9944 1551
rect 9964 1531 9976 1551
rect 8231 1457 8243 1477
rect 8263 1457 8275 1477
rect 9932 1489 9976 1531
rect 10026 1551 10068 1589
rect 10026 1531 10040 1551
rect 10060 1531 10068 1551
rect 10026 1489 10068 1531
rect 10150 1551 10194 1589
rect 10150 1531 10162 1551
rect 10182 1531 10194 1551
rect 10150 1489 10194 1531
rect 10244 1551 10286 1589
rect 10244 1531 10258 1551
rect 10278 1531 10286 1551
rect 10244 1489 10286 1531
rect 10360 1551 10402 1589
rect 10360 1531 10368 1551
rect 10388 1531 10402 1551
rect 10360 1489 10402 1531
rect 10452 1558 10497 1589
rect 10452 1551 10496 1558
rect 10452 1531 10464 1551
rect 10484 1531 10496 1551
rect 14296 1564 14340 1602
rect 10452 1489 10496 1531
rect 12088 1489 12132 1531
rect 8231 1419 8275 1457
rect 294 1300 338 1338
rect 294 1280 306 1300
rect 326 1280 338 1300
rect 294 1238 338 1280
rect 388 1300 430 1338
rect 388 1280 402 1300
rect 422 1280 430 1300
rect 388 1238 430 1280
rect 512 1300 556 1338
rect 512 1280 524 1300
rect 544 1280 556 1300
rect 512 1238 556 1280
rect 606 1300 648 1338
rect 606 1280 620 1300
rect 640 1280 648 1300
rect 606 1238 648 1280
rect 722 1300 764 1338
rect 722 1280 730 1300
rect 750 1280 764 1300
rect 722 1238 764 1280
rect 814 1307 859 1338
rect 814 1300 858 1307
rect 814 1280 826 1300
rect 846 1280 858 1300
rect 814 1238 858 1280
rect 12088 1469 12100 1489
rect 12120 1469 12132 1489
rect 12088 1462 12132 1469
rect 12087 1431 12132 1462
rect 12182 1489 12224 1531
rect 12182 1469 12196 1489
rect 12216 1469 12224 1489
rect 12182 1431 12224 1469
rect 12298 1489 12340 1531
rect 12298 1469 12306 1489
rect 12326 1469 12340 1489
rect 12298 1431 12340 1469
rect 12390 1489 12434 1531
rect 12390 1469 12402 1489
rect 12422 1469 12434 1489
rect 12390 1431 12434 1469
rect 12516 1489 12558 1531
rect 12516 1469 12524 1489
rect 12544 1469 12558 1489
rect 12516 1431 12558 1469
rect 12608 1489 12652 1531
rect 14296 1544 14308 1564
rect 14328 1544 14340 1564
rect 12608 1469 12620 1489
rect 12640 1469 12652 1489
rect 14296 1502 14340 1544
rect 14390 1564 14432 1602
rect 14390 1544 14404 1564
rect 14424 1544 14432 1564
rect 14390 1502 14432 1544
rect 14514 1564 14558 1602
rect 14514 1544 14526 1564
rect 14546 1544 14558 1564
rect 14514 1502 14558 1544
rect 14608 1564 14650 1602
rect 14608 1544 14622 1564
rect 14642 1544 14650 1564
rect 14608 1502 14650 1544
rect 14724 1564 14766 1602
rect 14724 1544 14732 1564
rect 14752 1544 14766 1564
rect 14724 1502 14766 1544
rect 14816 1571 14861 1602
rect 14816 1564 14860 1571
rect 14816 1544 14828 1564
rect 14848 1544 14860 1564
rect 14816 1502 14860 1544
rect 16452 1502 16496 1544
rect 12608 1431 12652 1469
rect 4658 1313 4702 1351
rect 4658 1293 4670 1313
rect 4690 1293 4702 1313
rect 2550 1236 2594 1278
rect 2550 1216 2562 1236
rect 2582 1216 2594 1236
rect 2550 1209 2594 1216
rect 2549 1178 2594 1209
rect 2644 1236 2686 1278
rect 2644 1216 2658 1236
rect 2678 1216 2686 1236
rect 2644 1178 2686 1216
rect 2760 1236 2802 1278
rect 2760 1216 2768 1236
rect 2788 1216 2802 1236
rect 2760 1178 2802 1216
rect 2852 1236 2896 1278
rect 2852 1216 2864 1236
rect 2884 1216 2896 1236
rect 2852 1178 2896 1216
rect 2978 1236 3020 1278
rect 2978 1216 2986 1236
rect 3006 1216 3020 1236
rect 2978 1178 3020 1216
rect 3070 1236 3114 1278
rect 4658 1251 4702 1293
rect 4752 1313 4794 1351
rect 4752 1293 4766 1313
rect 4786 1293 4794 1313
rect 4752 1251 4794 1293
rect 4876 1313 4920 1351
rect 4876 1293 4888 1313
rect 4908 1293 4920 1313
rect 4876 1251 4920 1293
rect 4970 1313 5012 1351
rect 4970 1293 4984 1313
rect 5004 1293 5012 1313
rect 4970 1251 5012 1293
rect 5086 1313 5128 1351
rect 5086 1293 5094 1313
rect 5114 1293 5128 1313
rect 5086 1251 5128 1293
rect 5178 1320 5223 1351
rect 5178 1313 5222 1320
rect 5178 1293 5190 1313
rect 5210 1293 5222 1313
rect 5178 1251 5222 1293
rect 16452 1482 16464 1502
rect 16484 1482 16496 1502
rect 16452 1475 16496 1482
rect 16451 1444 16496 1475
rect 16546 1502 16588 1544
rect 16546 1482 16560 1502
rect 16580 1482 16588 1502
rect 16546 1444 16588 1482
rect 16662 1502 16704 1544
rect 16662 1482 16670 1502
rect 16690 1482 16704 1502
rect 16662 1444 16704 1482
rect 16754 1502 16798 1544
rect 16754 1482 16766 1502
rect 16786 1482 16798 1502
rect 16754 1444 16798 1482
rect 16880 1502 16922 1544
rect 16880 1482 16888 1502
rect 16908 1482 16922 1502
rect 16880 1444 16922 1482
rect 16972 1502 17016 1544
rect 16972 1482 16984 1502
rect 17004 1482 17016 1502
rect 16972 1444 17016 1482
rect 9035 1325 9079 1363
rect 9035 1305 9047 1325
rect 9067 1305 9079 1325
rect 3070 1216 3082 1236
rect 3102 1216 3114 1236
rect 3070 1178 3114 1216
rect 1092 1116 1136 1154
rect 1092 1096 1104 1116
rect 1124 1096 1136 1116
rect 1092 1054 1136 1096
rect 1186 1116 1228 1154
rect 1186 1096 1200 1116
rect 1220 1096 1228 1116
rect 1186 1054 1228 1096
rect 1310 1116 1354 1154
rect 1310 1096 1322 1116
rect 1342 1096 1354 1116
rect 1310 1054 1354 1096
rect 1404 1116 1446 1154
rect 1404 1096 1418 1116
rect 1438 1096 1446 1116
rect 1404 1054 1446 1096
rect 1520 1116 1562 1154
rect 1520 1096 1528 1116
rect 1548 1096 1562 1116
rect 1520 1054 1562 1096
rect 1612 1123 1657 1154
rect 1612 1116 1656 1123
rect 1612 1096 1624 1116
rect 1644 1096 1656 1116
rect 1612 1054 1656 1096
rect 6914 1249 6958 1291
rect 6914 1229 6926 1249
rect 6946 1229 6958 1249
rect 6914 1222 6958 1229
rect 6913 1191 6958 1222
rect 7008 1249 7050 1291
rect 7008 1229 7022 1249
rect 7042 1229 7050 1249
rect 7008 1191 7050 1229
rect 7124 1249 7166 1291
rect 7124 1229 7132 1249
rect 7152 1229 7166 1249
rect 7124 1191 7166 1229
rect 7216 1249 7260 1291
rect 7216 1229 7228 1249
rect 7248 1229 7260 1249
rect 7216 1191 7260 1229
rect 7342 1249 7384 1291
rect 7342 1229 7350 1249
rect 7370 1229 7384 1249
rect 7342 1191 7384 1229
rect 7434 1249 7478 1291
rect 9035 1263 9079 1305
rect 9129 1325 9171 1363
rect 9129 1305 9143 1325
rect 9163 1305 9171 1325
rect 9129 1263 9171 1305
rect 9253 1325 9297 1363
rect 9253 1305 9265 1325
rect 9285 1305 9297 1325
rect 9253 1263 9297 1305
rect 9347 1325 9389 1363
rect 9347 1305 9361 1325
rect 9381 1305 9389 1325
rect 9347 1263 9389 1305
rect 9463 1325 9505 1363
rect 9463 1305 9471 1325
rect 9491 1305 9505 1325
rect 9463 1263 9505 1305
rect 9555 1332 9600 1363
rect 9555 1325 9599 1332
rect 9555 1305 9567 1325
rect 9587 1305 9599 1325
rect 9555 1263 9599 1305
rect 13399 1338 13443 1376
rect 13399 1318 13411 1338
rect 13431 1318 13443 1338
rect 7434 1229 7446 1249
rect 7466 1229 7478 1249
rect 7434 1191 7478 1229
rect 5456 1129 5500 1167
rect 5456 1109 5468 1129
rect 5488 1109 5500 1129
rect 3348 1052 3392 1094
rect 3348 1032 3360 1052
rect 3380 1032 3392 1052
rect 3348 1025 3392 1032
rect 3347 994 3392 1025
rect 3442 1052 3484 1094
rect 3442 1032 3456 1052
rect 3476 1032 3484 1052
rect 3442 994 3484 1032
rect 3558 1052 3600 1094
rect 3558 1032 3566 1052
rect 3586 1032 3600 1052
rect 3558 994 3600 1032
rect 3650 1052 3694 1094
rect 3650 1032 3662 1052
rect 3682 1032 3694 1052
rect 3650 994 3694 1032
rect 3776 1052 3818 1094
rect 3776 1032 3784 1052
rect 3804 1032 3818 1052
rect 3776 994 3818 1032
rect 3868 1052 3912 1094
rect 5456 1067 5500 1109
rect 5550 1129 5592 1167
rect 5550 1109 5564 1129
rect 5584 1109 5592 1129
rect 5550 1067 5592 1109
rect 5674 1129 5718 1167
rect 5674 1109 5686 1129
rect 5706 1109 5718 1129
rect 5674 1067 5718 1109
rect 5768 1129 5810 1167
rect 5768 1109 5782 1129
rect 5802 1109 5810 1129
rect 5768 1067 5810 1109
rect 5884 1129 5926 1167
rect 5884 1109 5892 1129
rect 5912 1109 5926 1129
rect 5884 1067 5926 1109
rect 5976 1136 6021 1167
rect 5976 1129 6020 1136
rect 5976 1109 5988 1129
rect 6008 1109 6020 1129
rect 5976 1067 6020 1109
rect 11291 1261 11335 1303
rect 11291 1241 11303 1261
rect 11323 1241 11335 1261
rect 11291 1234 11335 1241
rect 11290 1203 11335 1234
rect 11385 1261 11427 1303
rect 11385 1241 11399 1261
rect 11419 1241 11427 1261
rect 11385 1203 11427 1241
rect 11501 1261 11543 1303
rect 11501 1241 11509 1261
rect 11529 1241 11543 1261
rect 11501 1203 11543 1241
rect 11593 1261 11637 1303
rect 11593 1241 11605 1261
rect 11625 1241 11637 1261
rect 11593 1203 11637 1241
rect 11719 1261 11761 1303
rect 11719 1241 11727 1261
rect 11747 1241 11761 1261
rect 11719 1203 11761 1241
rect 11811 1261 11855 1303
rect 13399 1276 13443 1318
rect 13493 1338 13535 1376
rect 13493 1318 13507 1338
rect 13527 1318 13535 1338
rect 13493 1276 13535 1318
rect 13617 1338 13661 1376
rect 13617 1318 13629 1338
rect 13649 1318 13661 1338
rect 13617 1276 13661 1318
rect 13711 1338 13753 1376
rect 13711 1318 13725 1338
rect 13745 1318 13753 1338
rect 13711 1276 13753 1318
rect 13827 1338 13869 1376
rect 13827 1318 13835 1338
rect 13855 1318 13869 1338
rect 13827 1276 13869 1318
rect 13919 1345 13964 1376
rect 13919 1338 13963 1345
rect 13919 1318 13931 1338
rect 13951 1318 13963 1338
rect 13919 1276 13963 1318
rect 11811 1241 11823 1261
rect 11843 1241 11855 1261
rect 11811 1203 11855 1241
rect 9833 1141 9877 1179
rect 9833 1121 9845 1141
rect 9865 1121 9877 1141
rect 3868 1032 3880 1052
rect 3900 1032 3912 1052
rect 3868 994 3912 1032
rect 7712 1065 7756 1107
rect 7712 1045 7724 1065
rect 7744 1045 7756 1065
rect 7712 1038 7756 1045
rect 7711 1007 7756 1038
rect 7806 1065 7848 1107
rect 7806 1045 7820 1065
rect 7840 1045 7848 1065
rect 7806 1007 7848 1045
rect 7922 1065 7964 1107
rect 7922 1045 7930 1065
rect 7950 1045 7964 1065
rect 7922 1007 7964 1045
rect 8014 1065 8058 1107
rect 8014 1045 8026 1065
rect 8046 1045 8058 1065
rect 8014 1007 8058 1045
rect 8140 1065 8182 1107
rect 8140 1045 8148 1065
rect 8168 1045 8182 1065
rect 8140 1007 8182 1045
rect 8232 1065 8276 1107
rect 9833 1079 9877 1121
rect 9927 1141 9969 1179
rect 9927 1121 9941 1141
rect 9961 1121 9969 1141
rect 9927 1079 9969 1121
rect 10051 1141 10095 1179
rect 10051 1121 10063 1141
rect 10083 1121 10095 1141
rect 10051 1079 10095 1121
rect 10145 1141 10187 1179
rect 10145 1121 10159 1141
rect 10179 1121 10187 1141
rect 10145 1079 10187 1121
rect 10261 1141 10303 1179
rect 10261 1121 10269 1141
rect 10289 1121 10303 1141
rect 10261 1079 10303 1121
rect 10353 1148 10398 1179
rect 10353 1141 10397 1148
rect 10353 1121 10365 1141
rect 10385 1121 10397 1141
rect 10353 1079 10397 1121
rect 15655 1274 15699 1316
rect 15655 1254 15667 1274
rect 15687 1254 15699 1274
rect 15655 1247 15699 1254
rect 15654 1216 15699 1247
rect 15749 1274 15791 1316
rect 15749 1254 15763 1274
rect 15783 1254 15791 1274
rect 15749 1216 15791 1254
rect 15865 1274 15907 1316
rect 15865 1254 15873 1274
rect 15893 1254 15907 1274
rect 15865 1216 15907 1254
rect 15957 1274 16001 1316
rect 15957 1254 15969 1274
rect 15989 1254 16001 1274
rect 15957 1216 16001 1254
rect 16083 1274 16125 1316
rect 16083 1254 16091 1274
rect 16111 1254 16125 1274
rect 16083 1216 16125 1254
rect 16175 1274 16219 1316
rect 16175 1254 16187 1274
rect 16207 1254 16219 1274
rect 16175 1216 16219 1254
rect 14197 1154 14241 1192
rect 14197 1134 14209 1154
rect 14229 1134 14241 1154
rect 8232 1045 8244 1065
rect 8264 1045 8276 1065
rect 8232 1007 8276 1045
rect 12089 1077 12133 1119
rect 12089 1057 12101 1077
rect 12121 1057 12133 1077
rect 12089 1050 12133 1057
rect 12088 1019 12133 1050
rect 12183 1077 12225 1119
rect 12183 1057 12197 1077
rect 12217 1057 12225 1077
rect 12183 1019 12225 1057
rect 12299 1077 12341 1119
rect 12299 1057 12307 1077
rect 12327 1057 12341 1077
rect 12299 1019 12341 1057
rect 12391 1077 12435 1119
rect 12391 1057 12403 1077
rect 12423 1057 12435 1077
rect 12391 1019 12435 1057
rect 12517 1077 12559 1119
rect 12517 1057 12525 1077
rect 12545 1057 12559 1077
rect 12517 1019 12559 1057
rect 12609 1077 12653 1119
rect 14197 1092 14241 1134
rect 14291 1154 14333 1192
rect 14291 1134 14305 1154
rect 14325 1134 14333 1154
rect 14291 1092 14333 1134
rect 14415 1154 14459 1192
rect 14415 1134 14427 1154
rect 14447 1134 14459 1154
rect 14415 1092 14459 1134
rect 14509 1154 14551 1192
rect 14509 1134 14523 1154
rect 14543 1134 14551 1154
rect 14509 1092 14551 1134
rect 14625 1154 14667 1192
rect 14625 1134 14633 1154
rect 14653 1134 14667 1154
rect 14625 1092 14667 1134
rect 14717 1161 14762 1192
rect 14717 1154 14761 1161
rect 14717 1134 14729 1154
rect 14749 1134 14761 1154
rect 14717 1092 14761 1134
rect 12609 1057 12621 1077
rect 12641 1057 12653 1077
rect 12609 1019 12653 1057
rect 16453 1090 16497 1132
rect 16453 1070 16465 1090
rect 16485 1070 16497 1090
rect 16453 1063 16497 1070
rect 16452 1032 16497 1063
rect 16547 1090 16589 1132
rect 16547 1070 16561 1090
rect 16581 1070 16589 1090
rect 16547 1032 16589 1070
rect 16663 1090 16705 1132
rect 16663 1070 16671 1090
rect 16691 1070 16705 1090
rect 16663 1032 16705 1070
rect 16755 1090 16799 1132
rect 16755 1070 16767 1090
rect 16787 1070 16799 1090
rect 16755 1032 16799 1070
rect 16881 1090 16923 1132
rect 16881 1070 16889 1090
rect 16909 1070 16923 1090
rect 16881 1032 16923 1070
rect 16973 1090 17017 1132
rect 16973 1070 16985 1090
rect 17005 1070 17017 1090
rect 16973 1032 17017 1070
rect 295 888 339 926
rect 295 868 307 888
rect 327 868 339 888
rect 295 826 339 868
rect 389 888 431 926
rect 389 868 403 888
rect 423 868 431 888
rect 389 826 431 868
rect 513 888 557 926
rect 513 868 525 888
rect 545 868 557 888
rect 513 826 557 868
rect 607 888 649 926
rect 607 868 621 888
rect 641 868 649 888
rect 607 826 649 868
rect 723 888 765 926
rect 723 868 731 888
rect 751 868 765 888
rect 723 826 765 868
rect 815 895 860 926
rect 815 888 859 895
rect 815 868 827 888
rect 847 868 859 888
rect 815 826 859 868
rect 4659 901 4703 939
rect 4659 881 4671 901
rect 4691 881 4703 901
rect 4659 839 4703 881
rect 4753 901 4795 939
rect 4753 881 4767 901
rect 4787 881 4795 901
rect 4753 839 4795 881
rect 4877 901 4921 939
rect 4877 881 4889 901
rect 4909 881 4921 901
rect 4877 839 4921 881
rect 4971 901 5013 939
rect 4971 881 4985 901
rect 5005 881 5013 901
rect 4971 839 5013 881
rect 5087 901 5129 939
rect 5087 881 5095 901
rect 5115 881 5129 901
rect 5087 839 5129 881
rect 5179 908 5224 939
rect 5179 901 5223 908
rect 5179 881 5191 901
rect 5211 881 5223 901
rect 5179 839 5223 881
rect 9036 913 9080 951
rect 9036 893 9048 913
rect 9068 893 9080 913
rect 9036 851 9080 893
rect 9130 913 9172 951
rect 9130 893 9144 913
rect 9164 893 9172 913
rect 9130 851 9172 893
rect 9254 913 9298 951
rect 9254 893 9266 913
rect 9286 893 9298 913
rect 9254 851 9298 893
rect 9348 913 9390 951
rect 9348 893 9362 913
rect 9382 893 9390 913
rect 9348 851 9390 893
rect 9464 913 9506 951
rect 9464 893 9472 913
rect 9492 893 9506 913
rect 9464 851 9506 893
rect 9556 920 9601 951
rect 9556 913 9600 920
rect 9556 893 9568 913
rect 9588 893 9600 913
rect 9556 851 9600 893
rect 13400 926 13444 964
rect 13400 906 13412 926
rect 13432 906 13444 926
rect 13400 864 13444 906
rect 13494 926 13536 964
rect 13494 906 13508 926
rect 13528 906 13536 926
rect 13494 864 13536 906
rect 13618 926 13662 964
rect 13618 906 13630 926
rect 13650 906 13662 926
rect 13618 864 13662 906
rect 13712 926 13754 964
rect 13712 906 13726 926
rect 13746 906 13754 926
rect 13712 864 13754 906
rect 13828 926 13870 964
rect 13828 906 13836 926
rect 13856 906 13870 926
rect 13828 864 13870 906
rect 13920 933 13965 964
rect 13920 926 13964 933
rect 13920 906 13932 926
rect 13952 906 13964 926
rect 13920 864 13964 906
rect 1508 312 1552 350
rect 1508 292 1520 312
rect 1540 292 1552 312
rect 1508 250 1552 292
rect 1602 312 1644 350
rect 1602 292 1616 312
rect 1636 292 1644 312
rect 1602 250 1644 292
rect 1726 312 1770 350
rect 1726 292 1738 312
rect 1758 292 1770 312
rect 1726 250 1770 292
rect 1820 312 1862 350
rect 1820 292 1834 312
rect 1854 292 1862 312
rect 1820 250 1862 292
rect 1936 312 1978 350
rect 1936 292 1944 312
rect 1964 292 1978 312
rect 1936 250 1978 292
rect 2028 319 2073 350
rect 5872 325 5916 363
rect 2028 312 2072 319
rect 2028 292 2040 312
rect 2060 292 2072 312
rect 2028 250 2072 292
rect 5872 305 5884 325
rect 5904 305 5916 325
rect 3997 238 4041 276
rect 3997 218 4009 238
rect 4029 218 4041 238
rect 3997 176 4041 218
rect 4091 238 4133 276
rect 4091 218 4105 238
rect 4125 218 4133 238
rect 4091 176 4133 218
rect 4215 238 4259 276
rect 4215 218 4227 238
rect 4247 218 4259 238
rect 4215 176 4259 218
rect 4309 238 4351 276
rect 4309 218 4323 238
rect 4343 218 4351 238
rect 4309 176 4351 218
rect 4425 238 4467 276
rect 4425 218 4433 238
rect 4453 218 4467 238
rect 4425 176 4467 218
rect 4517 245 4562 276
rect 5872 263 5916 305
rect 5966 325 6008 363
rect 5966 305 5980 325
rect 6000 305 6008 325
rect 5966 263 6008 305
rect 6090 325 6134 363
rect 6090 305 6102 325
rect 6122 305 6134 325
rect 6090 263 6134 305
rect 6184 325 6226 363
rect 6184 305 6198 325
rect 6218 305 6226 325
rect 6184 263 6226 305
rect 6300 325 6342 363
rect 6300 305 6308 325
rect 6328 305 6342 325
rect 6300 263 6342 305
rect 6392 332 6437 363
rect 10249 337 10293 375
rect 6392 325 6436 332
rect 6392 305 6404 325
rect 6424 305 6436 325
rect 10249 317 10261 337
rect 10281 317 10293 337
rect 6392 263 6436 305
rect 4517 238 4561 245
rect 4517 218 4529 238
rect 4549 218 4561 238
rect 4517 176 4561 218
rect 8445 262 8489 300
rect 8445 242 8457 262
rect 8477 242 8489 262
rect 8445 200 8489 242
rect 8539 262 8581 300
rect 8539 242 8553 262
rect 8573 242 8581 262
rect 8539 200 8581 242
rect 8663 262 8707 300
rect 8663 242 8675 262
rect 8695 242 8707 262
rect 8663 200 8707 242
rect 8757 262 8799 300
rect 8757 242 8771 262
rect 8791 242 8799 262
rect 8757 200 8799 242
rect 8873 262 8915 300
rect 8873 242 8881 262
rect 8901 242 8915 262
rect 8873 200 8915 242
rect 8965 269 9010 300
rect 10249 275 10293 317
rect 10343 337 10385 375
rect 10343 317 10357 337
rect 10377 317 10385 337
rect 10343 275 10385 317
rect 10467 337 10511 375
rect 10467 317 10479 337
rect 10499 317 10511 337
rect 10467 275 10511 317
rect 10561 337 10603 375
rect 10561 317 10575 337
rect 10595 317 10603 337
rect 10561 275 10603 317
rect 10677 337 10719 375
rect 10677 317 10685 337
rect 10705 317 10719 337
rect 10677 275 10719 317
rect 10769 344 10814 375
rect 14613 350 14657 388
rect 10769 337 10813 344
rect 10769 317 10781 337
rect 10801 317 10813 337
rect 10769 275 10813 317
rect 14613 330 14625 350
rect 14645 330 14657 350
rect 8965 262 9009 269
rect 8965 242 8977 262
rect 8997 242 9009 262
rect 8965 200 9009 242
rect 12738 263 12782 301
rect 12738 243 12750 263
rect 12770 243 12782 263
rect 12738 201 12782 243
rect 12832 263 12874 301
rect 12832 243 12846 263
rect 12866 243 12874 263
rect 12832 201 12874 243
rect 12956 263 13000 301
rect 12956 243 12968 263
rect 12988 243 13000 263
rect 12956 201 13000 243
rect 13050 263 13092 301
rect 13050 243 13064 263
rect 13084 243 13092 263
rect 13050 201 13092 243
rect 13166 263 13208 301
rect 13166 243 13174 263
rect 13194 243 13208 263
rect 13166 201 13208 243
rect 13258 270 13303 301
rect 14613 288 14657 330
rect 14707 350 14749 388
rect 14707 330 14721 350
rect 14741 330 14749 350
rect 14707 288 14749 330
rect 14831 350 14875 388
rect 14831 330 14843 350
rect 14863 330 14875 350
rect 14831 288 14875 330
rect 14925 350 14967 388
rect 14925 330 14939 350
rect 14959 330 14967 350
rect 14925 288 14967 330
rect 15041 350 15083 388
rect 15041 330 15049 350
rect 15069 330 15083 350
rect 15041 288 15083 330
rect 15133 357 15178 388
rect 15133 350 15177 357
rect 15133 330 15145 350
rect 15165 330 15177 350
rect 15133 288 15177 330
rect 13258 263 13302 270
rect 13258 243 13270 263
rect 13290 243 13302 263
rect 13258 201 13302 243
<< ndiffc >>
rect 3480 8719 3500 8739
rect 3583 8715 3603 8735
rect 3691 8715 3711 8735
rect 3794 8719 3814 8739
rect 3909 8715 3929 8735
rect 4012 8719 4032 8739
rect 4199 8726 4217 8744
rect 263 8664 281 8682
rect 7844 8732 7864 8752
rect 7947 8728 7967 8748
rect 8055 8728 8075 8748
rect 8158 8732 8178 8752
rect 8273 8728 8293 8748
rect 8376 8732 8396 8752
rect 8563 8739 8581 8757
rect 4627 8677 4645 8695
rect 261 8565 279 8583
rect 4197 8627 4215 8645
rect 12221 8744 12241 8764
rect 12324 8740 12344 8760
rect 12432 8740 12452 8760
rect 12535 8744 12555 8764
rect 12650 8740 12670 8760
rect 12753 8744 12773 8764
rect 12940 8751 12958 8769
rect 9004 8689 9022 8707
rect 4625 8578 4643 8596
rect 2683 8491 2703 8511
rect 2786 8487 2806 8507
rect 2894 8487 2914 8507
rect 2997 8491 3017 8511
rect 3112 8487 3132 8507
rect 8561 8640 8579 8658
rect 16585 8757 16605 8777
rect 16688 8753 16708 8773
rect 16796 8753 16816 8773
rect 16899 8757 16919 8777
rect 17014 8753 17034 8773
rect 17117 8757 17137 8777
rect 17304 8764 17322 8782
rect 13368 8702 13386 8720
rect 9002 8590 9020 8608
rect 3215 8491 3235 8511
rect 4192 8508 4210 8526
rect 7047 8504 7067 8524
rect 7150 8500 7170 8520
rect 7258 8500 7278 8520
rect 7361 8504 7381 8524
rect 7476 8500 7496 8520
rect 12938 8652 12956 8670
rect 13366 8603 13384 8621
rect 7579 8504 7599 8524
rect 8556 8521 8574 8539
rect 11424 8516 11444 8536
rect 11527 8512 11547 8532
rect 11635 8512 11655 8532
rect 11738 8516 11758 8536
rect 11853 8512 11873 8532
rect 17302 8665 17320 8683
rect 11956 8516 11976 8536
rect 12933 8533 12951 8551
rect 15788 8529 15808 8549
rect 15891 8525 15911 8545
rect 15999 8525 16019 8545
rect 16102 8529 16122 8549
rect 16217 8525 16237 8545
rect 16320 8529 16340 8549
rect 17297 8546 17315 8564
rect 4190 8409 4208 8427
rect 258 8340 276 8358
rect 8554 8422 8572 8440
rect 3481 8307 3501 8327
rect 256 8241 274 8259
rect 427 8257 447 8277
rect 530 8261 550 8281
rect 645 8257 665 8277
rect 748 8261 768 8281
rect 856 8261 876 8281
rect 3584 8303 3604 8323
rect 3692 8303 3712 8323
rect 3795 8307 3815 8327
rect 3910 8303 3930 8323
rect 4013 8307 4033 8327
rect 4186 8325 4204 8343
rect 4622 8353 4640 8371
rect 959 8257 979 8277
rect 12931 8434 12949 8452
rect 7845 8320 7865 8340
rect 4184 8226 4202 8244
rect 4620 8254 4638 8272
rect 4791 8270 4811 8290
rect 4894 8274 4914 8294
rect 5009 8270 5029 8290
rect 5112 8274 5132 8294
rect 5220 8274 5240 8294
rect 7948 8316 7968 8336
rect 8056 8316 8076 8336
rect 8159 8320 8179 8340
rect 8274 8316 8294 8336
rect 8377 8320 8397 8340
rect 8550 8338 8568 8356
rect 8999 8365 9017 8383
rect 5323 8270 5343 8290
rect 252 8157 270 8175
rect 17295 8447 17313 8465
rect 12222 8332 12242 8352
rect 8548 8239 8566 8257
rect 8997 8266 9015 8284
rect 9168 8282 9188 8302
rect 9271 8286 9291 8306
rect 9386 8282 9406 8302
rect 9489 8286 9509 8306
rect 9597 8286 9617 8306
rect 12325 8328 12345 8348
rect 12433 8328 12453 8348
rect 12536 8332 12556 8352
rect 12651 8328 12671 8348
rect 12754 8332 12774 8352
rect 12927 8350 12945 8368
rect 13363 8378 13381 8396
rect 9700 8282 9720 8302
rect 4616 8170 4634 8188
rect 250 8058 268 8076
rect 1225 8073 1245 8093
rect 1328 8077 1348 8097
rect 1443 8073 1463 8093
rect 1546 8077 1566 8097
rect 1654 8077 1674 8097
rect 1757 8073 1777 8093
rect 2584 8081 2604 8101
rect 2687 8077 2707 8097
rect 2795 8077 2815 8097
rect 2898 8081 2918 8101
rect 3013 8077 3033 8097
rect 16586 8345 16606 8365
rect 12925 8251 12943 8269
rect 13361 8279 13379 8297
rect 13532 8295 13552 8315
rect 13635 8299 13655 8319
rect 13750 8295 13770 8315
rect 13853 8299 13873 8319
rect 13961 8299 13981 8319
rect 16689 8341 16709 8361
rect 16797 8341 16817 8361
rect 16900 8345 16920 8365
rect 17015 8341 17035 8361
rect 17118 8345 17138 8365
rect 17291 8363 17309 8381
rect 14064 8295 14084 8315
rect 8993 8182 9011 8200
rect 3116 8081 3136 8101
rect 4614 8071 4632 8089
rect 5589 8086 5609 8106
rect 245 7939 263 7957
rect 5692 8090 5712 8110
rect 5807 8086 5827 8106
rect 5910 8090 5930 8110
rect 6018 8090 6038 8110
rect 6121 8086 6141 8106
rect 6948 8094 6968 8114
rect 7051 8090 7071 8110
rect 7159 8090 7179 8110
rect 7262 8094 7282 8114
rect 7377 8090 7397 8110
rect 17289 8264 17307 8282
rect 13357 8195 13375 8213
rect 7480 8094 7500 8114
rect 4181 8001 4199 8019
rect 4609 7952 4627 7970
rect 8991 8083 9009 8101
rect 9966 8098 9986 8118
rect 10069 8102 10089 8122
rect 10184 8098 10204 8118
rect 10287 8102 10307 8122
rect 10395 8102 10415 8122
rect 10498 8098 10518 8118
rect 11325 8106 11345 8126
rect 11428 8102 11448 8122
rect 11536 8102 11556 8122
rect 11639 8106 11659 8126
rect 11754 8102 11774 8122
rect 11857 8106 11877 8126
rect 13355 8096 13373 8114
rect 14330 8111 14350 8131
rect 8545 8014 8563 8032
rect 4179 7902 4197 7920
rect 243 7840 261 7858
rect 428 7845 448 7865
rect 531 7849 551 7869
rect 646 7845 666 7865
rect 749 7849 769 7869
rect 857 7849 877 7869
rect 960 7845 980 7865
rect 8986 7964 9004 7982
rect 14433 8115 14453 8135
rect 14548 8111 14568 8131
rect 14651 8115 14671 8135
rect 14759 8115 14779 8135
rect 14862 8111 14882 8131
rect 15689 8119 15709 8139
rect 15792 8115 15812 8135
rect 15900 8115 15920 8135
rect 16003 8119 16023 8139
rect 16118 8115 16138 8135
rect 16221 8119 16241 8139
rect 12922 8026 12940 8044
rect 8543 7915 8561 7933
rect 4607 7853 4625 7871
rect 4792 7858 4812 7878
rect 4895 7862 4915 7882
rect 5010 7858 5030 7878
rect 5113 7862 5133 7882
rect 5221 7862 5241 7882
rect 5324 7858 5344 7878
rect 13350 7977 13368 7995
rect 17286 8039 17304 8057
rect 12920 7927 12938 7945
rect 8984 7865 9002 7883
rect 9169 7870 9189 7890
rect 9272 7874 9292 7894
rect 9387 7870 9407 7890
rect 9490 7874 9510 7894
rect 9598 7874 9618 7894
rect 9701 7870 9721 7890
rect 17284 7940 17302 7958
rect 13348 7878 13366 7896
rect 13533 7883 13553 7903
rect 13636 7887 13656 7907
rect 13751 7883 13771 7903
rect 13854 7887 13874 7907
rect 13962 7887 13982 7907
rect 14065 7883 14085 7903
rect 3463 7701 3483 7721
rect 3566 7697 3586 7717
rect 3674 7697 3694 7717
rect 3777 7701 3797 7721
rect 3892 7697 3912 7717
rect 3995 7701 4015 7721
rect 4182 7708 4200 7726
rect 246 7646 264 7664
rect 7827 7714 7847 7734
rect 7930 7710 7950 7730
rect 8038 7710 8058 7730
rect 8141 7714 8161 7734
rect 8256 7710 8276 7730
rect 8359 7714 8379 7734
rect 8546 7721 8564 7739
rect 4610 7659 4628 7677
rect 244 7547 262 7565
rect 4180 7609 4198 7627
rect 12204 7726 12224 7746
rect 12307 7722 12327 7742
rect 12415 7722 12435 7742
rect 12518 7726 12538 7746
rect 12633 7722 12653 7742
rect 12736 7726 12756 7746
rect 12923 7733 12941 7751
rect 8987 7671 9005 7689
rect 4608 7560 4626 7578
rect 1307 7465 1327 7485
rect 1410 7469 1430 7489
rect 1525 7465 1545 7485
rect 1628 7469 1648 7489
rect 1736 7469 1756 7489
rect 1839 7465 1859 7485
rect 2666 7473 2686 7493
rect 2769 7469 2789 7489
rect 2877 7469 2897 7489
rect 2980 7473 3000 7493
rect 3095 7469 3115 7489
rect 8544 7622 8562 7640
rect 16568 7739 16588 7759
rect 16671 7735 16691 7755
rect 16779 7735 16799 7755
rect 16882 7739 16902 7759
rect 16997 7735 17017 7755
rect 17100 7739 17120 7759
rect 17287 7746 17305 7764
rect 13351 7684 13369 7702
rect 8985 7572 9003 7590
rect 3198 7473 3218 7493
rect 4175 7490 4193 7508
rect 5671 7478 5691 7498
rect 5774 7482 5794 7502
rect 5889 7478 5909 7498
rect 5992 7482 6012 7502
rect 6100 7482 6120 7502
rect 6203 7478 6223 7498
rect 7030 7486 7050 7506
rect 7133 7482 7153 7502
rect 7241 7482 7261 7502
rect 7344 7486 7364 7506
rect 7459 7482 7479 7502
rect 7562 7486 7582 7506
rect 8539 7503 8557 7521
rect 12921 7634 12939 7652
rect 13349 7585 13367 7603
rect 10048 7490 10068 7510
rect 4173 7391 4191 7409
rect 241 7322 259 7340
rect 10151 7494 10171 7514
rect 10266 7490 10286 7510
rect 10369 7494 10389 7514
rect 10477 7494 10497 7514
rect 10580 7490 10600 7510
rect 11407 7498 11427 7518
rect 11510 7494 11530 7514
rect 11618 7494 11638 7514
rect 11721 7498 11741 7518
rect 11836 7494 11856 7514
rect 17285 7647 17303 7665
rect 11939 7498 11959 7518
rect 12916 7515 12934 7533
rect 14412 7503 14432 7523
rect 8537 7404 8555 7422
rect 3464 7289 3484 7309
rect 239 7223 257 7241
rect 410 7239 430 7259
rect 513 7243 533 7263
rect 628 7239 648 7259
rect 731 7243 751 7263
rect 839 7243 859 7263
rect 3567 7285 3587 7305
rect 3675 7285 3695 7305
rect 3778 7289 3798 7309
rect 3893 7285 3913 7305
rect 3996 7289 4016 7309
rect 4169 7307 4187 7325
rect 4605 7335 4623 7353
rect 942 7239 962 7259
rect 14515 7507 14535 7527
rect 14630 7503 14650 7523
rect 14733 7507 14753 7527
rect 14841 7507 14861 7527
rect 14944 7503 14964 7523
rect 15771 7511 15791 7531
rect 15874 7507 15894 7527
rect 15982 7507 16002 7527
rect 16085 7511 16105 7531
rect 16200 7507 16220 7527
rect 16303 7511 16323 7531
rect 17280 7528 17298 7546
rect 12914 7416 12932 7434
rect 7828 7302 7848 7322
rect 4167 7208 4185 7226
rect 4603 7236 4621 7254
rect 4774 7252 4794 7272
rect 4877 7256 4897 7276
rect 4992 7252 5012 7272
rect 5095 7256 5115 7276
rect 5203 7256 5223 7276
rect 7931 7298 7951 7318
rect 8039 7298 8059 7318
rect 8142 7302 8162 7322
rect 8257 7298 8277 7318
rect 8360 7302 8380 7322
rect 8533 7320 8551 7338
rect 8982 7347 9000 7365
rect 5306 7252 5326 7272
rect 235 7139 253 7157
rect 17278 7429 17296 7447
rect 12205 7314 12225 7334
rect 8531 7221 8549 7239
rect 8980 7248 8998 7266
rect 9151 7264 9171 7284
rect 9254 7268 9274 7288
rect 9369 7264 9389 7284
rect 9472 7268 9492 7288
rect 9580 7268 9600 7288
rect 12308 7310 12328 7330
rect 12416 7310 12436 7330
rect 12519 7314 12539 7334
rect 12634 7310 12654 7330
rect 12737 7314 12757 7334
rect 12910 7332 12928 7350
rect 13346 7360 13364 7378
rect 9683 7264 9703 7284
rect 4599 7152 4617 7170
rect 233 7040 251 7058
rect 1208 7055 1228 7075
rect 1311 7059 1331 7079
rect 1426 7055 1446 7075
rect 1529 7059 1549 7079
rect 1637 7059 1657 7079
rect 1740 7055 1760 7075
rect 2501 7065 2521 7085
rect 2604 7061 2624 7081
rect 2712 7061 2732 7081
rect 2815 7065 2835 7085
rect 2930 7061 2950 7081
rect 16569 7327 16589 7347
rect 12908 7233 12926 7251
rect 13344 7261 13362 7279
rect 13515 7277 13535 7297
rect 13618 7281 13638 7301
rect 13733 7277 13753 7297
rect 13836 7281 13856 7301
rect 13944 7281 13964 7301
rect 16672 7323 16692 7343
rect 16780 7323 16800 7343
rect 16883 7327 16903 7347
rect 16998 7323 17018 7343
rect 17101 7327 17121 7347
rect 17274 7345 17292 7363
rect 14047 7277 14067 7297
rect 8976 7164 8994 7182
rect 3033 7065 3053 7085
rect 228 6921 246 6939
rect 4597 7053 4615 7071
rect 5572 7068 5592 7088
rect 5675 7072 5695 7092
rect 5790 7068 5810 7088
rect 5893 7072 5913 7092
rect 6001 7072 6021 7092
rect 6104 7068 6124 7088
rect 6865 7078 6885 7098
rect 6968 7074 6988 7094
rect 7076 7074 7096 7094
rect 7179 7078 7199 7098
rect 7294 7074 7314 7094
rect 17272 7246 17290 7264
rect 13340 7177 13358 7195
rect 7397 7078 7417 7098
rect 4164 6983 4182 7001
rect 4592 6934 4610 6952
rect 8974 7065 8992 7083
rect 9949 7080 9969 7100
rect 10052 7084 10072 7104
rect 10167 7080 10187 7100
rect 10270 7084 10290 7104
rect 10378 7084 10398 7104
rect 10481 7080 10501 7100
rect 11242 7090 11262 7110
rect 11345 7086 11365 7106
rect 11453 7086 11473 7106
rect 11556 7090 11576 7110
rect 11671 7086 11691 7106
rect 11774 7090 11794 7110
rect 8528 6996 8546 7014
rect 4162 6884 4180 6902
rect 226 6822 244 6840
rect 411 6827 431 6847
rect 514 6831 534 6851
rect 629 6827 649 6847
rect 732 6831 752 6851
rect 840 6831 860 6851
rect 943 6827 963 6847
rect 8969 6946 8987 6964
rect 13338 7078 13356 7096
rect 14313 7093 14333 7113
rect 14416 7097 14436 7117
rect 14531 7093 14551 7113
rect 14634 7097 14654 7117
rect 14742 7097 14762 7117
rect 14845 7093 14865 7113
rect 15606 7103 15626 7123
rect 15709 7099 15729 7119
rect 15817 7099 15837 7119
rect 15920 7103 15940 7123
rect 16035 7099 16055 7119
rect 16138 7103 16158 7123
rect 12905 7008 12923 7026
rect 8526 6897 8544 6915
rect 4590 6835 4608 6853
rect 4775 6840 4795 6860
rect 4878 6844 4898 6864
rect 4993 6840 5013 6860
rect 5096 6844 5116 6864
rect 5204 6844 5224 6864
rect 5307 6840 5327 6860
rect 13333 6959 13351 6977
rect 17269 7021 17287 7039
rect 12903 6909 12921 6927
rect 8967 6847 8985 6865
rect 9152 6852 9172 6872
rect 9255 6856 9275 6876
rect 9370 6852 9390 6872
rect 9473 6856 9493 6876
rect 9581 6856 9601 6876
rect 9684 6852 9704 6872
rect 17267 6922 17285 6940
rect 13331 6860 13349 6878
rect 13516 6865 13536 6885
rect 13619 6869 13639 6889
rect 13734 6865 13754 6885
rect 13837 6869 13857 6889
rect 13945 6869 13965 6889
rect 14048 6865 14068 6885
rect 3443 6683 3463 6703
rect 3546 6679 3566 6699
rect 3654 6679 3674 6699
rect 3757 6683 3777 6703
rect 3872 6679 3892 6699
rect 3975 6683 3995 6703
rect 4162 6690 4180 6708
rect 226 6628 244 6646
rect 7807 6696 7827 6716
rect 7910 6692 7930 6712
rect 8018 6692 8038 6712
rect 8121 6696 8141 6716
rect 8236 6692 8256 6712
rect 8339 6696 8359 6716
rect 8526 6703 8544 6721
rect 4590 6641 4608 6659
rect 224 6529 242 6547
rect 4160 6591 4178 6609
rect 12184 6708 12204 6728
rect 12287 6704 12307 6724
rect 12395 6704 12415 6724
rect 12498 6708 12518 6728
rect 12613 6704 12633 6724
rect 12716 6708 12736 6728
rect 12903 6715 12921 6733
rect 8967 6653 8985 6671
rect 4588 6542 4606 6560
rect 1353 6445 1373 6465
rect 1456 6449 1476 6469
rect 1571 6445 1591 6465
rect 1674 6449 1694 6469
rect 1782 6449 1802 6469
rect 1885 6445 1905 6465
rect 2646 6455 2666 6475
rect 2749 6451 2769 6471
rect 2857 6451 2877 6471
rect 2960 6455 2980 6475
rect 3075 6451 3095 6471
rect 3178 6455 3198 6475
rect 4155 6472 4173 6490
rect 8524 6604 8542 6622
rect 16548 6721 16568 6741
rect 16651 6717 16671 6737
rect 16759 6717 16779 6737
rect 16862 6721 16882 6741
rect 16977 6717 16997 6737
rect 17080 6721 17100 6741
rect 17267 6728 17285 6746
rect 13331 6666 13349 6684
rect 8965 6554 8983 6572
rect 5717 6458 5737 6478
rect 5820 6462 5840 6482
rect 5935 6458 5955 6478
rect 6038 6462 6058 6482
rect 6146 6462 6166 6482
rect 6249 6458 6269 6478
rect 7010 6468 7030 6488
rect 7113 6464 7133 6484
rect 7221 6464 7241 6484
rect 7324 6468 7344 6488
rect 7439 6464 7459 6484
rect 7542 6468 7562 6488
rect 8519 6485 8537 6503
rect 12901 6616 12919 6634
rect 13329 6567 13347 6585
rect 10094 6470 10114 6490
rect 4153 6373 4171 6391
rect 221 6304 239 6322
rect 10197 6474 10217 6494
rect 10312 6470 10332 6490
rect 10415 6474 10435 6494
rect 10523 6474 10543 6494
rect 10626 6470 10646 6490
rect 11387 6480 11407 6500
rect 11490 6476 11510 6496
rect 11598 6476 11618 6496
rect 11701 6480 11721 6500
rect 11816 6476 11836 6496
rect 11919 6480 11939 6500
rect 12896 6497 12914 6515
rect 17265 6629 17283 6647
rect 14458 6483 14478 6503
rect 8517 6386 8535 6404
rect 3444 6271 3464 6291
rect 219 6205 237 6223
rect 390 6221 410 6241
rect 493 6225 513 6245
rect 608 6221 628 6241
rect 711 6225 731 6245
rect 819 6225 839 6245
rect 3547 6267 3567 6287
rect 3655 6267 3675 6287
rect 3758 6271 3778 6291
rect 3873 6267 3893 6287
rect 3976 6271 3996 6291
rect 4149 6289 4167 6307
rect 4585 6317 4603 6335
rect 922 6221 942 6241
rect 14561 6487 14581 6507
rect 14676 6483 14696 6503
rect 14779 6487 14799 6507
rect 14887 6487 14907 6507
rect 14990 6483 15010 6503
rect 15751 6493 15771 6513
rect 15854 6489 15874 6509
rect 15962 6489 15982 6509
rect 16065 6493 16085 6513
rect 16180 6489 16200 6509
rect 16283 6493 16303 6513
rect 17260 6510 17278 6528
rect 12894 6398 12912 6416
rect 7808 6284 7828 6304
rect 4147 6190 4165 6208
rect 4583 6218 4601 6236
rect 4754 6234 4774 6254
rect 4857 6238 4877 6258
rect 4972 6234 4992 6254
rect 5075 6238 5095 6258
rect 5183 6238 5203 6258
rect 7911 6280 7931 6300
rect 8019 6280 8039 6300
rect 8122 6284 8142 6304
rect 8237 6280 8257 6300
rect 8340 6284 8360 6304
rect 8513 6302 8531 6320
rect 8962 6329 8980 6347
rect 5286 6234 5306 6254
rect 215 6121 233 6139
rect 17258 6411 17276 6429
rect 12185 6296 12205 6316
rect 8511 6203 8529 6221
rect 8960 6230 8978 6248
rect 9131 6246 9151 6266
rect 9234 6250 9254 6270
rect 9349 6246 9369 6266
rect 9452 6250 9472 6270
rect 9560 6250 9580 6270
rect 12288 6292 12308 6312
rect 12396 6292 12416 6312
rect 12499 6296 12519 6316
rect 12614 6292 12634 6312
rect 12717 6296 12737 6316
rect 12890 6314 12908 6332
rect 13326 6342 13344 6360
rect 9663 6246 9683 6266
rect 4579 6134 4597 6152
rect 213 6022 231 6040
rect 1188 6037 1208 6057
rect 1291 6041 1311 6061
rect 1406 6037 1426 6057
rect 1509 6041 1529 6061
rect 1617 6041 1637 6061
rect 1720 6037 1740 6057
rect 2547 6045 2567 6065
rect 2650 6041 2670 6061
rect 2758 6041 2778 6061
rect 2861 6045 2881 6065
rect 2976 6041 2996 6061
rect 16549 6309 16569 6329
rect 12888 6215 12906 6233
rect 13324 6243 13342 6261
rect 13495 6259 13515 6279
rect 13598 6263 13618 6283
rect 13713 6259 13733 6279
rect 13816 6263 13836 6283
rect 13924 6263 13944 6283
rect 16652 6305 16672 6325
rect 16760 6305 16780 6325
rect 16863 6309 16883 6329
rect 16978 6305 16998 6325
rect 17081 6309 17101 6329
rect 17254 6327 17272 6345
rect 14027 6259 14047 6279
rect 8956 6146 8974 6164
rect 3079 6045 3099 6065
rect 4577 6035 4595 6053
rect 5552 6050 5572 6070
rect 208 5903 226 5921
rect 5655 6054 5675 6074
rect 5770 6050 5790 6070
rect 5873 6054 5893 6074
rect 5981 6054 6001 6074
rect 6084 6050 6104 6070
rect 6911 6058 6931 6078
rect 7014 6054 7034 6074
rect 7122 6054 7142 6074
rect 7225 6058 7245 6078
rect 7340 6054 7360 6074
rect 17252 6228 17270 6246
rect 13320 6159 13338 6177
rect 7443 6058 7463 6078
rect 4144 5965 4162 5983
rect 4572 5916 4590 5934
rect 8954 6047 8972 6065
rect 9929 6062 9949 6082
rect 10032 6066 10052 6086
rect 10147 6062 10167 6082
rect 10250 6066 10270 6086
rect 10358 6066 10378 6086
rect 10461 6062 10481 6082
rect 11288 6070 11308 6090
rect 11391 6066 11411 6086
rect 11499 6066 11519 6086
rect 11602 6070 11622 6090
rect 11717 6066 11737 6086
rect 11820 6070 11840 6090
rect 13318 6060 13336 6078
rect 14293 6075 14313 6095
rect 8508 5978 8526 5996
rect 4142 5866 4160 5884
rect 206 5804 224 5822
rect 391 5809 411 5829
rect 494 5813 514 5833
rect 609 5809 629 5829
rect 712 5813 732 5833
rect 820 5813 840 5833
rect 923 5809 943 5829
rect 8949 5928 8967 5946
rect 14396 6079 14416 6099
rect 14511 6075 14531 6095
rect 14614 6079 14634 6099
rect 14722 6079 14742 6099
rect 14825 6075 14845 6095
rect 15652 6083 15672 6103
rect 15755 6079 15775 6099
rect 15863 6079 15883 6099
rect 15966 6083 15986 6103
rect 16081 6079 16101 6099
rect 16184 6083 16204 6103
rect 12885 5990 12903 6008
rect 8506 5879 8524 5897
rect 4570 5817 4588 5835
rect 4755 5822 4775 5842
rect 4858 5826 4878 5846
rect 4973 5822 4993 5842
rect 5076 5826 5096 5846
rect 5184 5826 5204 5846
rect 5287 5822 5307 5842
rect 13313 5941 13331 5959
rect 17249 6003 17267 6021
rect 12883 5891 12901 5909
rect 8947 5829 8965 5847
rect 9132 5834 9152 5854
rect 9235 5838 9255 5858
rect 9350 5834 9370 5854
rect 9453 5838 9473 5858
rect 9561 5838 9581 5858
rect 9664 5834 9684 5854
rect 17247 5904 17265 5922
rect 13311 5842 13329 5860
rect 13496 5847 13516 5867
rect 13599 5851 13619 5871
rect 13714 5847 13734 5867
rect 13817 5851 13837 5871
rect 13925 5851 13945 5871
rect 14028 5847 14048 5867
rect 3426 5665 3446 5685
rect 3529 5661 3549 5681
rect 3637 5661 3657 5681
rect 3740 5665 3760 5685
rect 3855 5661 3875 5681
rect 3958 5665 3978 5685
rect 4145 5672 4163 5690
rect 209 5610 227 5628
rect 7790 5678 7810 5698
rect 7893 5674 7913 5694
rect 8001 5674 8021 5694
rect 8104 5678 8124 5698
rect 8219 5674 8239 5694
rect 8322 5678 8342 5698
rect 8509 5685 8527 5703
rect 4573 5623 4591 5641
rect 207 5511 225 5529
rect 4143 5573 4161 5591
rect 12167 5690 12187 5710
rect 12270 5686 12290 5706
rect 12378 5686 12398 5706
rect 12481 5690 12501 5710
rect 12596 5686 12616 5706
rect 12699 5690 12719 5710
rect 12886 5697 12904 5715
rect 8950 5635 8968 5653
rect 4571 5524 4589 5542
rect 1270 5429 1290 5449
rect 1373 5433 1393 5453
rect 1488 5429 1508 5449
rect 1591 5433 1611 5453
rect 1699 5433 1719 5453
rect 1802 5429 1822 5449
rect 2629 5437 2649 5457
rect 2732 5433 2752 5453
rect 2840 5433 2860 5453
rect 2943 5437 2963 5457
rect 3058 5433 3078 5453
rect 8507 5586 8525 5604
rect 16531 5703 16551 5723
rect 16634 5699 16654 5719
rect 16742 5699 16762 5719
rect 16845 5703 16865 5723
rect 16960 5699 16980 5719
rect 17063 5703 17083 5723
rect 17250 5710 17268 5728
rect 13314 5648 13332 5666
rect 8948 5536 8966 5554
rect 3161 5437 3181 5457
rect 4138 5454 4156 5472
rect 5634 5442 5654 5462
rect 5737 5446 5757 5466
rect 5852 5442 5872 5462
rect 5955 5446 5975 5466
rect 6063 5446 6083 5466
rect 6166 5442 6186 5462
rect 6993 5450 7013 5470
rect 7096 5446 7116 5466
rect 7204 5446 7224 5466
rect 7307 5450 7327 5470
rect 7422 5446 7442 5466
rect 7525 5450 7545 5470
rect 8502 5467 8520 5485
rect 12884 5598 12902 5616
rect 13312 5549 13330 5567
rect 10011 5454 10031 5474
rect 4136 5355 4154 5373
rect 204 5286 222 5304
rect 10114 5458 10134 5478
rect 10229 5454 10249 5474
rect 10332 5458 10352 5478
rect 10440 5458 10460 5478
rect 10543 5454 10563 5474
rect 11370 5462 11390 5482
rect 11473 5458 11493 5478
rect 11581 5458 11601 5478
rect 11684 5462 11704 5482
rect 11799 5458 11819 5478
rect 17248 5611 17266 5629
rect 11902 5462 11922 5482
rect 12879 5479 12897 5497
rect 14375 5467 14395 5487
rect 8500 5368 8518 5386
rect 3427 5253 3447 5273
rect 202 5187 220 5205
rect 373 5203 393 5223
rect 476 5207 496 5227
rect 591 5203 611 5223
rect 694 5207 714 5227
rect 802 5207 822 5227
rect 3530 5249 3550 5269
rect 3638 5249 3658 5269
rect 3741 5253 3761 5273
rect 3856 5249 3876 5269
rect 3959 5253 3979 5273
rect 4132 5271 4150 5289
rect 4568 5299 4586 5317
rect 905 5203 925 5223
rect 14478 5471 14498 5491
rect 14593 5467 14613 5487
rect 14696 5471 14716 5491
rect 14804 5471 14824 5491
rect 14907 5467 14927 5487
rect 15734 5475 15754 5495
rect 15837 5471 15857 5491
rect 15945 5471 15965 5491
rect 16048 5475 16068 5495
rect 16163 5471 16183 5491
rect 16266 5475 16286 5495
rect 17243 5492 17261 5510
rect 12877 5380 12895 5398
rect 7791 5266 7811 5286
rect 4130 5172 4148 5190
rect 4566 5200 4584 5218
rect 4737 5216 4757 5236
rect 4840 5220 4860 5240
rect 4955 5216 4975 5236
rect 5058 5220 5078 5240
rect 5166 5220 5186 5240
rect 7894 5262 7914 5282
rect 8002 5262 8022 5282
rect 8105 5266 8125 5286
rect 8220 5262 8240 5282
rect 8323 5266 8343 5286
rect 8496 5284 8514 5302
rect 8945 5311 8963 5329
rect 5269 5216 5289 5236
rect 198 5103 216 5121
rect 17241 5393 17259 5411
rect 12168 5278 12188 5298
rect 8494 5185 8512 5203
rect 8943 5212 8961 5230
rect 9114 5228 9134 5248
rect 9217 5232 9237 5252
rect 9332 5228 9352 5248
rect 9435 5232 9455 5252
rect 9543 5232 9563 5252
rect 12271 5274 12291 5294
rect 12379 5274 12399 5294
rect 12482 5278 12502 5298
rect 12597 5274 12617 5294
rect 12700 5278 12720 5298
rect 12873 5296 12891 5314
rect 13309 5324 13327 5342
rect 9646 5228 9666 5248
rect 4562 5116 4580 5134
rect 196 5004 214 5022
rect 1171 5019 1191 5039
rect 1274 5023 1294 5043
rect 1389 5019 1409 5039
rect 1492 5023 1512 5043
rect 1600 5023 1620 5043
rect 1703 5019 1723 5039
rect 2325 5031 2345 5051
rect 2428 5027 2448 5047
rect 2536 5027 2556 5047
rect 2639 5031 2659 5051
rect 2754 5027 2774 5047
rect 16532 5291 16552 5311
rect 12871 5197 12889 5215
rect 13307 5225 13325 5243
rect 13478 5241 13498 5261
rect 13581 5245 13601 5265
rect 13696 5241 13716 5261
rect 13799 5245 13819 5265
rect 13907 5245 13927 5265
rect 16635 5287 16655 5307
rect 16743 5287 16763 5307
rect 16846 5291 16866 5311
rect 16961 5287 16981 5307
rect 17064 5291 17084 5311
rect 17237 5309 17255 5327
rect 14010 5241 14030 5261
rect 8939 5128 8957 5146
rect 2857 5031 2877 5051
rect 191 4885 209 4903
rect 4560 5017 4578 5035
rect 5535 5032 5555 5052
rect 5638 5036 5658 5056
rect 5753 5032 5773 5052
rect 5856 5036 5876 5056
rect 5964 5036 5984 5056
rect 6067 5032 6087 5052
rect 6689 5044 6709 5064
rect 6792 5040 6812 5060
rect 6900 5040 6920 5060
rect 7003 5044 7023 5064
rect 7118 5040 7138 5060
rect 17235 5210 17253 5228
rect 13303 5141 13321 5159
rect 7221 5044 7241 5064
rect 4127 4947 4145 4965
rect 4555 4898 4573 4916
rect 8937 5029 8955 5047
rect 9912 5044 9932 5064
rect 10015 5048 10035 5068
rect 10130 5044 10150 5064
rect 10233 5048 10253 5068
rect 10341 5048 10361 5068
rect 10444 5044 10464 5064
rect 11066 5056 11086 5076
rect 11169 5052 11189 5072
rect 11277 5052 11297 5072
rect 11380 5056 11400 5076
rect 11495 5052 11515 5072
rect 11598 5056 11618 5076
rect 8491 4960 8509 4978
rect 4125 4848 4143 4866
rect 189 4786 207 4804
rect 374 4791 394 4811
rect 477 4795 497 4815
rect 592 4791 612 4811
rect 695 4795 715 4815
rect 803 4795 823 4815
rect 906 4791 926 4811
rect 8932 4910 8950 4928
rect 13301 5042 13319 5060
rect 14276 5057 14296 5077
rect 14379 5061 14399 5081
rect 14494 5057 14514 5077
rect 14597 5061 14617 5081
rect 14705 5061 14725 5081
rect 14808 5057 14828 5077
rect 15430 5069 15450 5089
rect 15533 5065 15553 5085
rect 15641 5065 15661 5085
rect 15744 5069 15764 5089
rect 15859 5065 15879 5085
rect 15962 5069 15982 5089
rect 12868 4972 12886 4990
rect 8489 4861 8507 4879
rect 4553 4799 4571 4817
rect 4738 4804 4758 4824
rect 4841 4808 4861 4828
rect 4956 4804 4976 4824
rect 5059 4808 5079 4828
rect 5167 4808 5187 4828
rect 5270 4804 5290 4824
rect 13296 4923 13314 4941
rect 17232 4985 17250 5003
rect 12866 4873 12884 4891
rect 8930 4811 8948 4829
rect 9115 4816 9135 4836
rect 9218 4820 9238 4840
rect 9333 4816 9353 4836
rect 9436 4820 9456 4840
rect 9544 4820 9564 4840
rect 9647 4816 9667 4836
rect 17230 4886 17248 4904
rect 13294 4824 13312 4842
rect 13479 4829 13499 4849
rect 13582 4833 13602 4853
rect 13697 4829 13717 4849
rect 13800 4833 13820 4853
rect 13908 4833 13928 4853
rect 14011 4829 14031 4849
rect 3407 4647 3427 4667
rect 3510 4643 3530 4663
rect 3618 4643 3638 4663
rect 3721 4647 3741 4667
rect 3836 4643 3856 4663
rect 3939 4647 3959 4667
rect 4126 4654 4144 4672
rect 190 4592 208 4610
rect 7771 4660 7791 4680
rect 7874 4656 7894 4676
rect 7982 4656 8002 4676
rect 8085 4660 8105 4680
rect 8200 4656 8220 4676
rect 8303 4660 8323 4680
rect 8490 4667 8508 4685
rect 4554 4605 4572 4623
rect 188 4493 206 4511
rect 4124 4555 4142 4573
rect 12148 4672 12168 4692
rect 12251 4668 12271 4688
rect 12359 4668 12379 4688
rect 12462 4672 12482 4692
rect 12577 4668 12597 4688
rect 12680 4672 12700 4692
rect 12867 4679 12885 4697
rect 8931 4617 8949 4635
rect 4552 4506 4570 4524
rect 1456 4407 1476 4427
rect 1559 4411 1579 4431
rect 1674 4407 1694 4427
rect 1777 4411 1797 4431
rect 1885 4411 1905 4431
rect 1988 4407 2008 4427
rect 2610 4419 2630 4439
rect 2713 4415 2733 4435
rect 2821 4415 2841 4435
rect 2924 4419 2944 4439
rect 3039 4415 3059 4435
rect 3142 4419 3162 4439
rect 4119 4436 4137 4454
rect 8488 4568 8506 4586
rect 16512 4685 16532 4705
rect 16615 4681 16635 4701
rect 16723 4681 16743 4701
rect 16826 4685 16846 4705
rect 16941 4681 16961 4701
rect 17044 4685 17064 4705
rect 17231 4692 17249 4710
rect 13295 4630 13313 4648
rect 8929 4518 8947 4536
rect 5820 4420 5840 4440
rect 5923 4424 5943 4444
rect 6038 4420 6058 4440
rect 6141 4424 6161 4444
rect 6249 4424 6269 4444
rect 6352 4420 6372 4440
rect 6974 4432 6994 4452
rect 7077 4428 7097 4448
rect 7185 4428 7205 4448
rect 7288 4432 7308 4452
rect 7403 4428 7423 4448
rect 7506 4432 7526 4452
rect 8483 4449 8501 4467
rect 12865 4580 12883 4598
rect 13293 4531 13311 4549
rect 10197 4432 10217 4452
rect 4117 4337 4135 4355
rect 185 4268 203 4286
rect 10300 4436 10320 4456
rect 10415 4432 10435 4452
rect 10518 4436 10538 4456
rect 10626 4436 10646 4456
rect 10729 4432 10749 4452
rect 11351 4444 11371 4464
rect 11454 4440 11474 4460
rect 11562 4440 11582 4460
rect 11665 4444 11685 4464
rect 11780 4440 11800 4460
rect 11883 4444 11903 4464
rect 12860 4461 12878 4479
rect 17229 4593 17247 4611
rect 14561 4445 14581 4465
rect 8481 4350 8499 4368
rect 3408 4235 3428 4255
rect 183 4169 201 4187
rect 354 4185 374 4205
rect 457 4189 477 4209
rect 572 4185 592 4205
rect 675 4189 695 4209
rect 783 4189 803 4209
rect 3511 4231 3531 4251
rect 3619 4231 3639 4251
rect 3722 4235 3742 4255
rect 3837 4231 3857 4251
rect 3940 4235 3960 4255
rect 4113 4253 4131 4271
rect 4549 4281 4567 4299
rect 886 4185 906 4205
rect 14664 4449 14684 4469
rect 14779 4445 14799 4465
rect 14882 4449 14902 4469
rect 14990 4449 15010 4469
rect 15093 4445 15113 4465
rect 15715 4457 15735 4477
rect 15818 4453 15838 4473
rect 15926 4453 15946 4473
rect 16029 4457 16049 4477
rect 16144 4453 16164 4473
rect 16247 4457 16267 4477
rect 17224 4474 17242 4492
rect 12858 4362 12876 4380
rect 7772 4248 7792 4268
rect 4111 4154 4129 4172
rect 4547 4182 4565 4200
rect 4718 4198 4738 4218
rect 4821 4202 4841 4222
rect 4936 4198 4956 4218
rect 5039 4202 5059 4222
rect 5147 4202 5167 4222
rect 7875 4244 7895 4264
rect 7983 4244 8003 4264
rect 8086 4248 8106 4268
rect 8201 4244 8221 4264
rect 8304 4248 8324 4268
rect 8477 4266 8495 4284
rect 8926 4293 8944 4311
rect 5250 4198 5270 4218
rect 179 4085 197 4103
rect 17222 4375 17240 4393
rect 12149 4260 12169 4280
rect 8475 4167 8493 4185
rect 8924 4194 8942 4212
rect 9095 4210 9115 4230
rect 9198 4214 9218 4234
rect 9313 4210 9333 4230
rect 9416 4214 9436 4234
rect 9524 4214 9544 4234
rect 12252 4256 12272 4276
rect 12360 4256 12380 4276
rect 12463 4260 12483 4280
rect 12578 4256 12598 4276
rect 12681 4260 12701 4280
rect 12854 4278 12872 4296
rect 13290 4306 13308 4324
rect 9627 4210 9647 4230
rect 4543 4098 4561 4116
rect 177 3986 195 4004
rect 1152 4001 1172 4021
rect 1255 4005 1275 4025
rect 1370 4001 1390 4021
rect 1473 4005 1493 4025
rect 1581 4005 1601 4025
rect 1684 4001 1704 4021
rect 2511 4009 2531 4029
rect 2614 4005 2634 4025
rect 2722 4005 2742 4025
rect 2825 4009 2845 4029
rect 2940 4005 2960 4025
rect 16513 4273 16533 4293
rect 12852 4179 12870 4197
rect 13288 4207 13306 4225
rect 13459 4223 13479 4243
rect 13562 4227 13582 4247
rect 13677 4223 13697 4243
rect 13780 4227 13800 4247
rect 13888 4227 13908 4247
rect 16616 4269 16636 4289
rect 16724 4269 16744 4289
rect 16827 4273 16847 4293
rect 16942 4269 16962 4289
rect 17045 4273 17065 4293
rect 17218 4291 17236 4309
rect 13991 4223 14011 4243
rect 8920 4110 8938 4128
rect 3043 4009 3063 4029
rect 4541 3999 4559 4017
rect 5516 4014 5536 4034
rect 172 3867 190 3885
rect 5619 4018 5639 4038
rect 5734 4014 5754 4034
rect 5837 4018 5857 4038
rect 5945 4018 5965 4038
rect 6048 4014 6068 4034
rect 6875 4022 6895 4042
rect 6978 4018 6998 4038
rect 7086 4018 7106 4038
rect 7189 4022 7209 4042
rect 7304 4018 7324 4038
rect 17216 4192 17234 4210
rect 13284 4123 13302 4141
rect 7407 4022 7427 4042
rect 4108 3929 4126 3947
rect 4536 3880 4554 3898
rect 8918 4011 8936 4029
rect 9893 4026 9913 4046
rect 9996 4030 10016 4050
rect 10111 4026 10131 4046
rect 10214 4030 10234 4050
rect 10322 4030 10342 4050
rect 10425 4026 10445 4046
rect 11252 4034 11272 4054
rect 11355 4030 11375 4050
rect 11463 4030 11483 4050
rect 11566 4034 11586 4054
rect 11681 4030 11701 4050
rect 11784 4034 11804 4054
rect 13282 4024 13300 4042
rect 14257 4039 14277 4059
rect 8472 3942 8490 3960
rect 4106 3830 4124 3848
rect 170 3768 188 3786
rect 355 3773 375 3793
rect 458 3777 478 3797
rect 573 3773 593 3793
rect 676 3777 696 3797
rect 784 3777 804 3797
rect 887 3773 907 3793
rect 8913 3892 8931 3910
rect 14360 4043 14380 4063
rect 14475 4039 14495 4059
rect 14578 4043 14598 4063
rect 14686 4043 14706 4063
rect 14789 4039 14809 4059
rect 15616 4047 15636 4067
rect 15719 4043 15739 4063
rect 15827 4043 15847 4063
rect 15930 4047 15950 4067
rect 16045 4043 16065 4063
rect 16148 4047 16168 4067
rect 12849 3954 12867 3972
rect 8470 3843 8488 3861
rect 4534 3781 4552 3799
rect 4719 3786 4739 3806
rect 4822 3790 4842 3810
rect 4937 3786 4957 3806
rect 5040 3790 5060 3810
rect 5148 3790 5168 3810
rect 5251 3786 5271 3806
rect 13277 3905 13295 3923
rect 17213 3967 17231 3985
rect 12847 3855 12865 3873
rect 8911 3793 8929 3811
rect 9096 3798 9116 3818
rect 9199 3802 9219 3822
rect 9314 3798 9334 3818
rect 9417 3802 9437 3822
rect 9525 3802 9545 3822
rect 9628 3798 9648 3818
rect 17211 3868 17229 3886
rect 13275 3806 13293 3824
rect 13460 3811 13480 3831
rect 13563 3815 13583 3835
rect 13678 3811 13698 3831
rect 13781 3815 13801 3835
rect 13889 3815 13909 3835
rect 13992 3811 14012 3831
rect 3390 3629 3410 3649
rect 3493 3625 3513 3645
rect 3601 3625 3621 3645
rect 3704 3629 3724 3649
rect 3819 3625 3839 3645
rect 3922 3629 3942 3649
rect 4109 3636 4127 3654
rect 173 3574 191 3592
rect 7754 3642 7774 3662
rect 7857 3638 7877 3658
rect 7965 3638 7985 3658
rect 8068 3642 8088 3662
rect 8183 3638 8203 3658
rect 8286 3642 8306 3662
rect 8473 3649 8491 3667
rect 4537 3587 4555 3605
rect 171 3475 189 3493
rect 4107 3537 4125 3555
rect 12131 3654 12151 3674
rect 12234 3650 12254 3670
rect 12342 3650 12362 3670
rect 12445 3654 12465 3674
rect 12560 3650 12580 3670
rect 12663 3654 12683 3674
rect 12850 3661 12868 3679
rect 8914 3599 8932 3617
rect 4535 3488 4553 3506
rect 1234 3393 1254 3413
rect 1337 3397 1357 3417
rect 1452 3393 1472 3413
rect 1555 3397 1575 3417
rect 1663 3397 1683 3417
rect 1766 3393 1786 3413
rect 2593 3401 2613 3421
rect 2696 3397 2716 3417
rect 2804 3397 2824 3417
rect 2907 3401 2927 3421
rect 3022 3397 3042 3417
rect 8471 3550 8489 3568
rect 16495 3667 16515 3687
rect 16598 3663 16618 3683
rect 16706 3663 16726 3683
rect 16809 3667 16829 3687
rect 16924 3663 16944 3683
rect 17027 3667 17047 3687
rect 17214 3674 17232 3692
rect 13278 3612 13296 3630
rect 8912 3500 8930 3518
rect 3125 3401 3145 3421
rect 4102 3418 4120 3436
rect 5598 3406 5618 3426
rect 5701 3410 5721 3430
rect 5816 3406 5836 3426
rect 5919 3410 5939 3430
rect 6027 3410 6047 3430
rect 6130 3406 6150 3426
rect 6957 3414 6977 3434
rect 7060 3410 7080 3430
rect 7168 3410 7188 3430
rect 7271 3414 7291 3434
rect 7386 3410 7406 3430
rect 7489 3414 7509 3434
rect 8466 3431 8484 3449
rect 12848 3562 12866 3580
rect 13276 3513 13294 3531
rect 9975 3418 9995 3438
rect 4100 3319 4118 3337
rect 168 3250 186 3268
rect 10078 3422 10098 3442
rect 10193 3418 10213 3438
rect 10296 3422 10316 3442
rect 10404 3422 10424 3442
rect 10507 3418 10527 3438
rect 11334 3426 11354 3446
rect 11437 3422 11457 3442
rect 11545 3422 11565 3442
rect 11648 3426 11668 3446
rect 11763 3422 11783 3442
rect 17212 3575 17230 3593
rect 11866 3426 11886 3446
rect 12843 3443 12861 3461
rect 14339 3431 14359 3451
rect 8464 3332 8482 3350
rect 3391 3217 3411 3237
rect 166 3151 184 3169
rect 337 3167 357 3187
rect 440 3171 460 3191
rect 555 3167 575 3187
rect 658 3171 678 3191
rect 766 3171 786 3191
rect 3494 3213 3514 3233
rect 3602 3213 3622 3233
rect 3705 3217 3725 3237
rect 3820 3213 3840 3233
rect 3923 3217 3943 3237
rect 4096 3235 4114 3253
rect 4532 3263 4550 3281
rect 869 3167 889 3187
rect 14442 3435 14462 3455
rect 14557 3431 14577 3451
rect 14660 3435 14680 3455
rect 14768 3435 14788 3455
rect 14871 3431 14891 3451
rect 15698 3439 15718 3459
rect 15801 3435 15821 3455
rect 15909 3435 15929 3455
rect 16012 3439 16032 3459
rect 16127 3435 16147 3455
rect 16230 3439 16250 3459
rect 17207 3456 17225 3474
rect 12841 3344 12859 3362
rect 7755 3230 7775 3250
rect 4094 3136 4112 3154
rect 4530 3164 4548 3182
rect 4701 3180 4721 3200
rect 4804 3184 4824 3204
rect 4919 3180 4939 3200
rect 5022 3184 5042 3204
rect 5130 3184 5150 3204
rect 7858 3226 7878 3246
rect 7966 3226 7986 3246
rect 8069 3230 8089 3250
rect 8184 3226 8204 3246
rect 8287 3230 8307 3250
rect 8460 3248 8478 3266
rect 8909 3275 8927 3293
rect 5233 3180 5253 3200
rect 162 3067 180 3085
rect 17205 3357 17223 3375
rect 12132 3242 12152 3262
rect 8458 3149 8476 3167
rect 8907 3176 8925 3194
rect 9078 3192 9098 3212
rect 9181 3196 9201 3216
rect 9296 3192 9316 3212
rect 9399 3196 9419 3216
rect 9507 3196 9527 3216
rect 12235 3238 12255 3258
rect 12343 3238 12363 3258
rect 12446 3242 12466 3262
rect 12561 3238 12581 3258
rect 12664 3242 12684 3262
rect 12837 3260 12855 3278
rect 13273 3288 13291 3306
rect 9610 3192 9630 3212
rect 4526 3080 4544 3098
rect 160 2968 178 2986
rect 1135 2983 1155 3003
rect 1238 2987 1258 3007
rect 1353 2983 1373 3003
rect 1456 2987 1476 3007
rect 1564 2987 1584 3007
rect 1667 2983 1687 3003
rect 2428 2993 2448 3013
rect 2531 2989 2551 3009
rect 2639 2989 2659 3009
rect 2742 2993 2762 3013
rect 2857 2989 2877 3009
rect 16496 3255 16516 3275
rect 12835 3161 12853 3179
rect 13271 3189 13289 3207
rect 13442 3205 13462 3225
rect 13545 3209 13565 3229
rect 13660 3205 13680 3225
rect 13763 3209 13783 3229
rect 13871 3209 13891 3229
rect 16599 3251 16619 3271
rect 16707 3251 16727 3271
rect 16810 3255 16830 3275
rect 16925 3251 16945 3271
rect 17028 3255 17048 3275
rect 17201 3273 17219 3291
rect 13974 3205 13994 3225
rect 8903 3092 8921 3110
rect 2960 2993 2980 3013
rect 155 2849 173 2867
rect 4524 2981 4542 2999
rect 5499 2996 5519 3016
rect 5602 3000 5622 3020
rect 5717 2996 5737 3016
rect 5820 3000 5840 3020
rect 5928 3000 5948 3020
rect 6031 2996 6051 3016
rect 6792 3006 6812 3026
rect 6895 3002 6915 3022
rect 7003 3002 7023 3022
rect 7106 3006 7126 3026
rect 7221 3002 7241 3022
rect 17199 3174 17217 3192
rect 13267 3105 13285 3123
rect 7324 3006 7344 3026
rect 4091 2911 4109 2929
rect 4519 2862 4537 2880
rect 8901 2993 8919 3011
rect 9876 3008 9896 3028
rect 9979 3012 9999 3032
rect 10094 3008 10114 3028
rect 10197 3012 10217 3032
rect 10305 3012 10325 3032
rect 10408 3008 10428 3028
rect 11169 3018 11189 3038
rect 11272 3014 11292 3034
rect 11380 3014 11400 3034
rect 11483 3018 11503 3038
rect 11598 3014 11618 3034
rect 11701 3018 11721 3038
rect 8455 2924 8473 2942
rect 4089 2812 4107 2830
rect 153 2750 171 2768
rect 338 2755 358 2775
rect 441 2759 461 2779
rect 556 2755 576 2775
rect 659 2759 679 2779
rect 767 2759 787 2779
rect 870 2755 890 2775
rect 8896 2874 8914 2892
rect 13265 3006 13283 3024
rect 14240 3021 14260 3041
rect 14343 3025 14363 3045
rect 14458 3021 14478 3041
rect 14561 3025 14581 3045
rect 14669 3025 14689 3045
rect 14772 3021 14792 3041
rect 15533 3031 15553 3051
rect 15636 3027 15656 3047
rect 15744 3027 15764 3047
rect 15847 3031 15867 3051
rect 15962 3027 15982 3047
rect 16065 3031 16085 3051
rect 12832 2936 12850 2954
rect 8453 2825 8471 2843
rect 4517 2763 4535 2781
rect 4702 2768 4722 2788
rect 4805 2772 4825 2792
rect 4920 2768 4940 2788
rect 5023 2772 5043 2792
rect 5131 2772 5151 2792
rect 5234 2768 5254 2788
rect 13260 2887 13278 2905
rect 17196 2949 17214 2967
rect 12830 2837 12848 2855
rect 8894 2775 8912 2793
rect 9079 2780 9099 2800
rect 9182 2784 9202 2804
rect 9297 2780 9317 2800
rect 9400 2784 9420 2804
rect 9508 2784 9528 2804
rect 9611 2780 9631 2800
rect 17194 2850 17212 2868
rect 13258 2788 13276 2806
rect 13443 2793 13463 2813
rect 13546 2797 13566 2817
rect 13661 2793 13681 2813
rect 13764 2797 13784 2817
rect 13872 2797 13892 2817
rect 13975 2793 13995 2813
rect 3370 2611 3390 2631
rect 3473 2607 3493 2627
rect 3581 2607 3601 2627
rect 3684 2611 3704 2631
rect 3799 2607 3819 2627
rect 3902 2611 3922 2631
rect 4089 2618 4107 2636
rect 153 2556 171 2574
rect 7734 2624 7754 2644
rect 7837 2620 7857 2640
rect 7945 2620 7965 2640
rect 8048 2624 8068 2644
rect 8163 2620 8183 2640
rect 8266 2624 8286 2644
rect 8453 2631 8471 2649
rect 4517 2569 4535 2587
rect 151 2457 169 2475
rect 4087 2519 4105 2537
rect 12111 2636 12131 2656
rect 12214 2632 12234 2652
rect 12322 2632 12342 2652
rect 12425 2636 12445 2656
rect 12540 2632 12560 2652
rect 12643 2636 12663 2656
rect 12830 2643 12848 2661
rect 8894 2581 8912 2599
rect 4515 2470 4533 2488
rect 1280 2373 1300 2393
rect 1383 2377 1403 2397
rect 1498 2373 1518 2393
rect 1601 2377 1621 2397
rect 1709 2377 1729 2397
rect 1812 2373 1832 2393
rect 2573 2383 2593 2403
rect 2676 2379 2696 2399
rect 2784 2379 2804 2399
rect 2887 2383 2907 2403
rect 3002 2379 3022 2399
rect 3105 2383 3125 2403
rect 4082 2400 4100 2418
rect 8451 2532 8469 2550
rect 16475 2649 16495 2669
rect 16578 2645 16598 2665
rect 16686 2645 16706 2665
rect 16789 2649 16809 2669
rect 16904 2645 16924 2665
rect 17007 2649 17027 2669
rect 17194 2656 17212 2674
rect 13258 2594 13276 2612
rect 8892 2482 8910 2500
rect 5644 2386 5664 2406
rect 5747 2390 5767 2410
rect 5862 2386 5882 2406
rect 5965 2390 5985 2410
rect 6073 2390 6093 2410
rect 6176 2386 6196 2406
rect 6937 2396 6957 2416
rect 7040 2392 7060 2412
rect 7148 2392 7168 2412
rect 7251 2396 7271 2416
rect 7366 2392 7386 2412
rect 7469 2396 7489 2416
rect 8446 2413 8464 2431
rect 12828 2544 12846 2562
rect 13256 2495 13274 2513
rect 10021 2398 10041 2418
rect 4080 2301 4098 2319
rect 148 2232 166 2250
rect 10124 2402 10144 2422
rect 10239 2398 10259 2418
rect 10342 2402 10362 2422
rect 10450 2402 10470 2422
rect 10553 2398 10573 2418
rect 11314 2408 11334 2428
rect 11417 2404 11437 2424
rect 11525 2404 11545 2424
rect 11628 2408 11648 2428
rect 11743 2404 11763 2424
rect 11846 2408 11866 2428
rect 12823 2425 12841 2443
rect 17192 2557 17210 2575
rect 14385 2411 14405 2431
rect 8444 2314 8462 2332
rect 3371 2199 3391 2219
rect 146 2133 164 2151
rect 317 2149 337 2169
rect 420 2153 440 2173
rect 535 2149 555 2169
rect 638 2153 658 2173
rect 746 2153 766 2173
rect 3474 2195 3494 2215
rect 3582 2195 3602 2215
rect 3685 2199 3705 2219
rect 3800 2195 3820 2215
rect 3903 2199 3923 2219
rect 4076 2217 4094 2235
rect 4512 2245 4530 2263
rect 849 2149 869 2169
rect 14488 2415 14508 2435
rect 14603 2411 14623 2431
rect 14706 2415 14726 2435
rect 14814 2415 14834 2435
rect 14917 2411 14937 2431
rect 15678 2421 15698 2441
rect 15781 2417 15801 2437
rect 15889 2417 15909 2437
rect 15992 2421 16012 2441
rect 16107 2417 16127 2437
rect 16210 2421 16230 2441
rect 17187 2438 17205 2456
rect 12821 2326 12839 2344
rect 7735 2212 7755 2232
rect 4074 2118 4092 2136
rect 4510 2146 4528 2164
rect 4681 2162 4701 2182
rect 4784 2166 4804 2186
rect 4899 2162 4919 2182
rect 5002 2166 5022 2186
rect 5110 2166 5130 2186
rect 7838 2208 7858 2228
rect 7946 2208 7966 2228
rect 8049 2212 8069 2232
rect 8164 2208 8184 2228
rect 8267 2212 8287 2232
rect 8440 2230 8458 2248
rect 8889 2257 8907 2275
rect 5213 2162 5233 2182
rect 142 2049 160 2067
rect 17185 2339 17203 2357
rect 12112 2224 12132 2244
rect 8438 2131 8456 2149
rect 8887 2158 8905 2176
rect 9058 2174 9078 2194
rect 9161 2178 9181 2198
rect 9276 2174 9296 2194
rect 9379 2178 9399 2198
rect 9487 2178 9507 2198
rect 12215 2220 12235 2240
rect 12323 2220 12343 2240
rect 12426 2224 12446 2244
rect 12541 2220 12561 2240
rect 12644 2224 12664 2244
rect 12817 2242 12835 2260
rect 13253 2270 13271 2288
rect 9590 2174 9610 2194
rect 4506 2062 4524 2080
rect 140 1950 158 1968
rect 1115 1965 1135 1985
rect 1218 1969 1238 1989
rect 1333 1965 1353 1985
rect 1436 1969 1456 1989
rect 1544 1969 1564 1989
rect 1647 1965 1667 1985
rect 2474 1973 2494 1993
rect 2577 1969 2597 1989
rect 2685 1969 2705 1989
rect 2788 1973 2808 1993
rect 2903 1969 2923 1989
rect 16476 2237 16496 2257
rect 12815 2143 12833 2161
rect 13251 2171 13269 2189
rect 13422 2187 13442 2207
rect 13525 2191 13545 2211
rect 13640 2187 13660 2207
rect 13743 2191 13763 2211
rect 13851 2191 13871 2211
rect 16579 2233 16599 2253
rect 16687 2233 16707 2253
rect 16790 2237 16810 2257
rect 16905 2233 16925 2253
rect 17008 2237 17028 2257
rect 17181 2255 17199 2273
rect 13954 2187 13974 2207
rect 8883 2074 8901 2092
rect 3006 1973 3026 1993
rect 4504 1963 4522 1981
rect 5479 1978 5499 1998
rect 135 1831 153 1849
rect 5582 1982 5602 2002
rect 5697 1978 5717 1998
rect 5800 1982 5820 2002
rect 5908 1982 5928 2002
rect 6011 1978 6031 1998
rect 6838 1986 6858 2006
rect 6941 1982 6961 2002
rect 7049 1982 7069 2002
rect 7152 1986 7172 2006
rect 7267 1982 7287 2002
rect 17179 2156 17197 2174
rect 13247 2087 13265 2105
rect 7370 1986 7390 2006
rect 4071 1893 4089 1911
rect 4499 1844 4517 1862
rect 8881 1975 8899 1993
rect 9856 1990 9876 2010
rect 9959 1994 9979 2014
rect 10074 1990 10094 2010
rect 10177 1994 10197 2014
rect 10285 1994 10305 2014
rect 10388 1990 10408 2010
rect 11215 1998 11235 2018
rect 11318 1994 11338 2014
rect 11426 1994 11446 2014
rect 11529 1998 11549 2018
rect 11644 1994 11664 2014
rect 11747 1998 11767 2018
rect 13245 1988 13263 2006
rect 14220 2003 14240 2023
rect 8435 1906 8453 1924
rect 4069 1794 4087 1812
rect 133 1732 151 1750
rect 318 1737 338 1757
rect 421 1741 441 1761
rect 536 1737 556 1757
rect 639 1741 659 1761
rect 747 1741 767 1761
rect 850 1737 870 1757
rect 8876 1856 8894 1874
rect 14323 2007 14343 2027
rect 14438 2003 14458 2023
rect 14541 2007 14561 2027
rect 14649 2007 14669 2027
rect 14752 2003 14772 2023
rect 15579 2011 15599 2031
rect 15682 2007 15702 2027
rect 15790 2007 15810 2027
rect 15893 2011 15913 2031
rect 16008 2007 16028 2027
rect 16111 2011 16131 2031
rect 12812 1918 12830 1936
rect 8433 1807 8451 1825
rect 4497 1745 4515 1763
rect 4682 1750 4702 1770
rect 4785 1754 4805 1774
rect 4900 1750 4920 1770
rect 5003 1754 5023 1774
rect 5111 1754 5131 1774
rect 5214 1750 5234 1770
rect 13240 1869 13258 1887
rect 17176 1931 17194 1949
rect 12810 1819 12828 1837
rect 8874 1757 8892 1775
rect 9059 1762 9079 1782
rect 9162 1766 9182 1786
rect 9277 1762 9297 1782
rect 9380 1766 9400 1786
rect 9488 1766 9508 1786
rect 9591 1762 9611 1782
rect 17174 1832 17192 1850
rect 13238 1770 13256 1788
rect 13423 1775 13443 1795
rect 13526 1779 13546 1799
rect 13641 1775 13661 1795
rect 13744 1779 13764 1799
rect 13852 1779 13872 1799
rect 13955 1775 13975 1795
rect 3353 1593 3373 1613
rect 3456 1589 3476 1609
rect 3564 1589 3584 1609
rect 3667 1593 3687 1613
rect 3782 1589 3802 1609
rect 3885 1593 3905 1613
rect 4072 1600 4090 1618
rect 136 1538 154 1556
rect 7717 1606 7737 1626
rect 7820 1602 7840 1622
rect 7928 1602 7948 1622
rect 8031 1606 8051 1626
rect 8146 1602 8166 1622
rect 8249 1606 8269 1626
rect 8436 1613 8454 1631
rect 4500 1551 4518 1569
rect 134 1439 152 1457
rect 4070 1501 4088 1519
rect 12094 1618 12114 1638
rect 12197 1614 12217 1634
rect 12305 1614 12325 1634
rect 12408 1618 12428 1638
rect 12523 1614 12543 1634
rect 12626 1618 12646 1638
rect 12813 1625 12831 1643
rect 8877 1563 8895 1581
rect 4498 1452 4516 1470
rect 1197 1357 1217 1377
rect 1300 1361 1320 1381
rect 1415 1357 1435 1377
rect 1518 1361 1538 1381
rect 1626 1361 1646 1381
rect 1729 1357 1749 1377
rect 2556 1365 2576 1385
rect 2659 1361 2679 1381
rect 2767 1361 2787 1381
rect 2870 1365 2890 1385
rect 2985 1361 3005 1381
rect 8434 1514 8452 1532
rect 16458 1631 16478 1651
rect 16561 1627 16581 1647
rect 16669 1627 16689 1647
rect 16772 1631 16792 1651
rect 16887 1627 16907 1647
rect 16990 1631 17010 1651
rect 17177 1638 17195 1656
rect 13241 1576 13259 1594
rect 8875 1464 8893 1482
rect 3088 1365 3108 1385
rect 4065 1382 4083 1400
rect 5561 1370 5581 1390
rect 5664 1374 5684 1394
rect 5779 1370 5799 1390
rect 5882 1374 5902 1394
rect 5990 1374 6010 1394
rect 6093 1370 6113 1390
rect 6920 1378 6940 1398
rect 7023 1374 7043 1394
rect 7131 1374 7151 1394
rect 7234 1378 7254 1398
rect 7349 1374 7369 1394
rect 7452 1378 7472 1398
rect 8429 1395 8447 1413
rect 12811 1526 12829 1544
rect 13239 1477 13257 1495
rect 9938 1382 9958 1402
rect 4063 1283 4081 1301
rect 131 1214 149 1232
rect 10041 1386 10061 1406
rect 10156 1382 10176 1402
rect 10259 1386 10279 1406
rect 10367 1386 10387 1406
rect 10470 1382 10490 1402
rect 11297 1390 11317 1410
rect 11400 1386 11420 1406
rect 11508 1386 11528 1406
rect 11611 1390 11631 1410
rect 11726 1386 11746 1406
rect 17175 1539 17193 1557
rect 11829 1390 11849 1410
rect 12806 1407 12824 1425
rect 14302 1395 14322 1415
rect 8427 1296 8445 1314
rect 3354 1181 3374 1201
rect 129 1115 147 1133
rect 300 1131 320 1151
rect 403 1135 423 1155
rect 518 1131 538 1151
rect 621 1135 641 1155
rect 729 1135 749 1155
rect 3457 1177 3477 1197
rect 3565 1177 3585 1197
rect 3668 1181 3688 1201
rect 3783 1177 3803 1197
rect 3886 1181 3906 1201
rect 4059 1199 4077 1217
rect 4495 1227 4513 1245
rect 832 1131 852 1151
rect 14405 1399 14425 1419
rect 14520 1395 14540 1415
rect 14623 1399 14643 1419
rect 14731 1399 14751 1419
rect 14834 1395 14854 1415
rect 15661 1403 15681 1423
rect 15764 1399 15784 1419
rect 15872 1399 15892 1419
rect 15975 1403 15995 1423
rect 16090 1399 16110 1419
rect 16193 1403 16213 1423
rect 17170 1420 17188 1438
rect 12804 1308 12822 1326
rect 7718 1194 7738 1214
rect 4057 1100 4075 1118
rect 4493 1128 4511 1146
rect 4664 1144 4684 1164
rect 4767 1148 4787 1168
rect 4882 1144 4902 1164
rect 4985 1148 5005 1168
rect 5093 1148 5113 1168
rect 7821 1190 7841 1210
rect 7929 1190 7949 1210
rect 8032 1194 8052 1214
rect 8147 1190 8167 1210
rect 8250 1194 8270 1214
rect 8423 1212 8441 1230
rect 8872 1239 8890 1257
rect 5196 1144 5216 1164
rect 125 1031 143 1049
rect 17168 1321 17186 1339
rect 12095 1206 12115 1226
rect 8421 1113 8439 1131
rect 8870 1140 8888 1158
rect 9041 1156 9061 1176
rect 9144 1160 9164 1180
rect 9259 1156 9279 1176
rect 9362 1160 9382 1180
rect 9470 1160 9490 1180
rect 12198 1202 12218 1222
rect 12306 1202 12326 1222
rect 12409 1206 12429 1226
rect 12524 1202 12544 1222
rect 12627 1206 12647 1226
rect 12800 1224 12818 1242
rect 13236 1252 13254 1270
rect 9573 1156 9593 1176
rect 4489 1044 4507 1062
rect 16459 1219 16479 1239
rect 12798 1125 12816 1143
rect 13234 1153 13252 1171
rect 13405 1169 13425 1189
rect 13508 1173 13528 1193
rect 13623 1169 13643 1189
rect 13726 1173 13746 1193
rect 13834 1173 13854 1193
rect 16562 1215 16582 1235
rect 16670 1215 16690 1235
rect 16773 1219 16793 1239
rect 16888 1215 16908 1235
rect 16991 1219 17011 1239
rect 17164 1237 17182 1255
rect 13937 1169 13957 1189
rect 8866 1056 8884 1074
rect 17162 1138 17180 1156
rect 13230 1069 13248 1087
rect 123 932 141 950
rect 1098 947 1118 967
rect 1201 951 1221 971
rect 1316 947 1336 967
rect 1419 951 1439 971
rect 1527 951 1547 971
rect 1630 947 1650 967
rect 4487 945 4505 963
rect 5462 960 5482 980
rect 118 813 136 831
rect 5565 964 5585 984
rect 5680 960 5700 980
rect 5783 964 5803 984
rect 5891 964 5911 984
rect 5994 960 6014 980
rect 8864 957 8882 975
rect 9839 972 9859 992
rect 4054 875 4072 893
rect 4482 826 4500 844
rect 9942 976 9962 996
rect 10057 972 10077 992
rect 10160 976 10180 996
rect 10268 976 10288 996
rect 10371 972 10391 992
rect 13228 970 13246 988
rect 14203 985 14223 1005
rect 8418 888 8436 906
rect 4052 776 4070 794
rect 116 714 134 732
rect 301 719 321 739
rect 404 723 424 743
rect 519 719 539 739
rect 622 723 642 743
rect 730 723 750 743
rect 833 719 853 739
rect 8859 838 8877 856
rect 14306 989 14326 1009
rect 14421 985 14441 1005
rect 14524 989 14544 1009
rect 14632 989 14652 1009
rect 14735 985 14755 1005
rect 12795 900 12813 918
rect 8416 789 8434 807
rect 4480 727 4498 745
rect 4665 732 4685 752
rect 4768 736 4788 756
rect 4883 732 4903 752
rect 4986 736 5006 756
rect 5094 736 5114 756
rect 5197 732 5217 752
rect 13223 851 13241 869
rect 17159 913 17177 931
rect 12793 801 12811 819
rect 8857 739 8875 757
rect 9042 744 9062 764
rect 9145 748 9165 768
rect 9260 744 9280 764
rect 9363 748 9383 768
rect 9471 748 9491 768
rect 9574 744 9594 764
rect 17157 814 17175 832
rect 13221 752 13239 770
rect 13406 757 13426 777
rect 13509 761 13529 781
rect 13624 757 13644 777
rect 13727 761 13747 781
rect 13835 761 13855 781
rect 13938 757 13958 777
rect 1514 143 1534 163
rect 1617 147 1637 167
rect 1732 143 1752 163
rect 1835 147 1855 167
rect 1943 147 1963 167
rect 2046 143 2066 163
rect 5878 156 5898 176
rect 5981 160 6001 180
rect 6096 156 6116 176
rect 6199 160 6219 180
rect 6307 160 6327 180
rect 6410 156 6430 176
rect 10255 168 10275 188
rect 10358 172 10378 192
rect 10473 168 10493 188
rect 10576 172 10596 192
rect 10684 172 10704 192
rect 10787 168 10807 188
rect 14619 181 14639 201
rect 14722 185 14742 205
rect 14837 181 14857 201
rect 14940 185 14960 205
rect 15048 185 15068 205
rect 15151 181 15171 201
rect 4003 69 4023 89
rect 4106 73 4126 93
rect 4221 69 4241 89
rect 4324 73 4344 93
rect 4432 73 4452 93
rect 4535 69 4555 89
rect 8451 93 8471 113
rect 8554 97 8574 117
rect 8669 93 8689 113
rect 8772 97 8792 117
rect 8880 97 8900 117
rect 8983 93 9003 113
rect 12744 94 12764 114
rect 12847 98 12867 118
rect 12962 94 12982 114
rect 13065 98 13085 118
rect 13173 98 13193 118
rect 13276 94 13296 114
<< pdiffc >>
rect 3486 8570 3506 8590
rect 3582 8570 3602 8590
rect 3692 8570 3712 8590
rect 3788 8570 3808 8590
rect 3910 8570 3930 8590
rect 4006 8570 4026 8590
rect 7850 8583 7870 8603
rect 7946 8583 7966 8603
rect 8056 8583 8076 8603
rect 8152 8583 8172 8603
rect 8274 8583 8294 8603
rect 8370 8583 8390 8603
rect 12227 8595 12247 8615
rect 12323 8595 12343 8615
rect 12433 8595 12453 8615
rect 12529 8595 12549 8615
rect 12651 8595 12671 8615
rect 12747 8595 12767 8615
rect 16591 8608 16611 8628
rect 16687 8608 16707 8628
rect 16797 8608 16817 8628
rect 16893 8608 16913 8628
rect 17015 8608 17035 8628
rect 17111 8608 17131 8628
rect 433 8406 453 8426
rect 529 8406 549 8426
rect 651 8406 671 8426
rect 747 8406 767 8426
rect 857 8406 877 8426
rect 953 8406 973 8426
rect 4797 8419 4817 8439
rect 2689 8342 2709 8362
rect 2785 8342 2805 8362
rect 2895 8342 2915 8362
rect 2991 8342 3011 8362
rect 3113 8342 3133 8362
rect 4893 8419 4913 8439
rect 5015 8419 5035 8439
rect 5111 8419 5131 8439
rect 5221 8419 5241 8439
rect 5317 8419 5337 8439
rect 9174 8431 9194 8451
rect 3209 8342 3229 8362
rect 1231 8222 1251 8242
rect 1327 8222 1347 8242
rect 1449 8222 1469 8242
rect 1545 8222 1565 8242
rect 1655 8222 1675 8242
rect 1751 8222 1771 8242
rect 7053 8355 7073 8375
rect 7149 8355 7169 8375
rect 7259 8355 7279 8375
rect 7355 8355 7375 8375
rect 7477 8355 7497 8375
rect 9270 8431 9290 8451
rect 9392 8431 9412 8451
rect 9488 8431 9508 8451
rect 9598 8431 9618 8451
rect 9694 8431 9714 8451
rect 13538 8444 13558 8464
rect 7573 8355 7593 8375
rect 5595 8235 5615 8255
rect 3487 8158 3507 8178
rect 3583 8158 3603 8178
rect 3693 8158 3713 8178
rect 3789 8158 3809 8178
rect 3911 8158 3931 8178
rect 5691 8235 5711 8255
rect 5813 8235 5833 8255
rect 5909 8235 5929 8255
rect 6019 8235 6039 8255
rect 6115 8235 6135 8255
rect 11430 8367 11450 8387
rect 11526 8367 11546 8387
rect 11636 8367 11656 8387
rect 11732 8367 11752 8387
rect 11854 8367 11874 8387
rect 13634 8444 13654 8464
rect 13756 8444 13776 8464
rect 13852 8444 13872 8464
rect 13962 8444 13982 8464
rect 14058 8444 14078 8464
rect 11950 8367 11970 8387
rect 9972 8247 9992 8267
rect 4007 8158 4027 8178
rect 7851 8171 7871 8191
rect 7947 8171 7967 8191
rect 8057 8171 8077 8191
rect 8153 8171 8173 8191
rect 8275 8171 8295 8191
rect 10068 8247 10088 8267
rect 10190 8247 10210 8267
rect 10286 8247 10306 8267
rect 10396 8247 10416 8267
rect 10492 8247 10512 8267
rect 15794 8380 15814 8400
rect 15890 8380 15910 8400
rect 16000 8380 16020 8400
rect 16096 8380 16116 8400
rect 16218 8380 16238 8400
rect 16314 8380 16334 8400
rect 14336 8260 14356 8280
rect 8371 8171 8391 8191
rect 434 7994 454 8014
rect 530 7994 550 8014
rect 652 7994 672 8014
rect 748 7994 768 8014
rect 858 7994 878 8014
rect 954 7994 974 8014
rect 12228 8183 12248 8203
rect 12324 8183 12344 8203
rect 12434 8183 12454 8203
rect 12530 8183 12550 8203
rect 12652 8183 12672 8203
rect 14432 8260 14452 8280
rect 14554 8260 14574 8280
rect 14650 8260 14670 8280
rect 14760 8260 14780 8280
rect 14856 8260 14876 8280
rect 12748 8183 12768 8203
rect 2590 7932 2610 7952
rect 2686 7932 2706 7952
rect 2796 7932 2816 7952
rect 2892 7932 2912 7952
rect 3014 7932 3034 7952
rect 4798 8007 4818 8027
rect 3110 7932 3130 7952
rect 4894 8007 4914 8027
rect 5016 8007 5036 8027
rect 5112 8007 5132 8027
rect 5222 8007 5242 8027
rect 5318 8007 5338 8027
rect 16592 8196 16612 8216
rect 16688 8196 16708 8216
rect 16798 8196 16818 8216
rect 16894 8196 16914 8216
rect 17016 8196 17036 8216
rect 17112 8196 17132 8216
rect 6954 7945 6974 7965
rect 7050 7945 7070 7965
rect 7160 7945 7180 7965
rect 7256 7945 7276 7965
rect 7378 7945 7398 7965
rect 9175 8019 9195 8039
rect 7474 7945 7494 7965
rect 9271 8019 9291 8039
rect 9393 8019 9413 8039
rect 9489 8019 9509 8039
rect 9599 8019 9619 8039
rect 9695 8019 9715 8039
rect 11331 7957 11351 7977
rect 11427 7957 11447 7977
rect 11537 7957 11557 7977
rect 11633 7957 11653 7977
rect 11755 7957 11775 7977
rect 13539 8032 13559 8052
rect 11851 7957 11871 7977
rect 13635 8032 13655 8052
rect 13757 8032 13777 8052
rect 13853 8032 13873 8052
rect 13963 8032 13983 8052
rect 14059 8032 14079 8052
rect 15695 7970 15715 7990
rect 15791 7970 15811 7990
rect 15901 7970 15921 7990
rect 15997 7970 16017 7990
rect 16119 7970 16139 7990
rect 16215 7970 16235 7990
rect 1313 7614 1333 7634
rect 1409 7614 1429 7634
rect 1531 7614 1551 7634
rect 1627 7614 1647 7634
rect 1737 7614 1757 7634
rect 1833 7614 1853 7634
rect 3469 7552 3489 7572
rect 3565 7552 3585 7572
rect 3675 7552 3695 7572
rect 3771 7552 3791 7572
rect 3893 7552 3913 7572
rect 5677 7627 5697 7647
rect 3989 7552 4009 7572
rect 5773 7627 5793 7647
rect 5895 7627 5915 7647
rect 5991 7627 6011 7647
rect 6101 7627 6121 7647
rect 6197 7627 6217 7647
rect 7833 7565 7853 7585
rect 7929 7565 7949 7585
rect 8039 7565 8059 7585
rect 8135 7565 8155 7585
rect 8257 7565 8277 7585
rect 10054 7639 10074 7659
rect 8353 7565 8373 7585
rect 10150 7639 10170 7659
rect 10272 7639 10292 7659
rect 10368 7639 10388 7659
rect 10478 7639 10498 7659
rect 10574 7639 10594 7659
rect 416 7388 436 7408
rect 512 7388 532 7408
rect 634 7388 654 7408
rect 730 7388 750 7408
rect 840 7388 860 7408
rect 936 7388 956 7408
rect 12210 7577 12230 7597
rect 12306 7577 12326 7597
rect 12416 7577 12436 7597
rect 12512 7577 12532 7597
rect 12634 7577 12654 7597
rect 14418 7652 14438 7672
rect 12730 7577 12750 7597
rect 14514 7652 14534 7672
rect 14636 7652 14656 7672
rect 14732 7652 14752 7672
rect 14842 7652 14862 7672
rect 14938 7652 14958 7672
rect 4780 7401 4800 7421
rect 2672 7324 2692 7344
rect 2768 7324 2788 7344
rect 2878 7324 2898 7344
rect 2974 7324 2994 7344
rect 3096 7324 3116 7344
rect 4876 7401 4896 7421
rect 4998 7401 5018 7421
rect 5094 7401 5114 7421
rect 5204 7401 5224 7421
rect 5300 7401 5320 7421
rect 16574 7590 16594 7610
rect 16670 7590 16690 7610
rect 16780 7590 16800 7610
rect 16876 7590 16896 7610
rect 16998 7590 17018 7610
rect 17094 7590 17114 7610
rect 9157 7413 9177 7433
rect 3192 7324 3212 7344
rect 1214 7204 1234 7224
rect 1310 7204 1330 7224
rect 1432 7204 1452 7224
rect 1528 7204 1548 7224
rect 1638 7204 1658 7224
rect 1734 7204 1754 7224
rect 7036 7337 7056 7357
rect 7132 7337 7152 7357
rect 7242 7337 7262 7357
rect 7338 7337 7358 7357
rect 7460 7337 7480 7357
rect 9253 7413 9273 7433
rect 9375 7413 9395 7433
rect 9471 7413 9491 7433
rect 9581 7413 9601 7433
rect 9677 7413 9697 7433
rect 13521 7426 13541 7446
rect 7556 7337 7576 7357
rect 5578 7217 5598 7237
rect 3470 7140 3490 7160
rect 3566 7140 3586 7160
rect 3676 7140 3696 7160
rect 3772 7140 3792 7160
rect 3894 7140 3914 7160
rect 5674 7217 5694 7237
rect 5796 7217 5816 7237
rect 5892 7217 5912 7237
rect 6002 7217 6022 7237
rect 6098 7217 6118 7237
rect 11413 7349 11433 7369
rect 11509 7349 11529 7369
rect 11619 7349 11639 7369
rect 11715 7349 11735 7369
rect 11837 7349 11857 7369
rect 13617 7426 13637 7446
rect 13739 7426 13759 7446
rect 13835 7426 13855 7446
rect 13945 7426 13965 7446
rect 14041 7426 14061 7446
rect 11933 7349 11953 7369
rect 9955 7229 9975 7249
rect 3990 7140 4010 7160
rect 7834 7153 7854 7173
rect 7930 7153 7950 7173
rect 8040 7153 8060 7173
rect 8136 7153 8156 7173
rect 8258 7153 8278 7173
rect 10051 7229 10071 7249
rect 10173 7229 10193 7249
rect 10269 7229 10289 7249
rect 10379 7229 10399 7249
rect 10475 7229 10495 7249
rect 15777 7362 15797 7382
rect 15873 7362 15893 7382
rect 15983 7362 16003 7382
rect 16079 7362 16099 7382
rect 16201 7362 16221 7382
rect 16297 7362 16317 7382
rect 14319 7242 14339 7262
rect 8354 7153 8374 7173
rect 417 6976 437 6996
rect 513 6976 533 6996
rect 635 6976 655 6996
rect 731 6976 751 6996
rect 841 6976 861 6996
rect 937 6976 957 6996
rect 12211 7165 12231 7185
rect 12307 7165 12327 7185
rect 12417 7165 12437 7185
rect 12513 7165 12533 7185
rect 12635 7165 12655 7185
rect 14415 7242 14435 7262
rect 14537 7242 14557 7262
rect 14633 7242 14653 7262
rect 14743 7242 14763 7262
rect 14839 7242 14859 7262
rect 12731 7165 12751 7185
rect 2507 6916 2527 6936
rect 2603 6916 2623 6936
rect 2713 6916 2733 6936
rect 2809 6916 2829 6936
rect 2931 6916 2951 6936
rect 4781 6989 4801 7009
rect 3027 6916 3047 6936
rect 4877 6989 4897 7009
rect 4999 6989 5019 7009
rect 5095 6989 5115 7009
rect 5205 6989 5225 7009
rect 5301 6989 5321 7009
rect 16575 7178 16595 7198
rect 16671 7178 16691 7198
rect 16781 7178 16801 7198
rect 16877 7178 16897 7198
rect 16999 7178 17019 7198
rect 17095 7178 17115 7198
rect 6871 6929 6891 6949
rect 6967 6929 6987 6949
rect 7077 6929 7097 6949
rect 7173 6929 7193 6949
rect 7295 6929 7315 6949
rect 9158 7001 9178 7021
rect 7391 6929 7411 6949
rect 9254 7001 9274 7021
rect 9376 7001 9396 7021
rect 9472 7001 9492 7021
rect 9582 7001 9602 7021
rect 9678 7001 9698 7021
rect 11248 6941 11268 6961
rect 11344 6941 11364 6961
rect 11454 6941 11474 6961
rect 11550 6941 11570 6961
rect 11672 6941 11692 6961
rect 13522 7014 13542 7034
rect 11768 6941 11788 6961
rect 13618 7014 13638 7034
rect 13740 7014 13760 7034
rect 13836 7014 13856 7034
rect 13946 7014 13966 7034
rect 14042 7014 14062 7034
rect 15612 6954 15632 6974
rect 15708 6954 15728 6974
rect 15818 6954 15838 6974
rect 15914 6954 15934 6974
rect 16036 6954 16056 6974
rect 16132 6954 16152 6974
rect 1359 6594 1379 6614
rect 1455 6594 1475 6614
rect 1577 6594 1597 6614
rect 1673 6594 1693 6614
rect 1783 6594 1803 6614
rect 1879 6594 1899 6614
rect 3449 6534 3469 6554
rect 3545 6534 3565 6554
rect 3655 6534 3675 6554
rect 3751 6534 3771 6554
rect 3873 6534 3893 6554
rect 5723 6607 5743 6627
rect 3969 6534 3989 6554
rect 5819 6607 5839 6627
rect 5941 6607 5961 6627
rect 6037 6607 6057 6627
rect 6147 6607 6167 6627
rect 6243 6607 6263 6627
rect 7813 6547 7833 6567
rect 7909 6547 7929 6567
rect 8019 6547 8039 6567
rect 8115 6547 8135 6567
rect 8237 6547 8257 6567
rect 10100 6619 10120 6639
rect 8333 6547 8353 6567
rect 10196 6619 10216 6639
rect 10318 6619 10338 6639
rect 10414 6619 10434 6639
rect 10524 6619 10544 6639
rect 10620 6619 10640 6639
rect 396 6370 416 6390
rect 492 6370 512 6390
rect 614 6370 634 6390
rect 710 6370 730 6390
rect 820 6370 840 6390
rect 916 6370 936 6390
rect 12190 6559 12210 6579
rect 12286 6559 12306 6579
rect 12396 6559 12416 6579
rect 12492 6559 12512 6579
rect 12614 6559 12634 6579
rect 14464 6632 14484 6652
rect 12710 6559 12730 6579
rect 14560 6632 14580 6652
rect 14682 6632 14702 6652
rect 14778 6632 14798 6652
rect 14888 6632 14908 6652
rect 14984 6632 15004 6652
rect 4760 6383 4780 6403
rect 2652 6306 2672 6326
rect 2748 6306 2768 6326
rect 2858 6306 2878 6326
rect 2954 6306 2974 6326
rect 3076 6306 3096 6326
rect 4856 6383 4876 6403
rect 4978 6383 4998 6403
rect 5074 6383 5094 6403
rect 5184 6383 5204 6403
rect 5280 6383 5300 6403
rect 16554 6572 16574 6592
rect 16650 6572 16670 6592
rect 16760 6572 16780 6592
rect 16856 6572 16876 6592
rect 16978 6572 16998 6592
rect 17074 6572 17094 6592
rect 9137 6395 9157 6415
rect 3172 6306 3192 6326
rect 1194 6186 1214 6206
rect 1290 6186 1310 6206
rect 1412 6186 1432 6206
rect 1508 6186 1528 6206
rect 1618 6186 1638 6206
rect 1714 6186 1734 6206
rect 7016 6319 7036 6339
rect 7112 6319 7132 6339
rect 7222 6319 7242 6339
rect 7318 6319 7338 6339
rect 7440 6319 7460 6339
rect 9233 6395 9253 6415
rect 9355 6395 9375 6415
rect 9451 6395 9471 6415
rect 9561 6395 9581 6415
rect 9657 6395 9677 6415
rect 13501 6408 13521 6428
rect 7536 6319 7556 6339
rect 5558 6199 5578 6219
rect 3450 6122 3470 6142
rect 3546 6122 3566 6142
rect 3656 6122 3676 6142
rect 3752 6122 3772 6142
rect 3874 6122 3894 6142
rect 5654 6199 5674 6219
rect 5776 6199 5796 6219
rect 5872 6199 5892 6219
rect 5982 6199 6002 6219
rect 6078 6199 6098 6219
rect 11393 6331 11413 6351
rect 11489 6331 11509 6351
rect 11599 6331 11619 6351
rect 11695 6331 11715 6351
rect 11817 6331 11837 6351
rect 13597 6408 13617 6428
rect 13719 6408 13739 6428
rect 13815 6408 13835 6428
rect 13925 6408 13945 6428
rect 14021 6408 14041 6428
rect 11913 6331 11933 6351
rect 9935 6211 9955 6231
rect 3970 6122 3990 6142
rect 7814 6135 7834 6155
rect 7910 6135 7930 6155
rect 8020 6135 8040 6155
rect 8116 6135 8136 6155
rect 8238 6135 8258 6155
rect 10031 6211 10051 6231
rect 10153 6211 10173 6231
rect 10249 6211 10269 6231
rect 10359 6211 10379 6231
rect 10455 6211 10475 6231
rect 15757 6344 15777 6364
rect 15853 6344 15873 6364
rect 15963 6344 15983 6364
rect 16059 6344 16079 6364
rect 16181 6344 16201 6364
rect 16277 6344 16297 6364
rect 14299 6224 14319 6244
rect 8334 6135 8354 6155
rect 397 5958 417 5978
rect 493 5958 513 5978
rect 615 5958 635 5978
rect 711 5958 731 5978
rect 821 5958 841 5978
rect 917 5958 937 5978
rect 12191 6147 12211 6167
rect 12287 6147 12307 6167
rect 12397 6147 12417 6167
rect 12493 6147 12513 6167
rect 12615 6147 12635 6167
rect 14395 6224 14415 6244
rect 14517 6224 14537 6244
rect 14613 6224 14633 6244
rect 14723 6224 14743 6244
rect 14819 6224 14839 6244
rect 12711 6147 12731 6167
rect 2553 5896 2573 5916
rect 2649 5896 2669 5916
rect 2759 5896 2779 5916
rect 2855 5896 2875 5916
rect 2977 5896 2997 5916
rect 4761 5971 4781 5991
rect 3073 5896 3093 5916
rect 4857 5971 4877 5991
rect 4979 5971 4999 5991
rect 5075 5971 5095 5991
rect 5185 5971 5205 5991
rect 5281 5971 5301 5991
rect 16555 6160 16575 6180
rect 16651 6160 16671 6180
rect 16761 6160 16781 6180
rect 16857 6160 16877 6180
rect 16979 6160 16999 6180
rect 17075 6160 17095 6180
rect 6917 5909 6937 5929
rect 7013 5909 7033 5929
rect 7123 5909 7143 5929
rect 7219 5909 7239 5929
rect 7341 5909 7361 5929
rect 9138 5983 9158 6003
rect 7437 5909 7457 5929
rect 9234 5983 9254 6003
rect 9356 5983 9376 6003
rect 9452 5983 9472 6003
rect 9562 5983 9582 6003
rect 9658 5983 9678 6003
rect 11294 5921 11314 5941
rect 11390 5921 11410 5941
rect 11500 5921 11520 5941
rect 11596 5921 11616 5941
rect 11718 5921 11738 5941
rect 13502 5996 13522 6016
rect 11814 5921 11834 5941
rect 13598 5996 13618 6016
rect 13720 5996 13740 6016
rect 13816 5996 13836 6016
rect 13926 5996 13946 6016
rect 14022 5996 14042 6016
rect 15658 5934 15678 5954
rect 15754 5934 15774 5954
rect 15864 5934 15884 5954
rect 15960 5934 15980 5954
rect 16082 5934 16102 5954
rect 16178 5934 16198 5954
rect 1276 5578 1296 5598
rect 1372 5578 1392 5598
rect 1494 5578 1514 5598
rect 1590 5578 1610 5598
rect 1700 5578 1720 5598
rect 1796 5578 1816 5598
rect 3432 5516 3452 5536
rect 3528 5516 3548 5536
rect 3638 5516 3658 5536
rect 3734 5516 3754 5536
rect 3856 5516 3876 5536
rect 5640 5591 5660 5611
rect 3952 5516 3972 5536
rect 5736 5591 5756 5611
rect 5858 5591 5878 5611
rect 5954 5591 5974 5611
rect 6064 5591 6084 5611
rect 6160 5591 6180 5611
rect 7796 5529 7816 5549
rect 7892 5529 7912 5549
rect 8002 5529 8022 5549
rect 8098 5529 8118 5549
rect 8220 5529 8240 5549
rect 10017 5603 10037 5623
rect 8316 5529 8336 5549
rect 10113 5603 10133 5623
rect 10235 5603 10255 5623
rect 10331 5603 10351 5623
rect 10441 5603 10461 5623
rect 10537 5603 10557 5623
rect 379 5352 399 5372
rect 475 5352 495 5372
rect 597 5352 617 5372
rect 693 5352 713 5372
rect 803 5352 823 5372
rect 899 5352 919 5372
rect 12173 5541 12193 5561
rect 12269 5541 12289 5561
rect 12379 5541 12399 5561
rect 12475 5541 12495 5561
rect 12597 5541 12617 5561
rect 14381 5616 14401 5636
rect 12693 5541 12713 5561
rect 14477 5616 14497 5636
rect 14599 5616 14619 5636
rect 14695 5616 14715 5636
rect 14805 5616 14825 5636
rect 14901 5616 14921 5636
rect 4743 5365 4763 5385
rect 2635 5288 2655 5308
rect 2731 5288 2751 5308
rect 2841 5288 2861 5308
rect 2937 5288 2957 5308
rect 3059 5288 3079 5308
rect 4839 5365 4859 5385
rect 4961 5365 4981 5385
rect 5057 5365 5077 5385
rect 5167 5365 5187 5385
rect 5263 5365 5283 5385
rect 16537 5554 16557 5574
rect 16633 5554 16653 5574
rect 16743 5554 16763 5574
rect 16839 5554 16859 5574
rect 16961 5554 16981 5574
rect 17057 5554 17077 5574
rect 9120 5377 9140 5397
rect 3155 5288 3175 5308
rect 1177 5168 1197 5188
rect 1273 5168 1293 5188
rect 1395 5168 1415 5188
rect 1491 5168 1511 5188
rect 1601 5168 1621 5188
rect 1697 5168 1717 5188
rect 6999 5301 7019 5321
rect 7095 5301 7115 5321
rect 7205 5301 7225 5321
rect 7301 5301 7321 5321
rect 7423 5301 7443 5321
rect 9216 5377 9236 5397
rect 9338 5377 9358 5397
rect 9434 5377 9454 5397
rect 9544 5377 9564 5397
rect 9640 5377 9660 5397
rect 13484 5390 13504 5410
rect 7519 5301 7539 5321
rect 5541 5181 5561 5201
rect 3433 5104 3453 5124
rect 3529 5104 3549 5124
rect 3639 5104 3659 5124
rect 3735 5104 3755 5124
rect 3857 5104 3877 5124
rect 5637 5181 5657 5201
rect 5759 5181 5779 5201
rect 5855 5181 5875 5201
rect 5965 5181 5985 5201
rect 6061 5181 6081 5201
rect 11376 5313 11396 5333
rect 11472 5313 11492 5333
rect 11582 5313 11602 5333
rect 11678 5313 11698 5333
rect 11800 5313 11820 5333
rect 13580 5390 13600 5410
rect 13702 5390 13722 5410
rect 13798 5390 13818 5410
rect 13908 5390 13928 5410
rect 14004 5390 14024 5410
rect 11896 5313 11916 5333
rect 9918 5193 9938 5213
rect 3953 5104 3973 5124
rect 7797 5117 7817 5137
rect 7893 5117 7913 5137
rect 8003 5117 8023 5137
rect 8099 5117 8119 5137
rect 8221 5117 8241 5137
rect 10014 5193 10034 5213
rect 10136 5193 10156 5213
rect 10232 5193 10252 5213
rect 10342 5193 10362 5213
rect 10438 5193 10458 5213
rect 15740 5326 15760 5346
rect 15836 5326 15856 5346
rect 15946 5326 15966 5346
rect 16042 5326 16062 5346
rect 16164 5326 16184 5346
rect 16260 5326 16280 5346
rect 14282 5206 14302 5226
rect 8317 5117 8337 5137
rect 380 4940 400 4960
rect 476 4940 496 4960
rect 598 4940 618 4960
rect 694 4940 714 4960
rect 804 4940 824 4960
rect 900 4940 920 4960
rect 12174 5129 12194 5149
rect 12270 5129 12290 5149
rect 12380 5129 12400 5149
rect 12476 5129 12496 5149
rect 12598 5129 12618 5149
rect 14378 5206 14398 5226
rect 14500 5206 14520 5226
rect 14596 5206 14616 5226
rect 14706 5206 14726 5226
rect 14802 5206 14822 5226
rect 12694 5129 12714 5149
rect 2331 4882 2351 4902
rect 2427 4882 2447 4902
rect 2537 4882 2557 4902
rect 2633 4882 2653 4902
rect 2755 4882 2775 4902
rect 4744 4953 4764 4973
rect 2851 4882 2871 4902
rect 4840 4953 4860 4973
rect 4962 4953 4982 4973
rect 5058 4953 5078 4973
rect 5168 4953 5188 4973
rect 5264 4953 5284 4973
rect 16538 5142 16558 5162
rect 16634 5142 16654 5162
rect 16744 5142 16764 5162
rect 16840 5142 16860 5162
rect 16962 5142 16982 5162
rect 17058 5142 17078 5162
rect 6695 4895 6715 4915
rect 6791 4895 6811 4915
rect 6901 4895 6921 4915
rect 6997 4895 7017 4915
rect 7119 4895 7139 4915
rect 9121 4965 9141 4985
rect 7215 4895 7235 4915
rect 9217 4965 9237 4985
rect 9339 4965 9359 4985
rect 9435 4965 9455 4985
rect 9545 4965 9565 4985
rect 9641 4965 9661 4985
rect 11072 4907 11092 4927
rect 11168 4907 11188 4927
rect 11278 4907 11298 4927
rect 11374 4907 11394 4927
rect 11496 4907 11516 4927
rect 13485 4978 13505 4998
rect 11592 4907 11612 4927
rect 13581 4978 13601 4998
rect 13703 4978 13723 4998
rect 13799 4978 13819 4998
rect 13909 4978 13929 4998
rect 14005 4978 14025 4998
rect 15436 4920 15456 4940
rect 15532 4920 15552 4940
rect 15642 4920 15662 4940
rect 15738 4920 15758 4940
rect 15860 4920 15880 4940
rect 15956 4920 15976 4940
rect 1462 4556 1482 4576
rect 1558 4556 1578 4576
rect 1680 4556 1700 4576
rect 1776 4556 1796 4576
rect 1886 4556 1906 4576
rect 1982 4556 2002 4576
rect 3413 4498 3433 4518
rect 3509 4498 3529 4518
rect 3619 4498 3639 4518
rect 3715 4498 3735 4518
rect 3837 4498 3857 4518
rect 5826 4569 5846 4589
rect 3933 4498 3953 4518
rect 5922 4569 5942 4589
rect 6044 4569 6064 4589
rect 6140 4569 6160 4589
rect 6250 4569 6270 4589
rect 6346 4569 6366 4589
rect 7777 4511 7797 4531
rect 7873 4511 7893 4531
rect 7983 4511 8003 4531
rect 8079 4511 8099 4531
rect 8201 4511 8221 4531
rect 10203 4581 10223 4601
rect 8297 4511 8317 4531
rect 10299 4581 10319 4601
rect 10421 4581 10441 4601
rect 10517 4581 10537 4601
rect 10627 4581 10647 4601
rect 10723 4581 10743 4601
rect 360 4334 380 4354
rect 456 4334 476 4354
rect 578 4334 598 4354
rect 674 4334 694 4354
rect 784 4334 804 4354
rect 880 4334 900 4354
rect 12154 4523 12174 4543
rect 12250 4523 12270 4543
rect 12360 4523 12380 4543
rect 12456 4523 12476 4543
rect 12578 4523 12598 4543
rect 14567 4594 14587 4614
rect 12674 4523 12694 4543
rect 14663 4594 14683 4614
rect 14785 4594 14805 4614
rect 14881 4594 14901 4614
rect 14991 4594 15011 4614
rect 15087 4594 15107 4614
rect 4724 4347 4744 4367
rect 2616 4270 2636 4290
rect 2712 4270 2732 4290
rect 2822 4270 2842 4290
rect 2918 4270 2938 4290
rect 3040 4270 3060 4290
rect 4820 4347 4840 4367
rect 4942 4347 4962 4367
rect 5038 4347 5058 4367
rect 5148 4347 5168 4367
rect 5244 4347 5264 4367
rect 16518 4536 16538 4556
rect 16614 4536 16634 4556
rect 16724 4536 16744 4556
rect 16820 4536 16840 4556
rect 16942 4536 16962 4556
rect 17038 4536 17058 4556
rect 9101 4359 9121 4379
rect 3136 4270 3156 4290
rect 1158 4150 1178 4170
rect 1254 4150 1274 4170
rect 1376 4150 1396 4170
rect 1472 4150 1492 4170
rect 1582 4150 1602 4170
rect 1678 4150 1698 4170
rect 6980 4283 7000 4303
rect 7076 4283 7096 4303
rect 7186 4283 7206 4303
rect 7282 4283 7302 4303
rect 7404 4283 7424 4303
rect 9197 4359 9217 4379
rect 9319 4359 9339 4379
rect 9415 4359 9435 4379
rect 9525 4359 9545 4379
rect 9621 4359 9641 4379
rect 13465 4372 13485 4392
rect 7500 4283 7520 4303
rect 5522 4163 5542 4183
rect 3414 4086 3434 4106
rect 3510 4086 3530 4106
rect 3620 4086 3640 4106
rect 3716 4086 3736 4106
rect 3838 4086 3858 4106
rect 5618 4163 5638 4183
rect 5740 4163 5760 4183
rect 5836 4163 5856 4183
rect 5946 4163 5966 4183
rect 6042 4163 6062 4183
rect 11357 4295 11377 4315
rect 11453 4295 11473 4315
rect 11563 4295 11583 4315
rect 11659 4295 11679 4315
rect 11781 4295 11801 4315
rect 13561 4372 13581 4392
rect 13683 4372 13703 4392
rect 13779 4372 13799 4392
rect 13889 4372 13909 4392
rect 13985 4372 14005 4392
rect 11877 4295 11897 4315
rect 9899 4175 9919 4195
rect 3934 4086 3954 4106
rect 7778 4099 7798 4119
rect 7874 4099 7894 4119
rect 7984 4099 8004 4119
rect 8080 4099 8100 4119
rect 8202 4099 8222 4119
rect 9995 4175 10015 4195
rect 10117 4175 10137 4195
rect 10213 4175 10233 4195
rect 10323 4175 10343 4195
rect 10419 4175 10439 4195
rect 15721 4308 15741 4328
rect 15817 4308 15837 4328
rect 15927 4308 15947 4328
rect 16023 4308 16043 4328
rect 16145 4308 16165 4328
rect 16241 4308 16261 4328
rect 14263 4188 14283 4208
rect 8298 4099 8318 4119
rect 361 3922 381 3942
rect 457 3922 477 3942
rect 579 3922 599 3942
rect 675 3922 695 3942
rect 785 3922 805 3942
rect 881 3922 901 3942
rect 12155 4111 12175 4131
rect 12251 4111 12271 4131
rect 12361 4111 12381 4131
rect 12457 4111 12477 4131
rect 12579 4111 12599 4131
rect 14359 4188 14379 4208
rect 14481 4188 14501 4208
rect 14577 4188 14597 4208
rect 14687 4188 14707 4208
rect 14783 4188 14803 4208
rect 12675 4111 12695 4131
rect 2517 3860 2537 3880
rect 2613 3860 2633 3880
rect 2723 3860 2743 3880
rect 2819 3860 2839 3880
rect 2941 3860 2961 3880
rect 4725 3935 4745 3955
rect 3037 3860 3057 3880
rect 4821 3935 4841 3955
rect 4943 3935 4963 3955
rect 5039 3935 5059 3955
rect 5149 3935 5169 3955
rect 5245 3935 5265 3955
rect 16519 4124 16539 4144
rect 16615 4124 16635 4144
rect 16725 4124 16745 4144
rect 16821 4124 16841 4144
rect 16943 4124 16963 4144
rect 17039 4124 17059 4144
rect 6881 3873 6901 3893
rect 6977 3873 6997 3893
rect 7087 3873 7107 3893
rect 7183 3873 7203 3893
rect 7305 3873 7325 3893
rect 9102 3947 9122 3967
rect 7401 3873 7421 3893
rect 9198 3947 9218 3967
rect 9320 3947 9340 3967
rect 9416 3947 9436 3967
rect 9526 3947 9546 3967
rect 9622 3947 9642 3967
rect 11258 3885 11278 3905
rect 11354 3885 11374 3905
rect 11464 3885 11484 3905
rect 11560 3885 11580 3905
rect 11682 3885 11702 3905
rect 13466 3960 13486 3980
rect 11778 3885 11798 3905
rect 13562 3960 13582 3980
rect 13684 3960 13704 3980
rect 13780 3960 13800 3980
rect 13890 3960 13910 3980
rect 13986 3960 14006 3980
rect 15622 3898 15642 3918
rect 15718 3898 15738 3918
rect 15828 3898 15848 3918
rect 15924 3898 15944 3918
rect 16046 3898 16066 3918
rect 16142 3898 16162 3918
rect 1240 3542 1260 3562
rect 1336 3542 1356 3562
rect 1458 3542 1478 3562
rect 1554 3542 1574 3562
rect 1664 3542 1684 3562
rect 1760 3542 1780 3562
rect 3396 3480 3416 3500
rect 3492 3480 3512 3500
rect 3602 3480 3622 3500
rect 3698 3480 3718 3500
rect 3820 3480 3840 3500
rect 5604 3555 5624 3575
rect 3916 3480 3936 3500
rect 5700 3555 5720 3575
rect 5822 3555 5842 3575
rect 5918 3555 5938 3575
rect 6028 3555 6048 3575
rect 6124 3555 6144 3575
rect 7760 3493 7780 3513
rect 7856 3493 7876 3513
rect 7966 3493 7986 3513
rect 8062 3493 8082 3513
rect 8184 3493 8204 3513
rect 9981 3567 10001 3587
rect 8280 3493 8300 3513
rect 10077 3567 10097 3587
rect 10199 3567 10219 3587
rect 10295 3567 10315 3587
rect 10405 3567 10425 3587
rect 10501 3567 10521 3587
rect 343 3316 363 3336
rect 439 3316 459 3336
rect 561 3316 581 3336
rect 657 3316 677 3336
rect 767 3316 787 3336
rect 863 3316 883 3336
rect 12137 3505 12157 3525
rect 12233 3505 12253 3525
rect 12343 3505 12363 3525
rect 12439 3505 12459 3525
rect 12561 3505 12581 3525
rect 14345 3580 14365 3600
rect 12657 3505 12677 3525
rect 14441 3580 14461 3600
rect 14563 3580 14583 3600
rect 14659 3580 14679 3600
rect 14769 3580 14789 3600
rect 14865 3580 14885 3600
rect 4707 3329 4727 3349
rect 2599 3252 2619 3272
rect 2695 3252 2715 3272
rect 2805 3252 2825 3272
rect 2901 3252 2921 3272
rect 3023 3252 3043 3272
rect 4803 3329 4823 3349
rect 4925 3329 4945 3349
rect 5021 3329 5041 3349
rect 5131 3329 5151 3349
rect 5227 3329 5247 3349
rect 16501 3518 16521 3538
rect 16597 3518 16617 3538
rect 16707 3518 16727 3538
rect 16803 3518 16823 3538
rect 16925 3518 16945 3538
rect 17021 3518 17041 3538
rect 9084 3341 9104 3361
rect 3119 3252 3139 3272
rect 1141 3132 1161 3152
rect 1237 3132 1257 3152
rect 1359 3132 1379 3152
rect 1455 3132 1475 3152
rect 1565 3132 1585 3152
rect 1661 3132 1681 3152
rect 6963 3265 6983 3285
rect 7059 3265 7079 3285
rect 7169 3265 7189 3285
rect 7265 3265 7285 3285
rect 7387 3265 7407 3285
rect 9180 3341 9200 3361
rect 9302 3341 9322 3361
rect 9398 3341 9418 3361
rect 9508 3341 9528 3361
rect 9604 3341 9624 3361
rect 13448 3354 13468 3374
rect 7483 3265 7503 3285
rect 5505 3145 5525 3165
rect 3397 3068 3417 3088
rect 3493 3068 3513 3088
rect 3603 3068 3623 3088
rect 3699 3068 3719 3088
rect 3821 3068 3841 3088
rect 5601 3145 5621 3165
rect 5723 3145 5743 3165
rect 5819 3145 5839 3165
rect 5929 3145 5949 3165
rect 6025 3145 6045 3165
rect 11340 3277 11360 3297
rect 11436 3277 11456 3297
rect 11546 3277 11566 3297
rect 11642 3277 11662 3297
rect 11764 3277 11784 3297
rect 13544 3354 13564 3374
rect 13666 3354 13686 3374
rect 13762 3354 13782 3374
rect 13872 3354 13892 3374
rect 13968 3354 13988 3374
rect 11860 3277 11880 3297
rect 9882 3157 9902 3177
rect 3917 3068 3937 3088
rect 7761 3081 7781 3101
rect 7857 3081 7877 3101
rect 7967 3081 7987 3101
rect 8063 3081 8083 3101
rect 8185 3081 8205 3101
rect 9978 3157 9998 3177
rect 10100 3157 10120 3177
rect 10196 3157 10216 3177
rect 10306 3157 10326 3177
rect 10402 3157 10422 3177
rect 15704 3290 15724 3310
rect 15800 3290 15820 3310
rect 15910 3290 15930 3310
rect 16006 3290 16026 3310
rect 16128 3290 16148 3310
rect 16224 3290 16244 3310
rect 14246 3170 14266 3190
rect 8281 3081 8301 3101
rect 344 2904 364 2924
rect 440 2904 460 2924
rect 562 2904 582 2924
rect 658 2904 678 2924
rect 768 2904 788 2924
rect 864 2904 884 2924
rect 12138 3093 12158 3113
rect 12234 3093 12254 3113
rect 12344 3093 12364 3113
rect 12440 3093 12460 3113
rect 12562 3093 12582 3113
rect 14342 3170 14362 3190
rect 14464 3170 14484 3190
rect 14560 3170 14580 3190
rect 14670 3170 14690 3190
rect 14766 3170 14786 3190
rect 12658 3093 12678 3113
rect 2434 2844 2454 2864
rect 2530 2844 2550 2864
rect 2640 2844 2660 2864
rect 2736 2844 2756 2864
rect 2858 2844 2878 2864
rect 4708 2917 4728 2937
rect 2954 2844 2974 2864
rect 4804 2917 4824 2937
rect 4926 2917 4946 2937
rect 5022 2917 5042 2937
rect 5132 2917 5152 2937
rect 5228 2917 5248 2937
rect 16502 3106 16522 3126
rect 16598 3106 16618 3126
rect 16708 3106 16728 3126
rect 16804 3106 16824 3126
rect 16926 3106 16946 3126
rect 17022 3106 17042 3126
rect 6798 2857 6818 2877
rect 6894 2857 6914 2877
rect 7004 2857 7024 2877
rect 7100 2857 7120 2877
rect 7222 2857 7242 2877
rect 9085 2929 9105 2949
rect 7318 2857 7338 2877
rect 9181 2929 9201 2949
rect 9303 2929 9323 2949
rect 9399 2929 9419 2949
rect 9509 2929 9529 2949
rect 9605 2929 9625 2949
rect 11175 2869 11195 2889
rect 11271 2869 11291 2889
rect 11381 2869 11401 2889
rect 11477 2869 11497 2889
rect 11599 2869 11619 2889
rect 13449 2942 13469 2962
rect 11695 2869 11715 2889
rect 13545 2942 13565 2962
rect 13667 2942 13687 2962
rect 13763 2942 13783 2962
rect 13873 2942 13893 2962
rect 13969 2942 13989 2962
rect 15539 2882 15559 2902
rect 15635 2882 15655 2902
rect 15745 2882 15765 2902
rect 15841 2882 15861 2902
rect 15963 2882 15983 2902
rect 16059 2882 16079 2902
rect 1286 2522 1306 2542
rect 1382 2522 1402 2542
rect 1504 2522 1524 2542
rect 1600 2522 1620 2542
rect 1710 2522 1730 2542
rect 1806 2522 1826 2542
rect 3376 2462 3396 2482
rect 3472 2462 3492 2482
rect 3582 2462 3602 2482
rect 3678 2462 3698 2482
rect 3800 2462 3820 2482
rect 5650 2535 5670 2555
rect 3896 2462 3916 2482
rect 5746 2535 5766 2555
rect 5868 2535 5888 2555
rect 5964 2535 5984 2555
rect 6074 2535 6094 2555
rect 6170 2535 6190 2555
rect 7740 2475 7760 2495
rect 7836 2475 7856 2495
rect 7946 2475 7966 2495
rect 8042 2475 8062 2495
rect 8164 2475 8184 2495
rect 10027 2547 10047 2567
rect 8260 2475 8280 2495
rect 10123 2547 10143 2567
rect 10245 2547 10265 2567
rect 10341 2547 10361 2567
rect 10451 2547 10471 2567
rect 10547 2547 10567 2567
rect 323 2298 343 2318
rect 419 2298 439 2318
rect 541 2298 561 2318
rect 637 2298 657 2318
rect 747 2298 767 2318
rect 843 2298 863 2318
rect 12117 2487 12137 2507
rect 12213 2487 12233 2507
rect 12323 2487 12343 2507
rect 12419 2487 12439 2507
rect 12541 2487 12561 2507
rect 14391 2560 14411 2580
rect 12637 2487 12657 2507
rect 14487 2560 14507 2580
rect 14609 2560 14629 2580
rect 14705 2560 14725 2580
rect 14815 2560 14835 2580
rect 14911 2560 14931 2580
rect 4687 2311 4707 2331
rect 2579 2234 2599 2254
rect 2675 2234 2695 2254
rect 2785 2234 2805 2254
rect 2881 2234 2901 2254
rect 3003 2234 3023 2254
rect 4783 2311 4803 2331
rect 4905 2311 4925 2331
rect 5001 2311 5021 2331
rect 5111 2311 5131 2331
rect 5207 2311 5227 2331
rect 16481 2500 16501 2520
rect 16577 2500 16597 2520
rect 16687 2500 16707 2520
rect 16783 2500 16803 2520
rect 16905 2500 16925 2520
rect 17001 2500 17021 2520
rect 9064 2323 9084 2343
rect 3099 2234 3119 2254
rect 1121 2114 1141 2134
rect 1217 2114 1237 2134
rect 1339 2114 1359 2134
rect 1435 2114 1455 2134
rect 1545 2114 1565 2134
rect 1641 2114 1661 2134
rect 6943 2247 6963 2267
rect 7039 2247 7059 2267
rect 7149 2247 7169 2267
rect 7245 2247 7265 2267
rect 7367 2247 7387 2267
rect 9160 2323 9180 2343
rect 9282 2323 9302 2343
rect 9378 2323 9398 2343
rect 9488 2323 9508 2343
rect 9584 2323 9604 2343
rect 13428 2336 13448 2356
rect 7463 2247 7483 2267
rect 5485 2127 5505 2147
rect 3377 2050 3397 2070
rect 3473 2050 3493 2070
rect 3583 2050 3603 2070
rect 3679 2050 3699 2070
rect 3801 2050 3821 2070
rect 5581 2127 5601 2147
rect 5703 2127 5723 2147
rect 5799 2127 5819 2147
rect 5909 2127 5929 2147
rect 6005 2127 6025 2147
rect 11320 2259 11340 2279
rect 11416 2259 11436 2279
rect 11526 2259 11546 2279
rect 11622 2259 11642 2279
rect 11744 2259 11764 2279
rect 13524 2336 13544 2356
rect 13646 2336 13666 2356
rect 13742 2336 13762 2356
rect 13852 2336 13872 2356
rect 13948 2336 13968 2356
rect 11840 2259 11860 2279
rect 9862 2139 9882 2159
rect 3897 2050 3917 2070
rect 7741 2063 7761 2083
rect 7837 2063 7857 2083
rect 7947 2063 7967 2083
rect 8043 2063 8063 2083
rect 8165 2063 8185 2083
rect 9958 2139 9978 2159
rect 10080 2139 10100 2159
rect 10176 2139 10196 2159
rect 10286 2139 10306 2159
rect 10382 2139 10402 2159
rect 15684 2272 15704 2292
rect 15780 2272 15800 2292
rect 15890 2272 15910 2292
rect 15986 2272 16006 2292
rect 16108 2272 16128 2292
rect 16204 2272 16224 2292
rect 14226 2152 14246 2172
rect 8261 2063 8281 2083
rect 324 1886 344 1906
rect 420 1886 440 1906
rect 542 1886 562 1906
rect 638 1886 658 1906
rect 748 1886 768 1906
rect 844 1886 864 1906
rect 12118 2075 12138 2095
rect 12214 2075 12234 2095
rect 12324 2075 12344 2095
rect 12420 2075 12440 2095
rect 12542 2075 12562 2095
rect 14322 2152 14342 2172
rect 14444 2152 14464 2172
rect 14540 2152 14560 2172
rect 14650 2152 14670 2172
rect 14746 2152 14766 2172
rect 12638 2075 12658 2095
rect 2480 1824 2500 1844
rect 2576 1824 2596 1844
rect 2686 1824 2706 1844
rect 2782 1824 2802 1844
rect 2904 1824 2924 1844
rect 4688 1899 4708 1919
rect 3000 1824 3020 1844
rect 4784 1899 4804 1919
rect 4906 1899 4926 1919
rect 5002 1899 5022 1919
rect 5112 1899 5132 1919
rect 5208 1899 5228 1919
rect 16482 2088 16502 2108
rect 16578 2088 16598 2108
rect 16688 2088 16708 2108
rect 16784 2088 16804 2108
rect 16906 2088 16926 2108
rect 17002 2088 17022 2108
rect 6844 1837 6864 1857
rect 6940 1837 6960 1857
rect 7050 1837 7070 1857
rect 7146 1837 7166 1857
rect 7268 1837 7288 1857
rect 9065 1911 9085 1931
rect 7364 1837 7384 1857
rect 9161 1911 9181 1931
rect 9283 1911 9303 1931
rect 9379 1911 9399 1931
rect 9489 1911 9509 1931
rect 9585 1911 9605 1931
rect 11221 1849 11241 1869
rect 11317 1849 11337 1869
rect 11427 1849 11447 1869
rect 11523 1849 11543 1869
rect 11645 1849 11665 1869
rect 13429 1924 13449 1944
rect 11741 1849 11761 1869
rect 13525 1924 13545 1944
rect 13647 1924 13667 1944
rect 13743 1924 13763 1944
rect 13853 1924 13873 1944
rect 13949 1924 13969 1944
rect 15585 1862 15605 1882
rect 15681 1862 15701 1882
rect 15791 1862 15811 1882
rect 15887 1862 15907 1882
rect 16009 1862 16029 1882
rect 16105 1862 16125 1882
rect 1203 1506 1223 1526
rect 1299 1506 1319 1526
rect 1421 1506 1441 1526
rect 1517 1506 1537 1526
rect 1627 1506 1647 1526
rect 1723 1506 1743 1526
rect 3359 1444 3379 1464
rect 3455 1444 3475 1464
rect 3565 1444 3585 1464
rect 3661 1444 3681 1464
rect 3783 1444 3803 1464
rect 5567 1519 5587 1539
rect 3879 1444 3899 1464
rect 5663 1519 5683 1539
rect 5785 1519 5805 1539
rect 5881 1519 5901 1539
rect 5991 1519 6011 1539
rect 6087 1519 6107 1539
rect 7723 1457 7743 1477
rect 7819 1457 7839 1477
rect 7929 1457 7949 1477
rect 8025 1457 8045 1477
rect 8147 1457 8167 1477
rect 9944 1531 9964 1551
rect 8243 1457 8263 1477
rect 10040 1531 10060 1551
rect 10162 1531 10182 1551
rect 10258 1531 10278 1551
rect 10368 1531 10388 1551
rect 10464 1531 10484 1551
rect 306 1280 326 1300
rect 402 1280 422 1300
rect 524 1280 544 1300
rect 620 1280 640 1300
rect 730 1280 750 1300
rect 826 1280 846 1300
rect 12100 1469 12120 1489
rect 12196 1469 12216 1489
rect 12306 1469 12326 1489
rect 12402 1469 12422 1489
rect 12524 1469 12544 1489
rect 14308 1544 14328 1564
rect 12620 1469 12640 1489
rect 14404 1544 14424 1564
rect 14526 1544 14546 1564
rect 14622 1544 14642 1564
rect 14732 1544 14752 1564
rect 14828 1544 14848 1564
rect 4670 1293 4690 1313
rect 2562 1216 2582 1236
rect 2658 1216 2678 1236
rect 2768 1216 2788 1236
rect 2864 1216 2884 1236
rect 2986 1216 3006 1236
rect 4766 1293 4786 1313
rect 4888 1293 4908 1313
rect 4984 1293 5004 1313
rect 5094 1293 5114 1313
rect 5190 1293 5210 1313
rect 16464 1482 16484 1502
rect 16560 1482 16580 1502
rect 16670 1482 16690 1502
rect 16766 1482 16786 1502
rect 16888 1482 16908 1502
rect 16984 1482 17004 1502
rect 9047 1305 9067 1325
rect 3082 1216 3102 1236
rect 1104 1096 1124 1116
rect 1200 1096 1220 1116
rect 1322 1096 1342 1116
rect 1418 1096 1438 1116
rect 1528 1096 1548 1116
rect 1624 1096 1644 1116
rect 6926 1229 6946 1249
rect 7022 1229 7042 1249
rect 7132 1229 7152 1249
rect 7228 1229 7248 1249
rect 7350 1229 7370 1249
rect 9143 1305 9163 1325
rect 9265 1305 9285 1325
rect 9361 1305 9381 1325
rect 9471 1305 9491 1325
rect 9567 1305 9587 1325
rect 13411 1318 13431 1338
rect 7446 1229 7466 1249
rect 5468 1109 5488 1129
rect 3360 1032 3380 1052
rect 3456 1032 3476 1052
rect 3566 1032 3586 1052
rect 3662 1032 3682 1052
rect 3784 1032 3804 1052
rect 5564 1109 5584 1129
rect 5686 1109 5706 1129
rect 5782 1109 5802 1129
rect 5892 1109 5912 1129
rect 5988 1109 6008 1129
rect 11303 1241 11323 1261
rect 11399 1241 11419 1261
rect 11509 1241 11529 1261
rect 11605 1241 11625 1261
rect 11727 1241 11747 1261
rect 13507 1318 13527 1338
rect 13629 1318 13649 1338
rect 13725 1318 13745 1338
rect 13835 1318 13855 1338
rect 13931 1318 13951 1338
rect 11823 1241 11843 1261
rect 9845 1121 9865 1141
rect 3880 1032 3900 1052
rect 7724 1045 7744 1065
rect 7820 1045 7840 1065
rect 7930 1045 7950 1065
rect 8026 1045 8046 1065
rect 8148 1045 8168 1065
rect 9941 1121 9961 1141
rect 10063 1121 10083 1141
rect 10159 1121 10179 1141
rect 10269 1121 10289 1141
rect 10365 1121 10385 1141
rect 15667 1254 15687 1274
rect 15763 1254 15783 1274
rect 15873 1254 15893 1274
rect 15969 1254 15989 1274
rect 16091 1254 16111 1274
rect 16187 1254 16207 1274
rect 14209 1134 14229 1154
rect 8244 1045 8264 1065
rect 12101 1057 12121 1077
rect 12197 1057 12217 1077
rect 12307 1057 12327 1077
rect 12403 1057 12423 1077
rect 12525 1057 12545 1077
rect 14305 1134 14325 1154
rect 14427 1134 14447 1154
rect 14523 1134 14543 1154
rect 14633 1134 14653 1154
rect 14729 1134 14749 1154
rect 12621 1057 12641 1077
rect 16465 1070 16485 1090
rect 16561 1070 16581 1090
rect 16671 1070 16691 1090
rect 16767 1070 16787 1090
rect 16889 1070 16909 1090
rect 16985 1070 17005 1090
rect 307 868 327 888
rect 403 868 423 888
rect 525 868 545 888
rect 621 868 641 888
rect 731 868 751 888
rect 827 868 847 888
rect 4671 881 4691 901
rect 4767 881 4787 901
rect 4889 881 4909 901
rect 4985 881 5005 901
rect 5095 881 5115 901
rect 5191 881 5211 901
rect 9048 893 9068 913
rect 9144 893 9164 913
rect 9266 893 9286 913
rect 9362 893 9382 913
rect 9472 893 9492 913
rect 9568 893 9588 913
rect 13412 906 13432 926
rect 13508 906 13528 926
rect 13630 906 13650 926
rect 13726 906 13746 926
rect 13836 906 13856 926
rect 13932 906 13952 926
rect 1520 292 1540 312
rect 1616 292 1636 312
rect 1738 292 1758 312
rect 1834 292 1854 312
rect 1944 292 1964 312
rect 2040 292 2060 312
rect 5884 305 5904 325
rect 4009 218 4029 238
rect 4105 218 4125 238
rect 4227 218 4247 238
rect 4323 218 4343 238
rect 4433 218 4453 238
rect 5980 305 6000 325
rect 6102 305 6122 325
rect 6198 305 6218 325
rect 6308 305 6328 325
rect 6404 305 6424 325
rect 10261 317 10281 337
rect 4529 218 4549 238
rect 8457 242 8477 262
rect 8553 242 8573 262
rect 8675 242 8695 262
rect 8771 242 8791 262
rect 8881 242 8901 262
rect 10357 317 10377 337
rect 10479 317 10499 337
rect 10575 317 10595 337
rect 10685 317 10705 337
rect 10781 317 10801 337
rect 14625 330 14645 350
rect 8977 242 8997 262
rect 12750 243 12770 263
rect 12846 243 12866 263
rect 12968 243 12988 263
rect 13064 243 13084 263
rect 13174 243 13194 263
rect 14721 330 14741 350
rect 14843 330 14863 350
rect 14939 330 14959 350
rect 15049 330 15069 350
rect 15145 330 15165 350
rect 13270 243 13290 263
<< poly >>
rect 3518 8751 3568 8767
rect 3726 8751 3776 8767
rect 3944 8751 3994 8767
rect 7882 8764 7932 8780
rect 8090 8764 8140 8780
rect 8308 8764 8358 8780
rect 12259 8776 12309 8792
rect 12467 8776 12517 8792
rect 12685 8776 12735 8792
rect 16623 8789 16673 8805
rect 16831 8789 16881 8805
rect 17049 8789 17099 8805
rect 3518 8679 3568 8709
rect 3518 8659 3525 8679
rect 3545 8659 3568 8679
rect 3518 8632 3568 8659
rect 3726 8677 3776 8709
rect 3726 8657 3743 8677
rect 3763 8657 3776 8677
rect 3726 8632 3776 8657
rect 3944 8680 3994 8709
rect 3944 8660 3961 8680
rect 3981 8660 3994 8680
rect 3944 8632 3994 8660
rect 7882 8692 7932 8722
rect 7882 8672 7889 8692
rect 7909 8672 7932 8692
rect 2721 8523 2771 8539
rect 2929 8523 2979 8539
rect 3147 8523 3197 8539
rect 7882 8645 7932 8672
rect 8090 8690 8140 8722
rect 8090 8670 8107 8690
rect 8127 8670 8140 8690
rect 8090 8645 8140 8670
rect 8308 8693 8358 8722
rect 8308 8673 8325 8693
rect 8345 8673 8358 8693
rect 8308 8645 8358 8673
rect 12259 8704 12309 8734
rect 12259 8684 12266 8704
rect 12286 8684 12309 8704
rect 3518 8519 3568 8532
rect 3726 8519 3776 8532
rect 3944 8519 3994 8532
rect 7085 8536 7135 8552
rect 7293 8536 7343 8552
rect 7511 8536 7561 8552
rect 12259 8657 12309 8684
rect 12467 8702 12517 8734
rect 12467 8682 12484 8702
rect 12504 8682 12517 8702
rect 12467 8657 12517 8682
rect 12685 8705 12735 8734
rect 12685 8685 12702 8705
rect 12722 8685 12735 8705
rect 12685 8657 12735 8685
rect 16623 8717 16673 8747
rect 16623 8697 16630 8717
rect 16650 8697 16673 8717
rect 7882 8532 7932 8545
rect 8090 8532 8140 8545
rect 8308 8532 8358 8545
rect 11462 8548 11512 8564
rect 11670 8548 11720 8564
rect 11888 8548 11938 8564
rect 16623 8670 16673 8697
rect 16831 8715 16881 8747
rect 16831 8695 16848 8715
rect 16868 8695 16881 8715
rect 16831 8670 16881 8695
rect 17049 8718 17099 8747
rect 17049 8698 17066 8718
rect 17086 8698 17099 8718
rect 17049 8670 17099 8698
rect 12259 8544 12309 8557
rect 12467 8544 12517 8557
rect 12685 8544 12735 8557
rect 15826 8561 15876 8577
rect 16034 8561 16084 8577
rect 16252 8561 16302 8577
rect 16623 8557 16673 8570
rect 16831 8557 16881 8570
rect 17049 8557 17099 8570
rect 465 8464 515 8477
rect 683 8464 733 8477
rect 891 8464 941 8477
rect 2721 8451 2771 8481
rect 2721 8431 2728 8451
rect 2748 8431 2771 8451
rect 2721 8404 2771 8431
rect 2929 8449 2979 8481
rect 2929 8429 2946 8449
rect 2966 8429 2979 8449
rect 2929 8404 2979 8429
rect 3147 8452 3197 8481
rect 3147 8432 3164 8452
rect 3184 8432 3197 8452
rect 4829 8477 4879 8490
rect 5047 8477 5097 8490
rect 5255 8477 5305 8490
rect 3147 8404 3197 8432
rect 465 8336 515 8364
rect 465 8316 478 8336
rect 498 8316 515 8336
rect 465 8287 515 8316
rect 683 8339 733 8364
rect 683 8319 696 8339
rect 716 8319 733 8339
rect 683 8287 733 8319
rect 891 8337 941 8364
rect 891 8317 914 8337
rect 934 8317 941 8337
rect 891 8287 941 8317
rect 7085 8464 7135 8494
rect 7085 8444 7092 8464
rect 7112 8444 7135 8464
rect 7085 8417 7135 8444
rect 7293 8462 7343 8494
rect 7293 8442 7310 8462
rect 7330 8442 7343 8462
rect 7293 8417 7343 8442
rect 7511 8465 7561 8494
rect 7511 8445 7528 8465
rect 7548 8445 7561 8465
rect 9206 8489 9256 8502
rect 9424 8489 9474 8502
rect 9632 8489 9682 8502
rect 7511 8417 7561 8445
rect 3519 8339 3569 8355
rect 3727 8339 3777 8355
rect 3945 8339 3995 8355
rect 1263 8280 1313 8293
rect 1481 8280 1531 8293
rect 1689 8280 1739 8293
rect 2721 8291 2771 8304
rect 2929 8291 2979 8304
rect 3147 8291 3197 8304
rect 4829 8349 4879 8377
rect 465 8229 515 8245
rect 683 8229 733 8245
rect 891 8229 941 8245
rect 3519 8267 3569 8297
rect 3519 8247 3526 8267
rect 3546 8247 3569 8267
rect 3519 8220 3569 8247
rect 3727 8265 3777 8297
rect 3727 8245 3744 8265
rect 3764 8245 3777 8265
rect 3727 8220 3777 8245
rect 3945 8268 3995 8297
rect 3945 8248 3962 8268
rect 3982 8248 3995 8268
rect 4829 8329 4842 8349
rect 4862 8329 4879 8349
rect 4829 8300 4879 8329
rect 5047 8352 5097 8377
rect 5047 8332 5060 8352
rect 5080 8332 5097 8352
rect 5047 8300 5097 8332
rect 5255 8350 5305 8377
rect 5255 8330 5278 8350
rect 5298 8330 5305 8350
rect 5255 8300 5305 8330
rect 11462 8476 11512 8506
rect 11462 8456 11469 8476
rect 11489 8456 11512 8476
rect 11462 8429 11512 8456
rect 11670 8474 11720 8506
rect 11670 8454 11687 8474
rect 11707 8454 11720 8474
rect 11670 8429 11720 8454
rect 11888 8477 11938 8506
rect 11888 8457 11905 8477
rect 11925 8457 11938 8477
rect 13570 8502 13620 8515
rect 13788 8502 13838 8515
rect 13996 8502 14046 8515
rect 11888 8429 11938 8457
rect 7883 8352 7933 8368
rect 8091 8352 8141 8368
rect 8309 8352 8359 8368
rect 3945 8220 3995 8248
rect 5627 8293 5677 8306
rect 5845 8293 5895 8306
rect 6053 8293 6103 8306
rect 7085 8304 7135 8317
rect 7293 8304 7343 8317
rect 7511 8304 7561 8317
rect 9206 8361 9256 8389
rect 4829 8242 4879 8258
rect 5047 8242 5097 8258
rect 5255 8242 5305 8258
rect 1263 8152 1313 8180
rect 1263 8132 1276 8152
rect 1296 8132 1313 8152
rect 1263 8103 1313 8132
rect 1481 8155 1531 8180
rect 1481 8135 1494 8155
rect 1514 8135 1531 8155
rect 1481 8103 1531 8135
rect 1689 8153 1739 8180
rect 1689 8133 1712 8153
rect 1732 8133 1739 8153
rect 1689 8103 1739 8133
rect 2622 8113 2672 8129
rect 2830 8113 2880 8129
rect 3048 8113 3098 8129
rect 7883 8280 7933 8310
rect 7883 8260 7890 8280
rect 7910 8260 7933 8280
rect 7883 8233 7933 8260
rect 8091 8278 8141 8310
rect 8091 8258 8108 8278
rect 8128 8258 8141 8278
rect 8091 8233 8141 8258
rect 8309 8281 8359 8310
rect 8309 8261 8326 8281
rect 8346 8261 8359 8281
rect 9206 8341 9219 8361
rect 9239 8341 9256 8361
rect 9206 8312 9256 8341
rect 9424 8364 9474 8389
rect 9424 8344 9437 8364
rect 9457 8344 9474 8364
rect 9424 8312 9474 8344
rect 9632 8362 9682 8389
rect 9632 8342 9655 8362
rect 9675 8342 9682 8362
rect 9632 8312 9682 8342
rect 15826 8489 15876 8519
rect 15826 8469 15833 8489
rect 15853 8469 15876 8489
rect 15826 8442 15876 8469
rect 16034 8487 16084 8519
rect 16034 8467 16051 8487
rect 16071 8467 16084 8487
rect 16034 8442 16084 8467
rect 16252 8490 16302 8519
rect 16252 8470 16269 8490
rect 16289 8470 16302 8490
rect 16252 8442 16302 8470
rect 12260 8364 12310 8380
rect 12468 8364 12518 8380
rect 12686 8364 12736 8380
rect 8309 8233 8359 8261
rect 10004 8305 10054 8318
rect 10222 8305 10272 8318
rect 10430 8305 10480 8318
rect 11462 8316 11512 8329
rect 11670 8316 11720 8329
rect 11888 8316 11938 8329
rect 13570 8374 13620 8402
rect 9206 8254 9256 8270
rect 9424 8254 9474 8270
rect 9632 8254 9682 8270
rect 5627 8165 5677 8193
rect 466 8052 516 8065
rect 684 8052 734 8065
rect 892 8052 942 8065
rect 3519 8107 3569 8120
rect 3727 8107 3777 8120
rect 3945 8107 3995 8120
rect 5627 8145 5640 8165
rect 5660 8145 5677 8165
rect 5627 8116 5677 8145
rect 5845 8168 5895 8193
rect 5845 8148 5858 8168
rect 5878 8148 5895 8168
rect 5845 8116 5895 8148
rect 6053 8166 6103 8193
rect 6053 8146 6076 8166
rect 6096 8146 6103 8166
rect 6053 8116 6103 8146
rect 6986 8126 7036 8142
rect 7194 8126 7244 8142
rect 7412 8126 7462 8142
rect 12260 8292 12310 8322
rect 12260 8272 12267 8292
rect 12287 8272 12310 8292
rect 12260 8245 12310 8272
rect 12468 8290 12518 8322
rect 12468 8270 12485 8290
rect 12505 8270 12518 8290
rect 12468 8245 12518 8270
rect 12686 8293 12736 8322
rect 12686 8273 12703 8293
rect 12723 8273 12736 8293
rect 13570 8354 13583 8374
rect 13603 8354 13620 8374
rect 13570 8325 13620 8354
rect 13788 8377 13838 8402
rect 13788 8357 13801 8377
rect 13821 8357 13838 8377
rect 13788 8325 13838 8357
rect 13996 8375 14046 8402
rect 13996 8355 14019 8375
rect 14039 8355 14046 8375
rect 13996 8325 14046 8355
rect 16624 8377 16674 8393
rect 16832 8377 16882 8393
rect 17050 8377 17100 8393
rect 12686 8245 12736 8273
rect 14368 8318 14418 8331
rect 14586 8318 14636 8331
rect 14794 8318 14844 8331
rect 15826 8329 15876 8342
rect 16034 8329 16084 8342
rect 16252 8329 16302 8342
rect 13570 8267 13620 8283
rect 13788 8267 13838 8283
rect 13996 8267 14046 8283
rect 10004 8177 10054 8205
rect 1263 8045 1313 8061
rect 1481 8045 1531 8061
rect 1689 8045 1739 8061
rect 2622 8041 2672 8071
rect 2622 8021 2629 8041
rect 2649 8021 2672 8041
rect 2622 7994 2672 8021
rect 2830 8039 2880 8071
rect 2830 8019 2847 8039
rect 2867 8019 2880 8039
rect 2830 7994 2880 8019
rect 3048 8042 3098 8071
rect 4830 8065 4880 8078
rect 5048 8065 5098 8078
rect 5256 8065 5306 8078
rect 7883 8120 7933 8133
rect 8091 8120 8141 8133
rect 8309 8120 8359 8133
rect 10004 8157 10017 8177
rect 10037 8157 10054 8177
rect 10004 8128 10054 8157
rect 10222 8180 10272 8205
rect 10222 8160 10235 8180
rect 10255 8160 10272 8180
rect 10222 8128 10272 8160
rect 10430 8178 10480 8205
rect 10430 8158 10453 8178
rect 10473 8158 10480 8178
rect 10430 8128 10480 8158
rect 11363 8138 11413 8154
rect 11571 8138 11621 8154
rect 11789 8138 11839 8154
rect 16624 8305 16674 8335
rect 16624 8285 16631 8305
rect 16651 8285 16674 8305
rect 16624 8258 16674 8285
rect 16832 8303 16882 8335
rect 16832 8283 16849 8303
rect 16869 8283 16882 8303
rect 16832 8258 16882 8283
rect 17050 8306 17100 8335
rect 17050 8286 17067 8306
rect 17087 8286 17100 8306
rect 17050 8258 17100 8286
rect 14368 8190 14418 8218
rect 3048 8022 3065 8042
rect 3085 8022 3098 8042
rect 3048 7994 3098 8022
rect 466 7924 516 7952
rect 466 7904 479 7924
rect 499 7904 516 7924
rect 466 7875 516 7904
rect 684 7927 734 7952
rect 684 7907 697 7927
rect 717 7907 734 7927
rect 684 7875 734 7907
rect 892 7925 942 7952
rect 892 7905 915 7925
rect 935 7905 942 7925
rect 892 7875 942 7905
rect 5627 8058 5677 8074
rect 5845 8058 5895 8074
rect 6053 8058 6103 8074
rect 6986 8054 7036 8084
rect 6986 8034 6993 8054
rect 7013 8034 7036 8054
rect 6986 8007 7036 8034
rect 7194 8052 7244 8084
rect 7194 8032 7211 8052
rect 7231 8032 7244 8052
rect 7194 8007 7244 8032
rect 7412 8055 7462 8084
rect 9207 8077 9257 8090
rect 9425 8077 9475 8090
rect 9633 8077 9683 8090
rect 12260 8132 12310 8145
rect 12468 8132 12518 8145
rect 12686 8132 12736 8145
rect 14368 8170 14381 8190
rect 14401 8170 14418 8190
rect 14368 8141 14418 8170
rect 14586 8193 14636 8218
rect 14586 8173 14599 8193
rect 14619 8173 14636 8193
rect 14586 8141 14636 8173
rect 14794 8191 14844 8218
rect 14794 8171 14817 8191
rect 14837 8171 14844 8191
rect 14794 8141 14844 8171
rect 15727 8151 15777 8167
rect 15935 8151 15985 8167
rect 16153 8151 16203 8167
rect 7412 8035 7429 8055
rect 7449 8035 7462 8055
rect 7412 8007 7462 8035
rect 4830 7937 4880 7965
rect 2622 7881 2672 7894
rect 2830 7881 2880 7894
rect 3048 7881 3098 7894
rect 4830 7917 4843 7937
rect 4863 7917 4880 7937
rect 4830 7888 4880 7917
rect 5048 7940 5098 7965
rect 5048 7920 5061 7940
rect 5081 7920 5098 7940
rect 5048 7888 5098 7920
rect 5256 7938 5306 7965
rect 5256 7918 5279 7938
rect 5299 7918 5306 7938
rect 5256 7888 5306 7918
rect 10004 8070 10054 8086
rect 10222 8070 10272 8086
rect 10430 8070 10480 8086
rect 11363 8066 11413 8096
rect 11363 8046 11370 8066
rect 11390 8046 11413 8066
rect 11363 8019 11413 8046
rect 11571 8064 11621 8096
rect 11571 8044 11588 8064
rect 11608 8044 11621 8064
rect 11571 8019 11621 8044
rect 11789 8067 11839 8096
rect 13571 8090 13621 8103
rect 13789 8090 13839 8103
rect 13997 8090 14047 8103
rect 16624 8145 16674 8158
rect 16832 8145 16882 8158
rect 17050 8145 17100 8158
rect 11789 8047 11806 8067
rect 11826 8047 11839 8067
rect 11789 8019 11839 8047
rect 9207 7949 9257 7977
rect 6986 7894 7036 7907
rect 7194 7894 7244 7907
rect 7412 7894 7462 7907
rect 9207 7929 9220 7949
rect 9240 7929 9257 7949
rect 9207 7900 9257 7929
rect 9425 7952 9475 7977
rect 9425 7932 9438 7952
rect 9458 7932 9475 7952
rect 9425 7900 9475 7932
rect 9633 7950 9683 7977
rect 9633 7930 9656 7950
rect 9676 7930 9683 7950
rect 9633 7900 9683 7930
rect 14368 8083 14418 8099
rect 14586 8083 14636 8099
rect 14794 8083 14844 8099
rect 15727 8079 15777 8109
rect 15727 8059 15734 8079
rect 15754 8059 15777 8079
rect 15727 8032 15777 8059
rect 15935 8077 15985 8109
rect 15935 8057 15952 8077
rect 15972 8057 15985 8077
rect 15935 8032 15985 8057
rect 16153 8080 16203 8109
rect 16153 8060 16170 8080
rect 16190 8060 16203 8080
rect 16153 8032 16203 8060
rect 13571 7962 13621 7990
rect 11363 7906 11413 7919
rect 11571 7906 11621 7919
rect 11789 7906 11839 7919
rect 13571 7942 13584 7962
rect 13604 7942 13621 7962
rect 13571 7913 13621 7942
rect 13789 7965 13839 7990
rect 13789 7945 13802 7965
rect 13822 7945 13839 7965
rect 13789 7913 13839 7945
rect 13997 7963 14047 7990
rect 13997 7943 14020 7963
rect 14040 7943 14047 7963
rect 13997 7913 14047 7943
rect 15727 7919 15777 7932
rect 15935 7919 15985 7932
rect 16153 7919 16203 7932
rect 466 7817 516 7833
rect 684 7817 734 7833
rect 892 7817 942 7833
rect 4830 7830 4880 7846
rect 5048 7830 5098 7846
rect 5256 7830 5306 7846
rect 9207 7842 9257 7858
rect 9425 7842 9475 7858
rect 9633 7842 9683 7858
rect 13571 7855 13621 7871
rect 13789 7855 13839 7871
rect 13997 7855 14047 7871
rect 3501 7733 3551 7749
rect 3709 7733 3759 7749
rect 3927 7733 3977 7749
rect 7865 7746 7915 7762
rect 8073 7746 8123 7762
rect 8291 7746 8341 7762
rect 12242 7758 12292 7774
rect 12450 7758 12500 7774
rect 12668 7758 12718 7774
rect 16606 7771 16656 7787
rect 16814 7771 16864 7787
rect 17032 7771 17082 7787
rect 1345 7672 1395 7685
rect 1563 7672 1613 7685
rect 1771 7672 1821 7685
rect 3501 7661 3551 7691
rect 3501 7641 3508 7661
rect 3528 7641 3551 7661
rect 3501 7614 3551 7641
rect 3709 7659 3759 7691
rect 3709 7639 3726 7659
rect 3746 7639 3759 7659
rect 3709 7614 3759 7639
rect 3927 7662 3977 7691
rect 3927 7642 3944 7662
rect 3964 7642 3977 7662
rect 5709 7685 5759 7698
rect 5927 7685 5977 7698
rect 6135 7685 6185 7698
rect 3927 7614 3977 7642
rect 1345 7544 1395 7572
rect 1345 7524 1358 7544
rect 1378 7524 1395 7544
rect 1345 7495 1395 7524
rect 1563 7547 1613 7572
rect 1563 7527 1576 7547
rect 1596 7527 1613 7547
rect 1563 7495 1613 7527
rect 1771 7545 1821 7572
rect 1771 7525 1794 7545
rect 1814 7525 1821 7545
rect 1771 7495 1821 7525
rect 2704 7505 2754 7521
rect 2912 7505 2962 7521
rect 3130 7505 3180 7521
rect 7865 7674 7915 7704
rect 7865 7654 7872 7674
rect 7892 7654 7915 7674
rect 7865 7627 7915 7654
rect 8073 7672 8123 7704
rect 8073 7652 8090 7672
rect 8110 7652 8123 7672
rect 8073 7627 8123 7652
rect 8291 7675 8341 7704
rect 8291 7655 8308 7675
rect 8328 7655 8341 7675
rect 10086 7697 10136 7710
rect 10304 7697 10354 7710
rect 10512 7697 10562 7710
rect 8291 7627 8341 7655
rect 5709 7557 5759 7585
rect 5709 7537 5722 7557
rect 5742 7537 5759 7557
rect 448 7446 498 7459
rect 666 7446 716 7459
rect 874 7446 924 7459
rect 3501 7501 3551 7514
rect 3709 7501 3759 7514
rect 3927 7501 3977 7514
rect 5709 7508 5759 7537
rect 5927 7560 5977 7585
rect 5927 7540 5940 7560
rect 5960 7540 5977 7560
rect 5927 7508 5977 7540
rect 6135 7558 6185 7585
rect 6135 7538 6158 7558
rect 6178 7538 6185 7558
rect 6135 7508 6185 7538
rect 7068 7518 7118 7534
rect 7276 7518 7326 7534
rect 7494 7518 7544 7534
rect 12242 7686 12292 7716
rect 12242 7666 12249 7686
rect 12269 7666 12292 7686
rect 12242 7639 12292 7666
rect 12450 7684 12500 7716
rect 12450 7664 12467 7684
rect 12487 7664 12500 7684
rect 12450 7639 12500 7664
rect 12668 7687 12718 7716
rect 12668 7667 12685 7687
rect 12705 7667 12718 7687
rect 14450 7710 14500 7723
rect 14668 7710 14718 7723
rect 14876 7710 14926 7723
rect 12668 7639 12718 7667
rect 10086 7569 10136 7597
rect 10086 7549 10099 7569
rect 10119 7549 10136 7569
rect 1345 7437 1395 7453
rect 1563 7437 1613 7453
rect 1771 7437 1821 7453
rect 2704 7433 2754 7463
rect 2704 7413 2711 7433
rect 2731 7413 2754 7433
rect 2704 7386 2754 7413
rect 2912 7431 2962 7463
rect 2912 7411 2929 7431
rect 2949 7411 2962 7431
rect 2912 7386 2962 7411
rect 3130 7434 3180 7463
rect 3130 7414 3147 7434
rect 3167 7414 3180 7434
rect 4812 7459 4862 7472
rect 5030 7459 5080 7472
rect 5238 7459 5288 7472
rect 7865 7514 7915 7527
rect 8073 7514 8123 7527
rect 8291 7514 8341 7527
rect 10086 7520 10136 7549
rect 10304 7572 10354 7597
rect 10304 7552 10317 7572
rect 10337 7552 10354 7572
rect 10304 7520 10354 7552
rect 10512 7570 10562 7597
rect 10512 7550 10535 7570
rect 10555 7550 10562 7570
rect 10512 7520 10562 7550
rect 11445 7530 11495 7546
rect 11653 7530 11703 7546
rect 11871 7530 11921 7546
rect 16606 7699 16656 7729
rect 16606 7679 16613 7699
rect 16633 7679 16656 7699
rect 16606 7652 16656 7679
rect 16814 7697 16864 7729
rect 16814 7677 16831 7697
rect 16851 7677 16864 7697
rect 16814 7652 16864 7677
rect 17032 7700 17082 7729
rect 17032 7680 17049 7700
rect 17069 7680 17082 7700
rect 17032 7652 17082 7680
rect 14450 7582 14500 7610
rect 14450 7562 14463 7582
rect 14483 7562 14500 7582
rect 3130 7386 3180 7414
rect 448 7318 498 7346
rect 448 7298 461 7318
rect 481 7298 498 7318
rect 448 7269 498 7298
rect 666 7321 716 7346
rect 666 7301 679 7321
rect 699 7301 716 7321
rect 666 7269 716 7301
rect 874 7319 924 7346
rect 874 7299 897 7319
rect 917 7299 924 7319
rect 874 7269 924 7299
rect 5709 7450 5759 7466
rect 5927 7450 5977 7466
rect 6135 7450 6185 7466
rect 7068 7446 7118 7476
rect 7068 7426 7075 7446
rect 7095 7426 7118 7446
rect 7068 7399 7118 7426
rect 7276 7444 7326 7476
rect 7276 7424 7293 7444
rect 7313 7424 7326 7444
rect 7276 7399 7326 7424
rect 7494 7447 7544 7476
rect 7494 7427 7511 7447
rect 7531 7427 7544 7447
rect 9189 7471 9239 7484
rect 9407 7471 9457 7484
rect 9615 7471 9665 7484
rect 12242 7526 12292 7539
rect 12450 7526 12500 7539
rect 12668 7526 12718 7539
rect 14450 7533 14500 7562
rect 14668 7585 14718 7610
rect 14668 7565 14681 7585
rect 14701 7565 14718 7585
rect 14668 7533 14718 7565
rect 14876 7583 14926 7610
rect 14876 7563 14899 7583
rect 14919 7563 14926 7583
rect 14876 7533 14926 7563
rect 15809 7543 15859 7559
rect 16017 7543 16067 7559
rect 16235 7543 16285 7559
rect 7494 7399 7544 7427
rect 3502 7321 3552 7337
rect 3710 7321 3760 7337
rect 3928 7321 3978 7337
rect 1246 7262 1296 7275
rect 1464 7262 1514 7275
rect 1672 7262 1722 7275
rect 2704 7273 2754 7286
rect 2912 7273 2962 7286
rect 3130 7273 3180 7286
rect 4812 7331 4862 7359
rect 448 7211 498 7227
rect 666 7211 716 7227
rect 874 7211 924 7227
rect 3502 7249 3552 7279
rect 3502 7229 3509 7249
rect 3529 7229 3552 7249
rect 3502 7202 3552 7229
rect 3710 7247 3760 7279
rect 3710 7227 3727 7247
rect 3747 7227 3760 7247
rect 3710 7202 3760 7227
rect 3928 7250 3978 7279
rect 3928 7230 3945 7250
rect 3965 7230 3978 7250
rect 4812 7311 4825 7331
rect 4845 7311 4862 7331
rect 4812 7282 4862 7311
rect 5030 7334 5080 7359
rect 5030 7314 5043 7334
rect 5063 7314 5080 7334
rect 5030 7282 5080 7314
rect 5238 7332 5288 7359
rect 5238 7312 5261 7332
rect 5281 7312 5288 7332
rect 5238 7282 5288 7312
rect 10086 7462 10136 7478
rect 10304 7462 10354 7478
rect 10512 7462 10562 7478
rect 11445 7458 11495 7488
rect 11445 7438 11452 7458
rect 11472 7438 11495 7458
rect 11445 7411 11495 7438
rect 11653 7456 11703 7488
rect 11653 7436 11670 7456
rect 11690 7436 11703 7456
rect 11653 7411 11703 7436
rect 11871 7459 11921 7488
rect 11871 7439 11888 7459
rect 11908 7439 11921 7459
rect 13553 7484 13603 7497
rect 13771 7484 13821 7497
rect 13979 7484 14029 7497
rect 16606 7539 16656 7552
rect 16814 7539 16864 7552
rect 17032 7539 17082 7552
rect 11871 7411 11921 7439
rect 7866 7334 7916 7350
rect 8074 7334 8124 7350
rect 8292 7334 8342 7350
rect 3928 7202 3978 7230
rect 5610 7275 5660 7288
rect 5828 7275 5878 7288
rect 6036 7275 6086 7288
rect 7068 7286 7118 7299
rect 7276 7286 7326 7299
rect 7494 7286 7544 7299
rect 9189 7343 9239 7371
rect 4812 7224 4862 7240
rect 5030 7224 5080 7240
rect 5238 7224 5288 7240
rect 1246 7134 1296 7162
rect 1246 7114 1259 7134
rect 1279 7114 1296 7134
rect 1246 7085 1296 7114
rect 1464 7137 1514 7162
rect 1464 7117 1477 7137
rect 1497 7117 1514 7137
rect 1464 7085 1514 7117
rect 1672 7135 1722 7162
rect 1672 7115 1695 7135
rect 1715 7115 1722 7135
rect 1672 7085 1722 7115
rect 2539 7097 2589 7113
rect 2747 7097 2797 7113
rect 2965 7097 3015 7113
rect 7866 7262 7916 7292
rect 7866 7242 7873 7262
rect 7893 7242 7916 7262
rect 7866 7215 7916 7242
rect 8074 7260 8124 7292
rect 8074 7240 8091 7260
rect 8111 7240 8124 7260
rect 8074 7215 8124 7240
rect 8292 7263 8342 7292
rect 8292 7243 8309 7263
rect 8329 7243 8342 7263
rect 9189 7323 9202 7343
rect 9222 7323 9239 7343
rect 9189 7294 9239 7323
rect 9407 7346 9457 7371
rect 9407 7326 9420 7346
rect 9440 7326 9457 7346
rect 9407 7294 9457 7326
rect 9615 7344 9665 7371
rect 9615 7324 9638 7344
rect 9658 7324 9665 7344
rect 9615 7294 9665 7324
rect 14450 7475 14500 7491
rect 14668 7475 14718 7491
rect 14876 7475 14926 7491
rect 15809 7471 15859 7501
rect 15809 7451 15816 7471
rect 15836 7451 15859 7471
rect 15809 7424 15859 7451
rect 16017 7469 16067 7501
rect 16017 7449 16034 7469
rect 16054 7449 16067 7469
rect 16017 7424 16067 7449
rect 16235 7472 16285 7501
rect 16235 7452 16252 7472
rect 16272 7452 16285 7472
rect 16235 7424 16285 7452
rect 12243 7346 12293 7362
rect 12451 7346 12501 7362
rect 12669 7346 12719 7362
rect 8292 7215 8342 7243
rect 9987 7287 10037 7300
rect 10205 7287 10255 7300
rect 10413 7287 10463 7300
rect 11445 7298 11495 7311
rect 11653 7298 11703 7311
rect 11871 7298 11921 7311
rect 13553 7356 13603 7384
rect 9189 7236 9239 7252
rect 9407 7236 9457 7252
rect 9615 7236 9665 7252
rect 5610 7147 5660 7175
rect 449 7034 499 7047
rect 667 7034 717 7047
rect 875 7034 925 7047
rect 3502 7089 3552 7102
rect 3710 7089 3760 7102
rect 3928 7089 3978 7102
rect 5610 7127 5623 7147
rect 5643 7127 5660 7147
rect 5610 7098 5660 7127
rect 5828 7150 5878 7175
rect 5828 7130 5841 7150
rect 5861 7130 5878 7150
rect 5828 7098 5878 7130
rect 6036 7148 6086 7175
rect 6036 7128 6059 7148
rect 6079 7128 6086 7148
rect 6036 7098 6086 7128
rect 6903 7110 6953 7126
rect 7111 7110 7161 7126
rect 7329 7110 7379 7126
rect 12243 7274 12293 7304
rect 12243 7254 12250 7274
rect 12270 7254 12293 7274
rect 12243 7227 12293 7254
rect 12451 7272 12501 7304
rect 12451 7252 12468 7272
rect 12488 7252 12501 7272
rect 12451 7227 12501 7252
rect 12669 7275 12719 7304
rect 12669 7255 12686 7275
rect 12706 7255 12719 7275
rect 13553 7336 13566 7356
rect 13586 7336 13603 7356
rect 13553 7307 13603 7336
rect 13771 7359 13821 7384
rect 13771 7339 13784 7359
rect 13804 7339 13821 7359
rect 13771 7307 13821 7339
rect 13979 7357 14029 7384
rect 13979 7337 14002 7357
rect 14022 7337 14029 7357
rect 13979 7307 14029 7337
rect 16607 7359 16657 7375
rect 16815 7359 16865 7375
rect 17033 7359 17083 7375
rect 12669 7227 12719 7255
rect 14351 7300 14401 7313
rect 14569 7300 14619 7313
rect 14777 7300 14827 7313
rect 15809 7311 15859 7324
rect 16017 7311 16067 7324
rect 16235 7311 16285 7324
rect 13553 7249 13603 7265
rect 13771 7249 13821 7265
rect 13979 7249 14029 7265
rect 9987 7159 10037 7187
rect 1246 7027 1296 7043
rect 1464 7027 1514 7043
rect 1672 7027 1722 7043
rect 2539 7025 2589 7055
rect 2539 7005 2546 7025
rect 2566 7005 2589 7025
rect 2539 6978 2589 7005
rect 2747 7023 2797 7055
rect 2747 7003 2764 7023
rect 2784 7003 2797 7023
rect 2747 6978 2797 7003
rect 2965 7026 3015 7055
rect 4813 7047 4863 7060
rect 5031 7047 5081 7060
rect 5239 7047 5289 7060
rect 7866 7102 7916 7115
rect 8074 7102 8124 7115
rect 8292 7102 8342 7115
rect 9987 7139 10000 7159
rect 10020 7139 10037 7159
rect 9987 7110 10037 7139
rect 10205 7162 10255 7187
rect 10205 7142 10218 7162
rect 10238 7142 10255 7162
rect 10205 7110 10255 7142
rect 10413 7160 10463 7187
rect 10413 7140 10436 7160
rect 10456 7140 10463 7160
rect 10413 7110 10463 7140
rect 11280 7122 11330 7138
rect 11488 7122 11538 7138
rect 11706 7122 11756 7138
rect 16607 7287 16657 7317
rect 16607 7267 16614 7287
rect 16634 7267 16657 7287
rect 16607 7240 16657 7267
rect 16815 7285 16865 7317
rect 16815 7265 16832 7285
rect 16852 7265 16865 7285
rect 16815 7240 16865 7265
rect 17033 7288 17083 7317
rect 17033 7268 17050 7288
rect 17070 7268 17083 7288
rect 17033 7240 17083 7268
rect 14351 7172 14401 7200
rect 2965 7006 2982 7026
rect 3002 7006 3015 7026
rect 2965 6978 3015 7006
rect 449 6906 499 6934
rect 449 6886 462 6906
rect 482 6886 499 6906
rect 449 6857 499 6886
rect 667 6909 717 6934
rect 667 6889 680 6909
rect 700 6889 717 6909
rect 667 6857 717 6889
rect 875 6907 925 6934
rect 875 6887 898 6907
rect 918 6887 925 6907
rect 875 6857 925 6887
rect 5610 7040 5660 7056
rect 5828 7040 5878 7056
rect 6036 7040 6086 7056
rect 6903 7038 6953 7068
rect 6903 7018 6910 7038
rect 6930 7018 6953 7038
rect 6903 6991 6953 7018
rect 7111 7036 7161 7068
rect 7111 7016 7128 7036
rect 7148 7016 7161 7036
rect 7111 6991 7161 7016
rect 7329 7039 7379 7068
rect 9190 7059 9240 7072
rect 9408 7059 9458 7072
rect 9616 7059 9666 7072
rect 12243 7114 12293 7127
rect 12451 7114 12501 7127
rect 12669 7114 12719 7127
rect 14351 7152 14364 7172
rect 14384 7152 14401 7172
rect 14351 7123 14401 7152
rect 14569 7175 14619 7200
rect 14569 7155 14582 7175
rect 14602 7155 14619 7175
rect 14569 7123 14619 7155
rect 14777 7173 14827 7200
rect 14777 7153 14800 7173
rect 14820 7153 14827 7173
rect 14777 7123 14827 7153
rect 15644 7135 15694 7151
rect 15852 7135 15902 7151
rect 16070 7135 16120 7151
rect 7329 7019 7346 7039
rect 7366 7019 7379 7039
rect 7329 6991 7379 7019
rect 4813 6919 4863 6947
rect 2539 6865 2589 6878
rect 2747 6865 2797 6878
rect 2965 6865 3015 6878
rect 4813 6899 4826 6919
rect 4846 6899 4863 6919
rect 4813 6870 4863 6899
rect 5031 6922 5081 6947
rect 5031 6902 5044 6922
rect 5064 6902 5081 6922
rect 5031 6870 5081 6902
rect 5239 6920 5289 6947
rect 5239 6900 5262 6920
rect 5282 6900 5289 6920
rect 5239 6870 5289 6900
rect 9987 7052 10037 7068
rect 10205 7052 10255 7068
rect 10413 7052 10463 7068
rect 11280 7050 11330 7080
rect 11280 7030 11287 7050
rect 11307 7030 11330 7050
rect 11280 7003 11330 7030
rect 11488 7048 11538 7080
rect 11488 7028 11505 7048
rect 11525 7028 11538 7048
rect 11488 7003 11538 7028
rect 11706 7051 11756 7080
rect 13554 7072 13604 7085
rect 13772 7072 13822 7085
rect 13980 7072 14030 7085
rect 16607 7127 16657 7140
rect 16815 7127 16865 7140
rect 17033 7127 17083 7140
rect 11706 7031 11723 7051
rect 11743 7031 11756 7051
rect 11706 7003 11756 7031
rect 9190 6931 9240 6959
rect 6903 6878 6953 6891
rect 7111 6878 7161 6891
rect 7329 6878 7379 6891
rect 9190 6911 9203 6931
rect 9223 6911 9240 6931
rect 9190 6882 9240 6911
rect 9408 6934 9458 6959
rect 9408 6914 9421 6934
rect 9441 6914 9458 6934
rect 9408 6882 9458 6914
rect 9616 6932 9666 6959
rect 9616 6912 9639 6932
rect 9659 6912 9666 6932
rect 9616 6882 9666 6912
rect 14351 7065 14401 7081
rect 14569 7065 14619 7081
rect 14777 7065 14827 7081
rect 15644 7063 15694 7093
rect 15644 7043 15651 7063
rect 15671 7043 15694 7063
rect 15644 7016 15694 7043
rect 15852 7061 15902 7093
rect 15852 7041 15869 7061
rect 15889 7041 15902 7061
rect 15852 7016 15902 7041
rect 16070 7064 16120 7093
rect 16070 7044 16087 7064
rect 16107 7044 16120 7064
rect 16070 7016 16120 7044
rect 13554 6944 13604 6972
rect 11280 6890 11330 6903
rect 11488 6890 11538 6903
rect 11706 6890 11756 6903
rect 13554 6924 13567 6944
rect 13587 6924 13604 6944
rect 13554 6895 13604 6924
rect 13772 6947 13822 6972
rect 13772 6927 13785 6947
rect 13805 6927 13822 6947
rect 13772 6895 13822 6927
rect 13980 6945 14030 6972
rect 13980 6925 14003 6945
rect 14023 6925 14030 6945
rect 13980 6895 14030 6925
rect 15644 6903 15694 6916
rect 15852 6903 15902 6916
rect 16070 6903 16120 6916
rect 449 6799 499 6815
rect 667 6799 717 6815
rect 875 6799 925 6815
rect 4813 6812 4863 6828
rect 5031 6812 5081 6828
rect 5239 6812 5289 6828
rect 9190 6824 9240 6840
rect 9408 6824 9458 6840
rect 9616 6824 9666 6840
rect 13554 6837 13604 6853
rect 13772 6837 13822 6853
rect 13980 6837 14030 6853
rect 3481 6715 3531 6731
rect 3689 6715 3739 6731
rect 3907 6715 3957 6731
rect 7845 6728 7895 6744
rect 8053 6728 8103 6744
rect 8271 6728 8321 6744
rect 12222 6740 12272 6756
rect 12430 6740 12480 6756
rect 12648 6740 12698 6756
rect 16586 6753 16636 6769
rect 16794 6753 16844 6769
rect 17012 6753 17062 6769
rect 1391 6652 1441 6665
rect 1609 6652 1659 6665
rect 1817 6652 1867 6665
rect 3481 6643 3531 6673
rect 3481 6623 3488 6643
rect 3508 6623 3531 6643
rect 3481 6596 3531 6623
rect 3689 6641 3739 6673
rect 3689 6621 3706 6641
rect 3726 6621 3739 6641
rect 3689 6596 3739 6621
rect 3907 6644 3957 6673
rect 3907 6624 3924 6644
rect 3944 6624 3957 6644
rect 5755 6665 5805 6678
rect 5973 6665 6023 6678
rect 6181 6665 6231 6678
rect 3907 6596 3957 6624
rect 1391 6524 1441 6552
rect 1391 6504 1404 6524
rect 1424 6504 1441 6524
rect 1391 6475 1441 6504
rect 1609 6527 1659 6552
rect 1609 6507 1622 6527
rect 1642 6507 1659 6527
rect 1609 6475 1659 6507
rect 1817 6525 1867 6552
rect 1817 6505 1840 6525
rect 1860 6505 1867 6525
rect 1817 6475 1867 6505
rect 2684 6487 2734 6503
rect 2892 6487 2942 6503
rect 3110 6487 3160 6503
rect 7845 6656 7895 6686
rect 7845 6636 7852 6656
rect 7872 6636 7895 6656
rect 7845 6609 7895 6636
rect 8053 6654 8103 6686
rect 8053 6634 8070 6654
rect 8090 6634 8103 6654
rect 8053 6609 8103 6634
rect 8271 6657 8321 6686
rect 8271 6637 8288 6657
rect 8308 6637 8321 6657
rect 10132 6677 10182 6690
rect 10350 6677 10400 6690
rect 10558 6677 10608 6690
rect 8271 6609 8321 6637
rect 5755 6537 5805 6565
rect 5755 6517 5768 6537
rect 5788 6517 5805 6537
rect 428 6428 478 6441
rect 646 6428 696 6441
rect 854 6428 904 6441
rect 3481 6483 3531 6496
rect 3689 6483 3739 6496
rect 3907 6483 3957 6496
rect 5755 6488 5805 6517
rect 5973 6540 6023 6565
rect 5973 6520 5986 6540
rect 6006 6520 6023 6540
rect 5973 6488 6023 6520
rect 6181 6538 6231 6565
rect 6181 6518 6204 6538
rect 6224 6518 6231 6538
rect 6181 6488 6231 6518
rect 7048 6500 7098 6516
rect 7256 6500 7306 6516
rect 7474 6500 7524 6516
rect 12222 6668 12272 6698
rect 12222 6648 12229 6668
rect 12249 6648 12272 6668
rect 12222 6621 12272 6648
rect 12430 6666 12480 6698
rect 12430 6646 12447 6666
rect 12467 6646 12480 6666
rect 12430 6621 12480 6646
rect 12648 6669 12698 6698
rect 12648 6649 12665 6669
rect 12685 6649 12698 6669
rect 14496 6690 14546 6703
rect 14714 6690 14764 6703
rect 14922 6690 14972 6703
rect 12648 6621 12698 6649
rect 10132 6549 10182 6577
rect 10132 6529 10145 6549
rect 10165 6529 10182 6549
rect 1391 6417 1441 6433
rect 1609 6417 1659 6433
rect 1817 6417 1867 6433
rect 2684 6415 2734 6445
rect 2684 6395 2691 6415
rect 2711 6395 2734 6415
rect 2684 6368 2734 6395
rect 2892 6413 2942 6445
rect 2892 6393 2909 6413
rect 2929 6393 2942 6413
rect 2892 6368 2942 6393
rect 3110 6416 3160 6445
rect 3110 6396 3127 6416
rect 3147 6396 3160 6416
rect 4792 6441 4842 6454
rect 5010 6441 5060 6454
rect 5218 6441 5268 6454
rect 7845 6496 7895 6509
rect 8053 6496 8103 6509
rect 8271 6496 8321 6509
rect 10132 6500 10182 6529
rect 10350 6552 10400 6577
rect 10350 6532 10363 6552
rect 10383 6532 10400 6552
rect 10350 6500 10400 6532
rect 10558 6550 10608 6577
rect 10558 6530 10581 6550
rect 10601 6530 10608 6550
rect 10558 6500 10608 6530
rect 11425 6512 11475 6528
rect 11633 6512 11683 6528
rect 11851 6512 11901 6528
rect 16586 6681 16636 6711
rect 16586 6661 16593 6681
rect 16613 6661 16636 6681
rect 16586 6634 16636 6661
rect 16794 6679 16844 6711
rect 16794 6659 16811 6679
rect 16831 6659 16844 6679
rect 16794 6634 16844 6659
rect 17012 6682 17062 6711
rect 17012 6662 17029 6682
rect 17049 6662 17062 6682
rect 17012 6634 17062 6662
rect 14496 6562 14546 6590
rect 14496 6542 14509 6562
rect 14529 6542 14546 6562
rect 3110 6368 3160 6396
rect 428 6300 478 6328
rect 428 6280 441 6300
rect 461 6280 478 6300
rect 428 6251 478 6280
rect 646 6303 696 6328
rect 646 6283 659 6303
rect 679 6283 696 6303
rect 646 6251 696 6283
rect 854 6301 904 6328
rect 854 6281 877 6301
rect 897 6281 904 6301
rect 854 6251 904 6281
rect 5755 6430 5805 6446
rect 5973 6430 6023 6446
rect 6181 6430 6231 6446
rect 7048 6428 7098 6458
rect 7048 6408 7055 6428
rect 7075 6408 7098 6428
rect 7048 6381 7098 6408
rect 7256 6426 7306 6458
rect 7256 6406 7273 6426
rect 7293 6406 7306 6426
rect 7256 6381 7306 6406
rect 7474 6429 7524 6458
rect 7474 6409 7491 6429
rect 7511 6409 7524 6429
rect 9169 6453 9219 6466
rect 9387 6453 9437 6466
rect 9595 6453 9645 6466
rect 12222 6508 12272 6521
rect 12430 6508 12480 6521
rect 12648 6508 12698 6521
rect 14496 6513 14546 6542
rect 14714 6565 14764 6590
rect 14714 6545 14727 6565
rect 14747 6545 14764 6565
rect 14714 6513 14764 6545
rect 14922 6563 14972 6590
rect 14922 6543 14945 6563
rect 14965 6543 14972 6563
rect 14922 6513 14972 6543
rect 15789 6525 15839 6541
rect 15997 6525 16047 6541
rect 16215 6525 16265 6541
rect 7474 6381 7524 6409
rect 3482 6303 3532 6319
rect 3690 6303 3740 6319
rect 3908 6303 3958 6319
rect 1226 6244 1276 6257
rect 1444 6244 1494 6257
rect 1652 6244 1702 6257
rect 2684 6255 2734 6268
rect 2892 6255 2942 6268
rect 3110 6255 3160 6268
rect 4792 6313 4842 6341
rect 428 6193 478 6209
rect 646 6193 696 6209
rect 854 6193 904 6209
rect 3482 6231 3532 6261
rect 3482 6211 3489 6231
rect 3509 6211 3532 6231
rect 3482 6184 3532 6211
rect 3690 6229 3740 6261
rect 3690 6209 3707 6229
rect 3727 6209 3740 6229
rect 3690 6184 3740 6209
rect 3908 6232 3958 6261
rect 3908 6212 3925 6232
rect 3945 6212 3958 6232
rect 4792 6293 4805 6313
rect 4825 6293 4842 6313
rect 4792 6264 4842 6293
rect 5010 6316 5060 6341
rect 5010 6296 5023 6316
rect 5043 6296 5060 6316
rect 5010 6264 5060 6296
rect 5218 6314 5268 6341
rect 5218 6294 5241 6314
rect 5261 6294 5268 6314
rect 5218 6264 5268 6294
rect 10132 6442 10182 6458
rect 10350 6442 10400 6458
rect 10558 6442 10608 6458
rect 11425 6440 11475 6470
rect 11425 6420 11432 6440
rect 11452 6420 11475 6440
rect 11425 6393 11475 6420
rect 11633 6438 11683 6470
rect 11633 6418 11650 6438
rect 11670 6418 11683 6438
rect 11633 6393 11683 6418
rect 11851 6441 11901 6470
rect 11851 6421 11868 6441
rect 11888 6421 11901 6441
rect 13533 6466 13583 6479
rect 13751 6466 13801 6479
rect 13959 6466 14009 6479
rect 16586 6521 16636 6534
rect 16794 6521 16844 6534
rect 17012 6521 17062 6534
rect 11851 6393 11901 6421
rect 7846 6316 7896 6332
rect 8054 6316 8104 6332
rect 8272 6316 8322 6332
rect 3908 6184 3958 6212
rect 5590 6257 5640 6270
rect 5808 6257 5858 6270
rect 6016 6257 6066 6270
rect 7048 6268 7098 6281
rect 7256 6268 7306 6281
rect 7474 6268 7524 6281
rect 9169 6325 9219 6353
rect 4792 6206 4842 6222
rect 5010 6206 5060 6222
rect 5218 6206 5268 6222
rect 1226 6116 1276 6144
rect 1226 6096 1239 6116
rect 1259 6096 1276 6116
rect 1226 6067 1276 6096
rect 1444 6119 1494 6144
rect 1444 6099 1457 6119
rect 1477 6099 1494 6119
rect 1444 6067 1494 6099
rect 1652 6117 1702 6144
rect 1652 6097 1675 6117
rect 1695 6097 1702 6117
rect 1652 6067 1702 6097
rect 2585 6077 2635 6093
rect 2793 6077 2843 6093
rect 3011 6077 3061 6093
rect 7846 6244 7896 6274
rect 7846 6224 7853 6244
rect 7873 6224 7896 6244
rect 7846 6197 7896 6224
rect 8054 6242 8104 6274
rect 8054 6222 8071 6242
rect 8091 6222 8104 6242
rect 8054 6197 8104 6222
rect 8272 6245 8322 6274
rect 8272 6225 8289 6245
rect 8309 6225 8322 6245
rect 9169 6305 9182 6325
rect 9202 6305 9219 6325
rect 9169 6276 9219 6305
rect 9387 6328 9437 6353
rect 9387 6308 9400 6328
rect 9420 6308 9437 6328
rect 9387 6276 9437 6308
rect 9595 6326 9645 6353
rect 9595 6306 9618 6326
rect 9638 6306 9645 6326
rect 9595 6276 9645 6306
rect 14496 6455 14546 6471
rect 14714 6455 14764 6471
rect 14922 6455 14972 6471
rect 15789 6453 15839 6483
rect 15789 6433 15796 6453
rect 15816 6433 15839 6453
rect 15789 6406 15839 6433
rect 15997 6451 16047 6483
rect 15997 6431 16014 6451
rect 16034 6431 16047 6451
rect 15997 6406 16047 6431
rect 16215 6454 16265 6483
rect 16215 6434 16232 6454
rect 16252 6434 16265 6454
rect 16215 6406 16265 6434
rect 12223 6328 12273 6344
rect 12431 6328 12481 6344
rect 12649 6328 12699 6344
rect 8272 6197 8322 6225
rect 9967 6269 10017 6282
rect 10185 6269 10235 6282
rect 10393 6269 10443 6282
rect 11425 6280 11475 6293
rect 11633 6280 11683 6293
rect 11851 6280 11901 6293
rect 13533 6338 13583 6366
rect 9169 6218 9219 6234
rect 9387 6218 9437 6234
rect 9595 6218 9645 6234
rect 5590 6129 5640 6157
rect 429 6016 479 6029
rect 647 6016 697 6029
rect 855 6016 905 6029
rect 3482 6071 3532 6084
rect 3690 6071 3740 6084
rect 3908 6071 3958 6084
rect 5590 6109 5603 6129
rect 5623 6109 5640 6129
rect 5590 6080 5640 6109
rect 5808 6132 5858 6157
rect 5808 6112 5821 6132
rect 5841 6112 5858 6132
rect 5808 6080 5858 6112
rect 6016 6130 6066 6157
rect 6016 6110 6039 6130
rect 6059 6110 6066 6130
rect 6016 6080 6066 6110
rect 6949 6090 6999 6106
rect 7157 6090 7207 6106
rect 7375 6090 7425 6106
rect 12223 6256 12273 6286
rect 12223 6236 12230 6256
rect 12250 6236 12273 6256
rect 12223 6209 12273 6236
rect 12431 6254 12481 6286
rect 12431 6234 12448 6254
rect 12468 6234 12481 6254
rect 12431 6209 12481 6234
rect 12649 6257 12699 6286
rect 12649 6237 12666 6257
rect 12686 6237 12699 6257
rect 13533 6318 13546 6338
rect 13566 6318 13583 6338
rect 13533 6289 13583 6318
rect 13751 6341 13801 6366
rect 13751 6321 13764 6341
rect 13784 6321 13801 6341
rect 13751 6289 13801 6321
rect 13959 6339 14009 6366
rect 13959 6319 13982 6339
rect 14002 6319 14009 6339
rect 13959 6289 14009 6319
rect 16587 6341 16637 6357
rect 16795 6341 16845 6357
rect 17013 6341 17063 6357
rect 12649 6209 12699 6237
rect 14331 6282 14381 6295
rect 14549 6282 14599 6295
rect 14757 6282 14807 6295
rect 15789 6293 15839 6306
rect 15997 6293 16047 6306
rect 16215 6293 16265 6306
rect 13533 6231 13583 6247
rect 13751 6231 13801 6247
rect 13959 6231 14009 6247
rect 9967 6141 10017 6169
rect 1226 6009 1276 6025
rect 1444 6009 1494 6025
rect 1652 6009 1702 6025
rect 2585 6005 2635 6035
rect 2585 5985 2592 6005
rect 2612 5985 2635 6005
rect 2585 5958 2635 5985
rect 2793 6003 2843 6035
rect 2793 5983 2810 6003
rect 2830 5983 2843 6003
rect 2793 5958 2843 5983
rect 3011 6006 3061 6035
rect 4793 6029 4843 6042
rect 5011 6029 5061 6042
rect 5219 6029 5269 6042
rect 7846 6084 7896 6097
rect 8054 6084 8104 6097
rect 8272 6084 8322 6097
rect 9967 6121 9980 6141
rect 10000 6121 10017 6141
rect 9967 6092 10017 6121
rect 10185 6144 10235 6169
rect 10185 6124 10198 6144
rect 10218 6124 10235 6144
rect 10185 6092 10235 6124
rect 10393 6142 10443 6169
rect 10393 6122 10416 6142
rect 10436 6122 10443 6142
rect 10393 6092 10443 6122
rect 11326 6102 11376 6118
rect 11534 6102 11584 6118
rect 11752 6102 11802 6118
rect 16587 6269 16637 6299
rect 16587 6249 16594 6269
rect 16614 6249 16637 6269
rect 16587 6222 16637 6249
rect 16795 6267 16845 6299
rect 16795 6247 16812 6267
rect 16832 6247 16845 6267
rect 16795 6222 16845 6247
rect 17013 6270 17063 6299
rect 17013 6250 17030 6270
rect 17050 6250 17063 6270
rect 17013 6222 17063 6250
rect 14331 6154 14381 6182
rect 3011 5986 3028 6006
rect 3048 5986 3061 6006
rect 3011 5958 3061 5986
rect 429 5888 479 5916
rect 429 5868 442 5888
rect 462 5868 479 5888
rect 429 5839 479 5868
rect 647 5891 697 5916
rect 647 5871 660 5891
rect 680 5871 697 5891
rect 647 5839 697 5871
rect 855 5889 905 5916
rect 855 5869 878 5889
rect 898 5869 905 5889
rect 855 5839 905 5869
rect 5590 6022 5640 6038
rect 5808 6022 5858 6038
rect 6016 6022 6066 6038
rect 6949 6018 6999 6048
rect 6949 5998 6956 6018
rect 6976 5998 6999 6018
rect 6949 5971 6999 5998
rect 7157 6016 7207 6048
rect 7157 5996 7174 6016
rect 7194 5996 7207 6016
rect 7157 5971 7207 5996
rect 7375 6019 7425 6048
rect 9170 6041 9220 6054
rect 9388 6041 9438 6054
rect 9596 6041 9646 6054
rect 12223 6096 12273 6109
rect 12431 6096 12481 6109
rect 12649 6096 12699 6109
rect 14331 6134 14344 6154
rect 14364 6134 14381 6154
rect 14331 6105 14381 6134
rect 14549 6157 14599 6182
rect 14549 6137 14562 6157
rect 14582 6137 14599 6157
rect 14549 6105 14599 6137
rect 14757 6155 14807 6182
rect 14757 6135 14780 6155
rect 14800 6135 14807 6155
rect 14757 6105 14807 6135
rect 15690 6115 15740 6131
rect 15898 6115 15948 6131
rect 16116 6115 16166 6131
rect 7375 5999 7392 6019
rect 7412 5999 7425 6019
rect 7375 5971 7425 5999
rect 4793 5901 4843 5929
rect 2585 5845 2635 5858
rect 2793 5845 2843 5858
rect 3011 5845 3061 5858
rect 4793 5881 4806 5901
rect 4826 5881 4843 5901
rect 4793 5852 4843 5881
rect 5011 5904 5061 5929
rect 5011 5884 5024 5904
rect 5044 5884 5061 5904
rect 5011 5852 5061 5884
rect 5219 5902 5269 5929
rect 5219 5882 5242 5902
rect 5262 5882 5269 5902
rect 5219 5852 5269 5882
rect 9967 6034 10017 6050
rect 10185 6034 10235 6050
rect 10393 6034 10443 6050
rect 11326 6030 11376 6060
rect 11326 6010 11333 6030
rect 11353 6010 11376 6030
rect 11326 5983 11376 6010
rect 11534 6028 11584 6060
rect 11534 6008 11551 6028
rect 11571 6008 11584 6028
rect 11534 5983 11584 6008
rect 11752 6031 11802 6060
rect 13534 6054 13584 6067
rect 13752 6054 13802 6067
rect 13960 6054 14010 6067
rect 16587 6109 16637 6122
rect 16795 6109 16845 6122
rect 17013 6109 17063 6122
rect 11752 6011 11769 6031
rect 11789 6011 11802 6031
rect 11752 5983 11802 6011
rect 9170 5913 9220 5941
rect 6949 5858 6999 5871
rect 7157 5858 7207 5871
rect 7375 5858 7425 5871
rect 9170 5893 9183 5913
rect 9203 5893 9220 5913
rect 9170 5864 9220 5893
rect 9388 5916 9438 5941
rect 9388 5896 9401 5916
rect 9421 5896 9438 5916
rect 9388 5864 9438 5896
rect 9596 5914 9646 5941
rect 9596 5894 9619 5914
rect 9639 5894 9646 5914
rect 9596 5864 9646 5894
rect 14331 6047 14381 6063
rect 14549 6047 14599 6063
rect 14757 6047 14807 6063
rect 15690 6043 15740 6073
rect 15690 6023 15697 6043
rect 15717 6023 15740 6043
rect 15690 5996 15740 6023
rect 15898 6041 15948 6073
rect 15898 6021 15915 6041
rect 15935 6021 15948 6041
rect 15898 5996 15948 6021
rect 16116 6044 16166 6073
rect 16116 6024 16133 6044
rect 16153 6024 16166 6044
rect 16116 5996 16166 6024
rect 13534 5926 13584 5954
rect 11326 5870 11376 5883
rect 11534 5870 11584 5883
rect 11752 5870 11802 5883
rect 13534 5906 13547 5926
rect 13567 5906 13584 5926
rect 13534 5877 13584 5906
rect 13752 5929 13802 5954
rect 13752 5909 13765 5929
rect 13785 5909 13802 5929
rect 13752 5877 13802 5909
rect 13960 5927 14010 5954
rect 13960 5907 13983 5927
rect 14003 5907 14010 5927
rect 13960 5877 14010 5907
rect 15690 5883 15740 5896
rect 15898 5883 15948 5896
rect 16116 5883 16166 5896
rect 429 5781 479 5797
rect 647 5781 697 5797
rect 855 5781 905 5797
rect 4793 5794 4843 5810
rect 5011 5794 5061 5810
rect 5219 5794 5269 5810
rect 9170 5806 9220 5822
rect 9388 5806 9438 5822
rect 9596 5806 9646 5822
rect 13534 5819 13584 5835
rect 13752 5819 13802 5835
rect 13960 5819 14010 5835
rect 3464 5697 3514 5713
rect 3672 5697 3722 5713
rect 3890 5697 3940 5713
rect 7828 5710 7878 5726
rect 8036 5710 8086 5726
rect 8254 5710 8304 5726
rect 12205 5722 12255 5738
rect 12413 5722 12463 5738
rect 12631 5722 12681 5738
rect 16569 5735 16619 5751
rect 16777 5735 16827 5751
rect 16995 5735 17045 5751
rect 1308 5636 1358 5649
rect 1526 5636 1576 5649
rect 1734 5636 1784 5649
rect 3464 5625 3514 5655
rect 3464 5605 3471 5625
rect 3491 5605 3514 5625
rect 3464 5578 3514 5605
rect 3672 5623 3722 5655
rect 3672 5603 3689 5623
rect 3709 5603 3722 5623
rect 3672 5578 3722 5603
rect 3890 5626 3940 5655
rect 3890 5606 3907 5626
rect 3927 5606 3940 5626
rect 5672 5649 5722 5662
rect 5890 5649 5940 5662
rect 6098 5649 6148 5662
rect 3890 5578 3940 5606
rect 1308 5508 1358 5536
rect 1308 5488 1321 5508
rect 1341 5488 1358 5508
rect 1308 5459 1358 5488
rect 1526 5511 1576 5536
rect 1526 5491 1539 5511
rect 1559 5491 1576 5511
rect 1526 5459 1576 5491
rect 1734 5509 1784 5536
rect 1734 5489 1757 5509
rect 1777 5489 1784 5509
rect 1734 5459 1784 5489
rect 2667 5469 2717 5485
rect 2875 5469 2925 5485
rect 3093 5469 3143 5485
rect 7828 5638 7878 5668
rect 7828 5618 7835 5638
rect 7855 5618 7878 5638
rect 7828 5591 7878 5618
rect 8036 5636 8086 5668
rect 8036 5616 8053 5636
rect 8073 5616 8086 5636
rect 8036 5591 8086 5616
rect 8254 5639 8304 5668
rect 8254 5619 8271 5639
rect 8291 5619 8304 5639
rect 10049 5661 10099 5674
rect 10267 5661 10317 5674
rect 10475 5661 10525 5674
rect 8254 5591 8304 5619
rect 5672 5521 5722 5549
rect 5672 5501 5685 5521
rect 5705 5501 5722 5521
rect 411 5410 461 5423
rect 629 5410 679 5423
rect 837 5410 887 5423
rect 3464 5465 3514 5478
rect 3672 5465 3722 5478
rect 3890 5465 3940 5478
rect 5672 5472 5722 5501
rect 5890 5524 5940 5549
rect 5890 5504 5903 5524
rect 5923 5504 5940 5524
rect 5890 5472 5940 5504
rect 6098 5522 6148 5549
rect 6098 5502 6121 5522
rect 6141 5502 6148 5522
rect 6098 5472 6148 5502
rect 7031 5482 7081 5498
rect 7239 5482 7289 5498
rect 7457 5482 7507 5498
rect 12205 5650 12255 5680
rect 12205 5630 12212 5650
rect 12232 5630 12255 5650
rect 12205 5603 12255 5630
rect 12413 5648 12463 5680
rect 12413 5628 12430 5648
rect 12450 5628 12463 5648
rect 12413 5603 12463 5628
rect 12631 5651 12681 5680
rect 12631 5631 12648 5651
rect 12668 5631 12681 5651
rect 14413 5674 14463 5687
rect 14631 5674 14681 5687
rect 14839 5674 14889 5687
rect 12631 5603 12681 5631
rect 10049 5533 10099 5561
rect 10049 5513 10062 5533
rect 10082 5513 10099 5533
rect 1308 5401 1358 5417
rect 1526 5401 1576 5417
rect 1734 5401 1784 5417
rect 2667 5397 2717 5427
rect 2667 5377 2674 5397
rect 2694 5377 2717 5397
rect 2667 5350 2717 5377
rect 2875 5395 2925 5427
rect 2875 5375 2892 5395
rect 2912 5375 2925 5395
rect 2875 5350 2925 5375
rect 3093 5398 3143 5427
rect 3093 5378 3110 5398
rect 3130 5378 3143 5398
rect 4775 5423 4825 5436
rect 4993 5423 5043 5436
rect 5201 5423 5251 5436
rect 7828 5478 7878 5491
rect 8036 5478 8086 5491
rect 8254 5478 8304 5491
rect 10049 5484 10099 5513
rect 10267 5536 10317 5561
rect 10267 5516 10280 5536
rect 10300 5516 10317 5536
rect 10267 5484 10317 5516
rect 10475 5534 10525 5561
rect 10475 5514 10498 5534
rect 10518 5514 10525 5534
rect 10475 5484 10525 5514
rect 11408 5494 11458 5510
rect 11616 5494 11666 5510
rect 11834 5494 11884 5510
rect 16569 5663 16619 5693
rect 16569 5643 16576 5663
rect 16596 5643 16619 5663
rect 16569 5616 16619 5643
rect 16777 5661 16827 5693
rect 16777 5641 16794 5661
rect 16814 5641 16827 5661
rect 16777 5616 16827 5641
rect 16995 5664 17045 5693
rect 16995 5644 17012 5664
rect 17032 5644 17045 5664
rect 16995 5616 17045 5644
rect 14413 5546 14463 5574
rect 14413 5526 14426 5546
rect 14446 5526 14463 5546
rect 3093 5350 3143 5378
rect 411 5282 461 5310
rect 411 5262 424 5282
rect 444 5262 461 5282
rect 411 5233 461 5262
rect 629 5285 679 5310
rect 629 5265 642 5285
rect 662 5265 679 5285
rect 629 5233 679 5265
rect 837 5283 887 5310
rect 837 5263 860 5283
rect 880 5263 887 5283
rect 837 5233 887 5263
rect 5672 5414 5722 5430
rect 5890 5414 5940 5430
rect 6098 5414 6148 5430
rect 7031 5410 7081 5440
rect 7031 5390 7038 5410
rect 7058 5390 7081 5410
rect 7031 5363 7081 5390
rect 7239 5408 7289 5440
rect 7239 5388 7256 5408
rect 7276 5388 7289 5408
rect 7239 5363 7289 5388
rect 7457 5411 7507 5440
rect 7457 5391 7474 5411
rect 7494 5391 7507 5411
rect 9152 5435 9202 5448
rect 9370 5435 9420 5448
rect 9578 5435 9628 5448
rect 12205 5490 12255 5503
rect 12413 5490 12463 5503
rect 12631 5490 12681 5503
rect 14413 5497 14463 5526
rect 14631 5549 14681 5574
rect 14631 5529 14644 5549
rect 14664 5529 14681 5549
rect 14631 5497 14681 5529
rect 14839 5547 14889 5574
rect 14839 5527 14862 5547
rect 14882 5527 14889 5547
rect 14839 5497 14889 5527
rect 15772 5507 15822 5523
rect 15980 5507 16030 5523
rect 16198 5507 16248 5523
rect 7457 5363 7507 5391
rect 3465 5285 3515 5301
rect 3673 5285 3723 5301
rect 3891 5285 3941 5301
rect 1209 5226 1259 5239
rect 1427 5226 1477 5239
rect 1635 5226 1685 5239
rect 2667 5237 2717 5250
rect 2875 5237 2925 5250
rect 3093 5237 3143 5250
rect 4775 5295 4825 5323
rect 411 5175 461 5191
rect 629 5175 679 5191
rect 837 5175 887 5191
rect 3465 5213 3515 5243
rect 3465 5193 3472 5213
rect 3492 5193 3515 5213
rect 3465 5166 3515 5193
rect 3673 5211 3723 5243
rect 3673 5191 3690 5211
rect 3710 5191 3723 5211
rect 3673 5166 3723 5191
rect 3891 5214 3941 5243
rect 3891 5194 3908 5214
rect 3928 5194 3941 5214
rect 4775 5275 4788 5295
rect 4808 5275 4825 5295
rect 4775 5246 4825 5275
rect 4993 5298 5043 5323
rect 4993 5278 5006 5298
rect 5026 5278 5043 5298
rect 4993 5246 5043 5278
rect 5201 5296 5251 5323
rect 5201 5276 5224 5296
rect 5244 5276 5251 5296
rect 5201 5246 5251 5276
rect 10049 5426 10099 5442
rect 10267 5426 10317 5442
rect 10475 5426 10525 5442
rect 11408 5422 11458 5452
rect 11408 5402 11415 5422
rect 11435 5402 11458 5422
rect 11408 5375 11458 5402
rect 11616 5420 11666 5452
rect 11616 5400 11633 5420
rect 11653 5400 11666 5420
rect 11616 5375 11666 5400
rect 11834 5423 11884 5452
rect 11834 5403 11851 5423
rect 11871 5403 11884 5423
rect 13516 5448 13566 5461
rect 13734 5448 13784 5461
rect 13942 5448 13992 5461
rect 16569 5503 16619 5516
rect 16777 5503 16827 5516
rect 16995 5503 17045 5516
rect 11834 5375 11884 5403
rect 7829 5298 7879 5314
rect 8037 5298 8087 5314
rect 8255 5298 8305 5314
rect 3891 5166 3941 5194
rect 5573 5239 5623 5252
rect 5791 5239 5841 5252
rect 5999 5239 6049 5252
rect 7031 5250 7081 5263
rect 7239 5250 7289 5263
rect 7457 5250 7507 5263
rect 9152 5307 9202 5335
rect 4775 5188 4825 5204
rect 4993 5188 5043 5204
rect 5201 5188 5251 5204
rect 1209 5098 1259 5126
rect 1209 5078 1222 5098
rect 1242 5078 1259 5098
rect 1209 5049 1259 5078
rect 1427 5101 1477 5126
rect 1427 5081 1440 5101
rect 1460 5081 1477 5101
rect 1427 5049 1477 5081
rect 1635 5099 1685 5126
rect 1635 5079 1658 5099
rect 1678 5079 1685 5099
rect 1635 5049 1685 5079
rect 2363 5063 2413 5079
rect 2571 5063 2621 5079
rect 2789 5063 2839 5079
rect 7829 5226 7879 5256
rect 7829 5206 7836 5226
rect 7856 5206 7879 5226
rect 7829 5179 7879 5206
rect 8037 5224 8087 5256
rect 8037 5204 8054 5224
rect 8074 5204 8087 5224
rect 8037 5179 8087 5204
rect 8255 5227 8305 5256
rect 8255 5207 8272 5227
rect 8292 5207 8305 5227
rect 9152 5287 9165 5307
rect 9185 5287 9202 5307
rect 9152 5258 9202 5287
rect 9370 5310 9420 5335
rect 9370 5290 9383 5310
rect 9403 5290 9420 5310
rect 9370 5258 9420 5290
rect 9578 5308 9628 5335
rect 9578 5288 9601 5308
rect 9621 5288 9628 5308
rect 9578 5258 9628 5288
rect 14413 5439 14463 5455
rect 14631 5439 14681 5455
rect 14839 5439 14889 5455
rect 15772 5435 15822 5465
rect 15772 5415 15779 5435
rect 15799 5415 15822 5435
rect 15772 5388 15822 5415
rect 15980 5433 16030 5465
rect 15980 5413 15997 5433
rect 16017 5413 16030 5433
rect 15980 5388 16030 5413
rect 16198 5436 16248 5465
rect 16198 5416 16215 5436
rect 16235 5416 16248 5436
rect 16198 5388 16248 5416
rect 12206 5310 12256 5326
rect 12414 5310 12464 5326
rect 12632 5310 12682 5326
rect 8255 5179 8305 5207
rect 9950 5251 10000 5264
rect 10168 5251 10218 5264
rect 10376 5251 10426 5264
rect 11408 5262 11458 5275
rect 11616 5262 11666 5275
rect 11834 5262 11884 5275
rect 13516 5320 13566 5348
rect 9152 5200 9202 5216
rect 9370 5200 9420 5216
rect 9578 5200 9628 5216
rect 5573 5111 5623 5139
rect 412 4998 462 5011
rect 630 4998 680 5011
rect 838 4998 888 5011
rect 3465 5053 3515 5066
rect 3673 5053 3723 5066
rect 3891 5053 3941 5066
rect 5573 5091 5586 5111
rect 5606 5091 5623 5111
rect 5573 5062 5623 5091
rect 5791 5114 5841 5139
rect 5791 5094 5804 5114
rect 5824 5094 5841 5114
rect 5791 5062 5841 5094
rect 5999 5112 6049 5139
rect 5999 5092 6022 5112
rect 6042 5092 6049 5112
rect 5999 5062 6049 5092
rect 6727 5076 6777 5092
rect 6935 5076 6985 5092
rect 7153 5076 7203 5092
rect 12206 5238 12256 5268
rect 12206 5218 12213 5238
rect 12233 5218 12256 5238
rect 12206 5191 12256 5218
rect 12414 5236 12464 5268
rect 12414 5216 12431 5236
rect 12451 5216 12464 5236
rect 12414 5191 12464 5216
rect 12632 5239 12682 5268
rect 12632 5219 12649 5239
rect 12669 5219 12682 5239
rect 13516 5300 13529 5320
rect 13549 5300 13566 5320
rect 13516 5271 13566 5300
rect 13734 5323 13784 5348
rect 13734 5303 13747 5323
rect 13767 5303 13784 5323
rect 13734 5271 13784 5303
rect 13942 5321 13992 5348
rect 13942 5301 13965 5321
rect 13985 5301 13992 5321
rect 13942 5271 13992 5301
rect 16570 5323 16620 5339
rect 16778 5323 16828 5339
rect 16996 5323 17046 5339
rect 12632 5191 12682 5219
rect 14314 5264 14364 5277
rect 14532 5264 14582 5277
rect 14740 5264 14790 5277
rect 15772 5275 15822 5288
rect 15980 5275 16030 5288
rect 16198 5275 16248 5288
rect 13516 5213 13566 5229
rect 13734 5213 13784 5229
rect 13942 5213 13992 5229
rect 9950 5123 10000 5151
rect 1209 4991 1259 5007
rect 1427 4991 1477 5007
rect 1635 4991 1685 5007
rect 2363 4991 2413 5021
rect 2363 4971 2370 4991
rect 2390 4971 2413 4991
rect 2363 4944 2413 4971
rect 2571 4989 2621 5021
rect 2571 4969 2588 4989
rect 2608 4969 2621 4989
rect 2571 4944 2621 4969
rect 2789 4992 2839 5021
rect 4776 5011 4826 5024
rect 4994 5011 5044 5024
rect 5202 5011 5252 5024
rect 7829 5066 7879 5079
rect 8037 5066 8087 5079
rect 8255 5066 8305 5079
rect 9950 5103 9963 5123
rect 9983 5103 10000 5123
rect 9950 5074 10000 5103
rect 10168 5126 10218 5151
rect 10168 5106 10181 5126
rect 10201 5106 10218 5126
rect 10168 5074 10218 5106
rect 10376 5124 10426 5151
rect 10376 5104 10399 5124
rect 10419 5104 10426 5124
rect 10376 5074 10426 5104
rect 11104 5088 11154 5104
rect 11312 5088 11362 5104
rect 11530 5088 11580 5104
rect 16570 5251 16620 5281
rect 16570 5231 16577 5251
rect 16597 5231 16620 5251
rect 16570 5204 16620 5231
rect 16778 5249 16828 5281
rect 16778 5229 16795 5249
rect 16815 5229 16828 5249
rect 16778 5204 16828 5229
rect 16996 5252 17046 5281
rect 16996 5232 17013 5252
rect 17033 5232 17046 5252
rect 16996 5204 17046 5232
rect 14314 5136 14364 5164
rect 2789 4972 2806 4992
rect 2826 4972 2839 4992
rect 2789 4944 2839 4972
rect 412 4870 462 4898
rect 412 4850 425 4870
rect 445 4850 462 4870
rect 412 4821 462 4850
rect 630 4873 680 4898
rect 630 4853 643 4873
rect 663 4853 680 4873
rect 630 4821 680 4853
rect 838 4871 888 4898
rect 838 4851 861 4871
rect 881 4851 888 4871
rect 838 4821 888 4851
rect 5573 5004 5623 5020
rect 5791 5004 5841 5020
rect 5999 5004 6049 5020
rect 6727 5004 6777 5034
rect 6727 4984 6734 5004
rect 6754 4984 6777 5004
rect 6727 4957 6777 4984
rect 6935 5002 6985 5034
rect 6935 4982 6952 5002
rect 6972 4982 6985 5002
rect 6935 4957 6985 4982
rect 7153 5005 7203 5034
rect 9153 5023 9203 5036
rect 9371 5023 9421 5036
rect 9579 5023 9629 5036
rect 12206 5078 12256 5091
rect 12414 5078 12464 5091
rect 12632 5078 12682 5091
rect 14314 5116 14327 5136
rect 14347 5116 14364 5136
rect 14314 5087 14364 5116
rect 14532 5139 14582 5164
rect 14532 5119 14545 5139
rect 14565 5119 14582 5139
rect 14532 5087 14582 5119
rect 14740 5137 14790 5164
rect 14740 5117 14763 5137
rect 14783 5117 14790 5137
rect 14740 5087 14790 5117
rect 15468 5101 15518 5117
rect 15676 5101 15726 5117
rect 15894 5101 15944 5117
rect 7153 4985 7170 5005
rect 7190 4985 7203 5005
rect 7153 4957 7203 4985
rect 4776 4883 4826 4911
rect 2363 4831 2413 4844
rect 2571 4831 2621 4844
rect 2789 4831 2839 4844
rect 4776 4863 4789 4883
rect 4809 4863 4826 4883
rect 4776 4834 4826 4863
rect 4994 4886 5044 4911
rect 4994 4866 5007 4886
rect 5027 4866 5044 4886
rect 4994 4834 5044 4866
rect 5202 4884 5252 4911
rect 5202 4864 5225 4884
rect 5245 4864 5252 4884
rect 5202 4834 5252 4864
rect 9950 5016 10000 5032
rect 10168 5016 10218 5032
rect 10376 5016 10426 5032
rect 11104 5016 11154 5046
rect 11104 4996 11111 5016
rect 11131 4996 11154 5016
rect 11104 4969 11154 4996
rect 11312 5014 11362 5046
rect 11312 4994 11329 5014
rect 11349 4994 11362 5014
rect 11312 4969 11362 4994
rect 11530 5017 11580 5046
rect 13517 5036 13567 5049
rect 13735 5036 13785 5049
rect 13943 5036 13993 5049
rect 16570 5091 16620 5104
rect 16778 5091 16828 5104
rect 16996 5091 17046 5104
rect 11530 4997 11547 5017
rect 11567 4997 11580 5017
rect 11530 4969 11580 4997
rect 9153 4895 9203 4923
rect 6727 4844 6777 4857
rect 6935 4844 6985 4857
rect 7153 4844 7203 4857
rect 9153 4875 9166 4895
rect 9186 4875 9203 4895
rect 9153 4846 9203 4875
rect 9371 4898 9421 4923
rect 9371 4878 9384 4898
rect 9404 4878 9421 4898
rect 9371 4846 9421 4878
rect 9579 4896 9629 4923
rect 9579 4876 9602 4896
rect 9622 4876 9629 4896
rect 9579 4846 9629 4876
rect 14314 5029 14364 5045
rect 14532 5029 14582 5045
rect 14740 5029 14790 5045
rect 15468 5029 15518 5059
rect 15468 5009 15475 5029
rect 15495 5009 15518 5029
rect 15468 4982 15518 5009
rect 15676 5027 15726 5059
rect 15676 5007 15693 5027
rect 15713 5007 15726 5027
rect 15676 4982 15726 5007
rect 15894 5030 15944 5059
rect 15894 5010 15911 5030
rect 15931 5010 15944 5030
rect 15894 4982 15944 5010
rect 13517 4908 13567 4936
rect 11104 4856 11154 4869
rect 11312 4856 11362 4869
rect 11530 4856 11580 4869
rect 13517 4888 13530 4908
rect 13550 4888 13567 4908
rect 13517 4859 13567 4888
rect 13735 4911 13785 4936
rect 13735 4891 13748 4911
rect 13768 4891 13785 4911
rect 13735 4859 13785 4891
rect 13943 4909 13993 4936
rect 13943 4889 13966 4909
rect 13986 4889 13993 4909
rect 13943 4859 13993 4889
rect 15468 4869 15518 4882
rect 15676 4869 15726 4882
rect 15894 4869 15944 4882
rect 412 4763 462 4779
rect 630 4763 680 4779
rect 838 4763 888 4779
rect 4776 4776 4826 4792
rect 4994 4776 5044 4792
rect 5202 4776 5252 4792
rect 9153 4788 9203 4804
rect 9371 4788 9421 4804
rect 9579 4788 9629 4804
rect 13517 4801 13567 4817
rect 13735 4801 13785 4817
rect 13943 4801 13993 4817
rect 3445 4679 3495 4695
rect 3653 4679 3703 4695
rect 3871 4679 3921 4695
rect 7809 4692 7859 4708
rect 8017 4692 8067 4708
rect 8235 4692 8285 4708
rect 12186 4704 12236 4720
rect 12394 4704 12444 4720
rect 12612 4704 12662 4720
rect 16550 4717 16600 4733
rect 16758 4717 16808 4733
rect 16976 4717 17026 4733
rect 1494 4614 1544 4627
rect 1712 4614 1762 4627
rect 1920 4614 1970 4627
rect 3445 4607 3495 4637
rect 3445 4587 3452 4607
rect 3472 4587 3495 4607
rect 3445 4560 3495 4587
rect 3653 4605 3703 4637
rect 3653 4585 3670 4605
rect 3690 4585 3703 4605
rect 3653 4560 3703 4585
rect 3871 4608 3921 4637
rect 3871 4588 3888 4608
rect 3908 4588 3921 4608
rect 5858 4627 5908 4640
rect 6076 4627 6126 4640
rect 6284 4627 6334 4640
rect 3871 4560 3921 4588
rect 1494 4486 1544 4514
rect 1494 4466 1507 4486
rect 1527 4466 1544 4486
rect 1494 4437 1544 4466
rect 1712 4489 1762 4514
rect 1712 4469 1725 4489
rect 1745 4469 1762 4489
rect 1712 4437 1762 4469
rect 1920 4487 1970 4514
rect 1920 4467 1943 4487
rect 1963 4467 1970 4487
rect 1920 4437 1970 4467
rect 2648 4451 2698 4467
rect 2856 4451 2906 4467
rect 3074 4451 3124 4467
rect 7809 4620 7859 4650
rect 7809 4600 7816 4620
rect 7836 4600 7859 4620
rect 7809 4573 7859 4600
rect 8017 4618 8067 4650
rect 8017 4598 8034 4618
rect 8054 4598 8067 4618
rect 8017 4573 8067 4598
rect 8235 4621 8285 4650
rect 8235 4601 8252 4621
rect 8272 4601 8285 4621
rect 10235 4639 10285 4652
rect 10453 4639 10503 4652
rect 10661 4639 10711 4652
rect 8235 4573 8285 4601
rect 5858 4499 5908 4527
rect 5858 4479 5871 4499
rect 5891 4479 5908 4499
rect 392 4392 442 4405
rect 610 4392 660 4405
rect 818 4392 868 4405
rect 3445 4447 3495 4460
rect 3653 4447 3703 4460
rect 3871 4447 3921 4460
rect 5858 4450 5908 4479
rect 6076 4502 6126 4527
rect 6076 4482 6089 4502
rect 6109 4482 6126 4502
rect 6076 4450 6126 4482
rect 6284 4500 6334 4527
rect 6284 4480 6307 4500
rect 6327 4480 6334 4500
rect 6284 4450 6334 4480
rect 7012 4464 7062 4480
rect 7220 4464 7270 4480
rect 7438 4464 7488 4480
rect 12186 4632 12236 4662
rect 12186 4612 12193 4632
rect 12213 4612 12236 4632
rect 12186 4585 12236 4612
rect 12394 4630 12444 4662
rect 12394 4610 12411 4630
rect 12431 4610 12444 4630
rect 12394 4585 12444 4610
rect 12612 4633 12662 4662
rect 12612 4613 12629 4633
rect 12649 4613 12662 4633
rect 14599 4652 14649 4665
rect 14817 4652 14867 4665
rect 15025 4652 15075 4665
rect 12612 4585 12662 4613
rect 10235 4511 10285 4539
rect 10235 4491 10248 4511
rect 10268 4491 10285 4511
rect 1494 4379 1544 4395
rect 1712 4379 1762 4395
rect 1920 4379 1970 4395
rect 2648 4379 2698 4409
rect 2648 4359 2655 4379
rect 2675 4359 2698 4379
rect 2648 4332 2698 4359
rect 2856 4377 2906 4409
rect 2856 4357 2873 4377
rect 2893 4357 2906 4377
rect 2856 4332 2906 4357
rect 3074 4380 3124 4409
rect 3074 4360 3091 4380
rect 3111 4360 3124 4380
rect 4756 4405 4806 4418
rect 4974 4405 5024 4418
rect 5182 4405 5232 4418
rect 7809 4460 7859 4473
rect 8017 4460 8067 4473
rect 8235 4460 8285 4473
rect 10235 4462 10285 4491
rect 10453 4514 10503 4539
rect 10453 4494 10466 4514
rect 10486 4494 10503 4514
rect 10453 4462 10503 4494
rect 10661 4512 10711 4539
rect 10661 4492 10684 4512
rect 10704 4492 10711 4512
rect 10661 4462 10711 4492
rect 11389 4476 11439 4492
rect 11597 4476 11647 4492
rect 11815 4476 11865 4492
rect 16550 4645 16600 4675
rect 16550 4625 16557 4645
rect 16577 4625 16600 4645
rect 16550 4598 16600 4625
rect 16758 4643 16808 4675
rect 16758 4623 16775 4643
rect 16795 4623 16808 4643
rect 16758 4598 16808 4623
rect 16976 4646 17026 4675
rect 16976 4626 16993 4646
rect 17013 4626 17026 4646
rect 16976 4598 17026 4626
rect 14599 4524 14649 4552
rect 14599 4504 14612 4524
rect 14632 4504 14649 4524
rect 3074 4332 3124 4360
rect 392 4264 442 4292
rect 392 4244 405 4264
rect 425 4244 442 4264
rect 392 4215 442 4244
rect 610 4267 660 4292
rect 610 4247 623 4267
rect 643 4247 660 4267
rect 610 4215 660 4247
rect 818 4265 868 4292
rect 818 4245 841 4265
rect 861 4245 868 4265
rect 818 4215 868 4245
rect 5858 4392 5908 4408
rect 6076 4392 6126 4408
rect 6284 4392 6334 4408
rect 7012 4392 7062 4422
rect 7012 4372 7019 4392
rect 7039 4372 7062 4392
rect 7012 4345 7062 4372
rect 7220 4390 7270 4422
rect 7220 4370 7237 4390
rect 7257 4370 7270 4390
rect 7220 4345 7270 4370
rect 7438 4393 7488 4422
rect 7438 4373 7455 4393
rect 7475 4373 7488 4393
rect 9133 4417 9183 4430
rect 9351 4417 9401 4430
rect 9559 4417 9609 4430
rect 12186 4472 12236 4485
rect 12394 4472 12444 4485
rect 12612 4472 12662 4485
rect 14599 4475 14649 4504
rect 14817 4527 14867 4552
rect 14817 4507 14830 4527
rect 14850 4507 14867 4527
rect 14817 4475 14867 4507
rect 15025 4525 15075 4552
rect 15025 4505 15048 4525
rect 15068 4505 15075 4525
rect 15025 4475 15075 4505
rect 15753 4489 15803 4505
rect 15961 4489 16011 4505
rect 16179 4489 16229 4505
rect 7438 4345 7488 4373
rect 3446 4267 3496 4283
rect 3654 4267 3704 4283
rect 3872 4267 3922 4283
rect 1190 4208 1240 4221
rect 1408 4208 1458 4221
rect 1616 4208 1666 4221
rect 2648 4219 2698 4232
rect 2856 4219 2906 4232
rect 3074 4219 3124 4232
rect 4756 4277 4806 4305
rect 392 4157 442 4173
rect 610 4157 660 4173
rect 818 4157 868 4173
rect 3446 4195 3496 4225
rect 3446 4175 3453 4195
rect 3473 4175 3496 4195
rect 3446 4148 3496 4175
rect 3654 4193 3704 4225
rect 3654 4173 3671 4193
rect 3691 4173 3704 4193
rect 3654 4148 3704 4173
rect 3872 4196 3922 4225
rect 3872 4176 3889 4196
rect 3909 4176 3922 4196
rect 4756 4257 4769 4277
rect 4789 4257 4806 4277
rect 4756 4228 4806 4257
rect 4974 4280 5024 4305
rect 4974 4260 4987 4280
rect 5007 4260 5024 4280
rect 4974 4228 5024 4260
rect 5182 4278 5232 4305
rect 5182 4258 5205 4278
rect 5225 4258 5232 4278
rect 5182 4228 5232 4258
rect 10235 4404 10285 4420
rect 10453 4404 10503 4420
rect 10661 4404 10711 4420
rect 11389 4404 11439 4434
rect 11389 4384 11396 4404
rect 11416 4384 11439 4404
rect 11389 4357 11439 4384
rect 11597 4402 11647 4434
rect 11597 4382 11614 4402
rect 11634 4382 11647 4402
rect 11597 4357 11647 4382
rect 11815 4405 11865 4434
rect 11815 4385 11832 4405
rect 11852 4385 11865 4405
rect 13497 4430 13547 4443
rect 13715 4430 13765 4443
rect 13923 4430 13973 4443
rect 16550 4485 16600 4498
rect 16758 4485 16808 4498
rect 16976 4485 17026 4498
rect 11815 4357 11865 4385
rect 7810 4280 7860 4296
rect 8018 4280 8068 4296
rect 8236 4280 8286 4296
rect 3872 4148 3922 4176
rect 5554 4221 5604 4234
rect 5772 4221 5822 4234
rect 5980 4221 6030 4234
rect 7012 4232 7062 4245
rect 7220 4232 7270 4245
rect 7438 4232 7488 4245
rect 9133 4289 9183 4317
rect 4756 4170 4806 4186
rect 4974 4170 5024 4186
rect 5182 4170 5232 4186
rect 1190 4080 1240 4108
rect 1190 4060 1203 4080
rect 1223 4060 1240 4080
rect 1190 4031 1240 4060
rect 1408 4083 1458 4108
rect 1408 4063 1421 4083
rect 1441 4063 1458 4083
rect 1408 4031 1458 4063
rect 1616 4081 1666 4108
rect 1616 4061 1639 4081
rect 1659 4061 1666 4081
rect 1616 4031 1666 4061
rect 2549 4041 2599 4057
rect 2757 4041 2807 4057
rect 2975 4041 3025 4057
rect 7810 4208 7860 4238
rect 7810 4188 7817 4208
rect 7837 4188 7860 4208
rect 7810 4161 7860 4188
rect 8018 4206 8068 4238
rect 8018 4186 8035 4206
rect 8055 4186 8068 4206
rect 8018 4161 8068 4186
rect 8236 4209 8286 4238
rect 8236 4189 8253 4209
rect 8273 4189 8286 4209
rect 9133 4269 9146 4289
rect 9166 4269 9183 4289
rect 9133 4240 9183 4269
rect 9351 4292 9401 4317
rect 9351 4272 9364 4292
rect 9384 4272 9401 4292
rect 9351 4240 9401 4272
rect 9559 4290 9609 4317
rect 9559 4270 9582 4290
rect 9602 4270 9609 4290
rect 9559 4240 9609 4270
rect 14599 4417 14649 4433
rect 14817 4417 14867 4433
rect 15025 4417 15075 4433
rect 15753 4417 15803 4447
rect 15753 4397 15760 4417
rect 15780 4397 15803 4417
rect 15753 4370 15803 4397
rect 15961 4415 16011 4447
rect 15961 4395 15978 4415
rect 15998 4395 16011 4415
rect 15961 4370 16011 4395
rect 16179 4418 16229 4447
rect 16179 4398 16196 4418
rect 16216 4398 16229 4418
rect 16179 4370 16229 4398
rect 12187 4292 12237 4308
rect 12395 4292 12445 4308
rect 12613 4292 12663 4308
rect 8236 4161 8286 4189
rect 9931 4233 9981 4246
rect 10149 4233 10199 4246
rect 10357 4233 10407 4246
rect 11389 4244 11439 4257
rect 11597 4244 11647 4257
rect 11815 4244 11865 4257
rect 13497 4302 13547 4330
rect 9133 4182 9183 4198
rect 9351 4182 9401 4198
rect 9559 4182 9609 4198
rect 5554 4093 5604 4121
rect 393 3980 443 3993
rect 611 3980 661 3993
rect 819 3980 869 3993
rect 3446 4035 3496 4048
rect 3654 4035 3704 4048
rect 3872 4035 3922 4048
rect 5554 4073 5567 4093
rect 5587 4073 5604 4093
rect 5554 4044 5604 4073
rect 5772 4096 5822 4121
rect 5772 4076 5785 4096
rect 5805 4076 5822 4096
rect 5772 4044 5822 4076
rect 5980 4094 6030 4121
rect 5980 4074 6003 4094
rect 6023 4074 6030 4094
rect 5980 4044 6030 4074
rect 6913 4054 6963 4070
rect 7121 4054 7171 4070
rect 7339 4054 7389 4070
rect 12187 4220 12237 4250
rect 12187 4200 12194 4220
rect 12214 4200 12237 4220
rect 12187 4173 12237 4200
rect 12395 4218 12445 4250
rect 12395 4198 12412 4218
rect 12432 4198 12445 4218
rect 12395 4173 12445 4198
rect 12613 4221 12663 4250
rect 12613 4201 12630 4221
rect 12650 4201 12663 4221
rect 13497 4282 13510 4302
rect 13530 4282 13547 4302
rect 13497 4253 13547 4282
rect 13715 4305 13765 4330
rect 13715 4285 13728 4305
rect 13748 4285 13765 4305
rect 13715 4253 13765 4285
rect 13923 4303 13973 4330
rect 13923 4283 13946 4303
rect 13966 4283 13973 4303
rect 13923 4253 13973 4283
rect 16551 4305 16601 4321
rect 16759 4305 16809 4321
rect 16977 4305 17027 4321
rect 12613 4173 12663 4201
rect 14295 4246 14345 4259
rect 14513 4246 14563 4259
rect 14721 4246 14771 4259
rect 15753 4257 15803 4270
rect 15961 4257 16011 4270
rect 16179 4257 16229 4270
rect 13497 4195 13547 4211
rect 13715 4195 13765 4211
rect 13923 4195 13973 4211
rect 9931 4105 9981 4133
rect 1190 3973 1240 3989
rect 1408 3973 1458 3989
rect 1616 3973 1666 3989
rect 2549 3969 2599 3999
rect 2549 3949 2556 3969
rect 2576 3949 2599 3969
rect 2549 3922 2599 3949
rect 2757 3967 2807 3999
rect 2757 3947 2774 3967
rect 2794 3947 2807 3967
rect 2757 3922 2807 3947
rect 2975 3970 3025 3999
rect 4757 3993 4807 4006
rect 4975 3993 5025 4006
rect 5183 3993 5233 4006
rect 7810 4048 7860 4061
rect 8018 4048 8068 4061
rect 8236 4048 8286 4061
rect 9931 4085 9944 4105
rect 9964 4085 9981 4105
rect 9931 4056 9981 4085
rect 10149 4108 10199 4133
rect 10149 4088 10162 4108
rect 10182 4088 10199 4108
rect 10149 4056 10199 4088
rect 10357 4106 10407 4133
rect 10357 4086 10380 4106
rect 10400 4086 10407 4106
rect 10357 4056 10407 4086
rect 11290 4066 11340 4082
rect 11498 4066 11548 4082
rect 11716 4066 11766 4082
rect 16551 4233 16601 4263
rect 16551 4213 16558 4233
rect 16578 4213 16601 4233
rect 16551 4186 16601 4213
rect 16759 4231 16809 4263
rect 16759 4211 16776 4231
rect 16796 4211 16809 4231
rect 16759 4186 16809 4211
rect 16977 4234 17027 4263
rect 16977 4214 16994 4234
rect 17014 4214 17027 4234
rect 16977 4186 17027 4214
rect 14295 4118 14345 4146
rect 2975 3950 2992 3970
rect 3012 3950 3025 3970
rect 2975 3922 3025 3950
rect 393 3852 443 3880
rect 393 3832 406 3852
rect 426 3832 443 3852
rect 393 3803 443 3832
rect 611 3855 661 3880
rect 611 3835 624 3855
rect 644 3835 661 3855
rect 611 3803 661 3835
rect 819 3853 869 3880
rect 819 3833 842 3853
rect 862 3833 869 3853
rect 819 3803 869 3833
rect 5554 3986 5604 4002
rect 5772 3986 5822 4002
rect 5980 3986 6030 4002
rect 6913 3982 6963 4012
rect 6913 3962 6920 3982
rect 6940 3962 6963 3982
rect 6913 3935 6963 3962
rect 7121 3980 7171 4012
rect 7121 3960 7138 3980
rect 7158 3960 7171 3980
rect 7121 3935 7171 3960
rect 7339 3983 7389 4012
rect 9134 4005 9184 4018
rect 9352 4005 9402 4018
rect 9560 4005 9610 4018
rect 12187 4060 12237 4073
rect 12395 4060 12445 4073
rect 12613 4060 12663 4073
rect 14295 4098 14308 4118
rect 14328 4098 14345 4118
rect 14295 4069 14345 4098
rect 14513 4121 14563 4146
rect 14513 4101 14526 4121
rect 14546 4101 14563 4121
rect 14513 4069 14563 4101
rect 14721 4119 14771 4146
rect 14721 4099 14744 4119
rect 14764 4099 14771 4119
rect 14721 4069 14771 4099
rect 15654 4079 15704 4095
rect 15862 4079 15912 4095
rect 16080 4079 16130 4095
rect 7339 3963 7356 3983
rect 7376 3963 7389 3983
rect 7339 3935 7389 3963
rect 4757 3865 4807 3893
rect 2549 3809 2599 3822
rect 2757 3809 2807 3822
rect 2975 3809 3025 3822
rect 4757 3845 4770 3865
rect 4790 3845 4807 3865
rect 4757 3816 4807 3845
rect 4975 3868 5025 3893
rect 4975 3848 4988 3868
rect 5008 3848 5025 3868
rect 4975 3816 5025 3848
rect 5183 3866 5233 3893
rect 5183 3846 5206 3866
rect 5226 3846 5233 3866
rect 5183 3816 5233 3846
rect 9931 3998 9981 4014
rect 10149 3998 10199 4014
rect 10357 3998 10407 4014
rect 11290 3994 11340 4024
rect 11290 3974 11297 3994
rect 11317 3974 11340 3994
rect 11290 3947 11340 3974
rect 11498 3992 11548 4024
rect 11498 3972 11515 3992
rect 11535 3972 11548 3992
rect 11498 3947 11548 3972
rect 11716 3995 11766 4024
rect 13498 4018 13548 4031
rect 13716 4018 13766 4031
rect 13924 4018 13974 4031
rect 16551 4073 16601 4086
rect 16759 4073 16809 4086
rect 16977 4073 17027 4086
rect 11716 3975 11733 3995
rect 11753 3975 11766 3995
rect 11716 3947 11766 3975
rect 9134 3877 9184 3905
rect 6913 3822 6963 3835
rect 7121 3822 7171 3835
rect 7339 3822 7389 3835
rect 9134 3857 9147 3877
rect 9167 3857 9184 3877
rect 9134 3828 9184 3857
rect 9352 3880 9402 3905
rect 9352 3860 9365 3880
rect 9385 3860 9402 3880
rect 9352 3828 9402 3860
rect 9560 3878 9610 3905
rect 9560 3858 9583 3878
rect 9603 3858 9610 3878
rect 9560 3828 9610 3858
rect 14295 4011 14345 4027
rect 14513 4011 14563 4027
rect 14721 4011 14771 4027
rect 15654 4007 15704 4037
rect 15654 3987 15661 4007
rect 15681 3987 15704 4007
rect 15654 3960 15704 3987
rect 15862 4005 15912 4037
rect 15862 3985 15879 4005
rect 15899 3985 15912 4005
rect 15862 3960 15912 3985
rect 16080 4008 16130 4037
rect 16080 3988 16097 4008
rect 16117 3988 16130 4008
rect 16080 3960 16130 3988
rect 13498 3890 13548 3918
rect 11290 3834 11340 3847
rect 11498 3834 11548 3847
rect 11716 3834 11766 3847
rect 13498 3870 13511 3890
rect 13531 3870 13548 3890
rect 13498 3841 13548 3870
rect 13716 3893 13766 3918
rect 13716 3873 13729 3893
rect 13749 3873 13766 3893
rect 13716 3841 13766 3873
rect 13924 3891 13974 3918
rect 13924 3871 13947 3891
rect 13967 3871 13974 3891
rect 13924 3841 13974 3871
rect 15654 3847 15704 3860
rect 15862 3847 15912 3860
rect 16080 3847 16130 3860
rect 393 3745 443 3761
rect 611 3745 661 3761
rect 819 3745 869 3761
rect 4757 3758 4807 3774
rect 4975 3758 5025 3774
rect 5183 3758 5233 3774
rect 9134 3770 9184 3786
rect 9352 3770 9402 3786
rect 9560 3770 9610 3786
rect 13498 3783 13548 3799
rect 13716 3783 13766 3799
rect 13924 3783 13974 3799
rect 3428 3661 3478 3677
rect 3636 3661 3686 3677
rect 3854 3661 3904 3677
rect 7792 3674 7842 3690
rect 8000 3674 8050 3690
rect 8218 3674 8268 3690
rect 12169 3686 12219 3702
rect 12377 3686 12427 3702
rect 12595 3686 12645 3702
rect 16533 3699 16583 3715
rect 16741 3699 16791 3715
rect 16959 3699 17009 3715
rect 1272 3600 1322 3613
rect 1490 3600 1540 3613
rect 1698 3600 1748 3613
rect 3428 3589 3478 3619
rect 3428 3569 3435 3589
rect 3455 3569 3478 3589
rect 3428 3542 3478 3569
rect 3636 3587 3686 3619
rect 3636 3567 3653 3587
rect 3673 3567 3686 3587
rect 3636 3542 3686 3567
rect 3854 3590 3904 3619
rect 3854 3570 3871 3590
rect 3891 3570 3904 3590
rect 5636 3613 5686 3626
rect 5854 3613 5904 3626
rect 6062 3613 6112 3626
rect 3854 3542 3904 3570
rect 1272 3472 1322 3500
rect 1272 3452 1285 3472
rect 1305 3452 1322 3472
rect 1272 3423 1322 3452
rect 1490 3475 1540 3500
rect 1490 3455 1503 3475
rect 1523 3455 1540 3475
rect 1490 3423 1540 3455
rect 1698 3473 1748 3500
rect 1698 3453 1721 3473
rect 1741 3453 1748 3473
rect 1698 3423 1748 3453
rect 2631 3433 2681 3449
rect 2839 3433 2889 3449
rect 3057 3433 3107 3449
rect 7792 3602 7842 3632
rect 7792 3582 7799 3602
rect 7819 3582 7842 3602
rect 7792 3555 7842 3582
rect 8000 3600 8050 3632
rect 8000 3580 8017 3600
rect 8037 3580 8050 3600
rect 8000 3555 8050 3580
rect 8218 3603 8268 3632
rect 8218 3583 8235 3603
rect 8255 3583 8268 3603
rect 10013 3625 10063 3638
rect 10231 3625 10281 3638
rect 10439 3625 10489 3638
rect 8218 3555 8268 3583
rect 5636 3485 5686 3513
rect 5636 3465 5649 3485
rect 5669 3465 5686 3485
rect 375 3374 425 3387
rect 593 3374 643 3387
rect 801 3374 851 3387
rect 3428 3429 3478 3442
rect 3636 3429 3686 3442
rect 3854 3429 3904 3442
rect 5636 3436 5686 3465
rect 5854 3488 5904 3513
rect 5854 3468 5867 3488
rect 5887 3468 5904 3488
rect 5854 3436 5904 3468
rect 6062 3486 6112 3513
rect 6062 3466 6085 3486
rect 6105 3466 6112 3486
rect 6062 3436 6112 3466
rect 6995 3446 7045 3462
rect 7203 3446 7253 3462
rect 7421 3446 7471 3462
rect 12169 3614 12219 3644
rect 12169 3594 12176 3614
rect 12196 3594 12219 3614
rect 12169 3567 12219 3594
rect 12377 3612 12427 3644
rect 12377 3592 12394 3612
rect 12414 3592 12427 3612
rect 12377 3567 12427 3592
rect 12595 3615 12645 3644
rect 12595 3595 12612 3615
rect 12632 3595 12645 3615
rect 14377 3638 14427 3651
rect 14595 3638 14645 3651
rect 14803 3638 14853 3651
rect 12595 3567 12645 3595
rect 10013 3497 10063 3525
rect 10013 3477 10026 3497
rect 10046 3477 10063 3497
rect 1272 3365 1322 3381
rect 1490 3365 1540 3381
rect 1698 3365 1748 3381
rect 2631 3361 2681 3391
rect 2631 3341 2638 3361
rect 2658 3341 2681 3361
rect 2631 3314 2681 3341
rect 2839 3359 2889 3391
rect 2839 3339 2856 3359
rect 2876 3339 2889 3359
rect 2839 3314 2889 3339
rect 3057 3362 3107 3391
rect 3057 3342 3074 3362
rect 3094 3342 3107 3362
rect 4739 3387 4789 3400
rect 4957 3387 5007 3400
rect 5165 3387 5215 3400
rect 7792 3442 7842 3455
rect 8000 3442 8050 3455
rect 8218 3442 8268 3455
rect 10013 3448 10063 3477
rect 10231 3500 10281 3525
rect 10231 3480 10244 3500
rect 10264 3480 10281 3500
rect 10231 3448 10281 3480
rect 10439 3498 10489 3525
rect 10439 3478 10462 3498
rect 10482 3478 10489 3498
rect 10439 3448 10489 3478
rect 11372 3458 11422 3474
rect 11580 3458 11630 3474
rect 11798 3458 11848 3474
rect 16533 3627 16583 3657
rect 16533 3607 16540 3627
rect 16560 3607 16583 3627
rect 16533 3580 16583 3607
rect 16741 3625 16791 3657
rect 16741 3605 16758 3625
rect 16778 3605 16791 3625
rect 16741 3580 16791 3605
rect 16959 3628 17009 3657
rect 16959 3608 16976 3628
rect 16996 3608 17009 3628
rect 16959 3580 17009 3608
rect 14377 3510 14427 3538
rect 14377 3490 14390 3510
rect 14410 3490 14427 3510
rect 3057 3314 3107 3342
rect 375 3246 425 3274
rect 375 3226 388 3246
rect 408 3226 425 3246
rect 375 3197 425 3226
rect 593 3249 643 3274
rect 593 3229 606 3249
rect 626 3229 643 3249
rect 593 3197 643 3229
rect 801 3247 851 3274
rect 801 3227 824 3247
rect 844 3227 851 3247
rect 801 3197 851 3227
rect 5636 3378 5686 3394
rect 5854 3378 5904 3394
rect 6062 3378 6112 3394
rect 6995 3374 7045 3404
rect 6995 3354 7002 3374
rect 7022 3354 7045 3374
rect 6995 3327 7045 3354
rect 7203 3372 7253 3404
rect 7203 3352 7220 3372
rect 7240 3352 7253 3372
rect 7203 3327 7253 3352
rect 7421 3375 7471 3404
rect 7421 3355 7438 3375
rect 7458 3355 7471 3375
rect 9116 3399 9166 3412
rect 9334 3399 9384 3412
rect 9542 3399 9592 3412
rect 12169 3454 12219 3467
rect 12377 3454 12427 3467
rect 12595 3454 12645 3467
rect 14377 3461 14427 3490
rect 14595 3513 14645 3538
rect 14595 3493 14608 3513
rect 14628 3493 14645 3513
rect 14595 3461 14645 3493
rect 14803 3511 14853 3538
rect 14803 3491 14826 3511
rect 14846 3491 14853 3511
rect 14803 3461 14853 3491
rect 15736 3471 15786 3487
rect 15944 3471 15994 3487
rect 16162 3471 16212 3487
rect 7421 3327 7471 3355
rect 3429 3249 3479 3265
rect 3637 3249 3687 3265
rect 3855 3249 3905 3265
rect 1173 3190 1223 3203
rect 1391 3190 1441 3203
rect 1599 3190 1649 3203
rect 2631 3201 2681 3214
rect 2839 3201 2889 3214
rect 3057 3201 3107 3214
rect 4739 3259 4789 3287
rect 375 3139 425 3155
rect 593 3139 643 3155
rect 801 3139 851 3155
rect 3429 3177 3479 3207
rect 3429 3157 3436 3177
rect 3456 3157 3479 3177
rect 3429 3130 3479 3157
rect 3637 3175 3687 3207
rect 3637 3155 3654 3175
rect 3674 3155 3687 3175
rect 3637 3130 3687 3155
rect 3855 3178 3905 3207
rect 3855 3158 3872 3178
rect 3892 3158 3905 3178
rect 4739 3239 4752 3259
rect 4772 3239 4789 3259
rect 4739 3210 4789 3239
rect 4957 3262 5007 3287
rect 4957 3242 4970 3262
rect 4990 3242 5007 3262
rect 4957 3210 5007 3242
rect 5165 3260 5215 3287
rect 5165 3240 5188 3260
rect 5208 3240 5215 3260
rect 5165 3210 5215 3240
rect 10013 3390 10063 3406
rect 10231 3390 10281 3406
rect 10439 3390 10489 3406
rect 11372 3386 11422 3416
rect 11372 3366 11379 3386
rect 11399 3366 11422 3386
rect 11372 3339 11422 3366
rect 11580 3384 11630 3416
rect 11580 3364 11597 3384
rect 11617 3364 11630 3384
rect 11580 3339 11630 3364
rect 11798 3387 11848 3416
rect 11798 3367 11815 3387
rect 11835 3367 11848 3387
rect 13480 3412 13530 3425
rect 13698 3412 13748 3425
rect 13906 3412 13956 3425
rect 16533 3467 16583 3480
rect 16741 3467 16791 3480
rect 16959 3467 17009 3480
rect 11798 3339 11848 3367
rect 7793 3262 7843 3278
rect 8001 3262 8051 3278
rect 8219 3262 8269 3278
rect 3855 3130 3905 3158
rect 5537 3203 5587 3216
rect 5755 3203 5805 3216
rect 5963 3203 6013 3216
rect 6995 3214 7045 3227
rect 7203 3214 7253 3227
rect 7421 3214 7471 3227
rect 9116 3271 9166 3299
rect 4739 3152 4789 3168
rect 4957 3152 5007 3168
rect 5165 3152 5215 3168
rect 1173 3062 1223 3090
rect 1173 3042 1186 3062
rect 1206 3042 1223 3062
rect 1173 3013 1223 3042
rect 1391 3065 1441 3090
rect 1391 3045 1404 3065
rect 1424 3045 1441 3065
rect 1391 3013 1441 3045
rect 1599 3063 1649 3090
rect 1599 3043 1622 3063
rect 1642 3043 1649 3063
rect 1599 3013 1649 3043
rect 2466 3025 2516 3041
rect 2674 3025 2724 3041
rect 2892 3025 2942 3041
rect 7793 3190 7843 3220
rect 7793 3170 7800 3190
rect 7820 3170 7843 3190
rect 7793 3143 7843 3170
rect 8001 3188 8051 3220
rect 8001 3168 8018 3188
rect 8038 3168 8051 3188
rect 8001 3143 8051 3168
rect 8219 3191 8269 3220
rect 8219 3171 8236 3191
rect 8256 3171 8269 3191
rect 9116 3251 9129 3271
rect 9149 3251 9166 3271
rect 9116 3222 9166 3251
rect 9334 3274 9384 3299
rect 9334 3254 9347 3274
rect 9367 3254 9384 3274
rect 9334 3222 9384 3254
rect 9542 3272 9592 3299
rect 9542 3252 9565 3272
rect 9585 3252 9592 3272
rect 9542 3222 9592 3252
rect 14377 3403 14427 3419
rect 14595 3403 14645 3419
rect 14803 3403 14853 3419
rect 15736 3399 15786 3429
rect 15736 3379 15743 3399
rect 15763 3379 15786 3399
rect 15736 3352 15786 3379
rect 15944 3397 15994 3429
rect 15944 3377 15961 3397
rect 15981 3377 15994 3397
rect 15944 3352 15994 3377
rect 16162 3400 16212 3429
rect 16162 3380 16179 3400
rect 16199 3380 16212 3400
rect 16162 3352 16212 3380
rect 12170 3274 12220 3290
rect 12378 3274 12428 3290
rect 12596 3274 12646 3290
rect 8219 3143 8269 3171
rect 9914 3215 9964 3228
rect 10132 3215 10182 3228
rect 10340 3215 10390 3228
rect 11372 3226 11422 3239
rect 11580 3226 11630 3239
rect 11798 3226 11848 3239
rect 13480 3284 13530 3312
rect 9116 3164 9166 3180
rect 9334 3164 9384 3180
rect 9542 3164 9592 3180
rect 5537 3075 5587 3103
rect 376 2962 426 2975
rect 594 2962 644 2975
rect 802 2962 852 2975
rect 3429 3017 3479 3030
rect 3637 3017 3687 3030
rect 3855 3017 3905 3030
rect 5537 3055 5550 3075
rect 5570 3055 5587 3075
rect 5537 3026 5587 3055
rect 5755 3078 5805 3103
rect 5755 3058 5768 3078
rect 5788 3058 5805 3078
rect 5755 3026 5805 3058
rect 5963 3076 6013 3103
rect 5963 3056 5986 3076
rect 6006 3056 6013 3076
rect 5963 3026 6013 3056
rect 6830 3038 6880 3054
rect 7038 3038 7088 3054
rect 7256 3038 7306 3054
rect 12170 3202 12220 3232
rect 12170 3182 12177 3202
rect 12197 3182 12220 3202
rect 12170 3155 12220 3182
rect 12378 3200 12428 3232
rect 12378 3180 12395 3200
rect 12415 3180 12428 3200
rect 12378 3155 12428 3180
rect 12596 3203 12646 3232
rect 12596 3183 12613 3203
rect 12633 3183 12646 3203
rect 13480 3264 13493 3284
rect 13513 3264 13530 3284
rect 13480 3235 13530 3264
rect 13698 3287 13748 3312
rect 13698 3267 13711 3287
rect 13731 3267 13748 3287
rect 13698 3235 13748 3267
rect 13906 3285 13956 3312
rect 13906 3265 13929 3285
rect 13949 3265 13956 3285
rect 13906 3235 13956 3265
rect 16534 3287 16584 3303
rect 16742 3287 16792 3303
rect 16960 3287 17010 3303
rect 12596 3155 12646 3183
rect 14278 3228 14328 3241
rect 14496 3228 14546 3241
rect 14704 3228 14754 3241
rect 15736 3239 15786 3252
rect 15944 3239 15994 3252
rect 16162 3239 16212 3252
rect 13480 3177 13530 3193
rect 13698 3177 13748 3193
rect 13906 3177 13956 3193
rect 9914 3087 9964 3115
rect 1173 2955 1223 2971
rect 1391 2955 1441 2971
rect 1599 2955 1649 2971
rect 2466 2953 2516 2983
rect 2466 2933 2473 2953
rect 2493 2933 2516 2953
rect 2466 2906 2516 2933
rect 2674 2951 2724 2983
rect 2674 2931 2691 2951
rect 2711 2931 2724 2951
rect 2674 2906 2724 2931
rect 2892 2954 2942 2983
rect 4740 2975 4790 2988
rect 4958 2975 5008 2988
rect 5166 2975 5216 2988
rect 7793 3030 7843 3043
rect 8001 3030 8051 3043
rect 8219 3030 8269 3043
rect 9914 3067 9927 3087
rect 9947 3067 9964 3087
rect 9914 3038 9964 3067
rect 10132 3090 10182 3115
rect 10132 3070 10145 3090
rect 10165 3070 10182 3090
rect 10132 3038 10182 3070
rect 10340 3088 10390 3115
rect 10340 3068 10363 3088
rect 10383 3068 10390 3088
rect 10340 3038 10390 3068
rect 11207 3050 11257 3066
rect 11415 3050 11465 3066
rect 11633 3050 11683 3066
rect 16534 3215 16584 3245
rect 16534 3195 16541 3215
rect 16561 3195 16584 3215
rect 16534 3168 16584 3195
rect 16742 3213 16792 3245
rect 16742 3193 16759 3213
rect 16779 3193 16792 3213
rect 16742 3168 16792 3193
rect 16960 3216 17010 3245
rect 16960 3196 16977 3216
rect 16997 3196 17010 3216
rect 16960 3168 17010 3196
rect 14278 3100 14328 3128
rect 2892 2934 2909 2954
rect 2929 2934 2942 2954
rect 2892 2906 2942 2934
rect 376 2834 426 2862
rect 376 2814 389 2834
rect 409 2814 426 2834
rect 376 2785 426 2814
rect 594 2837 644 2862
rect 594 2817 607 2837
rect 627 2817 644 2837
rect 594 2785 644 2817
rect 802 2835 852 2862
rect 802 2815 825 2835
rect 845 2815 852 2835
rect 802 2785 852 2815
rect 5537 2968 5587 2984
rect 5755 2968 5805 2984
rect 5963 2968 6013 2984
rect 6830 2966 6880 2996
rect 6830 2946 6837 2966
rect 6857 2946 6880 2966
rect 6830 2919 6880 2946
rect 7038 2964 7088 2996
rect 7038 2944 7055 2964
rect 7075 2944 7088 2964
rect 7038 2919 7088 2944
rect 7256 2967 7306 2996
rect 9117 2987 9167 3000
rect 9335 2987 9385 3000
rect 9543 2987 9593 3000
rect 12170 3042 12220 3055
rect 12378 3042 12428 3055
rect 12596 3042 12646 3055
rect 14278 3080 14291 3100
rect 14311 3080 14328 3100
rect 14278 3051 14328 3080
rect 14496 3103 14546 3128
rect 14496 3083 14509 3103
rect 14529 3083 14546 3103
rect 14496 3051 14546 3083
rect 14704 3101 14754 3128
rect 14704 3081 14727 3101
rect 14747 3081 14754 3101
rect 14704 3051 14754 3081
rect 15571 3063 15621 3079
rect 15779 3063 15829 3079
rect 15997 3063 16047 3079
rect 7256 2947 7273 2967
rect 7293 2947 7306 2967
rect 7256 2919 7306 2947
rect 4740 2847 4790 2875
rect 2466 2793 2516 2806
rect 2674 2793 2724 2806
rect 2892 2793 2942 2806
rect 4740 2827 4753 2847
rect 4773 2827 4790 2847
rect 4740 2798 4790 2827
rect 4958 2850 5008 2875
rect 4958 2830 4971 2850
rect 4991 2830 5008 2850
rect 4958 2798 5008 2830
rect 5166 2848 5216 2875
rect 5166 2828 5189 2848
rect 5209 2828 5216 2848
rect 5166 2798 5216 2828
rect 9914 2980 9964 2996
rect 10132 2980 10182 2996
rect 10340 2980 10390 2996
rect 11207 2978 11257 3008
rect 11207 2958 11214 2978
rect 11234 2958 11257 2978
rect 11207 2931 11257 2958
rect 11415 2976 11465 3008
rect 11415 2956 11432 2976
rect 11452 2956 11465 2976
rect 11415 2931 11465 2956
rect 11633 2979 11683 3008
rect 13481 3000 13531 3013
rect 13699 3000 13749 3013
rect 13907 3000 13957 3013
rect 16534 3055 16584 3068
rect 16742 3055 16792 3068
rect 16960 3055 17010 3068
rect 11633 2959 11650 2979
rect 11670 2959 11683 2979
rect 11633 2931 11683 2959
rect 9117 2859 9167 2887
rect 6830 2806 6880 2819
rect 7038 2806 7088 2819
rect 7256 2806 7306 2819
rect 9117 2839 9130 2859
rect 9150 2839 9167 2859
rect 9117 2810 9167 2839
rect 9335 2862 9385 2887
rect 9335 2842 9348 2862
rect 9368 2842 9385 2862
rect 9335 2810 9385 2842
rect 9543 2860 9593 2887
rect 9543 2840 9566 2860
rect 9586 2840 9593 2860
rect 9543 2810 9593 2840
rect 14278 2993 14328 3009
rect 14496 2993 14546 3009
rect 14704 2993 14754 3009
rect 15571 2991 15621 3021
rect 15571 2971 15578 2991
rect 15598 2971 15621 2991
rect 15571 2944 15621 2971
rect 15779 2989 15829 3021
rect 15779 2969 15796 2989
rect 15816 2969 15829 2989
rect 15779 2944 15829 2969
rect 15997 2992 16047 3021
rect 15997 2972 16014 2992
rect 16034 2972 16047 2992
rect 15997 2944 16047 2972
rect 13481 2872 13531 2900
rect 11207 2818 11257 2831
rect 11415 2818 11465 2831
rect 11633 2818 11683 2831
rect 13481 2852 13494 2872
rect 13514 2852 13531 2872
rect 13481 2823 13531 2852
rect 13699 2875 13749 2900
rect 13699 2855 13712 2875
rect 13732 2855 13749 2875
rect 13699 2823 13749 2855
rect 13907 2873 13957 2900
rect 13907 2853 13930 2873
rect 13950 2853 13957 2873
rect 13907 2823 13957 2853
rect 15571 2831 15621 2844
rect 15779 2831 15829 2844
rect 15997 2831 16047 2844
rect 376 2727 426 2743
rect 594 2727 644 2743
rect 802 2727 852 2743
rect 4740 2740 4790 2756
rect 4958 2740 5008 2756
rect 5166 2740 5216 2756
rect 9117 2752 9167 2768
rect 9335 2752 9385 2768
rect 9543 2752 9593 2768
rect 13481 2765 13531 2781
rect 13699 2765 13749 2781
rect 13907 2765 13957 2781
rect 3408 2643 3458 2659
rect 3616 2643 3666 2659
rect 3834 2643 3884 2659
rect 7772 2656 7822 2672
rect 7980 2656 8030 2672
rect 8198 2656 8248 2672
rect 12149 2668 12199 2684
rect 12357 2668 12407 2684
rect 12575 2668 12625 2684
rect 16513 2681 16563 2697
rect 16721 2681 16771 2697
rect 16939 2681 16989 2697
rect 1318 2580 1368 2593
rect 1536 2580 1586 2593
rect 1744 2580 1794 2593
rect 3408 2571 3458 2601
rect 3408 2551 3415 2571
rect 3435 2551 3458 2571
rect 3408 2524 3458 2551
rect 3616 2569 3666 2601
rect 3616 2549 3633 2569
rect 3653 2549 3666 2569
rect 3616 2524 3666 2549
rect 3834 2572 3884 2601
rect 3834 2552 3851 2572
rect 3871 2552 3884 2572
rect 5682 2593 5732 2606
rect 5900 2593 5950 2606
rect 6108 2593 6158 2606
rect 3834 2524 3884 2552
rect 1318 2452 1368 2480
rect 1318 2432 1331 2452
rect 1351 2432 1368 2452
rect 1318 2403 1368 2432
rect 1536 2455 1586 2480
rect 1536 2435 1549 2455
rect 1569 2435 1586 2455
rect 1536 2403 1586 2435
rect 1744 2453 1794 2480
rect 1744 2433 1767 2453
rect 1787 2433 1794 2453
rect 1744 2403 1794 2433
rect 2611 2415 2661 2431
rect 2819 2415 2869 2431
rect 3037 2415 3087 2431
rect 7772 2584 7822 2614
rect 7772 2564 7779 2584
rect 7799 2564 7822 2584
rect 7772 2537 7822 2564
rect 7980 2582 8030 2614
rect 7980 2562 7997 2582
rect 8017 2562 8030 2582
rect 7980 2537 8030 2562
rect 8198 2585 8248 2614
rect 8198 2565 8215 2585
rect 8235 2565 8248 2585
rect 10059 2605 10109 2618
rect 10277 2605 10327 2618
rect 10485 2605 10535 2618
rect 8198 2537 8248 2565
rect 5682 2465 5732 2493
rect 5682 2445 5695 2465
rect 5715 2445 5732 2465
rect 355 2356 405 2369
rect 573 2356 623 2369
rect 781 2356 831 2369
rect 3408 2411 3458 2424
rect 3616 2411 3666 2424
rect 3834 2411 3884 2424
rect 5682 2416 5732 2445
rect 5900 2468 5950 2493
rect 5900 2448 5913 2468
rect 5933 2448 5950 2468
rect 5900 2416 5950 2448
rect 6108 2466 6158 2493
rect 6108 2446 6131 2466
rect 6151 2446 6158 2466
rect 6108 2416 6158 2446
rect 6975 2428 7025 2444
rect 7183 2428 7233 2444
rect 7401 2428 7451 2444
rect 12149 2596 12199 2626
rect 12149 2576 12156 2596
rect 12176 2576 12199 2596
rect 12149 2549 12199 2576
rect 12357 2594 12407 2626
rect 12357 2574 12374 2594
rect 12394 2574 12407 2594
rect 12357 2549 12407 2574
rect 12575 2597 12625 2626
rect 12575 2577 12592 2597
rect 12612 2577 12625 2597
rect 14423 2618 14473 2631
rect 14641 2618 14691 2631
rect 14849 2618 14899 2631
rect 12575 2549 12625 2577
rect 10059 2477 10109 2505
rect 10059 2457 10072 2477
rect 10092 2457 10109 2477
rect 1318 2345 1368 2361
rect 1536 2345 1586 2361
rect 1744 2345 1794 2361
rect 2611 2343 2661 2373
rect 2611 2323 2618 2343
rect 2638 2323 2661 2343
rect 2611 2296 2661 2323
rect 2819 2341 2869 2373
rect 2819 2321 2836 2341
rect 2856 2321 2869 2341
rect 2819 2296 2869 2321
rect 3037 2344 3087 2373
rect 3037 2324 3054 2344
rect 3074 2324 3087 2344
rect 4719 2369 4769 2382
rect 4937 2369 4987 2382
rect 5145 2369 5195 2382
rect 7772 2424 7822 2437
rect 7980 2424 8030 2437
rect 8198 2424 8248 2437
rect 10059 2428 10109 2457
rect 10277 2480 10327 2505
rect 10277 2460 10290 2480
rect 10310 2460 10327 2480
rect 10277 2428 10327 2460
rect 10485 2478 10535 2505
rect 10485 2458 10508 2478
rect 10528 2458 10535 2478
rect 10485 2428 10535 2458
rect 11352 2440 11402 2456
rect 11560 2440 11610 2456
rect 11778 2440 11828 2456
rect 16513 2609 16563 2639
rect 16513 2589 16520 2609
rect 16540 2589 16563 2609
rect 16513 2562 16563 2589
rect 16721 2607 16771 2639
rect 16721 2587 16738 2607
rect 16758 2587 16771 2607
rect 16721 2562 16771 2587
rect 16939 2610 16989 2639
rect 16939 2590 16956 2610
rect 16976 2590 16989 2610
rect 16939 2562 16989 2590
rect 14423 2490 14473 2518
rect 14423 2470 14436 2490
rect 14456 2470 14473 2490
rect 3037 2296 3087 2324
rect 355 2228 405 2256
rect 355 2208 368 2228
rect 388 2208 405 2228
rect 355 2179 405 2208
rect 573 2231 623 2256
rect 573 2211 586 2231
rect 606 2211 623 2231
rect 573 2179 623 2211
rect 781 2229 831 2256
rect 781 2209 804 2229
rect 824 2209 831 2229
rect 781 2179 831 2209
rect 5682 2358 5732 2374
rect 5900 2358 5950 2374
rect 6108 2358 6158 2374
rect 6975 2356 7025 2386
rect 6975 2336 6982 2356
rect 7002 2336 7025 2356
rect 6975 2309 7025 2336
rect 7183 2354 7233 2386
rect 7183 2334 7200 2354
rect 7220 2334 7233 2354
rect 7183 2309 7233 2334
rect 7401 2357 7451 2386
rect 7401 2337 7418 2357
rect 7438 2337 7451 2357
rect 9096 2381 9146 2394
rect 9314 2381 9364 2394
rect 9522 2381 9572 2394
rect 12149 2436 12199 2449
rect 12357 2436 12407 2449
rect 12575 2436 12625 2449
rect 14423 2441 14473 2470
rect 14641 2493 14691 2518
rect 14641 2473 14654 2493
rect 14674 2473 14691 2493
rect 14641 2441 14691 2473
rect 14849 2491 14899 2518
rect 14849 2471 14872 2491
rect 14892 2471 14899 2491
rect 14849 2441 14899 2471
rect 15716 2453 15766 2469
rect 15924 2453 15974 2469
rect 16142 2453 16192 2469
rect 7401 2309 7451 2337
rect 3409 2231 3459 2247
rect 3617 2231 3667 2247
rect 3835 2231 3885 2247
rect 1153 2172 1203 2185
rect 1371 2172 1421 2185
rect 1579 2172 1629 2185
rect 2611 2183 2661 2196
rect 2819 2183 2869 2196
rect 3037 2183 3087 2196
rect 4719 2241 4769 2269
rect 355 2121 405 2137
rect 573 2121 623 2137
rect 781 2121 831 2137
rect 3409 2159 3459 2189
rect 3409 2139 3416 2159
rect 3436 2139 3459 2159
rect 3409 2112 3459 2139
rect 3617 2157 3667 2189
rect 3617 2137 3634 2157
rect 3654 2137 3667 2157
rect 3617 2112 3667 2137
rect 3835 2160 3885 2189
rect 3835 2140 3852 2160
rect 3872 2140 3885 2160
rect 4719 2221 4732 2241
rect 4752 2221 4769 2241
rect 4719 2192 4769 2221
rect 4937 2244 4987 2269
rect 4937 2224 4950 2244
rect 4970 2224 4987 2244
rect 4937 2192 4987 2224
rect 5145 2242 5195 2269
rect 5145 2222 5168 2242
rect 5188 2222 5195 2242
rect 5145 2192 5195 2222
rect 10059 2370 10109 2386
rect 10277 2370 10327 2386
rect 10485 2370 10535 2386
rect 11352 2368 11402 2398
rect 11352 2348 11359 2368
rect 11379 2348 11402 2368
rect 11352 2321 11402 2348
rect 11560 2366 11610 2398
rect 11560 2346 11577 2366
rect 11597 2346 11610 2366
rect 11560 2321 11610 2346
rect 11778 2369 11828 2398
rect 11778 2349 11795 2369
rect 11815 2349 11828 2369
rect 13460 2394 13510 2407
rect 13678 2394 13728 2407
rect 13886 2394 13936 2407
rect 16513 2449 16563 2462
rect 16721 2449 16771 2462
rect 16939 2449 16989 2462
rect 11778 2321 11828 2349
rect 7773 2244 7823 2260
rect 7981 2244 8031 2260
rect 8199 2244 8249 2260
rect 3835 2112 3885 2140
rect 5517 2185 5567 2198
rect 5735 2185 5785 2198
rect 5943 2185 5993 2198
rect 6975 2196 7025 2209
rect 7183 2196 7233 2209
rect 7401 2196 7451 2209
rect 9096 2253 9146 2281
rect 4719 2134 4769 2150
rect 4937 2134 4987 2150
rect 5145 2134 5195 2150
rect 1153 2044 1203 2072
rect 1153 2024 1166 2044
rect 1186 2024 1203 2044
rect 1153 1995 1203 2024
rect 1371 2047 1421 2072
rect 1371 2027 1384 2047
rect 1404 2027 1421 2047
rect 1371 1995 1421 2027
rect 1579 2045 1629 2072
rect 1579 2025 1602 2045
rect 1622 2025 1629 2045
rect 1579 1995 1629 2025
rect 2512 2005 2562 2021
rect 2720 2005 2770 2021
rect 2938 2005 2988 2021
rect 7773 2172 7823 2202
rect 7773 2152 7780 2172
rect 7800 2152 7823 2172
rect 7773 2125 7823 2152
rect 7981 2170 8031 2202
rect 7981 2150 7998 2170
rect 8018 2150 8031 2170
rect 7981 2125 8031 2150
rect 8199 2173 8249 2202
rect 8199 2153 8216 2173
rect 8236 2153 8249 2173
rect 9096 2233 9109 2253
rect 9129 2233 9146 2253
rect 9096 2204 9146 2233
rect 9314 2256 9364 2281
rect 9314 2236 9327 2256
rect 9347 2236 9364 2256
rect 9314 2204 9364 2236
rect 9522 2254 9572 2281
rect 9522 2234 9545 2254
rect 9565 2234 9572 2254
rect 9522 2204 9572 2234
rect 14423 2383 14473 2399
rect 14641 2383 14691 2399
rect 14849 2383 14899 2399
rect 15716 2381 15766 2411
rect 15716 2361 15723 2381
rect 15743 2361 15766 2381
rect 15716 2334 15766 2361
rect 15924 2379 15974 2411
rect 15924 2359 15941 2379
rect 15961 2359 15974 2379
rect 15924 2334 15974 2359
rect 16142 2382 16192 2411
rect 16142 2362 16159 2382
rect 16179 2362 16192 2382
rect 16142 2334 16192 2362
rect 12150 2256 12200 2272
rect 12358 2256 12408 2272
rect 12576 2256 12626 2272
rect 8199 2125 8249 2153
rect 9894 2197 9944 2210
rect 10112 2197 10162 2210
rect 10320 2197 10370 2210
rect 11352 2208 11402 2221
rect 11560 2208 11610 2221
rect 11778 2208 11828 2221
rect 13460 2266 13510 2294
rect 9096 2146 9146 2162
rect 9314 2146 9364 2162
rect 9522 2146 9572 2162
rect 5517 2057 5567 2085
rect 356 1944 406 1957
rect 574 1944 624 1957
rect 782 1944 832 1957
rect 3409 1999 3459 2012
rect 3617 1999 3667 2012
rect 3835 1999 3885 2012
rect 5517 2037 5530 2057
rect 5550 2037 5567 2057
rect 5517 2008 5567 2037
rect 5735 2060 5785 2085
rect 5735 2040 5748 2060
rect 5768 2040 5785 2060
rect 5735 2008 5785 2040
rect 5943 2058 5993 2085
rect 5943 2038 5966 2058
rect 5986 2038 5993 2058
rect 5943 2008 5993 2038
rect 6876 2018 6926 2034
rect 7084 2018 7134 2034
rect 7302 2018 7352 2034
rect 12150 2184 12200 2214
rect 12150 2164 12157 2184
rect 12177 2164 12200 2184
rect 12150 2137 12200 2164
rect 12358 2182 12408 2214
rect 12358 2162 12375 2182
rect 12395 2162 12408 2182
rect 12358 2137 12408 2162
rect 12576 2185 12626 2214
rect 12576 2165 12593 2185
rect 12613 2165 12626 2185
rect 13460 2246 13473 2266
rect 13493 2246 13510 2266
rect 13460 2217 13510 2246
rect 13678 2269 13728 2294
rect 13678 2249 13691 2269
rect 13711 2249 13728 2269
rect 13678 2217 13728 2249
rect 13886 2267 13936 2294
rect 13886 2247 13909 2267
rect 13929 2247 13936 2267
rect 13886 2217 13936 2247
rect 16514 2269 16564 2285
rect 16722 2269 16772 2285
rect 16940 2269 16990 2285
rect 12576 2137 12626 2165
rect 14258 2210 14308 2223
rect 14476 2210 14526 2223
rect 14684 2210 14734 2223
rect 15716 2221 15766 2234
rect 15924 2221 15974 2234
rect 16142 2221 16192 2234
rect 13460 2159 13510 2175
rect 13678 2159 13728 2175
rect 13886 2159 13936 2175
rect 9894 2069 9944 2097
rect 1153 1937 1203 1953
rect 1371 1937 1421 1953
rect 1579 1937 1629 1953
rect 2512 1933 2562 1963
rect 2512 1913 2519 1933
rect 2539 1913 2562 1933
rect 2512 1886 2562 1913
rect 2720 1931 2770 1963
rect 2720 1911 2737 1931
rect 2757 1911 2770 1931
rect 2720 1886 2770 1911
rect 2938 1934 2988 1963
rect 4720 1957 4770 1970
rect 4938 1957 4988 1970
rect 5146 1957 5196 1970
rect 7773 2012 7823 2025
rect 7981 2012 8031 2025
rect 8199 2012 8249 2025
rect 9894 2049 9907 2069
rect 9927 2049 9944 2069
rect 9894 2020 9944 2049
rect 10112 2072 10162 2097
rect 10112 2052 10125 2072
rect 10145 2052 10162 2072
rect 10112 2020 10162 2052
rect 10320 2070 10370 2097
rect 10320 2050 10343 2070
rect 10363 2050 10370 2070
rect 10320 2020 10370 2050
rect 11253 2030 11303 2046
rect 11461 2030 11511 2046
rect 11679 2030 11729 2046
rect 16514 2197 16564 2227
rect 16514 2177 16521 2197
rect 16541 2177 16564 2197
rect 16514 2150 16564 2177
rect 16722 2195 16772 2227
rect 16722 2175 16739 2195
rect 16759 2175 16772 2195
rect 16722 2150 16772 2175
rect 16940 2198 16990 2227
rect 16940 2178 16957 2198
rect 16977 2178 16990 2198
rect 16940 2150 16990 2178
rect 14258 2082 14308 2110
rect 2938 1914 2955 1934
rect 2975 1914 2988 1934
rect 2938 1886 2988 1914
rect 356 1816 406 1844
rect 356 1796 369 1816
rect 389 1796 406 1816
rect 356 1767 406 1796
rect 574 1819 624 1844
rect 574 1799 587 1819
rect 607 1799 624 1819
rect 574 1767 624 1799
rect 782 1817 832 1844
rect 782 1797 805 1817
rect 825 1797 832 1817
rect 782 1767 832 1797
rect 5517 1950 5567 1966
rect 5735 1950 5785 1966
rect 5943 1950 5993 1966
rect 6876 1946 6926 1976
rect 6876 1926 6883 1946
rect 6903 1926 6926 1946
rect 6876 1899 6926 1926
rect 7084 1944 7134 1976
rect 7084 1924 7101 1944
rect 7121 1924 7134 1944
rect 7084 1899 7134 1924
rect 7302 1947 7352 1976
rect 9097 1969 9147 1982
rect 9315 1969 9365 1982
rect 9523 1969 9573 1982
rect 12150 2024 12200 2037
rect 12358 2024 12408 2037
rect 12576 2024 12626 2037
rect 14258 2062 14271 2082
rect 14291 2062 14308 2082
rect 14258 2033 14308 2062
rect 14476 2085 14526 2110
rect 14476 2065 14489 2085
rect 14509 2065 14526 2085
rect 14476 2033 14526 2065
rect 14684 2083 14734 2110
rect 14684 2063 14707 2083
rect 14727 2063 14734 2083
rect 14684 2033 14734 2063
rect 15617 2043 15667 2059
rect 15825 2043 15875 2059
rect 16043 2043 16093 2059
rect 7302 1927 7319 1947
rect 7339 1927 7352 1947
rect 7302 1899 7352 1927
rect 4720 1829 4770 1857
rect 2512 1773 2562 1786
rect 2720 1773 2770 1786
rect 2938 1773 2988 1786
rect 4720 1809 4733 1829
rect 4753 1809 4770 1829
rect 4720 1780 4770 1809
rect 4938 1832 4988 1857
rect 4938 1812 4951 1832
rect 4971 1812 4988 1832
rect 4938 1780 4988 1812
rect 5146 1830 5196 1857
rect 5146 1810 5169 1830
rect 5189 1810 5196 1830
rect 5146 1780 5196 1810
rect 9894 1962 9944 1978
rect 10112 1962 10162 1978
rect 10320 1962 10370 1978
rect 11253 1958 11303 1988
rect 11253 1938 11260 1958
rect 11280 1938 11303 1958
rect 11253 1911 11303 1938
rect 11461 1956 11511 1988
rect 11461 1936 11478 1956
rect 11498 1936 11511 1956
rect 11461 1911 11511 1936
rect 11679 1959 11729 1988
rect 13461 1982 13511 1995
rect 13679 1982 13729 1995
rect 13887 1982 13937 1995
rect 16514 2037 16564 2050
rect 16722 2037 16772 2050
rect 16940 2037 16990 2050
rect 11679 1939 11696 1959
rect 11716 1939 11729 1959
rect 11679 1911 11729 1939
rect 9097 1841 9147 1869
rect 6876 1786 6926 1799
rect 7084 1786 7134 1799
rect 7302 1786 7352 1799
rect 9097 1821 9110 1841
rect 9130 1821 9147 1841
rect 9097 1792 9147 1821
rect 9315 1844 9365 1869
rect 9315 1824 9328 1844
rect 9348 1824 9365 1844
rect 9315 1792 9365 1824
rect 9523 1842 9573 1869
rect 9523 1822 9546 1842
rect 9566 1822 9573 1842
rect 9523 1792 9573 1822
rect 14258 1975 14308 1991
rect 14476 1975 14526 1991
rect 14684 1975 14734 1991
rect 15617 1971 15667 2001
rect 15617 1951 15624 1971
rect 15644 1951 15667 1971
rect 15617 1924 15667 1951
rect 15825 1969 15875 2001
rect 15825 1949 15842 1969
rect 15862 1949 15875 1969
rect 15825 1924 15875 1949
rect 16043 1972 16093 2001
rect 16043 1952 16060 1972
rect 16080 1952 16093 1972
rect 16043 1924 16093 1952
rect 13461 1854 13511 1882
rect 11253 1798 11303 1811
rect 11461 1798 11511 1811
rect 11679 1798 11729 1811
rect 13461 1834 13474 1854
rect 13494 1834 13511 1854
rect 13461 1805 13511 1834
rect 13679 1857 13729 1882
rect 13679 1837 13692 1857
rect 13712 1837 13729 1857
rect 13679 1805 13729 1837
rect 13887 1855 13937 1882
rect 13887 1835 13910 1855
rect 13930 1835 13937 1855
rect 13887 1805 13937 1835
rect 15617 1811 15667 1824
rect 15825 1811 15875 1824
rect 16043 1811 16093 1824
rect 356 1709 406 1725
rect 574 1709 624 1725
rect 782 1709 832 1725
rect 4720 1722 4770 1738
rect 4938 1722 4988 1738
rect 5146 1722 5196 1738
rect 9097 1734 9147 1750
rect 9315 1734 9365 1750
rect 9523 1734 9573 1750
rect 13461 1747 13511 1763
rect 13679 1747 13729 1763
rect 13887 1747 13937 1763
rect 3391 1625 3441 1641
rect 3599 1625 3649 1641
rect 3817 1625 3867 1641
rect 7755 1638 7805 1654
rect 7963 1638 8013 1654
rect 8181 1638 8231 1654
rect 12132 1650 12182 1666
rect 12340 1650 12390 1666
rect 12558 1650 12608 1666
rect 16496 1663 16546 1679
rect 16704 1663 16754 1679
rect 16922 1663 16972 1679
rect 1235 1564 1285 1577
rect 1453 1564 1503 1577
rect 1661 1564 1711 1577
rect 3391 1553 3441 1583
rect 3391 1533 3398 1553
rect 3418 1533 3441 1553
rect 3391 1506 3441 1533
rect 3599 1551 3649 1583
rect 3599 1531 3616 1551
rect 3636 1531 3649 1551
rect 3599 1506 3649 1531
rect 3817 1554 3867 1583
rect 3817 1534 3834 1554
rect 3854 1534 3867 1554
rect 5599 1577 5649 1590
rect 5817 1577 5867 1590
rect 6025 1577 6075 1590
rect 3817 1506 3867 1534
rect 1235 1436 1285 1464
rect 1235 1416 1248 1436
rect 1268 1416 1285 1436
rect 1235 1387 1285 1416
rect 1453 1439 1503 1464
rect 1453 1419 1466 1439
rect 1486 1419 1503 1439
rect 1453 1387 1503 1419
rect 1661 1437 1711 1464
rect 1661 1417 1684 1437
rect 1704 1417 1711 1437
rect 1661 1387 1711 1417
rect 2594 1397 2644 1413
rect 2802 1397 2852 1413
rect 3020 1397 3070 1413
rect 7755 1566 7805 1596
rect 7755 1546 7762 1566
rect 7782 1546 7805 1566
rect 7755 1519 7805 1546
rect 7963 1564 8013 1596
rect 7963 1544 7980 1564
rect 8000 1544 8013 1564
rect 7963 1519 8013 1544
rect 8181 1567 8231 1596
rect 8181 1547 8198 1567
rect 8218 1547 8231 1567
rect 9976 1589 10026 1602
rect 10194 1589 10244 1602
rect 10402 1589 10452 1602
rect 8181 1519 8231 1547
rect 5599 1449 5649 1477
rect 5599 1429 5612 1449
rect 5632 1429 5649 1449
rect 338 1338 388 1351
rect 556 1338 606 1351
rect 764 1338 814 1351
rect 3391 1393 3441 1406
rect 3599 1393 3649 1406
rect 3817 1393 3867 1406
rect 5599 1400 5649 1429
rect 5817 1452 5867 1477
rect 5817 1432 5830 1452
rect 5850 1432 5867 1452
rect 5817 1400 5867 1432
rect 6025 1450 6075 1477
rect 6025 1430 6048 1450
rect 6068 1430 6075 1450
rect 6025 1400 6075 1430
rect 6958 1410 7008 1426
rect 7166 1410 7216 1426
rect 7384 1410 7434 1426
rect 12132 1578 12182 1608
rect 12132 1558 12139 1578
rect 12159 1558 12182 1578
rect 12132 1531 12182 1558
rect 12340 1576 12390 1608
rect 12340 1556 12357 1576
rect 12377 1556 12390 1576
rect 12340 1531 12390 1556
rect 12558 1579 12608 1608
rect 12558 1559 12575 1579
rect 12595 1559 12608 1579
rect 14340 1602 14390 1615
rect 14558 1602 14608 1615
rect 14766 1602 14816 1615
rect 12558 1531 12608 1559
rect 9976 1461 10026 1489
rect 9976 1441 9989 1461
rect 10009 1441 10026 1461
rect 1235 1329 1285 1345
rect 1453 1329 1503 1345
rect 1661 1329 1711 1345
rect 2594 1325 2644 1355
rect 2594 1305 2601 1325
rect 2621 1305 2644 1325
rect 2594 1278 2644 1305
rect 2802 1323 2852 1355
rect 2802 1303 2819 1323
rect 2839 1303 2852 1323
rect 2802 1278 2852 1303
rect 3020 1326 3070 1355
rect 3020 1306 3037 1326
rect 3057 1306 3070 1326
rect 4702 1351 4752 1364
rect 4920 1351 4970 1364
rect 5128 1351 5178 1364
rect 7755 1406 7805 1419
rect 7963 1406 8013 1419
rect 8181 1406 8231 1419
rect 9976 1412 10026 1441
rect 10194 1464 10244 1489
rect 10194 1444 10207 1464
rect 10227 1444 10244 1464
rect 10194 1412 10244 1444
rect 10402 1462 10452 1489
rect 10402 1442 10425 1462
rect 10445 1442 10452 1462
rect 10402 1412 10452 1442
rect 11335 1422 11385 1438
rect 11543 1422 11593 1438
rect 11761 1422 11811 1438
rect 16496 1591 16546 1621
rect 16496 1571 16503 1591
rect 16523 1571 16546 1591
rect 16496 1544 16546 1571
rect 16704 1589 16754 1621
rect 16704 1569 16721 1589
rect 16741 1569 16754 1589
rect 16704 1544 16754 1569
rect 16922 1592 16972 1621
rect 16922 1572 16939 1592
rect 16959 1572 16972 1592
rect 16922 1544 16972 1572
rect 14340 1474 14390 1502
rect 14340 1454 14353 1474
rect 14373 1454 14390 1474
rect 3020 1278 3070 1306
rect 338 1210 388 1238
rect 338 1190 351 1210
rect 371 1190 388 1210
rect 338 1161 388 1190
rect 556 1213 606 1238
rect 556 1193 569 1213
rect 589 1193 606 1213
rect 556 1161 606 1193
rect 764 1211 814 1238
rect 764 1191 787 1211
rect 807 1191 814 1211
rect 764 1161 814 1191
rect 5599 1342 5649 1358
rect 5817 1342 5867 1358
rect 6025 1342 6075 1358
rect 6958 1338 7008 1368
rect 6958 1318 6965 1338
rect 6985 1318 7008 1338
rect 6958 1291 7008 1318
rect 7166 1336 7216 1368
rect 7166 1316 7183 1336
rect 7203 1316 7216 1336
rect 7166 1291 7216 1316
rect 7384 1339 7434 1368
rect 7384 1319 7401 1339
rect 7421 1319 7434 1339
rect 9079 1363 9129 1376
rect 9297 1363 9347 1376
rect 9505 1363 9555 1376
rect 12132 1418 12182 1431
rect 12340 1418 12390 1431
rect 12558 1418 12608 1431
rect 14340 1425 14390 1454
rect 14558 1477 14608 1502
rect 14558 1457 14571 1477
rect 14591 1457 14608 1477
rect 14558 1425 14608 1457
rect 14766 1475 14816 1502
rect 14766 1455 14789 1475
rect 14809 1455 14816 1475
rect 14766 1425 14816 1455
rect 15699 1435 15749 1451
rect 15907 1435 15957 1451
rect 16125 1435 16175 1451
rect 7384 1291 7434 1319
rect 3392 1213 3442 1229
rect 3600 1213 3650 1229
rect 3818 1213 3868 1229
rect 1136 1154 1186 1167
rect 1354 1154 1404 1167
rect 1562 1154 1612 1167
rect 2594 1165 2644 1178
rect 2802 1165 2852 1178
rect 3020 1165 3070 1178
rect 4702 1223 4752 1251
rect 338 1103 388 1119
rect 556 1103 606 1119
rect 764 1103 814 1119
rect 3392 1141 3442 1171
rect 3392 1121 3399 1141
rect 3419 1121 3442 1141
rect 3392 1094 3442 1121
rect 3600 1139 3650 1171
rect 3600 1119 3617 1139
rect 3637 1119 3650 1139
rect 3600 1094 3650 1119
rect 3818 1142 3868 1171
rect 3818 1122 3835 1142
rect 3855 1122 3868 1142
rect 4702 1203 4715 1223
rect 4735 1203 4752 1223
rect 4702 1174 4752 1203
rect 4920 1226 4970 1251
rect 4920 1206 4933 1226
rect 4953 1206 4970 1226
rect 4920 1174 4970 1206
rect 5128 1224 5178 1251
rect 5128 1204 5151 1224
rect 5171 1204 5178 1224
rect 5128 1174 5178 1204
rect 9976 1354 10026 1370
rect 10194 1354 10244 1370
rect 10402 1354 10452 1370
rect 11335 1350 11385 1380
rect 11335 1330 11342 1350
rect 11362 1330 11385 1350
rect 11335 1303 11385 1330
rect 11543 1348 11593 1380
rect 11543 1328 11560 1348
rect 11580 1328 11593 1348
rect 11543 1303 11593 1328
rect 11761 1351 11811 1380
rect 11761 1331 11778 1351
rect 11798 1331 11811 1351
rect 13443 1376 13493 1389
rect 13661 1376 13711 1389
rect 13869 1376 13919 1389
rect 16496 1431 16546 1444
rect 16704 1431 16754 1444
rect 16922 1431 16972 1444
rect 11761 1303 11811 1331
rect 7756 1226 7806 1242
rect 7964 1226 8014 1242
rect 8182 1226 8232 1242
rect 3818 1094 3868 1122
rect 5500 1167 5550 1180
rect 5718 1167 5768 1180
rect 5926 1167 5976 1180
rect 6958 1178 7008 1191
rect 7166 1178 7216 1191
rect 7384 1178 7434 1191
rect 9079 1235 9129 1263
rect 4702 1116 4752 1132
rect 4920 1116 4970 1132
rect 5128 1116 5178 1132
rect 1136 1026 1186 1054
rect 1136 1006 1149 1026
rect 1169 1006 1186 1026
rect 1136 977 1186 1006
rect 1354 1029 1404 1054
rect 1354 1009 1367 1029
rect 1387 1009 1404 1029
rect 1354 977 1404 1009
rect 1562 1027 1612 1054
rect 1562 1007 1585 1027
rect 1605 1007 1612 1027
rect 1562 977 1612 1007
rect 7756 1154 7806 1184
rect 7756 1134 7763 1154
rect 7783 1134 7806 1154
rect 7756 1107 7806 1134
rect 7964 1152 8014 1184
rect 7964 1132 7981 1152
rect 8001 1132 8014 1152
rect 7964 1107 8014 1132
rect 8182 1155 8232 1184
rect 8182 1135 8199 1155
rect 8219 1135 8232 1155
rect 9079 1215 9092 1235
rect 9112 1215 9129 1235
rect 9079 1186 9129 1215
rect 9297 1238 9347 1263
rect 9297 1218 9310 1238
rect 9330 1218 9347 1238
rect 9297 1186 9347 1218
rect 9505 1236 9555 1263
rect 9505 1216 9528 1236
rect 9548 1216 9555 1236
rect 9505 1186 9555 1216
rect 14340 1367 14390 1383
rect 14558 1367 14608 1383
rect 14766 1367 14816 1383
rect 15699 1363 15749 1393
rect 15699 1343 15706 1363
rect 15726 1343 15749 1363
rect 15699 1316 15749 1343
rect 15907 1361 15957 1393
rect 15907 1341 15924 1361
rect 15944 1341 15957 1361
rect 15907 1316 15957 1341
rect 16125 1364 16175 1393
rect 16125 1344 16142 1364
rect 16162 1344 16175 1364
rect 16125 1316 16175 1344
rect 12133 1238 12183 1254
rect 12341 1238 12391 1254
rect 12559 1238 12609 1254
rect 8182 1107 8232 1135
rect 9877 1179 9927 1192
rect 10095 1179 10145 1192
rect 10303 1179 10353 1192
rect 11335 1190 11385 1203
rect 11543 1190 11593 1203
rect 11761 1190 11811 1203
rect 13443 1248 13493 1276
rect 9079 1128 9129 1144
rect 9297 1128 9347 1144
rect 9505 1128 9555 1144
rect 5500 1039 5550 1067
rect 3392 981 3442 994
rect 3600 981 3650 994
rect 3818 981 3868 994
rect 5500 1019 5513 1039
rect 5533 1019 5550 1039
rect 5500 990 5550 1019
rect 5718 1042 5768 1067
rect 5718 1022 5731 1042
rect 5751 1022 5768 1042
rect 5718 990 5768 1022
rect 5926 1040 5976 1067
rect 5926 1020 5949 1040
rect 5969 1020 5976 1040
rect 5926 990 5976 1020
rect 12133 1166 12183 1196
rect 12133 1146 12140 1166
rect 12160 1146 12183 1166
rect 12133 1119 12183 1146
rect 12341 1164 12391 1196
rect 12341 1144 12358 1164
rect 12378 1144 12391 1164
rect 12341 1119 12391 1144
rect 12559 1167 12609 1196
rect 12559 1147 12576 1167
rect 12596 1147 12609 1167
rect 13443 1228 13456 1248
rect 13476 1228 13493 1248
rect 13443 1199 13493 1228
rect 13661 1251 13711 1276
rect 13661 1231 13674 1251
rect 13694 1231 13711 1251
rect 13661 1199 13711 1231
rect 13869 1249 13919 1276
rect 13869 1229 13892 1249
rect 13912 1229 13919 1249
rect 13869 1199 13919 1229
rect 16497 1251 16547 1267
rect 16705 1251 16755 1267
rect 16923 1251 16973 1267
rect 12559 1119 12609 1147
rect 14241 1192 14291 1205
rect 14459 1192 14509 1205
rect 14667 1192 14717 1205
rect 15699 1203 15749 1216
rect 15907 1203 15957 1216
rect 16125 1203 16175 1216
rect 13443 1141 13493 1157
rect 13661 1141 13711 1157
rect 13869 1141 13919 1157
rect 9877 1051 9927 1079
rect 7756 994 7806 1007
rect 7964 994 8014 1007
rect 8182 994 8232 1007
rect 9877 1031 9890 1051
rect 9910 1031 9927 1051
rect 9877 1002 9927 1031
rect 10095 1054 10145 1079
rect 10095 1034 10108 1054
rect 10128 1034 10145 1054
rect 10095 1002 10145 1034
rect 10303 1052 10353 1079
rect 10303 1032 10326 1052
rect 10346 1032 10353 1052
rect 10303 1002 10353 1032
rect 16497 1179 16547 1209
rect 16497 1159 16504 1179
rect 16524 1159 16547 1179
rect 16497 1132 16547 1159
rect 16705 1177 16755 1209
rect 16705 1157 16722 1177
rect 16742 1157 16755 1177
rect 16705 1132 16755 1157
rect 16923 1180 16973 1209
rect 16923 1160 16940 1180
rect 16960 1160 16973 1180
rect 16923 1132 16973 1160
rect 14241 1064 14291 1092
rect 12133 1006 12183 1019
rect 12341 1006 12391 1019
rect 12559 1006 12609 1019
rect 14241 1044 14254 1064
rect 14274 1044 14291 1064
rect 14241 1015 14291 1044
rect 14459 1067 14509 1092
rect 14459 1047 14472 1067
rect 14492 1047 14509 1067
rect 14459 1015 14509 1047
rect 14667 1065 14717 1092
rect 14667 1045 14690 1065
rect 14710 1045 14717 1065
rect 14667 1015 14717 1045
rect 16497 1019 16547 1032
rect 16705 1019 16755 1032
rect 16923 1019 16973 1032
rect 339 926 389 939
rect 557 926 607 939
rect 765 926 815 939
rect 1136 919 1186 935
rect 1354 919 1404 935
rect 1562 919 1612 935
rect 4703 939 4753 952
rect 4921 939 4971 952
rect 5129 939 5179 952
rect 339 798 389 826
rect 339 778 352 798
rect 372 778 389 798
rect 339 749 389 778
rect 557 801 607 826
rect 557 781 570 801
rect 590 781 607 801
rect 557 749 607 781
rect 765 799 815 826
rect 5500 932 5550 948
rect 5718 932 5768 948
rect 5926 932 5976 948
rect 9080 951 9130 964
rect 9298 951 9348 964
rect 9506 951 9556 964
rect 765 779 788 799
rect 808 779 815 799
rect 765 749 815 779
rect 4703 811 4753 839
rect 4703 791 4716 811
rect 4736 791 4753 811
rect 4703 762 4753 791
rect 4921 814 4971 839
rect 4921 794 4934 814
rect 4954 794 4971 814
rect 4921 762 4971 794
rect 5129 812 5179 839
rect 9877 944 9927 960
rect 10095 944 10145 960
rect 10303 944 10353 960
rect 13444 964 13494 977
rect 13662 964 13712 977
rect 13870 964 13920 977
rect 5129 792 5152 812
rect 5172 792 5179 812
rect 5129 762 5179 792
rect 9080 823 9130 851
rect 9080 803 9093 823
rect 9113 803 9130 823
rect 9080 774 9130 803
rect 9298 826 9348 851
rect 9298 806 9311 826
rect 9331 806 9348 826
rect 9298 774 9348 806
rect 9506 824 9556 851
rect 14241 957 14291 973
rect 14459 957 14509 973
rect 14667 957 14717 973
rect 9506 804 9529 824
rect 9549 804 9556 824
rect 9506 774 9556 804
rect 13444 836 13494 864
rect 13444 816 13457 836
rect 13477 816 13494 836
rect 13444 787 13494 816
rect 13662 839 13712 864
rect 13662 819 13675 839
rect 13695 819 13712 839
rect 13662 787 13712 819
rect 13870 837 13920 864
rect 13870 817 13893 837
rect 13913 817 13920 837
rect 13870 787 13920 817
rect 339 691 389 707
rect 557 691 607 707
rect 765 691 815 707
rect 4703 704 4753 720
rect 4921 704 4971 720
rect 5129 704 5179 720
rect 9080 716 9130 732
rect 9298 716 9348 732
rect 9506 716 9556 732
rect 13444 729 13494 745
rect 13662 729 13712 745
rect 13870 729 13920 745
rect 14657 388 14707 401
rect 14875 388 14925 401
rect 15083 388 15133 401
rect 5916 363 5966 376
rect 6134 363 6184 376
rect 6342 363 6392 376
rect 10293 375 10343 388
rect 10511 375 10561 388
rect 10719 375 10769 388
rect 1552 350 1602 363
rect 1770 350 1820 363
rect 1978 350 2028 363
rect 4041 276 4091 289
rect 4259 276 4309 289
rect 4467 276 4517 289
rect 1552 222 1602 250
rect 1552 202 1565 222
rect 1585 202 1602 222
rect 1552 173 1602 202
rect 1770 225 1820 250
rect 1770 205 1783 225
rect 1803 205 1820 225
rect 1770 173 1820 205
rect 1978 223 2028 250
rect 1978 203 2001 223
rect 2021 203 2028 223
rect 1978 173 2028 203
rect 8489 300 8539 313
rect 8707 300 8757 313
rect 8915 300 8965 313
rect 5916 235 5966 263
rect 5916 215 5929 235
rect 5949 215 5966 235
rect 5916 186 5966 215
rect 6134 238 6184 263
rect 6134 218 6147 238
rect 6167 218 6184 238
rect 6134 186 6184 218
rect 6342 236 6392 263
rect 6342 216 6365 236
rect 6385 216 6392 236
rect 6342 186 6392 216
rect 12782 301 12832 314
rect 13000 301 13050 314
rect 13208 301 13258 314
rect 10293 247 10343 275
rect 10293 227 10306 247
rect 10326 227 10343 247
rect 4041 148 4091 176
rect 1552 115 1602 131
rect 1770 115 1820 131
rect 1978 115 2028 131
rect 4041 128 4054 148
rect 4074 128 4091 148
rect 4041 99 4091 128
rect 4259 151 4309 176
rect 4259 131 4272 151
rect 4292 131 4309 151
rect 4259 99 4309 131
rect 4467 149 4517 176
rect 4467 129 4490 149
rect 4510 129 4517 149
rect 8489 172 8539 200
rect 8489 152 8502 172
rect 8522 152 8539 172
rect 4467 99 4517 129
rect 5916 128 5966 144
rect 6134 128 6184 144
rect 6342 128 6392 144
rect 8489 123 8539 152
rect 8707 175 8757 200
rect 8707 155 8720 175
rect 8740 155 8757 175
rect 8707 123 8757 155
rect 8915 173 8965 200
rect 10293 198 10343 227
rect 10511 250 10561 275
rect 10511 230 10524 250
rect 10544 230 10561 250
rect 10511 198 10561 230
rect 10719 248 10769 275
rect 10719 228 10742 248
rect 10762 228 10769 248
rect 10719 198 10769 228
rect 14657 260 14707 288
rect 14657 240 14670 260
rect 14690 240 14707 260
rect 14657 211 14707 240
rect 14875 263 14925 288
rect 14875 243 14888 263
rect 14908 243 14925 263
rect 14875 211 14925 243
rect 15083 261 15133 288
rect 15083 241 15106 261
rect 15126 241 15133 261
rect 15083 211 15133 241
rect 8915 153 8938 173
rect 8958 153 8965 173
rect 12782 173 12832 201
rect 8915 123 8965 153
rect 10293 140 10343 156
rect 10511 140 10561 156
rect 10719 140 10769 156
rect 12782 153 12795 173
rect 12815 153 12832 173
rect 12782 124 12832 153
rect 13000 176 13050 201
rect 13000 156 13013 176
rect 13033 156 13050 176
rect 13000 124 13050 156
rect 13208 174 13258 201
rect 13208 154 13231 174
rect 13251 154 13258 174
rect 13208 124 13258 154
rect 14657 153 14707 169
rect 14875 153 14925 169
rect 15083 153 15133 169
rect 8489 65 8539 81
rect 8707 65 8757 81
rect 8915 65 8965 81
rect 12782 66 12832 82
rect 13000 66 13050 82
rect 13208 66 13258 82
rect 4041 41 4091 57
rect 4259 41 4309 57
rect 4467 41 4517 57
<< polycont >>
rect 3525 8659 3545 8679
rect 3743 8657 3763 8677
rect 3961 8660 3981 8680
rect 7889 8672 7909 8692
rect 8107 8670 8127 8690
rect 8325 8673 8345 8693
rect 12266 8684 12286 8704
rect 12484 8682 12504 8702
rect 12702 8685 12722 8705
rect 16630 8697 16650 8717
rect 16848 8695 16868 8715
rect 17066 8698 17086 8718
rect 2728 8431 2748 8451
rect 2946 8429 2966 8449
rect 3164 8432 3184 8452
rect 478 8316 498 8336
rect 696 8319 716 8339
rect 914 8317 934 8337
rect 7092 8444 7112 8464
rect 7310 8442 7330 8462
rect 7528 8445 7548 8465
rect 3526 8247 3546 8267
rect 3744 8245 3764 8265
rect 3962 8248 3982 8268
rect 4842 8329 4862 8349
rect 5060 8332 5080 8352
rect 5278 8330 5298 8350
rect 11469 8456 11489 8476
rect 11687 8454 11707 8474
rect 11905 8457 11925 8477
rect 1276 8132 1296 8152
rect 1494 8135 1514 8155
rect 1712 8133 1732 8153
rect 7890 8260 7910 8280
rect 8108 8258 8128 8278
rect 8326 8261 8346 8281
rect 9219 8341 9239 8361
rect 9437 8344 9457 8364
rect 9655 8342 9675 8362
rect 15833 8469 15853 8489
rect 16051 8467 16071 8487
rect 16269 8470 16289 8490
rect 5640 8145 5660 8165
rect 5858 8148 5878 8168
rect 6076 8146 6096 8166
rect 12267 8272 12287 8292
rect 12485 8270 12505 8290
rect 12703 8273 12723 8293
rect 13583 8354 13603 8374
rect 13801 8357 13821 8377
rect 14019 8355 14039 8375
rect 2629 8021 2649 8041
rect 2847 8019 2867 8039
rect 10017 8157 10037 8177
rect 10235 8160 10255 8180
rect 10453 8158 10473 8178
rect 16631 8285 16651 8305
rect 16849 8283 16869 8303
rect 17067 8286 17087 8306
rect 3065 8022 3085 8042
rect 479 7904 499 7924
rect 697 7907 717 7927
rect 915 7905 935 7925
rect 6993 8034 7013 8054
rect 7211 8032 7231 8052
rect 14381 8170 14401 8190
rect 14599 8173 14619 8193
rect 14817 8171 14837 8191
rect 7429 8035 7449 8055
rect 4843 7917 4863 7937
rect 5061 7920 5081 7940
rect 5279 7918 5299 7938
rect 11370 8046 11390 8066
rect 11588 8044 11608 8064
rect 11806 8047 11826 8067
rect 9220 7929 9240 7949
rect 9438 7932 9458 7952
rect 9656 7930 9676 7950
rect 15734 8059 15754 8079
rect 15952 8057 15972 8077
rect 16170 8060 16190 8080
rect 13584 7942 13604 7962
rect 13802 7945 13822 7965
rect 14020 7943 14040 7963
rect 3508 7641 3528 7661
rect 3726 7639 3746 7659
rect 3944 7642 3964 7662
rect 1358 7524 1378 7544
rect 1576 7527 1596 7547
rect 1794 7525 1814 7545
rect 7872 7654 7892 7674
rect 8090 7652 8110 7672
rect 8308 7655 8328 7675
rect 5722 7537 5742 7557
rect 5940 7540 5960 7560
rect 6158 7538 6178 7558
rect 12249 7666 12269 7686
rect 12467 7664 12487 7684
rect 12685 7667 12705 7687
rect 10099 7549 10119 7569
rect 2711 7413 2731 7433
rect 2929 7411 2949 7431
rect 3147 7414 3167 7434
rect 10317 7552 10337 7572
rect 10535 7550 10555 7570
rect 16613 7679 16633 7699
rect 16831 7677 16851 7697
rect 17049 7680 17069 7700
rect 14463 7562 14483 7582
rect 461 7298 481 7318
rect 679 7301 699 7321
rect 897 7299 917 7319
rect 7075 7426 7095 7446
rect 7293 7424 7313 7444
rect 7511 7427 7531 7447
rect 14681 7565 14701 7585
rect 14899 7563 14919 7583
rect 3509 7229 3529 7249
rect 3727 7227 3747 7247
rect 3945 7230 3965 7250
rect 4825 7311 4845 7331
rect 5043 7314 5063 7334
rect 5261 7312 5281 7332
rect 11452 7438 11472 7458
rect 11670 7436 11690 7456
rect 11888 7439 11908 7459
rect 1259 7114 1279 7134
rect 1477 7117 1497 7137
rect 1695 7115 1715 7135
rect 7873 7242 7893 7262
rect 8091 7240 8111 7260
rect 8309 7243 8329 7263
rect 9202 7323 9222 7343
rect 9420 7326 9440 7346
rect 9638 7324 9658 7344
rect 15816 7451 15836 7471
rect 16034 7449 16054 7469
rect 16252 7452 16272 7472
rect 5623 7127 5643 7147
rect 5841 7130 5861 7150
rect 6059 7128 6079 7148
rect 12250 7254 12270 7274
rect 12468 7252 12488 7272
rect 12686 7255 12706 7275
rect 13566 7336 13586 7356
rect 13784 7339 13804 7359
rect 14002 7337 14022 7357
rect 2546 7005 2566 7025
rect 2764 7003 2784 7023
rect 10000 7139 10020 7159
rect 10218 7142 10238 7162
rect 10436 7140 10456 7160
rect 16614 7267 16634 7287
rect 16832 7265 16852 7285
rect 17050 7268 17070 7288
rect 2982 7006 3002 7026
rect 462 6886 482 6906
rect 680 6889 700 6909
rect 898 6887 918 6907
rect 6910 7018 6930 7038
rect 7128 7016 7148 7036
rect 14364 7152 14384 7172
rect 14582 7155 14602 7175
rect 14800 7153 14820 7173
rect 7346 7019 7366 7039
rect 4826 6899 4846 6919
rect 5044 6902 5064 6922
rect 5262 6900 5282 6920
rect 11287 7030 11307 7050
rect 11505 7028 11525 7048
rect 11723 7031 11743 7051
rect 9203 6911 9223 6931
rect 9421 6914 9441 6934
rect 9639 6912 9659 6932
rect 15651 7043 15671 7063
rect 15869 7041 15889 7061
rect 16087 7044 16107 7064
rect 13567 6924 13587 6944
rect 13785 6927 13805 6947
rect 14003 6925 14023 6945
rect 3488 6623 3508 6643
rect 3706 6621 3726 6641
rect 3924 6624 3944 6644
rect 1404 6504 1424 6524
rect 1622 6507 1642 6527
rect 1840 6505 1860 6525
rect 7852 6636 7872 6656
rect 8070 6634 8090 6654
rect 8288 6637 8308 6657
rect 5768 6517 5788 6537
rect 5986 6520 6006 6540
rect 6204 6518 6224 6538
rect 12229 6648 12249 6668
rect 12447 6646 12467 6666
rect 12665 6649 12685 6669
rect 10145 6529 10165 6549
rect 2691 6395 2711 6415
rect 2909 6393 2929 6413
rect 3127 6396 3147 6416
rect 10363 6532 10383 6552
rect 10581 6530 10601 6550
rect 16593 6661 16613 6681
rect 16811 6659 16831 6679
rect 17029 6662 17049 6682
rect 14509 6542 14529 6562
rect 441 6280 461 6300
rect 659 6283 679 6303
rect 877 6281 897 6301
rect 7055 6408 7075 6428
rect 7273 6406 7293 6426
rect 7491 6409 7511 6429
rect 14727 6545 14747 6565
rect 14945 6543 14965 6563
rect 3489 6211 3509 6231
rect 3707 6209 3727 6229
rect 3925 6212 3945 6232
rect 4805 6293 4825 6313
rect 5023 6296 5043 6316
rect 5241 6294 5261 6314
rect 11432 6420 11452 6440
rect 11650 6418 11670 6438
rect 11868 6421 11888 6441
rect 1239 6096 1259 6116
rect 1457 6099 1477 6119
rect 1675 6097 1695 6117
rect 7853 6224 7873 6244
rect 8071 6222 8091 6242
rect 8289 6225 8309 6245
rect 9182 6305 9202 6325
rect 9400 6308 9420 6328
rect 9618 6306 9638 6326
rect 15796 6433 15816 6453
rect 16014 6431 16034 6451
rect 16232 6434 16252 6454
rect 5603 6109 5623 6129
rect 5821 6112 5841 6132
rect 6039 6110 6059 6130
rect 12230 6236 12250 6256
rect 12448 6234 12468 6254
rect 12666 6237 12686 6257
rect 13546 6318 13566 6338
rect 13764 6321 13784 6341
rect 13982 6319 14002 6339
rect 2592 5985 2612 6005
rect 2810 5983 2830 6003
rect 9980 6121 10000 6141
rect 10198 6124 10218 6144
rect 10416 6122 10436 6142
rect 16594 6249 16614 6269
rect 16812 6247 16832 6267
rect 17030 6250 17050 6270
rect 3028 5986 3048 6006
rect 442 5868 462 5888
rect 660 5871 680 5891
rect 878 5869 898 5889
rect 6956 5998 6976 6018
rect 7174 5996 7194 6016
rect 14344 6134 14364 6154
rect 14562 6137 14582 6157
rect 14780 6135 14800 6155
rect 7392 5999 7412 6019
rect 4806 5881 4826 5901
rect 5024 5884 5044 5904
rect 5242 5882 5262 5902
rect 11333 6010 11353 6030
rect 11551 6008 11571 6028
rect 11769 6011 11789 6031
rect 9183 5893 9203 5913
rect 9401 5896 9421 5916
rect 9619 5894 9639 5914
rect 15697 6023 15717 6043
rect 15915 6021 15935 6041
rect 16133 6024 16153 6044
rect 13547 5906 13567 5926
rect 13765 5909 13785 5929
rect 13983 5907 14003 5927
rect 3471 5605 3491 5625
rect 3689 5603 3709 5623
rect 3907 5606 3927 5626
rect 1321 5488 1341 5508
rect 1539 5491 1559 5511
rect 1757 5489 1777 5509
rect 7835 5618 7855 5638
rect 8053 5616 8073 5636
rect 8271 5619 8291 5639
rect 5685 5501 5705 5521
rect 5903 5504 5923 5524
rect 6121 5502 6141 5522
rect 12212 5630 12232 5650
rect 12430 5628 12450 5648
rect 12648 5631 12668 5651
rect 10062 5513 10082 5533
rect 2674 5377 2694 5397
rect 2892 5375 2912 5395
rect 3110 5378 3130 5398
rect 10280 5516 10300 5536
rect 10498 5514 10518 5534
rect 16576 5643 16596 5663
rect 16794 5641 16814 5661
rect 17012 5644 17032 5664
rect 14426 5526 14446 5546
rect 424 5262 444 5282
rect 642 5265 662 5285
rect 860 5263 880 5283
rect 7038 5390 7058 5410
rect 7256 5388 7276 5408
rect 7474 5391 7494 5411
rect 14644 5529 14664 5549
rect 14862 5527 14882 5547
rect 3472 5193 3492 5213
rect 3690 5191 3710 5211
rect 3908 5194 3928 5214
rect 4788 5275 4808 5295
rect 5006 5278 5026 5298
rect 5224 5276 5244 5296
rect 11415 5402 11435 5422
rect 11633 5400 11653 5420
rect 11851 5403 11871 5423
rect 1222 5078 1242 5098
rect 1440 5081 1460 5101
rect 1658 5079 1678 5099
rect 7836 5206 7856 5226
rect 8054 5204 8074 5224
rect 8272 5207 8292 5227
rect 9165 5287 9185 5307
rect 9383 5290 9403 5310
rect 9601 5288 9621 5308
rect 15779 5415 15799 5435
rect 15997 5413 16017 5433
rect 16215 5416 16235 5436
rect 5586 5091 5606 5111
rect 5804 5094 5824 5114
rect 6022 5092 6042 5112
rect 12213 5218 12233 5238
rect 12431 5216 12451 5236
rect 12649 5219 12669 5239
rect 13529 5300 13549 5320
rect 13747 5303 13767 5323
rect 13965 5301 13985 5321
rect 2370 4971 2390 4991
rect 2588 4969 2608 4989
rect 9963 5103 9983 5123
rect 10181 5106 10201 5126
rect 10399 5104 10419 5124
rect 16577 5231 16597 5251
rect 16795 5229 16815 5249
rect 17013 5232 17033 5252
rect 2806 4972 2826 4992
rect 425 4850 445 4870
rect 643 4853 663 4873
rect 861 4851 881 4871
rect 6734 4984 6754 5004
rect 6952 4982 6972 5002
rect 14327 5116 14347 5136
rect 14545 5119 14565 5139
rect 14763 5117 14783 5137
rect 7170 4985 7190 5005
rect 4789 4863 4809 4883
rect 5007 4866 5027 4886
rect 5225 4864 5245 4884
rect 11111 4996 11131 5016
rect 11329 4994 11349 5014
rect 11547 4997 11567 5017
rect 9166 4875 9186 4895
rect 9384 4878 9404 4898
rect 9602 4876 9622 4896
rect 15475 5009 15495 5029
rect 15693 5007 15713 5027
rect 15911 5010 15931 5030
rect 13530 4888 13550 4908
rect 13748 4891 13768 4911
rect 13966 4889 13986 4909
rect 3452 4587 3472 4607
rect 3670 4585 3690 4605
rect 3888 4588 3908 4608
rect 1507 4466 1527 4486
rect 1725 4469 1745 4489
rect 1943 4467 1963 4487
rect 7816 4600 7836 4620
rect 8034 4598 8054 4618
rect 8252 4601 8272 4621
rect 5871 4479 5891 4499
rect 6089 4482 6109 4502
rect 6307 4480 6327 4500
rect 12193 4612 12213 4632
rect 12411 4610 12431 4630
rect 12629 4613 12649 4633
rect 10248 4491 10268 4511
rect 2655 4359 2675 4379
rect 2873 4357 2893 4377
rect 3091 4360 3111 4380
rect 10466 4494 10486 4514
rect 10684 4492 10704 4512
rect 16557 4625 16577 4645
rect 16775 4623 16795 4643
rect 16993 4626 17013 4646
rect 14612 4504 14632 4524
rect 405 4244 425 4264
rect 623 4247 643 4267
rect 841 4245 861 4265
rect 7019 4372 7039 4392
rect 7237 4370 7257 4390
rect 7455 4373 7475 4393
rect 14830 4507 14850 4527
rect 15048 4505 15068 4525
rect 3453 4175 3473 4195
rect 3671 4173 3691 4193
rect 3889 4176 3909 4196
rect 4769 4257 4789 4277
rect 4987 4260 5007 4280
rect 5205 4258 5225 4278
rect 11396 4384 11416 4404
rect 11614 4382 11634 4402
rect 11832 4385 11852 4405
rect 1203 4060 1223 4080
rect 1421 4063 1441 4083
rect 1639 4061 1659 4081
rect 7817 4188 7837 4208
rect 8035 4186 8055 4206
rect 8253 4189 8273 4209
rect 9146 4269 9166 4289
rect 9364 4272 9384 4292
rect 9582 4270 9602 4290
rect 15760 4397 15780 4417
rect 15978 4395 15998 4415
rect 16196 4398 16216 4418
rect 5567 4073 5587 4093
rect 5785 4076 5805 4096
rect 6003 4074 6023 4094
rect 12194 4200 12214 4220
rect 12412 4198 12432 4218
rect 12630 4201 12650 4221
rect 13510 4282 13530 4302
rect 13728 4285 13748 4305
rect 13946 4283 13966 4303
rect 2556 3949 2576 3969
rect 2774 3947 2794 3967
rect 9944 4085 9964 4105
rect 10162 4088 10182 4108
rect 10380 4086 10400 4106
rect 16558 4213 16578 4233
rect 16776 4211 16796 4231
rect 16994 4214 17014 4234
rect 2992 3950 3012 3970
rect 406 3832 426 3852
rect 624 3835 644 3855
rect 842 3833 862 3853
rect 6920 3962 6940 3982
rect 7138 3960 7158 3980
rect 14308 4098 14328 4118
rect 14526 4101 14546 4121
rect 14744 4099 14764 4119
rect 7356 3963 7376 3983
rect 4770 3845 4790 3865
rect 4988 3848 5008 3868
rect 5206 3846 5226 3866
rect 11297 3974 11317 3994
rect 11515 3972 11535 3992
rect 11733 3975 11753 3995
rect 9147 3857 9167 3877
rect 9365 3860 9385 3880
rect 9583 3858 9603 3878
rect 15661 3987 15681 4007
rect 15879 3985 15899 4005
rect 16097 3988 16117 4008
rect 13511 3870 13531 3890
rect 13729 3873 13749 3893
rect 13947 3871 13967 3891
rect 3435 3569 3455 3589
rect 3653 3567 3673 3587
rect 3871 3570 3891 3590
rect 1285 3452 1305 3472
rect 1503 3455 1523 3475
rect 1721 3453 1741 3473
rect 7799 3582 7819 3602
rect 8017 3580 8037 3600
rect 8235 3583 8255 3603
rect 5649 3465 5669 3485
rect 5867 3468 5887 3488
rect 6085 3466 6105 3486
rect 12176 3594 12196 3614
rect 12394 3592 12414 3612
rect 12612 3595 12632 3615
rect 10026 3477 10046 3497
rect 2638 3341 2658 3361
rect 2856 3339 2876 3359
rect 3074 3342 3094 3362
rect 10244 3480 10264 3500
rect 10462 3478 10482 3498
rect 16540 3607 16560 3627
rect 16758 3605 16778 3625
rect 16976 3608 16996 3628
rect 14390 3490 14410 3510
rect 388 3226 408 3246
rect 606 3229 626 3249
rect 824 3227 844 3247
rect 7002 3354 7022 3374
rect 7220 3352 7240 3372
rect 7438 3355 7458 3375
rect 14608 3493 14628 3513
rect 14826 3491 14846 3511
rect 3436 3157 3456 3177
rect 3654 3155 3674 3175
rect 3872 3158 3892 3178
rect 4752 3239 4772 3259
rect 4970 3242 4990 3262
rect 5188 3240 5208 3260
rect 11379 3366 11399 3386
rect 11597 3364 11617 3384
rect 11815 3367 11835 3387
rect 1186 3042 1206 3062
rect 1404 3045 1424 3065
rect 1622 3043 1642 3063
rect 7800 3170 7820 3190
rect 8018 3168 8038 3188
rect 8236 3171 8256 3191
rect 9129 3251 9149 3271
rect 9347 3254 9367 3274
rect 9565 3252 9585 3272
rect 15743 3379 15763 3399
rect 15961 3377 15981 3397
rect 16179 3380 16199 3400
rect 5550 3055 5570 3075
rect 5768 3058 5788 3078
rect 5986 3056 6006 3076
rect 12177 3182 12197 3202
rect 12395 3180 12415 3200
rect 12613 3183 12633 3203
rect 13493 3264 13513 3284
rect 13711 3267 13731 3287
rect 13929 3265 13949 3285
rect 2473 2933 2493 2953
rect 2691 2931 2711 2951
rect 9927 3067 9947 3087
rect 10145 3070 10165 3090
rect 10363 3068 10383 3088
rect 16541 3195 16561 3215
rect 16759 3193 16779 3213
rect 16977 3196 16997 3216
rect 2909 2934 2929 2954
rect 389 2814 409 2834
rect 607 2817 627 2837
rect 825 2815 845 2835
rect 6837 2946 6857 2966
rect 7055 2944 7075 2964
rect 14291 3080 14311 3100
rect 14509 3083 14529 3103
rect 14727 3081 14747 3101
rect 7273 2947 7293 2967
rect 4753 2827 4773 2847
rect 4971 2830 4991 2850
rect 5189 2828 5209 2848
rect 11214 2958 11234 2978
rect 11432 2956 11452 2976
rect 11650 2959 11670 2979
rect 9130 2839 9150 2859
rect 9348 2842 9368 2862
rect 9566 2840 9586 2860
rect 15578 2971 15598 2991
rect 15796 2969 15816 2989
rect 16014 2972 16034 2992
rect 13494 2852 13514 2872
rect 13712 2855 13732 2875
rect 13930 2853 13950 2873
rect 3415 2551 3435 2571
rect 3633 2549 3653 2569
rect 3851 2552 3871 2572
rect 1331 2432 1351 2452
rect 1549 2435 1569 2455
rect 1767 2433 1787 2453
rect 7779 2564 7799 2584
rect 7997 2562 8017 2582
rect 8215 2565 8235 2585
rect 5695 2445 5715 2465
rect 5913 2448 5933 2468
rect 6131 2446 6151 2466
rect 12156 2576 12176 2596
rect 12374 2574 12394 2594
rect 12592 2577 12612 2597
rect 10072 2457 10092 2477
rect 2618 2323 2638 2343
rect 2836 2321 2856 2341
rect 3054 2324 3074 2344
rect 10290 2460 10310 2480
rect 10508 2458 10528 2478
rect 16520 2589 16540 2609
rect 16738 2587 16758 2607
rect 16956 2590 16976 2610
rect 14436 2470 14456 2490
rect 368 2208 388 2228
rect 586 2211 606 2231
rect 804 2209 824 2229
rect 6982 2336 7002 2356
rect 7200 2334 7220 2354
rect 7418 2337 7438 2357
rect 14654 2473 14674 2493
rect 14872 2471 14892 2491
rect 3416 2139 3436 2159
rect 3634 2137 3654 2157
rect 3852 2140 3872 2160
rect 4732 2221 4752 2241
rect 4950 2224 4970 2244
rect 5168 2222 5188 2242
rect 11359 2348 11379 2368
rect 11577 2346 11597 2366
rect 11795 2349 11815 2369
rect 1166 2024 1186 2044
rect 1384 2027 1404 2047
rect 1602 2025 1622 2045
rect 7780 2152 7800 2172
rect 7998 2150 8018 2170
rect 8216 2153 8236 2173
rect 9109 2233 9129 2253
rect 9327 2236 9347 2256
rect 9545 2234 9565 2254
rect 15723 2361 15743 2381
rect 15941 2359 15961 2379
rect 16159 2362 16179 2382
rect 5530 2037 5550 2057
rect 5748 2040 5768 2060
rect 5966 2038 5986 2058
rect 12157 2164 12177 2184
rect 12375 2162 12395 2182
rect 12593 2165 12613 2185
rect 13473 2246 13493 2266
rect 13691 2249 13711 2269
rect 13909 2247 13929 2267
rect 2519 1913 2539 1933
rect 2737 1911 2757 1931
rect 9907 2049 9927 2069
rect 10125 2052 10145 2072
rect 10343 2050 10363 2070
rect 16521 2177 16541 2197
rect 16739 2175 16759 2195
rect 16957 2178 16977 2198
rect 2955 1914 2975 1934
rect 369 1796 389 1816
rect 587 1799 607 1819
rect 805 1797 825 1817
rect 6883 1926 6903 1946
rect 7101 1924 7121 1944
rect 14271 2062 14291 2082
rect 14489 2065 14509 2085
rect 14707 2063 14727 2083
rect 7319 1927 7339 1947
rect 4733 1809 4753 1829
rect 4951 1812 4971 1832
rect 5169 1810 5189 1830
rect 11260 1938 11280 1958
rect 11478 1936 11498 1956
rect 11696 1939 11716 1959
rect 9110 1821 9130 1841
rect 9328 1824 9348 1844
rect 9546 1822 9566 1842
rect 15624 1951 15644 1971
rect 15842 1949 15862 1969
rect 16060 1952 16080 1972
rect 13474 1834 13494 1854
rect 13692 1837 13712 1857
rect 13910 1835 13930 1855
rect 3398 1533 3418 1553
rect 3616 1531 3636 1551
rect 3834 1534 3854 1554
rect 1248 1416 1268 1436
rect 1466 1419 1486 1439
rect 1684 1417 1704 1437
rect 7762 1546 7782 1566
rect 7980 1544 8000 1564
rect 8198 1547 8218 1567
rect 5612 1429 5632 1449
rect 5830 1432 5850 1452
rect 6048 1430 6068 1450
rect 12139 1558 12159 1578
rect 12357 1556 12377 1576
rect 12575 1559 12595 1579
rect 9989 1441 10009 1461
rect 2601 1305 2621 1325
rect 2819 1303 2839 1323
rect 3037 1306 3057 1326
rect 10207 1444 10227 1464
rect 10425 1442 10445 1462
rect 16503 1571 16523 1591
rect 16721 1569 16741 1589
rect 16939 1572 16959 1592
rect 14353 1454 14373 1474
rect 351 1190 371 1210
rect 569 1193 589 1213
rect 787 1191 807 1211
rect 6965 1318 6985 1338
rect 7183 1316 7203 1336
rect 7401 1319 7421 1339
rect 14571 1457 14591 1477
rect 14789 1455 14809 1475
rect 3399 1121 3419 1141
rect 3617 1119 3637 1139
rect 3835 1122 3855 1142
rect 4715 1203 4735 1223
rect 4933 1206 4953 1226
rect 5151 1204 5171 1224
rect 11342 1330 11362 1350
rect 11560 1328 11580 1348
rect 11778 1331 11798 1351
rect 1149 1006 1169 1026
rect 1367 1009 1387 1029
rect 1585 1007 1605 1027
rect 7763 1134 7783 1154
rect 7981 1132 8001 1152
rect 8199 1135 8219 1155
rect 9092 1215 9112 1235
rect 9310 1218 9330 1238
rect 9528 1216 9548 1236
rect 15706 1343 15726 1363
rect 15924 1341 15944 1361
rect 16142 1344 16162 1364
rect 5513 1019 5533 1039
rect 5731 1022 5751 1042
rect 5949 1020 5969 1040
rect 12140 1146 12160 1166
rect 12358 1144 12378 1164
rect 12576 1147 12596 1167
rect 13456 1228 13476 1248
rect 13674 1231 13694 1251
rect 13892 1229 13912 1249
rect 9890 1031 9910 1051
rect 10108 1034 10128 1054
rect 10326 1032 10346 1052
rect 16504 1159 16524 1179
rect 16722 1157 16742 1177
rect 16940 1160 16960 1180
rect 14254 1044 14274 1064
rect 14472 1047 14492 1067
rect 14690 1045 14710 1065
rect 352 778 372 798
rect 570 781 590 801
rect 788 779 808 799
rect 4716 791 4736 811
rect 4934 794 4954 814
rect 5152 792 5172 812
rect 9093 803 9113 823
rect 9311 806 9331 826
rect 9529 804 9549 824
rect 13457 816 13477 836
rect 13675 819 13695 839
rect 13893 817 13913 837
rect 1565 202 1585 222
rect 1783 205 1803 225
rect 2001 203 2021 223
rect 5929 215 5949 235
rect 6147 218 6167 238
rect 6365 216 6385 236
rect 10306 227 10326 247
rect 4054 128 4074 148
rect 4272 131 4292 151
rect 4490 129 4510 149
rect 8502 152 8522 172
rect 8720 155 8740 175
rect 10524 230 10544 250
rect 10742 228 10762 248
rect 14670 240 14690 260
rect 14888 243 14908 263
rect 15106 241 15126 261
rect 8938 153 8958 173
rect 12795 153 12815 173
rect 13013 156 13033 176
rect 13231 154 13251 174
<< ndiffres >>
rect 4181 8744 4238 8763
rect 4181 8726 4199 8744
rect 4217 8741 4238 8744
rect 4217 8726 4332 8741
rect 240 8686 301 8702
rect 145 8682 301 8686
rect 145 8664 263 8682
rect 281 8664 301 8682
rect 145 8643 301 8664
rect 145 8642 245 8643
rect 146 8606 188 8642
rect 4181 8703 4332 8726
rect 8545 8757 8602 8776
rect 8545 8739 8563 8757
rect 8581 8754 8602 8757
rect 8581 8739 8696 8754
rect 4290 8667 4332 8703
rect 4604 8699 4665 8715
rect 4509 8695 4665 8699
rect 4509 8677 4627 8695
rect 4645 8677 4665 8695
rect 4233 8666 4333 8667
rect 4177 8645 4333 8666
rect 4509 8656 4665 8677
rect 4509 8655 4609 8656
rect 146 8583 297 8606
rect 146 8568 261 8583
rect 240 8565 261 8568
rect 279 8565 297 8583
rect 240 8546 297 8565
rect 4177 8627 4197 8645
rect 4215 8627 4333 8645
rect 4177 8623 4333 8627
rect 4177 8607 4238 8623
rect 4510 8619 4552 8655
rect 8545 8716 8696 8739
rect 12922 8769 12979 8788
rect 12922 8751 12940 8769
rect 12958 8766 12979 8769
rect 12958 8751 13073 8766
rect 8654 8680 8696 8716
rect 8981 8711 9042 8727
rect 8886 8707 9042 8711
rect 8886 8689 9004 8707
rect 9022 8689 9042 8707
rect 8597 8679 8697 8680
rect 8541 8658 8697 8679
rect 8886 8668 9042 8689
rect 8886 8667 8986 8668
rect 4510 8596 4661 8619
rect 4510 8581 4625 8596
rect 4604 8578 4625 8581
rect 4643 8578 4661 8596
rect 4604 8559 4661 8578
rect 4174 8526 4231 8545
rect 8541 8640 8561 8658
rect 8579 8640 8697 8658
rect 8541 8636 8697 8640
rect 8541 8620 8602 8636
rect 8887 8631 8929 8667
rect 12922 8728 13073 8751
rect 17286 8782 17343 8801
rect 17286 8764 17304 8782
rect 17322 8779 17343 8782
rect 17322 8764 17437 8779
rect 13031 8692 13073 8728
rect 13345 8724 13406 8740
rect 13250 8720 13406 8724
rect 13250 8702 13368 8720
rect 13386 8702 13406 8720
rect 12974 8691 13074 8692
rect 12918 8670 13074 8691
rect 13250 8681 13406 8702
rect 13250 8680 13350 8681
rect 8887 8608 9038 8631
rect 8887 8593 9002 8608
rect 8981 8590 9002 8593
rect 9020 8590 9038 8608
rect 8981 8571 9038 8590
rect 4174 8508 4192 8526
rect 4210 8523 4231 8526
rect 4210 8508 4325 8523
rect 4174 8485 4325 8508
rect 8538 8539 8595 8558
rect 12918 8652 12938 8670
rect 12956 8652 13074 8670
rect 12918 8648 13074 8652
rect 12918 8632 12979 8648
rect 13251 8644 13293 8680
rect 17286 8741 17437 8764
rect 17395 8705 17437 8741
rect 17338 8704 17438 8705
rect 17282 8683 17438 8704
rect 13251 8621 13402 8644
rect 13251 8606 13366 8621
rect 13345 8603 13366 8606
rect 13384 8603 13402 8621
rect 13345 8584 13402 8603
rect 8538 8521 8556 8539
rect 8574 8536 8595 8539
rect 8574 8521 8689 8536
rect 8538 8498 8689 8521
rect 12915 8551 12972 8570
rect 17282 8665 17302 8683
rect 17320 8665 17438 8683
rect 17282 8661 17438 8665
rect 17282 8645 17343 8661
rect 12915 8533 12933 8551
rect 12951 8548 12972 8551
rect 12951 8533 13066 8548
rect 12915 8510 13066 8533
rect 17279 8564 17336 8583
rect 17279 8546 17297 8564
rect 17315 8561 17336 8564
rect 17315 8546 17430 8561
rect 17279 8523 17430 8546
rect 235 8362 296 8378
rect 4283 8449 4325 8485
rect 4226 8448 4326 8449
rect 4170 8427 4326 8448
rect 4170 8409 4190 8427
rect 4208 8409 4326 8427
rect 4170 8405 4326 8409
rect 140 8358 296 8362
rect 140 8340 258 8358
rect 276 8340 296 8358
rect 140 8319 296 8340
rect 140 8318 240 8319
rect 141 8282 183 8318
rect 4170 8389 4231 8405
rect 4599 8375 4660 8391
rect 8647 8462 8689 8498
rect 8590 8461 8690 8462
rect 8534 8440 8690 8461
rect 8534 8422 8554 8440
rect 8572 8422 8690 8440
rect 8534 8418 8690 8422
rect 4504 8371 4660 8375
rect 4168 8343 4225 8362
rect 141 8259 292 8282
rect 141 8244 256 8259
rect 235 8241 256 8244
rect 274 8241 292 8259
rect 4168 8325 4186 8343
rect 4204 8340 4225 8343
rect 4504 8353 4622 8371
rect 4640 8353 4660 8371
rect 4204 8325 4319 8340
rect 4504 8332 4660 8353
rect 4504 8331 4604 8332
rect 4168 8302 4319 8325
rect 235 8222 292 8241
rect 229 8179 290 8195
rect 4277 8266 4319 8302
rect 4505 8295 4547 8331
rect 8534 8402 8595 8418
rect 8976 8387 9037 8403
rect 13024 8474 13066 8510
rect 12967 8473 13067 8474
rect 12911 8452 13067 8473
rect 12911 8434 12931 8452
rect 12949 8434 13067 8452
rect 12911 8430 13067 8434
rect 8881 8383 9037 8387
rect 8532 8356 8589 8375
rect 4505 8272 4656 8295
rect 4220 8265 4320 8266
rect 4164 8244 4320 8265
rect 4505 8257 4620 8272
rect 4164 8226 4184 8244
rect 4202 8226 4320 8244
rect 4599 8254 4620 8257
rect 4638 8254 4656 8272
rect 8532 8338 8550 8356
rect 8568 8353 8589 8356
rect 8881 8365 8999 8383
rect 9017 8365 9037 8383
rect 8568 8338 8683 8353
rect 8881 8344 9037 8365
rect 8881 8343 8981 8344
rect 8532 8315 8683 8338
rect 4599 8235 4656 8254
rect 4164 8222 4320 8226
rect 134 8175 290 8179
rect 134 8157 252 8175
rect 270 8157 290 8175
rect 134 8136 290 8157
rect 134 8135 234 8136
rect 135 8099 177 8135
rect 4164 8206 4225 8222
rect 4593 8192 4654 8208
rect 8641 8279 8683 8315
rect 8882 8307 8924 8343
rect 12911 8414 12972 8430
rect 13340 8400 13401 8416
rect 17388 8487 17430 8523
rect 17331 8486 17431 8487
rect 17275 8465 17431 8486
rect 17275 8447 17295 8465
rect 17313 8447 17431 8465
rect 17275 8443 17431 8447
rect 13245 8396 13401 8400
rect 12909 8368 12966 8387
rect 8882 8284 9033 8307
rect 8584 8278 8684 8279
rect 8528 8257 8684 8278
rect 8882 8269 8997 8284
rect 8528 8239 8548 8257
rect 8566 8239 8684 8257
rect 8976 8266 8997 8269
rect 9015 8266 9033 8284
rect 12909 8350 12927 8368
rect 12945 8365 12966 8368
rect 13245 8378 13363 8396
rect 13381 8378 13401 8396
rect 12945 8350 13060 8365
rect 13245 8357 13401 8378
rect 13245 8356 13345 8357
rect 12909 8327 13060 8350
rect 8976 8247 9033 8266
rect 8528 8235 8684 8239
rect 4498 8188 4654 8192
rect 4498 8170 4616 8188
rect 4634 8170 4654 8188
rect 4498 8149 4654 8170
rect 4498 8148 4598 8149
rect 135 8076 286 8099
rect 135 8061 250 8076
rect 229 8058 250 8061
rect 268 8058 286 8076
rect 229 8039 286 8058
rect 4499 8112 4541 8148
rect 8528 8219 8589 8235
rect 8970 8204 9031 8220
rect 13018 8291 13060 8327
rect 13246 8320 13288 8356
rect 17275 8427 17336 8443
rect 17273 8381 17330 8400
rect 13246 8297 13397 8320
rect 12961 8290 13061 8291
rect 12905 8269 13061 8290
rect 13246 8282 13361 8297
rect 12905 8251 12925 8269
rect 12943 8251 13061 8269
rect 13340 8279 13361 8282
rect 13379 8279 13397 8297
rect 17273 8363 17291 8381
rect 17309 8378 17330 8381
rect 17309 8363 17424 8378
rect 17273 8340 17424 8363
rect 13340 8260 13397 8279
rect 12905 8247 13061 8251
rect 8875 8200 9031 8204
rect 8875 8182 8993 8200
rect 9011 8182 9031 8200
rect 8875 8161 9031 8182
rect 8875 8160 8975 8161
rect 4499 8089 4650 8112
rect 4499 8074 4614 8089
rect 4593 8071 4614 8074
rect 4632 8071 4650 8089
rect 222 7961 283 7977
rect 127 7957 283 7961
rect 127 7939 245 7957
rect 263 7939 283 7957
rect 4593 8052 4650 8071
rect 8876 8124 8918 8160
rect 12905 8231 12966 8247
rect 13334 8217 13395 8233
rect 17382 8304 17424 8340
rect 17325 8303 17425 8304
rect 17269 8282 17425 8303
rect 17269 8264 17289 8282
rect 17307 8264 17425 8282
rect 17269 8260 17425 8264
rect 13239 8213 13395 8217
rect 13239 8195 13357 8213
rect 13375 8195 13395 8213
rect 13239 8174 13395 8195
rect 13239 8173 13339 8174
rect 8876 8101 9027 8124
rect 8876 8086 8991 8101
rect 4163 8019 4220 8038
rect 4163 8001 4181 8019
rect 4199 8016 4220 8019
rect 4199 8001 4314 8016
rect 127 7918 283 7939
rect 127 7917 227 7918
rect 128 7881 170 7917
rect 128 7858 279 7881
rect 4163 7978 4314 8001
rect 4272 7942 4314 7978
rect 4586 7974 4647 7990
rect 4491 7970 4647 7974
rect 4491 7952 4609 7970
rect 4627 7952 4647 7970
rect 8970 8083 8991 8086
rect 9009 8083 9027 8101
rect 8970 8064 9027 8083
rect 13240 8137 13282 8173
rect 17269 8244 17330 8260
rect 13240 8114 13391 8137
rect 13240 8099 13355 8114
rect 13334 8096 13355 8099
rect 13373 8096 13391 8114
rect 8527 8032 8584 8051
rect 8527 8014 8545 8032
rect 8563 8029 8584 8032
rect 8563 8014 8678 8029
rect 4215 7941 4315 7942
rect 4159 7920 4315 7941
rect 4491 7931 4647 7952
rect 4491 7930 4591 7931
rect 4159 7902 4179 7920
rect 4197 7902 4315 7920
rect 4159 7898 4315 7902
rect 4159 7882 4220 7898
rect 4492 7894 4534 7930
rect 128 7843 243 7858
rect 222 7840 243 7843
rect 261 7840 279 7858
rect 222 7821 279 7840
rect 4492 7871 4643 7894
rect 8527 7991 8678 8014
rect 8636 7955 8678 7991
rect 8963 7986 9024 8002
rect 8868 7982 9024 7986
rect 8868 7964 8986 7982
rect 9004 7964 9024 7982
rect 13334 8077 13391 8096
rect 12904 8044 12961 8063
rect 12904 8026 12922 8044
rect 12940 8041 12961 8044
rect 12940 8026 13055 8041
rect 8579 7954 8679 7955
rect 8523 7933 8679 7954
rect 8868 7943 9024 7964
rect 8868 7942 8968 7943
rect 8523 7915 8543 7933
rect 8561 7915 8679 7933
rect 8523 7911 8679 7915
rect 8523 7895 8584 7911
rect 8869 7906 8911 7942
rect 4492 7856 4607 7871
rect 4586 7853 4607 7856
rect 4625 7853 4643 7871
rect 4586 7834 4643 7853
rect 8869 7883 9020 7906
rect 12904 8003 13055 8026
rect 13013 7967 13055 8003
rect 13327 7999 13388 8015
rect 13232 7995 13388 7999
rect 13232 7977 13350 7995
rect 13368 7977 13388 7995
rect 17268 8057 17325 8076
rect 17268 8039 17286 8057
rect 17304 8054 17325 8057
rect 17304 8039 17419 8054
rect 12956 7966 13056 7967
rect 12900 7945 13056 7966
rect 13232 7956 13388 7977
rect 13232 7955 13332 7956
rect 12900 7927 12920 7945
rect 12938 7927 13056 7945
rect 12900 7923 13056 7927
rect 12900 7907 12961 7923
rect 13233 7919 13275 7955
rect 8869 7868 8984 7883
rect 8963 7865 8984 7868
rect 9002 7865 9020 7883
rect 8963 7846 9020 7865
rect 13233 7896 13384 7919
rect 17268 8016 17419 8039
rect 17377 7980 17419 8016
rect 17320 7979 17420 7980
rect 17264 7958 17420 7979
rect 17264 7940 17284 7958
rect 17302 7940 17420 7958
rect 17264 7936 17420 7940
rect 17264 7920 17325 7936
rect 13233 7881 13348 7896
rect 13327 7878 13348 7881
rect 13366 7878 13384 7896
rect 13327 7859 13384 7878
rect 4164 7726 4221 7745
rect 4164 7708 4182 7726
rect 4200 7723 4221 7726
rect 4200 7708 4315 7723
rect 223 7668 284 7684
rect 128 7664 284 7668
rect 128 7646 246 7664
rect 264 7646 284 7664
rect 128 7625 284 7646
rect 128 7624 228 7625
rect 129 7588 171 7624
rect 129 7565 280 7588
rect 4164 7685 4315 7708
rect 8528 7739 8585 7758
rect 8528 7721 8546 7739
rect 8564 7736 8585 7739
rect 8564 7721 8679 7736
rect 4273 7649 4315 7685
rect 4587 7681 4648 7697
rect 4492 7677 4648 7681
rect 4492 7659 4610 7677
rect 4628 7659 4648 7677
rect 4216 7648 4316 7649
rect 4160 7627 4316 7648
rect 4492 7638 4648 7659
rect 4492 7637 4592 7638
rect 129 7550 244 7565
rect 223 7547 244 7550
rect 262 7547 280 7565
rect 223 7528 280 7547
rect 4160 7609 4180 7627
rect 4198 7609 4316 7627
rect 4160 7605 4316 7609
rect 4160 7589 4221 7605
rect 4493 7601 4535 7637
rect 4493 7578 4644 7601
rect 8528 7698 8679 7721
rect 12905 7751 12962 7770
rect 12905 7733 12923 7751
rect 12941 7748 12962 7751
rect 12941 7733 13056 7748
rect 8637 7662 8679 7698
rect 8964 7693 9025 7709
rect 8869 7689 9025 7693
rect 8869 7671 8987 7689
rect 9005 7671 9025 7689
rect 8580 7661 8680 7662
rect 8524 7640 8680 7661
rect 8869 7650 9025 7671
rect 8869 7649 8969 7650
rect 4493 7563 4608 7578
rect 4587 7560 4608 7563
rect 4626 7560 4644 7578
rect 4587 7541 4644 7560
rect 4157 7508 4214 7527
rect 8524 7622 8544 7640
rect 8562 7622 8680 7640
rect 8524 7618 8680 7622
rect 8524 7602 8585 7618
rect 8870 7613 8912 7649
rect 8870 7590 9021 7613
rect 12905 7710 13056 7733
rect 17269 7764 17326 7783
rect 17269 7746 17287 7764
rect 17305 7761 17326 7764
rect 17305 7746 17420 7761
rect 13014 7674 13056 7710
rect 13328 7706 13389 7722
rect 13233 7702 13389 7706
rect 13233 7684 13351 7702
rect 13369 7684 13389 7702
rect 12957 7673 13057 7674
rect 12901 7652 13057 7673
rect 13233 7663 13389 7684
rect 13233 7662 13333 7663
rect 8870 7575 8985 7590
rect 8964 7572 8985 7575
rect 9003 7572 9021 7590
rect 8964 7553 9021 7572
rect 4157 7490 4175 7508
rect 4193 7505 4214 7508
rect 4193 7490 4308 7505
rect 4157 7467 4308 7490
rect 218 7344 279 7360
rect 4266 7431 4308 7467
rect 8521 7521 8578 7540
rect 8521 7503 8539 7521
rect 8557 7518 8578 7521
rect 12901 7634 12921 7652
rect 12939 7634 13057 7652
rect 12901 7630 13057 7634
rect 12901 7614 12962 7630
rect 13234 7626 13276 7662
rect 13234 7603 13385 7626
rect 17269 7723 17420 7746
rect 17378 7687 17420 7723
rect 17321 7686 17421 7687
rect 17265 7665 17421 7686
rect 13234 7588 13349 7603
rect 13328 7585 13349 7588
rect 13367 7585 13385 7603
rect 13328 7566 13385 7585
rect 8557 7503 8672 7518
rect 8521 7480 8672 7503
rect 4209 7430 4309 7431
rect 4153 7409 4309 7430
rect 4153 7391 4173 7409
rect 4191 7391 4309 7409
rect 4153 7387 4309 7391
rect 123 7340 279 7344
rect 123 7322 241 7340
rect 259 7322 279 7340
rect 123 7301 279 7322
rect 123 7300 223 7301
rect 124 7264 166 7300
rect 4153 7371 4214 7387
rect 4582 7357 4643 7373
rect 8630 7444 8672 7480
rect 12898 7533 12955 7552
rect 17265 7647 17285 7665
rect 17303 7647 17421 7665
rect 17265 7643 17421 7647
rect 17265 7627 17326 7643
rect 12898 7515 12916 7533
rect 12934 7530 12955 7533
rect 12934 7515 13049 7530
rect 12898 7492 13049 7515
rect 8573 7443 8673 7444
rect 8517 7422 8673 7443
rect 8517 7404 8537 7422
rect 8555 7404 8673 7422
rect 8517 7400 8673 7404
rect 4487 7353 4643 7357
rect 4151 7325 4208 7344
rect 124 7241 275 7264
rect 124 7226 239 7241
rect 218 7223 239 7226
rect 257 7223 275 7241
rect 4151 7307 4169 7325
rect 4187 7322 4208 7325
rect 4487 7335 4605 7353
rect 4623 7335 4643 7353
rect 4187 7307 4302 7322
rect 4487 7314 4643 7335
rect 4487 7313 4587 7314
rect 4151 7284 4302 7307
rect 218 7204 275 7223
rect 212 7161 273 7177
rect 4260 7248 4302 7284
rect 4488 7277 4530 7313
rect 8517 7384 8578 7400
rect 8959 7369 9020 7385
rect 13007 7456 13049 7492
rect 17262 7546 17319 7565
rect 17262 7528 17280 7546
rect 17298 7543 17319 7546
rect 17298 7528 17413 7543
rect 17262 7505 17413 7528
rect 12950 7455 13050 7456
rect 12894 7434 13050 7455
rect 12894 7416 12914 7434
rect 12932 7416 13050 7434
rect 12894 7412 13050 7416
rect 8864 7365 9020 7369
rect 8515 7338 8572 7357
rect 4488 7254 4639 7277
rect 4203 7247 4303 7248
rect 4147 7226 4303 7247
rect 4488 7239 4603 7254
rect 4147 7208 4167 7226
rect 4185 7208 4303 7226
rect 4582 7236 4603 7239
rect 4621 7236 4639 7254
rect 8515 7320 8533 7338
rect 8551 7335 8572 7338
rect 8864 7347 8982 7365
rect 9000 7347 9020 7365
rect 8551 7320 8666 7335
rect 8864 7326 9020 7347
rect 8864 7325 8964 7326
rect 8515 7297 8666 7320
rect 4582 7217 4639 7236
rect 4147 7204 4303 7208
rect 117 7157 273 7161
rect 117 7139 235 7157
rect 253 7139 273 7157
rect 117 7118 273 7139
rect 117 7117 217 7118
rect 118 7081 160 7117
rect 4147 7188 4208 7204
rect 4576 7174 4637 7190
rect 8624 7261 8666 7297
rect 8865 7289 8907 7325
rect 12894 7396 12955 7412
rect 13323 7382 13384 7398
rect 17371 7469 17413 7505
rect 17314 7468 17414 7469
rect 17258 7447 17414 7468
rect 17258 7429 17278 7447
rect 17296 7429 17414 7447
rect 17258 7425 17414 7429
rect 13228 7378 13384 7382
rect 12892 7350 12949 7369
rect 8865 7266 9016 7289
rect 8567 7260 8667 7261
rect 8511 7239 8667 7260
rect 8865 7251 8980 7266
rect 8511 7221 8531 7239
rect 8549 7221 8667 7239
rect 8959 7248 8980 7251
rect 8998 7248 9016 7266
rect 12892 7332 12910 7350
rect 12928 7347 12949 7350
rect 13228 7360 13346 7378
rect 13364 7360 13384 7378
rect 12928 7332 13043 7347
rect 13228 7339 13384 7360
rect 13228 7338 13328 7339
rect 12892 7309 13043 7332
rect 8959 7229 9016 7248
rect 8511 7217 8667 7221
rect 4481 7170 4637 7174
rect 4481 7152 4599 7170
rect 4617 7152 4637 7170
rect 4481 7131 4637 7152
rect 4481 7130 4581 7131
rect 118 7058 269 7081
rect 118 7043 233 7058
rect 212 7040 233 7043
rect 251 7040 269 7058
rect 212 7021 269 7040
rect 4482 7094 4524 7130
rect 8511 7201 8572 7217
rect 8953 7186 9014 7202
rect 13001 7273 13043 7309
rect 13229 7302 13271 7338
rect 17258 7409 17319 7425
rect 17256 7363 17313 7382
rect 13229 7279 13380 7302
rect 12944 7272 13044 7273
rect 12888 7251 13044 7272
rect 13229 7264 13344 7279
rect 12888 7233 12908 7251
rect 12926 7233 13044 7251
rect 13323 7261 13344 7264
rect 13362 7261 13380 7279
rect 17256 7345 17274 7363
rect 17292 7360 17313 7363
rect 17292 7345 17407 7360
rect 17256 7322 17407 7345
rect 13323 7242 13380 7261
rect 12888 7229 13044 7233
rect 8858 7182 9014 7186
rect 8858 7164 8976 7182
rect 8994 7164 9014 7182
rect 8858 7143 9014 7164
rect 8858 7142 8958 7143
rect 4482 7071 4633 7094
rect 4482 7056 4597 7071
rect 205 6943 266 6959
rect 110 6939 266 6943
rect 110 6921 228 6939
rect 246 6921 266 6939
rect 4576 7053 4597 7056
rect 4615 7053 4633 7071
rect 4576 7034 4633 7053
rect 8859 7106 8901 7142
rect 12888 7213 12949 7229
rect 13317 7199 13378 7215
rect 17365 7286 17407 7322
rect 17308 7285 17408 7286
rect 17252 7264 17408 7285
rect 17252 7246 17272 7264
rect 17290 7246 17408 7264
rect 17252 7242 17408 7246
rect 13222 7195 13378 7199
rect 13222 7177 13340 7195
rect 13358 7177 13378 7195
rect 13222 7156 13378 7177
rect 13222 7155 13322 7156
rect 8859 7083 9010 7106
rect 8859 7068 8974 7083
rect 4146 7001 4203 7020
rect 4146 6983 4164 7001
rect 4182 6998 4203 7001
rect 4182 6983 4297 6998
rect 110 6900 266 6921
rect 110 6899 210 6900
rect 111 6863 153 6899
rect 111 6840 262 6863
rect 4146 6960 4297 6983
rect 4255 6924 4297 6960
rect 4569 6956 4630 6972
rect 4474 6952 4630 6956
rect 4474 6934 4592 6952
rect 4610 6934 4630 6952
rect 8953 7065 8974 7068
rect 8992 7065 9010 7083
rect 8953 7046 9010 7065
rect 13223 7119 13265 7155
rect 17252 7226 17313 7242
rect 13223 7096 13374 7119
rect 13223 7081 13338 7096
rect 8510 7014 8567 7033
rect 8510 6996 8528 7014
rect 8546 7011 8567 7014
rect 8546 6996 8661 7011
rect 4198 6923 4298 6924
rect 4142 6902 4298 6923
rect 4474 6913 4630 6934
rect 4474 6912 4574 6913
rect 4142 6884 4162 6902
rect 4180 6884 4298 6902
rect 4142 6880 4298 6884
rect 4142 6864 4203 6880
rect 4475 6876 4517 6912
rect 111 6825 226 6840
rect 205 6822 226 6825
rect 244 6822 262 6840
rect 205 6803 262 6822
rect 4475 6853 4626 6876
rect 8510 6973 8661 6996
rect 8619 6937 8661 6973
rect 8946 6968 9007 6984
rect 8851 6964 9007 6968
rect 8851 6946 8969 6964
rect 8987 6946 9007 6964
rect 13317 7078 13338 7081
rect 13356 7078 13374 7096
rect 13317 7059 13374 7078
rect 12887 7026 12944 7045
rect 12887 7008 12905 7026
rect 12923 7023 12944 7026
rect 12923 7008 13038 7023
rect 8562 6936 8662 6937
rect 8506 6915 8662 6936
rect 8851 6925 9007 6946
rect 8851 6924 8951 6925
rect 8506 6897 8526 6915
rect 8544 6897 8662 6915
rect 8506 6893 8662 6897
rect 8506 6877 8567 6893
rect 8852 6888 8894 6924
rect 4475 6838 4590 6853
rect 4569 6835 4590 6838
rect 4608 6835 4626 6853
rect 4569 6816 4626 6835
rect 8852 6865 9003 6888
rect 12887 6985 13038 7008
rect 12996 6949 13038 6985
rect 13310 6981 13371 6997
rect 13215 6977 13371 6981
rect 13215 6959 13333 6977
rect 13351 6959 13371 6977
rect 17251 7039 17308 7058
rect 17251 7021 17269 7039
rect 17287 7036 17308 7039
rect 17287 7021 17402 7036
rect 12939 6948 13039 6949
rect 12883 6927 13039 6948
rect 13215 6938 13371 6959
rect 13215 6937 13315 6938
rect 12883 6909 12903 6927
rect 12921 6909 13039 6927
rect 12883 6905 13039 6909
rect 12883 6889 12944 6905
rect 13216 6901 13258 6937
rect 8852 6850 8967 6865
rect 8946 6847 8967 6850
rect 8985 6847 9003 6865
rect 8946 6828 9003 6847
rect 13216 6878 13367 6901
rect 17251 6998 17402 7021
rect 17360 6962 17402 6998
rect 17303 6961 17403 6962
rect 17247 6940 17403 6961
rect 17247 6922 17267 6940
rect 17285 6922 17403 6940
rect 17247 6918 17403 6922
rect 17247 6902 17308 6918
rect 13216 6863 13331 6878
rect 13310 6860 13331 6863
rect 13349 6860 13367 6878
rect 13310 6841 13367 6860
rect 4144 6708 4201 6727
rect 4144 6690 4162 6708
rect 4180 6705 4201 6708
rect 4180 6690 4295 6705
rect 203 6650 264 6666
rect 108 6646 264 6650
rect 108 6628 226 6646
rect 244 6628 264 6646
rect 108 6607 264 6628
rect 108 6606 208 6607
rect 109 6570 151 6606
rect 109 6547 260 6570
rect 4144 6667 4295 6690
rect 8508 6721 8565 6740
rect 8508 6703 8526 6721
rect 8544 6718 8565 6721
rect 8544 6703 8659 6718
rect 4253 6631 4295 6667
rect 4567 6663 4628 6679
rect 4472 6659 4628 6663
rect 4472 6641 4590 6659
rect 4608 6641 4628 6659
rect 4196 6630 4296 6631
rect 4140 6609 4296 6630
rect 4472 6620 4628 6641
rect 4472 6619 4572 6620
rect 109 6532 224 6547
rect 203 6529 224 6532
rect 242 6529 260 6547
rect 203 6510 260 6529
rect 4140 6591 4160 6609
rect 4178 6591 4296 6609
rect 4140 6587 4296 6591
rect 4140 6571 4201 6587
rect 4473 6583 4515 6619
rect 4473 6560 4624 6583
rect 8508 6680 8659 6703
rect 12885 6733 12942 6752
rect 12885 6715 12903 6733
rect 12921 6730 12942 6733
rect 12921 6715 13036 6730
rect 8617 6644 8659 6680
rect 8944 6675 9005 6691
rect 8849 6671 9005 6675
rect 8849 6653 8967 6671
rect 8985 6653 9005 6671
rect 8560 6643 8660 6644
rect 8504 6622 8660 6643
rect 8849 6632 9005 6653
rect 8849 6631 8949 6632
rect 4473 6545 4588 6560
rect 4567 6542 4588 6545
rect 4606 6542 4624 6560
rect 4567 6523 4624 6542
rect 4137 6490 4194 6509
rect 4137 6472 4155 6490
rect 4173 6487 4194 6490
rect 8504 6604 8524 6622
rect 8542 6604 8660 6622
rect 8504 6600 8660 6604
rect 8504 6584 8565 6600
rect 8850 6595 8892 6631
rect 8850 6572 9001 6595
rect 12885 6692 13036 6715
rect 17249 6746 17306 6765
rect 17249 6728 17267 6746
rect 17285 6743 17306 6746
rect 17285 6728 17400 6743
rect 12994 6656 13036 6692
rect 13308 6688 13369 6704
rect 13213 6684 13369 6688
rect 13213 6666 13331 6684
rect 13349 6666 13369 6684
rect 12937 6655 13037 6656
rect 12881 6634 13037 6655
rect 13213 6645 13369 6666
rect 13213 6644 13313 6645
rect 8850 6557 8965 6572
rect 8944 6554 8965 6557
rect 8983 6554 9001 6572
rect 8944 6535 9001 6554
rect 4173 6472 4288 6487
rect 4137 6449 4288 6472
rect 198 6326 259 6342
rect 4246 6413 4288 6449
rect 8501 6503 8558 6522
rect 8501 6485 8519 6503
rect 8537 6500 8558 6503
rect 12881 6616 12901 6634
rect 12919 6616 13037 6634
rect 12881 6612 13037 6616
rect 12881 6596 12942 6612
rect 13214 6608 13256 6644
rect 13214 6585 13365 6608
rect 17249 6705 17400 6728
rect 17358 6669 17400 6705
rect 17301 6668 17401 6669
rect 17245 6647 17401 6668
rect 13214 6570 13329 6585
rect 13308 6567 13329 6570
rect 13347 6567 13365 6585
rect 13308 6548 13365 6567
rect 8537 6485 8652 6500
rect 8501 6462 8652 6485
rect 4189 6412 4289 6413
rect 4133 6391 4289 6412
rect 4133 6373 4153 6391
rect 4171 6373 4289 6391
rect 4133 6369 4289 6373
rect 103 6322 259 6326
rect 103 6304 221 6322
rect 239 6304 259 6322
rect 103 6283 259 6304
rect 103 6282 203 6283
rect 104 6246 146 6282
rect 4133 6353 4194 6369
rect 4562 6339 4623 6355
rect 8610 6426 8652 6462
rect 12878 6515 12935 6534
rect 12878 6497 12896 6515
rect 12914 6512 12935 6515
rect 17245 6629 17265 6647
rect 17283 6629 17401 6647
rect 17245 6625 17401 6629
rect 17245 6609 17306 6625
rect 12914 6497 13029 6512
rect 12878 6474 13029 6497
rect 8553 6425 8653 6426
rect 8497 6404 8653 6425
rect 8497 6386 8517 6404
rect 8535 6386 8653 6404
rect 8497 6382 8653 6386
rect 4467 6335 4623 6339
rect 4131 6307 4188 6326
rect 104 6223 255 6246
rect 104 6208 219 6223
rect 198 6205 219 6208
rect 237 6205 255 6223
rect 4131 6289 4149 6307
rect 4167 6304 4188 6307
rect 4467 6317 4585 6335
rect 4603 6317 4623 6335
rect 4167 6289 4282 6304
rect 4467 6296 4623 6317
rect 4467 6295 4567 6296
rect 4131 6266 4282 6289
rect 198 6186 255 6205
rect 192 6143 253 6159
rect 4240 6230 4282 6266
rect 4468 6259 4510 6295
rect 8497 6366 8558 6382
rect 8939 6351 9000 6367
rect 12987 6438 13029 6474
rect 17242 6528 17299 6547
rect 17242 6510 17260 6528
rect 17278 6525 17299 6528
rect 17278 6510 17393 6525
rect 17242 6487 17393 6510
rect 12930 6437 13030 6438
rect 12874 6416 13030 6437
rect 12874 6398 12894 6416
rect 12912 6398 13030 6416
rect 12874 6394 13030 6398
rect 8844 6347 9000 6351
rect 8495 6320 8552 6339
rect 4468 6236 4619 6259
rect 4183 6229 4283 6230
rect 4127 6208 4283 6229
rect 4468 6221 4583 6236
rect 4127 6190 4147 6208
rect 4165 6190 4283 6208
rect 4562 6218 4583 6221
rect 4601 6218 4619 6236
rect 8495 6302 8513 6320
rect 8531 6317 8552 6320
rect 8844 6329 8962 6347
rect 8980 6329 9000 6347
rect 8531 6302 8646 6317
rect 8844 6308 9000 6329
rect 8844 6307 8944 6308
rect 8495 6279 8646 6302
rect 4562 6199 4619 6218
rect 4127 6186 4283 6190
rect 97 6139 253 6143
rect 97 6121 215 6139
rect 233 6121 253 6139
rect 97 6100 253 6121
rect 97 6099 197 6100
rect 98 6063 140 6099
rect 4127 6170 4188 6186
rect 4556 6156 4617 6172
rect 8604 6243 8646 6279
rect 8845 6271 8887 6307
rect 12874 6378 12935 6394
rect 13303 6364 13364 6380
rect 17351 6451 17393 6487
rect 17294 6450 17394 6451
rect 17238 6429 17394 6450
rect 17238 6411 17258 6429
rect 17276 6411 17394 6429
rect 17238 6407 17394 6411
rect 13208 6360 13364 6364
rect 12872 6332 12929 6351
rect 8845 6248 8996 6271
rect 8547 6242 8647 6243
rect 8491 6221 8647 6242
rect 8845 6233 8960 6248
rect 8491 6203 8511 6221
rect 8529 6203 8647 6221
rect 8939 6230 8960 6233
rect 8978 6230 8996 6248
rect 12872 6314 12890 6332
rect 12908 6329 12929 6332
rect 13208 6342 13326 6360
rect 13344 6342 13364 6360
rect 12908 6314 13023 6329
rect 13208 6321 13364 6342
rect 13208 6320 13308 6321
rect 12872 6291 13023 6314
rect 8939 6211 8996 6230
rect 8491 6199 8647 6203
rect 4461 6152 4617 6156
rect 4461 6134 4579 6152
rect 4597 6134 4617 6152
rect 4461 6113 4617 6134
rect 4461 6112 4561 6113
rect 98 6040 249 6063
rect 98 6025 213 6040
rect 192 6022 213 6025
rect 231 6022 249 6040
rect 192 6003 249 6022
rect 4462 6076 4504 6112
rect 8491 6183 8552 6199
rect 8933 6168 8994 6184
rect 12981 6255 13023 6291
rect 13209 6284 13251 6320
rect 17238 6391 17299 6407
rect 17236 6345 17293 6364
rect 13209 6261 13360 6284
rect 12924 6254 13024 6255
rect 12868 6233 13024 6254
rect 13209 6246 13324 6261
rect 12868 6215 12888 6233
rect 12906 6215 13024 6233
rect 13303 6243 13324 6246
rect 13342 6243 13360 6261
rect 17236 6327 17254 6345
rect 17272 6342 17293 6345
rect 17272 6327 17387 6342
rect 17236 6304 17387 6327
rect 13303 6224 13360 6243
rect 12868 6211 13024 6215
rect 8838 6164 8994 6168
rect 8838 6146 8956 6164
rect 8974 6146 8994 6164
rect 8838 6125 8994 6146
rect 8838 6124 8938 6125
rect 4462 6053 4613 6076
rect 4462 6038 4577 6053
rect 4556 6035 4577 6038
rect 4595 6035 4613 6053
rect 185 5925 246 5941
rect 90 5921 246 5925
rect 90 5903 208 5921
rect 226 5903 246 5921
rect 4556 6016 4613 6035
rect 8839 6088 8881 6124
rect 12868 6195 12929 6211
rect 13297 6181 13358 6197
rect 17345 6268 17387 6304
rect 17288 6267 17388 6268
rect 17232 6246 17388 6267
rect 17232 6228 17252 6246
rect 17270 6228 17388 6246
rect 17232 6224 17388 6228
rect 13202 6177 13358 6181
rect 13202 6159 13320 6177
rect 13338 6159 13358 6177
rect 13202 6138 13358 6159
rect 13202 6137 13302 6138
rect 8839 6065 8990 6088
rect 8839 6050 8954 6065
rect 4126 5983 4183 6002
rect 4126 5965 4144 5983
rect 4162 5980 4183 5983
rect 4162 5965 4277 5980
rect 90 5882 246 5903
rect 90 5881 190 5882
rect 91 5845 133 5881
rect 91 5822 242 5845
rect 4126 5942 4277 5965
rect 4235 5906 4277 5942
rect 4549 5938 4610 5954
rect 4454 5934 4610 5938
rect 4454 5916 4572 5934
rect 4590 5916 4610 5934
rect 8933 6047 8954 6050
rect 8972 6047 8990 6065
rect 8933 6028 8990 6047
rect 13203 6101 13245 6137
rect 17232 6208 17293 6224
rect 13203 6078 13354 6101
rect 13203 6063 13318 6078
rect 13297 6060 13318 6063
rect 13336 6060 13354 6078
rect 8490 5996 8547 6015
rect 8490 5978 8508 5996
rect 8526 5993 8547 5996
rect 8526 5978 8641 5993
rect 4178 5905 4278 5906
rect 4122 5884 4278 5905
rect 4454 5895 4610 5916
rect 4454 5894 4554 5895
rect 4122 5866 4142 5884
rect 4160 5866 4278 5884
rect 4122 5862 4278 5866
rect 4122 5846 4183 5862
rect 4455 5858 4497 5894
rect 91 5807 206 5822
rect 185 5804 206 5807
rect 224 5804 242 5822
rect 185 5785 242 5804
rect 4455 5835 4606 5858
rect 8490 5955 8641 5978
rect 8599 5919 8641 5955
rect 8926 5950 8987 5966
rect 8831 5946 8987 5950
rect 8831 5928 8949 5946
rect 8967 5928 8987 5946
rect 13297 6041 13354 6060
rect 12867 6008 12924 6027
rect 12867 5990 12885 6008
rect 12903 6005 12924 6008
rect 12903 5990 13018 6005
rect 8542 5918 8642 5919
rect 8486 5897 8642 5918
rect 8831 5907 8987 5928
rect 8831 5906 8931 5907
rect 8486 5879 8506 5897
rect 8524 5879 8642 5897
rect 8486 5875 8642 5879
rect 8486 5859 8547 5875
rect 8832 5870 8874 5906
rect 4455 5820 4570 5835
rect 4549 5817 4570 5820
rect 4588 5817 4606 5835
rect 4549 5798 4606 5817
rect 8832 5847 8983 5870
rect 12867 5967 13018 5990
rect 12976 5931 13018 5967
rect 13290 5963 13351 5979
rect 13195 5959 13351 5963
rect 13195 5941 13313 5959
rect 13331 5941 13351 5959
rect 17231 6021 17288 6040
rect 17231 6003 17249 6021
rect 17267 6018 17288 6021
rect 17267 6003 17382 6018
rect 12919 5930 13019 5931
rect 12863 5909 13019 5930
rect 13195 5920 13351 5941
rect 13195 5919 13295 5920
rect 12863 5891 12883 5909
rect 12901 5891 13019 5909
rect 12863 5887 13019 5891
rect 12863 5871 12924 5887
rect 13196 5883 13238 5919
rect 8832 5832 8947 5847
rect 8926 5829 8947 5832
rect 8965 5829 8983 5847
rect 8926 5810 8983 5829
rect 13196 5860 13347 5883
rect 17231 5980 17382 6003
rect 17340 5944 17382 5980
rect 17283 5943 17383 5944
rect 17227 5922 17383 5943
rect 17227 5904 17247 5922
rect 17265 5904 17383 5922
rect 17227 5900 17383 5904
rect 17227 5884 17288 5900
rect 13196 5845 13311 5860
rect 13290 5842 13311 5845
rect 13329 5842 13347 5860
rect 13290 5823 13347 5842
rect 4127 5690 4184 5709
rect 4127 5672 4145 5690
rect 4163 5687 4184 5690
rect 4163 5672 4278 5687
rect 186 5632 247 5648
rect 91 5628 247 5632
rect 91 5610 209 5628
rect 227 5610 247 5628
rect 91 5589 247 5610
rect 91 5588 191 5589
rect 92 5552 134 5588
rect 92 5529 243 5552
rect 4127 5649 4278 5672
rect 8491 5703 8548 5722
rect 8491 5685 8509 5703
rect 8527 5700 8548 5703
rect 8527 5685 8642 5700
rect 4236 5613 4278 5649
rect 4550 5645 4611 5661
rect 4455 5641 4611 5645
rect 4455 5623 4573 5641
rect 4591 5623 4611 5641
rect 4179 5612 4279 5613
rect 4123 5591 4279 5612
rect 4455 5602 4611 5623
rect 4455 5601 4555 5602
rect 92 5514 207 5529
rect 186 5511 207 5514
rect 225 5511 243 5529
rect 186 5492 243 5511
rect 4123 5573 4143 5591
rect 4161 5573 4279 5591
rect 4123 5569 4279 5573
rect 4123 5553 4184 5569
rect 4456 5565 4498 5601
rect 4456 5542 4607 5565
rect 8491 5662 8642 5685
rect 12868 5715 12925 5734
rect 12868 5697 12886 5715
rect 12904 5712 12925 5715
rect 12904 5697 13019 5712
rect 8600 5626 8642 5662
rect 8927 5657 8988 5673
rect 8832 5653 8988 5657
rect 8832 5635 8950 5653
rect 8968 5635 8988 5653
rect 8543 5625 8643 5626
rect 8487 5604 8643 5625
rect 8832 5614 8988 5635
rect 8832 5613 8932 5614
rect 4456 5527 4571 5542
rect 4550 5524 4571 5527
rect 4589 5524 4607 5542
rect 4550 5505 4607 5524
rect 4120 5472 4177 5491
rect 8487 5586 8507 5604
rect 8525 5586 8643 5604
rect 8487 5582 8643 5586
rect 8487 5566 8548 5582
rect 8833 5577 8875 5613
rect 8833 5554 8984 5577
rect 12868 5674 13019 5697
rect 17232 5728 17289 5747
rect 17232 5710 17250 5728
rect 17268 5725 17289 5728
rect 17268 5710 17383 5725
rect 12977 5638 13019 5674
rect 13291 5670 13352 5686
rect 13196 5666 13352 5670
rect 13196 5648 13314 5666
rect 13332 5648 13352 5666
rect 12920 5637 13020 5638
rect 12864 5616 13020 5637
rect 13196 5627 13352 5648
rect 13196 5626 13296 5627
rect 8833 5539 8948 5554
rect 8927 5536 8948 5539
rect 8966 5536 8984 5554
rect 8927 5517 8984 5536
rect 4120 5454 4138 5472
rect 4156 5469 4177 5472
rect 4156 5454 4271 5469
rect 4120 5431 4271 5454
rect 181 5308 242 5324
rect 4229 5395 4271 5431
rect 8484 5485 8541 5504
rect 8484 5467 8502 5485
rect 8520 5482 8541 5485
rect 12864 5598 12884 5616
rect 12902 5598 13020 5616
rect 12864 5594 13020 5598
rect 12864 5578 12925 5594
rect 13197 5590 13239 5626
rect 13197 5567 13348 5590
rect 17232 5687 17383 5710
rect 17341 5651 17383 5687
rect 17284 5650 17384 5651
rect 17228 5629 17384 5650
rect 13197 5552 13312 5567
rect 13291 5549 13312 5552
rect 13330 5549 13348 5567
rect 13291 5530 13348 5549
rect 8520 5467 8635 5482
rect 8484 5444 8635 5467
rect 4172 5394 4272 5395
rect 4116 5373 4272 5394
rect 4116 5355 4136 5373
rect 4154 5355 4272 5373
rect 4116 5351 4272 5355
rect 86 5304 242 5308
rect 86 5286 204 5304
rect 222 5286 242 5304
rect 86 5265 242 5286
rect 86 5264 186 5265
rect 87 5228 129 5264
rect 4116 5335 4177 5351
rect 4545 5321 4606 5337
rect 8593 5408 8635 5444
rect 12861 5497 12918 5516
rect 17228 5611 17248 5629
rect 17266 5611 17384 5629
rect 17228 5607 17384 5611
rect 17228 5591 17289 5607
rect 12861 5479 12879 5497
rect 12897 5494 12918 5497
rect 12897 5479 13012 5494
rect 12861 5456 13012 5479
rect 8536 5407 8636 5408
rect 8480 5386 8636 5407
rect 8480 5368 8500 5386
rect 8518 5368 8636 5386
rect 8480 5364 8636 5368
rect 4450 5317 4606 5321
rect 4114 5289 4171 5308
rect 87 5205 238 5228
rect 87 5190 202 5205
rect 181 5187 202 5190
rect 220 5187 238 5205
rect 4114 5271 4132 5289
rect 4150 5286 4171 5289
rect 4450 5299 4568 5317
rect 4586 5299 4606 5317
rect 4150 5271 4265 5286
rect 4450 5278 4606 5299
rect 4450 5277 4550 5278
rect 4114 5248 4265 5271
rect 181 5168 238 5187
rect 175 5125 236 5141
rect 4223 5212 4265 5248
rect 4451 5241 4493 5277
rect 8480 5348 8541 5364
rect 8922 5333 8983 5349
rect 12970 5420 13012 5456
rect 17225 5510 17282 5529
rect 17225 5492 17243 5510
rect 17261 5507 17282 5510
rect 17261 5492 17376 5507
rect 17225 5469 17376 5492
rect 12913 5419 13013 5420
rect 12857 5398 13013 5419
rect 12857 5380 12877 5398
rect 12895 5380 13013 5398
rect 12857 5376 13013 5380
rect 8827 5329 8983 5333
rect 8478 5302 8535 5321
rect 4451 5218 4602 5241
rect 4166 5211 4266 5212
rect 4110 5190 4266 5211
rect 4451 5203 4566 5218
rect 4110 5172 4130 5190
rect 4148 5172 4266 5190
rect 4545 5200 4566 5203
rect 4584 5200 4602 5218
rect 8478 5284 8496 5302
rect 8514 5299 8535 5302
rect 8827 5311 8945 5329
rect 8963 5311 8983 5329
rect 8514 5284 8629 5299
rect 8827 5290 8983 5311
rect 8827 5289 8927 5290
rect 8478 5261 8629 5284
rect 4545 5181 4602 5200
rect 4110 5168 4266 5172
rect 80 5121 236 5125
rect 80 5103 198 5121
rect 216 5103 236 5121
rect 80 5082 236 5103
rect 80 5081 180 5082
rect 81 5045 123 5081
rect 4110 5152 4171 5168
rect 4539 5138 4600 5154
rect 8587 5225 8629 5261
rect 8828 5253 8870 5289
rect 12857 5360 12918 5376
rect 13286 5346 13347 5362
rect 17334 5433 17376 5469
rect 17277 5432 17377 5433
rect 17221 5411 17377 5432
rect 17221 5393 17241 5411
rect 17259 5393 17377 5411
rect 17221 5389 17377 5393
rect 13191 5342 13347 5346
rect 12855 5314 12912 5333
rect 8828 5230 8979 5253
rect 8530 5224 8630 5225
rect 8474 5203 8630 5224
rect 8828 5215 8943 5230
rect 8474 5185 8494 5203
rect 8512 5185 8630 5203
rect 8922 5212 8943 5215
rect 8961 5212 8979 5230
rect 12855 5296 12873 5314
rect 12891 5311 12912 5314
rect 13191 5324 13309 5342
rect 13327 5324 13347 5342
rect 12891 5296 13006 5311
rect 13191 5303 13347 5324
rect 13191 5302 13291 5303
rect 12855 5273 13006 5296
rect 8922 5193 8979 5212
rect 8474 5181 8630 5185
rect 4444 5134 4600 5138
rect 4444 5116 4562 5134
rect 4580 5116 4600 5134
rect 4444 5095 4600 5116
rect 4444 5094 4544 5095
rect 81 5022 232 5045
rect 81 5007 196 5022
rect 175 5004 196 5007
rect 214 5004 232 5022
rect 175 4985 232 5004
rect 4445 5058 4487 5094
rect 8474 5165 8535 5181
rect 8916 5150 8977 5166
rect 12964 5237 13006 5273
rect 13192 5266 13234 5302
rect 17221 5373 17282 5389
rect 17219 5327 17276 5346
rect 13192 5243 13343 5266
rect 12907 5236 13007 5237
rect 12851 5215 13007 5236
rect 13192 5228 13307 5243
rect 12851 5197 12871 5215
rect 12889 5197 13007 5215
rect 13286 5225 13307 5228
rect 13325 5225 13343 5243
rect 17219 5309 17237 5327
rect 17255 5324 17276 5327
rect 17255 5309 17370 5324
rect 17219 5286 17370 5309
rect 13286 5206 13343 5225
rect 12851 5193 13007 5197
rect 8821 5146 8977 5150
rect 8821 5128 8939 5146
rect 8957 5128 8977 5146
rect 8821 5107 8977 5128
rect 8821 5106 8921 5107
rect 4445 5035 4596 5058
rect 168 4907 229 4923
rect 73 4903 229 4907
rect 73 4885 191 4903
rect 209 4885 229 4903
rect 4445 5020 4560 5035
rect 4539 5017 4560 5020
rect 4578 5017 4596 5035
rect 4539 4998 4596 5017
rect 8822 5070 8864 5106
rect 12851 5177 12912 5193
rect 13280 5163 13341 5179
rect 17328 5250 17370 5286
rect 17271 5249 17371 5250
rect 17215 5228 17371 5249
rect 17215 5210 17235 5228
rect 17253 5210 17371 5228
rect 17215 5206 17371 5210
rect 13185 5159 13341 5163
rect 13185 5141 13303 5159
rect 13321 5141 13341 5159
rect 13185 5120 13341 5141
rect 13185 5119 13285 5120
rect 8822 5047 8973 5070
rect 4109 4965 4166 4984
rect 4109 4947 4127 4965
rect 4145 4962 4166 4965
rect 4145 4947 4260 4962
rect 73 4864 229 4885
rect 73 4863 173 4864
rect 74 4827 116 4863
rect 74 4804 225 4827
rect 4109 4924 4260 4947
rect 4218 4888 4260 4924
rect 4532 4920 4593 4936
rect 4437 4916 4593 4920
rect 4437 4898 4555 4916
rect 4573 4898 4593 4916
rect 8822 5032 8937 5047
rect 8916 5029 8937 5032
rect 8955 5029 8973 5047
rect 8916 5010 8973 5029
rect 13186 5083 13228 5119
rect 17215 5190 17276 5206
rect 13186 5060 13337 5083
rect 8473 4978 8530 4997
rect 8473 4960 8491 4978
rect 8509 4975 8530 4978
rect 8509 4960 8624 4975
rect 4161 4887 4261 4888
rect 4105 4866 4261 4887
rect 4437 4877 4593 4898
rect 4437 4876 4537 4877
rect 4105 4848 4125 4866
rect 4143 4848 4261 4866
rect 4105 4844 4261 4848
rect 4105 4828 4166 4844
rect 4438 4840 4480 4876
rect 74 4789 189 4804
rect 168 4786 189 4789
rect 207 4786 225 4804
rect 168 4767 225 4786
rect 4438 4817 4589 4840
rect 8473 4937 8624 4960
rect 8582 4901 8624 4937
rect 8909 4932 8970 4948
rect 8814 4928 8970 4932
rect 8814 4910 8932 4928
rect 8950 4910 8970 4928
rect 13186 5045 13301 5060
rect 13280 5042 13301 5045
rect 13319 5042 13337 5060
rect 13280 5023 13337 5042
rect 12850 4990 12907 5009
rect 12850 4972 12868 4990
rect 12886 4987 12907 4990
rect 12886 4972 13001 4987
rect 8525 4900 8625 4901
rect 8469 4879 8625 4900
rect 8814 4889 8970 4910
rect 8814 4888 8914 4889
rect 8469 4861 8489 4879
rect 8507 4861 8625 4879
rect 8469 4857 8625 4861
rect 8469 4841 8530 4857
rect 8815 4852 8857 4888
rect 4438 4802 4553 4817
rect 4532 4799 4553 4802
rect 4571 4799 4589 4817
rect 4532 4780 4589 4799
rect 8815 4829 8966 4852
rect 12850 4949 13001 4972
rect 12959 4913 13001 4949
rect 13273 4945 13334 4961
rect 13178 4941 13334 4945
rect 13178 4923 13296 4941
rect 13314 4923 13334 4941
rect 17214 5003 17271 5022
rect 17214 4985 17232 5003
rect 17250 5000 17271 5003
rect 17250 4985 17365 5000
rect 12902 4912 13002 4913
rect 12846 4891 13002 4912
rect 13178 4902 13334 4923
rect 13178 4901 13278 4902
rect 12846 4873 12866 4891
rect 12884 4873 13002 4891
rect 12846 4869 13002 4873
rect 12846 4853 12907 4869
rect 13179 4865 13221 4901
rect 8815 4814 8930 4829
rect 8909 4811 8930 4814
rect 8948 4811 8966 4829
rect 8909 4792 8966 4811
rect 13179 4842 13330 4865
rect 17214 4962 17365 4985
rect 17323 4926 17365 4962
rect 17266 4925 17366 4926
rect 17210 4904 17366 4925
rect 17210 4886 17230 4904
rect 17248 4886 17366 4904
rect 17210 4882 17366 4886
rect 17210 4866 17271 4882
rect 13179 4827 13294 4842
rect 13273 4824 13294 4827
rect 13312 4824 13330 4842
rect 13273 4805 13330 4824
rect 4108 4672 4165 4691
rect 4108 4654 4126 4672
rect 4144 4669 4165 4672
rect 4144 4654 4259 4669
rect 167 4614 228 4630
rect 72 4610 228 4614
rect 72 4592 190 4610
rect 208 4592 228 4610
rect 72 4571 228 4592
rect 72 4570 172 4571
rect 73 4534 115 4570
rect 73 4511 224 4534
rect 4108 4631 4259 4654
rect 8472 4685 8529 4704
rect 8472 4667 8490 4685
rect 8508 4682 8529 4685
rect 8508 4667 8623 4682
rect 4217 4595 4259 4631
rect 4531 4627 4592 4643
rect 4436 4623 4592 4627
rect 4436 4605 4554 4623
rect 4572 4605 4592 4623
rect 4160 4594 4260 4595
rect 4104 4573 4260 4594
rect 4436 4584 4592 4605
rect 4436 4583 4536 4584
rect 73 4496 188 4511
rect 167 4493 188 4496
rect 206 4493 224 4511
rect 167 4474 224 4493
rect 4104 4555 4124 4573
rect 4142 4555 4260 4573
rect 4104 4551 4260 4555
rect 4104 4535 4165 4551
rect 4437 4547 4479 4583
rect 4437 4524 4588 4547
rect 8472 4644 8623 4667
rect 12849 4697 12906 4716
rect 12849 4679 12867 4697
rect 12885 4694 12906 4697
rect 12885 4679 13000 4694
rect 8581 4608 8623 4644
rect 8908 4639 8969 4655
rect 8813 4635 8969 4639
rect 8813 4617 8931 4635
rect 8949 4617 8969 4635
rect 8524 4607 8624 4608
rect 8468 4586 8624 4607
rect 8813 4596 8969 4617
rect 8813 4595 8913 4596
rect 4437 4509 4552 4524
rect 4531 4506 4552 4509
rect 4570 4506 4588 4524
rect 4531 4487 4588 4506
rect 4101 4454 4158 4473
rect 4101 4436 4119 4454
rect 4137 4451 4158 4454
rect 4137 4436 4252 4451
rect 8468 4568 8488 4586
rect 8506 4568 8624 4586
rect 8468 4564 8624 4568
rect 8468 4548 8529 4564
rect 8814 4559 8856 4595
rect 8814 4536 8965 4559
rect 12849 4656 13000 4679
rect 17213 4710 17270 4729
rect 17213 4692 17231 4710
rect 17249 4707 17270 4710
rect 17249 4692 17364 4707
rect 12958 4620 13000 4656
rect 13272 4652 13333 4668
rect 13177 4648 13333 4652
rect 13177 4630 13295 4648
rect 13313 4630 13333 4648
rect 12901 4619 13001 4620
rect 12845 4598 13001 4619
rect 13177 4609 13333 4630
rect 13177 4608 13277 4609
rect 8814 4521 8929 4536
rect 8908 4518 8929 4521
rect 8947 4518 8965 4536
rect 8908 4499 8965 4518
rect 4101 4413 4252 4436
rect 162 4290 223 4306
rect 4210 4377 4252 4413
rect 8465 4467 8522 4486
rect 8465 4449 8483 4467
rect 8501 4464 8522 4467
rect 8501 4449 8616 4464
rect 12845 4580 12865 4598
rect 12883 4580 13001 4598
rect 12845 4576 13001 4580
rect 12845 4560 12906 4576
rect 13178 4572 13220 4608
rect 13178 4549 13329 4572
rect 17213 4669 17364 4692
rect 17322 4633 17364 4669
rect 17265 4632 17365 4633
rect 17209 4611 17365 4632
rect 13178 4534 13293 4549
rect 13272 4531 13293 4534
rect 13311 4531 13329 4549
rect 13272 4512 13329 4531
rect 8465 4426 8616 4449
rect 4153 4376 4253 4377
rect 4097 4355 4253 4376
rect 4097 4337 4117 4355
rect 4135 4337 4253 4355
rect 4097 4333 4253 4337
rect 67 4286 223 4290
rect 67 4268 185 4286
rect 203 4268 223 4286
rect 67 4247 223 4268
rect 67 4246 167 4247
rect 68 4210 110 4246
rect 4097 4317 4158 4333
rect 4526 4303 4587 4319
rect 8574 4390 8616 4426
rect 12842 4479 12899 4498
rect 12842 4461 12860 4479
rect 12878 4476 12899 4479
rect 12878 4461 12993 4476
rect 17209 4593 17229 4611
rect 17247 4593 17365 4611
rect 17209 4589 17365 4593
rect 17209 4573 17270 4589
rect 12842 4438 12993 4461
rect 8517 4389 8617 4390
rect 8461 4368 8617 4389
rect 8461 4350 8481 4368
rect 8499 4350 8617 4368
rect 8461 4346 8617 4350
rect 4431 4299 4587 4303
rect 4095 4271 4152 4290
rect 68 4187 219 4210
rect 68 4172 183 4187
rect 162 4169 183 4172
rect 201 4169 219 4187
rect 4095 4253 4113 4271
rect 4131 4268 4152 4271
rect 4431 4281 4549 4299
rect 4567 4281 4587 4299
rect 4131 4253 4246 4268
rect 4431 4260 4587 4281
rect 4431 4259 4531 4260
rect 4095 4230 4246 4253
rect 162 4150 219 4169
rect 156 4107 217 4123
rect 4204 4194 4246 4230
rect 4432 4223 4474 4259
rect 8461 4330 8522 4346
rect 8903 4315 8964 4331
rect 12951 4402 12993 4438
rect 17206 4492 17263 4511
rect 17206 4474 17224 4492
rect 17242 4489 17263 4492
rect 17242 4474 17357 4489
rect 17206 4451 17357 4474
rect 12894 4401 12994 4402
rect 12838 4380 12994 4401
rect 12838 4362 12858 4380
rect 12876 4362 12994 4380
rect 12838 4358 12994 4362
rect 8808 4311 8964 4315
rect 8459 4284 8516 4303
rect 4432 4200 4583 4223
rect 4147 4193 4247 4194
rect 4091 4172 4247 4193
rect 4432 4185 4547 4200
rect 4091 4154 4111 4172
rect 4129 4154 4247 4172
rect 4526 4182 4547 4185
rect 4565 4182 4583 4200
rect 8459 4266 8477 4284
rect 8495 4281 8516 4284
rect 8808 4293 8926 4311
rect 8944 4293 8964 4311
rect 8495 4266 8610 4281
rect 8808 4272 8964 4293
rect 8808 4271 8908 4272
rect 8459 4243 8610 4266
rect 4526 4163 4583 4182
rect 4091 4150 4247 4154
rect 61 4103 217 4107
rect 61 4085 179 4103
rect 197 4085 217 4103
rect 61 4064 217 4085
rect 61 4063 161 4064
rect 62 4027 104 4063
rect 4091 4134 4152 4150
rect 4520 4120 4581 4136
rect 8568 4207 8610 4243
rect 8809 4235 8851 4271
rect 12838 4342 12899 4358
rect 13267 4328 13328 4344
rect 17315 4415 17357 4451
rect 17258 4414 17358 4415
rect 17202 4393 17358 4414
rect 17202 4375 17222 4393
rect 17240 4375 17358 4393
rect 17202 4371 17358 4375
rect 13172 4324 13328 4328
rect 12836 4296 12893 4315
rect 8809 4212 8960 4235
rect 8511 4206 8611 4207
rect 8455 4185 8611 4206
rect 8809 4197 8924 4212
rect 8455 4167 8475 4185
rect 8493 4167 8611 4185
rect 8903 4194 8924 4197
rect 8942 4194 8960 4212
rect 12836 4278 12854 4296
rect 12872 4293 12893 4296
rect 13172 4306 13290 4324
rect 13308 4306 13328 4324
rect 12872 4278 12987 4293
rect 13172 4285 13328 4306
rect 13172 4284 13272 4285
rect 12836 4255 12987 4278
rect 8903 4175 8960 4194
rect 8455 4163 8611 4167
rect 4425 4116 4581 4120
rect 4425 4098 4543 4116
rect 4561 4098 4581 4116
rect 4425 4077 4581 4098
rect 4425 4076 4525 4077
rect 62 4004 213 4027
rect 62 3989 177 4004
rect 156 3986 177 3989
rect 195 3986 213 4004
rect 156 3967 213 3986
rect 4426 4040 4468 4076
rect 8455 4147 8516 4163
rect 8897 4132 8958 4148
rect 12945 4219 12987 4255
rect 13173 4248 13215 4284
rect 17202 4355 17263 4371
rect 17200 4309 17257 4328
rect 13173 4225 13324 4248
rect 12888 4218 12988 4219
rect 12832 4197 12988 4218
rect 13173 4210 13288 4225
rect 12832 4179 12852 4197
rect 12870 4179 12988 4197
rect 13267 4207 13288 4210
rect 13306 4207 13324 4225
rect 17200 4291 17218 4309
rect 17236 4306 17257 4309
rect 17236 4291 17351 4306
rect 17200 4268 17351 4291
rect 13267 4188 13324 4207
rect 12832 4175 12988 4179
rect 8802 4128 8958 4132
rect 8802 4110 8920 4128
rect 8938 4110 8958 4128
rect 8802 4089 8958 4110
rect 8802 4088 8902 4089
rect 4426 4017 4577 4040
rect 4426 4002 4541 4017
rect 4520 3999 4541 4002
rect 4559 3999 4577 4017
rect 149 3889 210 3905
rect 54 3885 210 3889
rect 54 3867 172 3885
rect 190 3867 210 3885
rect 4520 3980 4577 3999
rect 8803 4052 8845 4088
rect 12832 4159 12893 4175
rect 13261 4145 13322 4161
rect 17309 4232 17351 4268
rect 17252 4231 17352 4232
rect 17196 4210 17352 4231
rect 17196 4192 17216 4210
rect 17234 4192 17352 4210
rect 17196 4188 17352 4192
rect 13166 4141 13322 4145
rect 13166 4123 13284 4141
rect 13302 4123 13322 4141
rect 13166 4102 13322 4123
rect 13166 4101 13266 4102
rect 8803 4029 8954 4052
rect 8803 4014 8918 4029
rect 4090 3947 4147 3966
rect 4090 3929 4108 3947
rect 4126 3944 4147 3947
rect 4126 3929 4241 3944
rect 54 3846 210 3867
rect 54 3845 154 3846
rect 55 3809 97 3845
rect 55 3786 206 3809
rect 4090 3906 4241 3929
rect 4199 3870 4241 3906
rect 4513 3902 4574 3918
rect 4418 3898 4574 3902
rect 4418 3880 4536 3898
rect 4554 3880 4574 3898
rect 8897 4011 8918 4014
rect 8936 4011 8954 4029
rect 8897 3992 8954 4011
rect 13167 4065 13209 4101
rect 17196 4172 17257 4188
rect 13167 4042 13318 4065
rect 13167 4027 13282 4042
rect 13261 4024 13282 4027
rect 13300 4024 13318 4042
rect 8454 3960 8511 3979
rect 8454 3942 8472 3960
rect 8490 3957 8511 3960
rect 8490 3942 8605 3957
rect 4142 3869 4242 3870
rect 4086 3848 4242 3869
rect 4418 3859 4574 3880
rect 4418 3858 4518 3859
rect 4086 3830 4106 3848
rect 4124 3830 4242 3848
rect 4086 3826 4242 3830
rect 4086 3810 4147 3826
rect 4419 3822 4461 3858
rect 55 3771 170 3786
rect 149 3768 170 3771
rect 188 3768 206 3786
rect 149 3749 206 3768
rect 4419 3799 4570 3822
rect 8454 3919 8605 3942
rect 8563 3883 8605 3919
rect 8890 3914 8951 3930
rect 8795 3910 8951 3914
rect 8795 3892 8913 3910
rect 8931 3892 8951 3910
rect 13261 4005 13318 4024
rect 12831 3972 12888 3991
rect 12831 3954 12849 3972
rect 12867 3969 12888 3972
rect 12867 3954 12982 3969
rect 8506 3882 8606 3883
rect 8450 3861 8606 3882
rect 8795 3871 8951 3892
rect 8795 3870 8895 3871
rect 8450 3843 8470 3861
rect 8488 3843 8606 3861
rect 8450 3839 8606 3843
rect 8450 3823 8511 3839
rect 8796 3834 8838 3870
rect 4419 3784 4534 3799
rect 4513 3781 4534 3784
rect 4552 3781 4570 3799
rect 4513 3762 4570 3781
rect 8796 3811 8947 3834
rect 12831 3931 12982 3954
rect 12940 3895 12982 3931
rect 13254 3927 13315 3943
rect 13159 3923 13315 3927
rect 13159 3905 13277 3923
rect 13295 3905 13315 3923
rect 17195 3985 17252 4004
rect 17195 3967 17213 3985
rect 17231 3982 17252 3985
rect 17231 3967 17346 3982
rect 12883 3894 12983 3895
rect 12827 3873 12983 3894
rect 13159 3884 13315 3905
rect 13159 3883 13259 3884
rect 12827 3855 12847 3873
rect 12865 3855 12983 3873
rect 12827 3851 12983 3855
rect 12827 3835 12888 3851
rect 13160 3847 13202 3883
rect 8796 3796 8911 3811
rect 8890 3793 8911 3796
rect 8929 3793 8947 3811
rect 8890 3774 8947 3793
rect 13160 3824 13311 3847
rect 17195 3944 17346 3967
rect 17304 3908 17346 3944
rect 17247 3907 17347 3908
rect 17191 3886 17347 3907
rect 17191 3868 17211 3886
rect 17229 3868 17347 3886
rect 17191 3864 17347 3868
rect 17191 3848 17252 3864
rect 13160 3809 13275 3824
rect 13254 3806 13275 3809
rect 13293 3806 13311 3824
rect 13254 3787 13311 3806
rect 4091 3654 4148 3673
rect 4091 3636 4109 3654
rect 4127 3651 4148 3654
rect 4127 3636 4242 3651
rect 150 3596 211 3612
rect 55 3592 211 3596
rect 55 3574 173 3592
rect 191 3574 211 3592
rect 55 3553 211 3574
rect 55 3552 155 3553
rect 56 3516 98 3552
rect 56 3493 207 3516
rect 4091 3613 4242 3636
rect 8455 3667 8512 3686
rect 8455 3649 8473 3667
rect 8491 3664 8512 3667
rect 8491 3649 8606 3664
rect 4200 3577 4242 3613
rect 4514 3609 4575 3625
rect 4419 3605 4575 3609
rect 4419 3587 4537 3605
rect 4555 3587 4575 3605
rect 4143 3576 4243 3577
rect 4087 3555 4243 3576
rect 4419 3566 4575 3587
rect 4419 3565 4519 3566
rect 56 3478 171 3493
rect 150 3475 171 3478
rect 189 3475 207 3493
rect 150 3456 207 3475
rect 4087 3537 4107 3555
rect 4125 3537 4243 3555
rect 4087 3533 4243 3537
rect 4087 3517 4148 3533
rect 4420 3529 4462 3565
rect 4420 3506 4571 3529
rect 8455 3626 8606 3649
rect 12832 3679 12889 3698
rect 12832 3661 12850 3679
rect 12868 3676 12889 3679
rect 12868 3661 12983 3676
rect 8564 3590 8606 3626
rect 8891 3621 8952 3637
rect 8796 3617 8952 3621
rect 8796 3599 8914 3617
rect 8932 3599 8952 3617
rect 8507 3589 8607 3590
rect 8451 3568 8607 3589
rect 8796 3578 8952 3599
rect 8796 3577 8896 3578
rect 4420 3491 4535 3506
rect 4514 3488 4535 3491
rect 4553 3488 4571 3506
rect 4514 3469 4571 3488
rect 4084 3436 4141 3455
rect 8451 3550 8471 3568
rect 8489 3550 8607 3568
rect 8451 3546 8607 3550
rect 8451 3530 8512 3546
rect 8797 3541 8839 3577
rect 8797 3518 8948 3541
rect 12832 3638 12983 3661
rect 17196 3692 17253 3711
rect 17196 3674 17214 3692
rect 17232 3689 17253 3692
rect 17232 3674 17347 3689
rect 12941 3602 12983 3638
rect 13255 3634 13316 3650
rect 13160 3630 13316 3634
rect 13160 3612 13278 3630
rect 13296 3612 13316 3630
rect 12884 3601 12984 3602
rect 12828 3580 12984 3601
rect 13160 3591 13316 3612
rect 13160 3590 13260 3591
rect 8797 3503 8912 3518
rect 8891 3500 8912 3503
rect 8930 3500 8948 3518
rect 8891 3481 8948 3500
rect 4084 3418 4102 3436
rect 4120 3433 4141 3436
rect 4120 3418 4235 3433
rect 4084 3395 4235 3418
rect 145 3272 206 3288
rect 4193 3359 4235 3395
rect 8448 3449 8505 3468
rect 8448 3431 8466 3449
rect 8484 3446 8505 3449
rect 12828 3562 12848 3580
rect 12866 3562 12984 3580
rect 12828 3558 12984 3562
rect 12828 3542 12889 3558
rect 13161 3554 13203 3590
rect 13161 3531 13312 3554
rect 17196 3651 17347 3674
rect 17305 3615 17347 3651
rect 17248 3614 17348 3615
rect 17192 3593 17348 3614
rect 13161 3516 13276 3531
rect 13255 3513 13276 3516
rect 13294 3513 13312 3531
rect 13255 3494 13312 3513
rect 8484 3431 8599 3446
rect 8448 3408 8599 3431
rect 4136 3358 4236 3359
rect 4080 3337 4236 3358
rect 4080 3319 4100 3337
rect 4118 3319 4236 3337
rect 4080 3315 4236 3319
rect 50 3268 206 3272
rect 50 3250 168 3268
rect 186 3250 206 3268
rect 50 3229 206 3250
rect 50 3228 150 3229
rect 51 3192 93 3228
rect 4080 3299 4141 3315
rect 4509 3285 4570 3301
rect 8557 3372 8599 3408
rect 12825 3461 12882 3480
rect 17192 3575 17212 3593
rect 17230 3575 17348 3593
rect 17192 3571 17348 3575
rect 17192 3555 17253 3571
rect 12825 3443 12843 3461
rect 12861 3458 12882 3461
rect 12861 3443 12976 3458
rect 12825 3420 12976 3443
rect 8500 3371 8600 3372
rect 8444 3350 8600 3371
rect 8444 3332 8464 3350
rect 8482 3332 8600 3350
rect 8444 3328 8600 3332
rect 4414 3281 4570 3285
rect 4078 3253 4135 3272
rect 51 3169 202 3192
rect 51 3154 166 3169
rect 145 3151 166 3154
rect 184 3151 202 3169
rect 4078 3235 4096 3253
rect 4114 3250 4135 3253
rect 4414 3263 4532 3281
rect 4550 3263 4570 3281
rect 4114 3235 4229 3250
rect 4414 3242 4570 3263
rect 4414 3241 4514 3242
rect 4078 3212 4229 3235
rect 145 3132 202 3151
rect 139 3089 200 3105
rect 4187 3176 4229 3212
rect 4415 3205 4457 3241
rect 8444 3312 8505 3328
rect 8886 3297 8947 3313
rect 12934 3384 12976 3420
rect 17189 3474 17246 3493
rect 17189 3456 17207 3474
rect 17225 3471 17246 3474
rect 17225 3456 17340 3471
rect 17189 3433 17340 3456
rect 12877 3383 12977 3384
rect 12821 3362 12977 3383
rect 12821 3344 12841 3362
rect 12859 3344 12977 3362
rect 12821 3340 12977 3344
rect 8791 3293 8947 3297
rect 8442 3266 8499 3285
rect 4415 3182 4566 3205
rect 4130 3175 4230 3176
rect 4074 3154 4230 3175
rect 4415 3167 4530 3182
rect 4074 3136 4094 3154
rect 4112 3136 4230 3154
rect 4509 3164 4530 3167
rect 4548 3164 4566 3182
rect 8442 3248 8460 3266
rect 8478 3263 8499 3266
rect 8791 3275 8909 3293
rect 8927 3275 8947 3293
rect 8478 3248 8593 3263
rect 8791 3254 8947 3275
rect 8791 3253 8891 3254
rect 8442 3225 8593 3248
rect 4509 3145 4566 3164
rect 4074 3132 4230 3136
rect 44 3085 200 3089
rect 44 3067 162 3085
rect 180 3067 200 3085
rect 44 3046 200 3067
rect 44 3045 144 3046
rect 45 3009 87 3045
rect 4074 3116 4135 3132
rect 4503 3102 4564 3118
rect 8551 3189 8593 3225
rect 8792 3217 8834 3253
rect 12821 3324 12882 3340
rect 13250 3310 13311 3326
rect 17298 3397 17340 3433
rect 17241 3396 17341 3397
rect 17185 3375 17341 3396
rect 17185 3357 17205 3375
rect 17223 3357 17341 3375
rect 17185 3353 17341 3357
rect 13155 3306 13311 3310
rect 12819 3278 12876 3297
rect 8792 3194 8943 3217
rect 8494 3188 8594 3189
rect 8438 3167 8594 3188
rect 8792 3179 8907 3194
rect 8438 3149 8458 3167
rect 8476 3149 8594 3167
rect 8886 3176 8907 3179
rect 8925 3176 8943 3194
rect 12819 3260 12837 3278
rect 12855 3275 12876 3278
rect 13155 3288 13273 3306
rect 13291 3288 13311 3306
rect 12855 3260 12970 3275
rect 13155 3267 13311 3288
rect 13155 3266 13255 3267
rect 12819 3237 12970 3260
rect 8886 3157 8943 3176
rect 8438 3145 8594 3149
rect 4408 3098 4564 3102
rect 4408 3080 4526 3098
rect 4544 3080 4564 3098
rect 4408 3059 4564 3080
rect 4408 3058 4508 3059
rect 45 2986 196 3009
rect 45 2971 160 2986
rect 139 2968 160 2971
rect 178 2968 196 2986
rect 139 2949 196 2968
rect 4409 3022 4451 3058
rect 8438 3129 8499 3145
rect 8880 3114 8941 3130
rect 12928 3201 12970 3237
rect 13156 3230 13198 3266
rect 17185 3337 17246 3353
rect 17183 3291 17240 3310
rect 13156 3207 13307 3230
rect 12871 3200 12971 3201
rect 12815 3179 12971 3200
rect 13156 3192 13271 3207
rect 12815 3161 12835 3179
rect 12853 3161 12971 3179
rect 13250 3189 13271 3192
rect 13289 3189 13307 3207
rect 17183 3273 17201 3291
rect 17219 3288 17240 3291
rect 17219 3273 17334 3288
rect 17183 3250 17334 3273
rect 13250 3170 13307 3189
rect 12815 3157 12971 3161
rect 8785 3110 8941 3114
rect 8785 3092 8903 3110
rect 8921 3092 8941 3110
rect 8785 3071 8941 3092
rect 8785 3070 8885 3071
rect 4409 2999 4560 3022
rect 4409 2984 4524 2999
rect 132 2871 193 2887
rect 37 2867 193 2871
rect 37 2849 155 2867
rect 173 2849 193 2867
rect 4503 2981 4524 2984
rect 4542 2981 4560 2999
rect 4503 2962 4560 2981
rect 8786 3034 8828 3070
rect 12815 3141 12876 3157
rect 13244 3127 13305 3143
rect 17292 3214 17334 3250
rect 17235 3213 17335 3214
rect 17179 3192 17335 3213
rect 17179 3174 17199 3192
rect 17217 3174 17335 3192
rect 17179 3170 17335 3174
rect 13149 3123 13305 3127
rect 13149 3105 13267 3123
rect 13285 3105 13305 3123
rect 13149 3084 13305 3105
rect 13149 3083 13249 3084
rect 8786 3011 8937 3034
rect 8786 2996 8901 3011
rect 4073 2929 4130 2948
rect 4073 2911 4091 2929
rect 4109 2926 4130 2929
rect 4109 2911 4224 2926
rect 37 2828 193 2849
rect 37 2827 137 2828
rect 38 2791 80 2827
rect 38 2768 189 2791
rect 4073 2888 4224 2911
rect 4182 2852 4224 2888
rect 4496 2884 4557 2900
rect 4401 2880 4557 2884
rect 4401 2862 4519 2880
rect 4537 2862 4557 2880
rect 8880 2993 8901 2996
rect 8919 2993 8937 3011
rect 8880 2974 8937 2993
rect 13150 3047 13192 3083
rect 17179 3154 17240 3170
rect 13150 3024 13301 3047
rect 13150 3009 13265 3024
rect 8437 2942 8494 2961
rect 8437 2924 8455 2942
rect 8473 2939 8494 2942
rect 8473 2924 8588 2939
rect 4125 2851 4225 2852
rect 4069 2830 4225 2851
rect 4401 2841 4557 2862
rect 4401 2840 4501 2841
rect 4069 2812 4089 2830
rect 4107 2812 4225 2830
rect 4069 2808 4225 2812
rect 4069 2792 4130 2808
rect 4402 2804 4444 2840
rect 38 2753 153 2768
rect 132 2750 153 2753
rect 171 2750 189 2768
rect 132 2731 189 2750
rect 4402 2781 4553 2804
rect 8437 2901 8588 2924
rect 8546 2865 8588 2901
rect 8873 2896 8934 2912
rect 8778 2892 8934 2896
rect 8778 2874 8896 2892
rect 8914 2874 8934 2892
rect 13244 3006 13265 3009
rect 13283 3006 13301 3024
rect 13244 2987 13301 3006
rect 12814 2954 12871 2973
rect 12814 2936 12832 2954
rect 12850 2951 12871 2954
rect 12850 2936 12965 2951
rect 8489 2864 8589 2865
rect 8433 2843 8589 2864
rect 8778 2853 8934 2874
rect 8778 2852 8878 2853
rect 8433 2825 8453 2843
rect 8471 2825 8589 2843
rect 8433 2821 8589 2825
rect 8433 2805 8494 2821
rect 8779 2816 8821 2852
rect 4402 2766 4517 2781
rect 4496 2763 4517 2766
rect 4535 2763 4553 2781
rect 4496 2744 4553 2763
rect 8779 2793 8930 2816
rect 12814 2913 12965 2936
rect 12923 2877 12965 2913
rect 13237 2909 13298 2925
rect 13142 2905 13298 2909
rect 13142 2887 13260 2905
rect 13278 2887 13298 2905
rect 17178 2967 17235 2986
rect 17178 2949 17196 2967
rect 17214 2964 17235 2967
rect 17214 2949 17329 2964
rect 12866 2876 12966 2877
rect 12810 2855 12966 2876
rect 13142 2866 13298 2887
rect 13142 2865 13242 2866
rect 12810 2837 12830 2855
rect 12848 2837 12966 2855
rect 12810 2833 12966 2837
rect 12810 2817 12871 2833
rect 13143 2829 13185 2865
rect 8779 2778 8894 2793
rect 8873 2775 8894 2778
rect 8912 2775 8930 2793
rect 8873 2756 8930 2775
rect 13143 2806 13294 2829
rect 17178 2926 17329 2949
rect 17287 2890 17329 2926
rect 17230 2889 17330 2890
rect 17174 2868 17330 2889
rect 17174 2850 17194 2868
rect 17212 2850 17330 2868
rect 17174 2846 17330 2850
rect 17174 2830 17235 2846
rect 13143 2791 13258 2806
rect 13237 2788 13258 2791
rect 13276 2788 13294 2806
rect 13237 2769 13294 2788
rect 4071 2636 4128 2655
rect 4071 2618 4089 2636
rect 4107 2633 4128 2636
rect 4107 2618 4222 2633
rect 130 2578 191 2594
rect 35 2574 191 2578
rect 35 2556 153 2574
rect 171 2556 191 2574
rect 35 2535 191 2556
rect 35 2534 135 2535
rect 36 2498 78 2534
rect 36 2475 187 2498
rect 4071 2595 4222 2618
rect 8435 2649 8492 2668
rect 8435 2631 8453 2649
rect 8471 2646 8492 2649
rect 8471 2631 8586 2646
rect 4180 2559 4222 2595
rect 4494 2591 4555 2607
rect 4399 2587 4555 2591
rect 4399 2569 4517 2587
rect 4535 2569 4555 2587
rect 4123 2558 4223 2559
rect 4067 2537 4223 2558
rect 4399 2548 4555 2569
rect 4399 2547 4499 2548
rect 36 2460 151 2475
rect 130 2457 151 2460
rect 169 2457 187 2475
rect 130 2438 187 2457
rect 4067 2519 4087 2537
rect 4105 2519 4223 2537
rect 4067 2515 4223 2519
rect 4067 2499 4128 2515
rect 4400 2511 4442 2547
rect 4400 2488 4551 2511
rect 8435 2608 8586 2631
rect 12812 2661 12869 2680
rect 12812 2643 12830 2661
rect 12848 2658 12869 2661
rect 12848 2643 12963 2658
rect 8544 2572 8586 2608
rect 8871 2603 8932 2619
rect 8776 2599 8932 2603
rect 8776 2581 8894 2599
rect 8912 2581 8932 2599
rect 8487 2571 8587 2572
rect 8431 2550 8587 2571
rect 8776 2560 8932 2581
rect 8776 2559 8876 2560
rect 4400 2473 4515 2488
rect 4494 2470 4515 2473
rect 4533 2470 4551 2488
rect 4494 2451 4551 2470
rect 4064 2418 4121 2437
rect 4064 2400 4082 2418
rect 4100 2415 4121 2418
rect 8431 2532 8451 2550
rect 8469 2532 8587 2550
rect 8431 2528 8587 2532
rect 8431 2512 8492 2528
rect 8777 2523 8819 2559
rect 8777 2500 8928 2523
rect 12812 2620 12963 2643
rect 17176 2674 17233 2693
rect 17176 2656 17194 2674
rect 17212 2671 17233 2674
rect 17212 2656 17327 2671
rect 12921 2584 12963 2620
rect 13235 2616 13296 2632
rect 13140 2612 13296 2616
rect 13140 2594 13258 2612
rect 13276 2594 13296 2612
rect 12864 2583 12964 2584
rect 12808 2562 12964 2583
rect 13140 2573 13296 2594
rect 13140 2572 13240 2573
rect 8777 2485 8892 2500
rect 8871 2482 8892 2485
rect 8910 2482 8928 2500
rect 8871 2463 8928 2482
rect 4100 2400 4215 2415
rect 4064 2377 4215 2400
rect 125 2254 186 2270
rect 4173 2341 4215 2377
rect 8428 2431 8485 2450
rect 8428 2413 8446 2431
rect 8464 2428 8485 2431
rect 12808 2544 12828 2562
rect 12846 2544 12964 2562
rect 12808 2540 12964 2544
rect 12808 2524 12869 2540
rect 13141 2536 13183 2572
rect 13141 2513 13292 2536
rect 17176 2633 17327 2656
rect 17285 2597 17327 2633
rect 17228 2596 17328 2597
rect 17172 2575 17328 2596
rect 13141 2498 13256 2513
rect 13235 2495 13256 2498
rect 13274 2495 13292 2513
rect 13235 2476 13292 2495
rect 8464 2413 8579 2428
rect 8428 2390 8579 2413
rect 4116 2340 4216 2341
rect 4060 2319 4216 2340
rect 4060 2301 4080 2319
rect 4098 2301 4216 2319
rect 4060 2297 4216 2301
rect 30 2250 186 2254
rect 30 2232 148 2250
rect 166 2232 186 2250
rect 30 2211 186 2232
rect 30 2210 130 2211
rect 31 2174 73 2210
rect 4060 2281 4121 2297
rect 4489 2267 4550 2283
rect 8537 2354 8579 2390
rect 12805 2443 12862 2462
rect 12805 2425 12823 2443
rect 12841 2440 12862 2443
rect 17172 2557 17192 2575
rect 17210 2557 17328 2575
rect 17172 2553 17328 2557
rect 17172 2537 17233 2553
rect 12841 2425 12956 2440
rect 12805 2402 12956 2425
rect 8480 2353 8580 2354
rect 8424 2332 8580 2353
rect 8424 2314 8444 2332
rect 8462 2314 8580 2332
rect 8424 2310 8580 2314
rect 4394 2263 4550 2267
rect 4058 2235 4115 2254
rect 31 2151 182 2174
rect 31 2136 146 2151
rect 125 2133 146 2136
rect 164 2133 182 2151
rect 4058 2217 4076 2235
rect 4094 2232 4115 2235
rect 4394 2245 4512 2263
rect 4530 2245 4550 2263
rect 4094 2217 4209 2232
rect 4394 2224 4550 2245
rect 4394 2223 4494 2224
rect 4058 2194 4209 2217
rect 125 2114 182 2133
rect 119 2071 180 2087
rect 4167 2158 4209 2194
rect 4395 2187 4437 2223
rect 8424 2294 8485 2310
rect 8866 2279 8927 2295
rect 12914 2366 12956 2402
rect 17169 2456 17226 2475
rect 17169 2438 17187 2456
rect 17205 2453 17226 2456
rect 17205 2438 17320 2453
rect 17169 2415 17320 2438
rect 12857 2365 12957 2366
rect 12801 2344 12957 2365
rect 12801 2326 12821 2344
rect 12839 2326 12957 2344
rect 12801 2322 12957 2326
rect 8771 2275 8927 2279
rect 8422 2248 8479 2267
rect 4395 2164 4546 2187
rect 4110 2157 4210 2158
rect 4054 2136 4210 2157
rect 4395 2149 4510 2164
rect 4054 2118 4074 2136
rect 4092 2118 4210 2136
rect 4489 2146 4510 2149
rect 4528 2146 4546 2164
rect 8422 2230 8440 2248
rect 8458 2245 8479 2248
rect 8771 2257 8889 2275
rect 8907 2257 8927 2275
rect 8458 2230 8573 2245
rect 8771 2236 8927 2257
rect 8771 2235 8871 2236
rect 8422 2207 8573 2230
rect 4489 2127 4546 2146
rect 4054 2114 4210 2118
rect 24 2067 180 2071
rect 24 2049 142 2067
rect 160 2049 180 2067
rect 24 2028 180 2049
rect 24 2027 124 2028
rect 25 1991 67 2027
rect 4054 2098 4115 2114
rect 4483 2084 4544 2100
rect 8531 2171 8573 2207
rect 8772 2199 8814 2235
rect 12801 2306 12862 2322
rect 13230 2292 13291 2308
rect 17278 2379 17320 2415
rect 17221 2378 17321 2379
rect 17165 2357 17321 2378
rect 17165 2339 17185 2357
rect 17203 2339 17321 2357
rect 17165 2335 17321 2339
rect 13135 2288 13291 2292
rect 12799 2260 12856 2279
rect 8772 2176 8923 2199
rect 8474 2170 8574 2171
rect 8418 2149 8574 2170
rect 8772 2161 8887 2176
rect 8418 2131 8438 2149
rect 8456 2131 8574 2149
rect 8866 2158 8887 2161
rect 8905 2158 8923 2176
rect 12799 2242 12817 2260
rect 12835 2257 12856 2260
rect 13135 2270 13253 2288
rect 13271 2270 13291 2288
rect 12835 2242 12950 2257
rect 13135 2249 13291 2270
rect 13135 2248 13235 2249
rect 12799 2219 12950 2242
rect 8866 2139 8923 2158
rect 8418 2127 8574 2131
rect 4388 2080 4544 2084
rect 4388 2062 4506 2080
rect 4524 2062 4544 2080
rect 4388 2041 4544 2062
rect 4388 2040 4488 2041
rect 25 1968 176 1991
rect 25 1953 140 1968
rect 119 1950 140 1953
rect 158 1950 176 1968
rect 119 1931 176 1950
rect 4389 2004 4431 2040
rect 8418 2111 8479 2127
rect 8860 2096 8921 2112
rect 12908 2183 12950 2219
rect 13136 2212 13178 2248
rect 17165 2319 17226 2335
rect 17163 2273 17220 2292
rect 13136 2189 13287 2212
rect 12851 2182 12951 2183
rect 12795 2161 12951 2182
rect 13136 2174 13251 2189
rect 12795 2143 12815 2161
rect 12833 2143 12951 2161
rect 13230 2171 13251 2174
rect 13269 2171 13287 2189
rect 17163 2255 17181 2273
rect 17199 2270 17220 2273
rect 17199 2255 17314 2270
rect 17163 2232 17314 2255
rect 13230 2152 13287 2171
rect 12795 2139 12951 2143
rect 8765 2092 8921 2096
rect 8765 2074 8883 2092
rect 8901 2074 8921 2092
rect 8765 2053 8921 2074
rect 8765 2052 8865 2053
rect 4389 1981 4540 2004
rect 4389 1966 4504 1981
rect 4483 1963 4504 1966
rect 4522 1963 4540 1981
rect 112 1853 173 1869
rect 17 1849 173 1853
rect 17 1831 135 1849
rect 153 1831 173 1849
rect 4483 1944 4540 1963
rect 8766 2016 8808 2052
rect 12795 2123 12856 2139
rect 13224 2109 13285 2125
rect 17272 2196 17314 2232
rect 17215 2195 17315 2196
rect 17159 2174 17315 2195
rect 17159 2156 17179 2174
rect 17197 2156 17315 2174
rect 17159 2152 17315 2156
rect 13129 2105 13285 2109
rect 13129 2087 13247 2105
rect 13265 2087 13285 2105
rect 13129 2066 13285 2087
rect 13129 2065 13229 2066
rect 8766 1993 8917 2016
rect 8766 1978 8881 1993
rect 4053 1911 4110 1930
rect 4053 1893 4071 1911
rect 4089 1908 4110 1911
rect 4089 1893 4204 1908
rect 17 1810 173 1831
rect 17 1809 117 1810
rect 18 1773 60 1809
rect 18 1750 169 1773
rect 4053 1870 4204 1893
rect 4162 1834 4204 1870
rect 4476 1866 4537 1882
rect 4381 1862 4537 1866
rect 4381 1844 4499 1862
rect 4517 1844 4537 1862
rect 8860 1975 8881 1978
rect 8899 1975 8917 1993
rect 8860 1956 8917 1975
rect 13130 2029 13172 2065
rect 17159 2136 17220 2152
rect 13130 2006 13281 2029
rect 13130 1991 13245 2006
rect 13224 1988 13245 1991
rect 13263 1988 13281 2006
rect 8417 1924 8474 1943
rect 8417 1906 8435 1924
rect 8453 1921 8474 1924
rect 8453 1906 8568 1921
rect 4105 1833 4205 1834
rect 4049 1812 4205 1833
rect 4381 1823 4537 1844
rect 4381 1822 4481 1823
rect 4049 1794 4069 1812
rect 4087 1794 4205 1812
rect 4049 1790 4205 1794
rect 4049 1774 4110 1790
rect 4382 1786 4424 1822
rect 18 1735 133 1750
rect 112 1732 133 1735
rect 151 1732 169 1750
rect 112 1713 169 1732
rect 4382 1763 4533 1786
rect 8417 1883 8568 1906
rect 8526 1847 8568 1883
rect 8853 1878 8914 1894
rect 8758 1874 8914 1878
rect 8758 1856 8876 1874
rect 8894 1856 8914 1874
rect 13224 1969 13281 1988
rect 12794 1936 12851 1955
rect 12794 1918 12812 1936
rect 12830 1933 12851 1936
rect 12830 1918 12945 1933
rect 8469 1846 8569 1847
rect 8413 1825 8569 1846
rect 8758 1835 8914 1856
rect 8758 1834 8858 1835
rect 8413 1807 8433 1825
rect 8451 1807 8569 1825
rect 8413 1803 8569 1807
rect 8413 1787 8474 1803
rect 8759 1798 8801 1834
rect 4382 1748 4497 1763
rect 4476 1745 4497 1748
rect 4515 1745 4533 1763
rect 4476 1726 4533 1745
rect 8759 1775 8910 1798
rect 12794 1895 12945 1918
rect 12903 1859 12945 1895
rect 13217 1891 13278 1907
rect 13122 1887 13278 1891
rect 13122 1869 13240 1887
rect 13258 1869 13278 1887
rect 17158 1949 17215 1968
rect 17158 1931 17176 1949
rect 17194 1946 17215 1949
rect 17194 1931 17309 1946
rect 12846 1858 12946 1859
rect 12790 1837 12946 1858
rect 13122 1848 13278 1869
rect 13122 1847 13222 1848
rect 12790 1819 12810 1837
rect 12828 1819 12946 1837
rect 12790 1815 12946 1819
rect 12790 1799 12851 1815
rect 13123 1811 13165 1847
rect 8759 1760 8874 1775
rect 8853 1757 8874 1760
rect 8892 1757 8910 1775
rect 8853 1738 8910 1757
rect 13123 1788 13274 1811
rect 17158 1908 17309 1931
rect 17267 1872 17309 1908
rect 17210 1871 17310 1872
rect 17154 1850 17310 1871
rect 17154 1832 17174 1850
rect 17192 1832 17310 1850
rect 17154 1828 17310 1832
rect 17154 1812 17215 1828
rect 13123 1773 13238 1788
rect 13217 1770 13238 1773
rect 13256 1770 13274 1788
rect 13217 1751 13274 1770
rect 4054 1618 4111 1637
rect 4054 1600 4072 1618
rect 4090 1615 4111 1618
rect 4090 1600 4205 1615
rect 113 1560 174 1576
rect 18 1556 174 1560
rect 18 1538 136 1556
rect 154 1538 174 1556
rect 18 1517 174 1538
rect 18 1516 118 1517
rect 19 1480 61 1516
rect 19 1457 170 1480
rect 4054 1577 4205 1600
rect 8418 1631 8475 1650
rect 8418 1613 8436 1631
rect 8454 1628 8475 1631
rect 8454 1613 8569 1628
rect 4163 1541 4205 1577
rect 4477 1573 4538 1589
rect 4382 1569 4538 1573
rect 4382 1551 4500 1569
rect 4518 1551 4538 1569
rect 4106 1540 4206 1541
rect 4050 1519 4206 1540
rect 4382 1530 4538 1551
rect 4382 1529 4482 1530
rect 19 1442 134 1457
rect 113 1439 134 1442
rect 152 1439 170 1457
rect 113 1420 170 1439
rect 4050 1501 4070 1519
rect 4088 1501 4206 1519
rect 4050 1497 4206 1501
rect 4050 1481 4111 1497
rect 4383 1493 4425 1529
rect 4383 1470 4534 1493
rect 8418 1590 8569 1613
rect 12795 1643 12852 1662
rect 12795 1625 12813 1643
rect 12831 1640 12852 1643
rect 12831 1625 12946 1640
rect 8527 1554 8569 1590
rect 8854 1585 8915 1601
rect 8759 1581 8915 1585
rect 8759 1563 8877 1581
rect 8895 1563 8915 1581
rect 8470 1553 8570 1554
rect 8414 1532 8570 1553
rect 8759 1542 8915 1563
rect 8759 1541 8859 1542
rect 4383 1455 4498 1470
rect 4477 1452 4498 1455
rect 4516 1452 4534 1470
rect 4477 1433 4534 1452
rect 4047 1400 4104 1419
rect 8414 1514 8434 1532
rect 8452 1514 8570 1532
rect 8414 1510 8570 1514
rect 8414 1494 8475 1510
rect 8760 1505 8802 1541
rect 8760 1482 8911 1505
rect 12795 1602 12946 1625
rect 17159 1656 17216 1675
rect 17159 1638 17177 1656
rect 17195 1653 17216 1656
rect 17195 1638 17310 1653
rect 12904 1566 12946 1602
rect 13218 1598 13279 1614
rect 13123 1594 13279 1598
rect 13123 1576 13241 1594
rect 13259 1576 13279 1594
rect 12847 1565 12947 1566
rect 12791 1544 12947 1565
rect 13123 1555 13279 1576
rect 13123 1554 13223 1555
rect 8760 1467 8875 1482
rect 8854 1464 8875 1467
rect 8893 1464 8911 1482
rect 8854 1445 8911 1464
rect 4047 1382 4065 1400
rect 4083 1397 4104 1400
rect 4083 1382 4198 1397
rect 4047 1359 4198 1382
rect 108 1236 169 1252
rect 4156 1323 4198 1359
rect 8411 1413 8468 1432
rect 8411 1395 8429 1413
rect 8447 1410 8468 1413
rect 12791 1526 12811 1544
rect 12829 1526 12947 1544
rect 12791 1522 12947 1526
rect 12791 1506 12852 1522
rect 13124 1518 13166 1554
rect 13124 1495 13275 1518
rect 17159 1615 17310 1638
rect 17268 1579 17310 1615
rect 17211 1578 17311 1579
rect 17155 1557 17311 1578
rect 13124 1480 13239 1495
rect 13218 1477 13239 1480
rect 13257 1477 13275 1495
rect 13218 1458 13275 1477
rect 8447 1395 8562 1410
rect 8411 1372 8562 1395
rect 4099 1322 4199 1323
rect 4043 1301 4199 1322
rect 4043 1283 4063 1301
rect 4081 1283 4199 1301
rect 4043 1279 4199 1283
rect 13 1232 169 1236
rect 13 1214 131 1232
rect 149 1214 169 1232
rect 13 1193 169 1214
rect 13 1192 113 1193
rect 14 1156 56 1192
rect 4043 1263 4104 1279
rect 4472 1249 4533 1265
rect 8520 1336 8562 1372
rect 12788 1425 12845 1444
rect 17155 1539 17175 1557
rect 17193 1539 17311 1557
rect 17155 1535 17311 1539
rect 17155 1519 17216 1535
rect 12788 1407 12806 1425
rect 12824 1422 12845 1425
rect 12824 1407 12939 1422
rect 12788 1384 12939 1407
rect 8463 1335 8563 1336
rect 8407 1314 8563 1335
rect 8407 1296 8427 1314
rect 8445 1296 8563 1314
rect 8407 1292 8563 1296
rect 4377 1245 4533 1249
rect 4041 1217 4098 1236
rect 14 1133 165 1156
rect 14 1118 129 1133
rect 108 1115 129 1118
rect 147 1115 165 1133
rect 4041 1199 4059 1217
rect 4077 1214 4098 1217
rect 4377 1227 4495 1245
rect 4513 1227 4533 1245
rect 4077 1199 4192 1214
rect 4377 1206 4533 1227
rect 4377 1205 4477 1206
rect 4041 1176 4192 1199
rect 108 1096 165 1115
rect 102 1053 163 1069
rect 4150 1140 4192 1176
rect 4378 1169 4420 1205
rect 8407 1276 8468 1292
rect 8849 1261 8910 1277
rect 12897 1348 12939 1384
rect 17152 1438 17209 1457
rect 17152 1420 17170 1438
rect 17188 1435 17209 1438
rect 17188 1420 17303 1435
rect 17152 1397 17303 1420
rect 12840 1347 12940 1348
rect 12784 1326 12940 1347
rect 12784 1308 12804 1326
rect 12822 1308 12940 1326
rect 12784 1304 12940 1308
rect 8754 1257 8910 1261
rect 8405 1230 8462 1249
rect 4378 1146 4529 1169
rect 4093 1139 4193 1140
rect 4037 1118 4193 1139
rect 4378 1131 4493 1146
rect 4037 1100 4057 1118
rect 4075 1100 4193 1118
rect 4472 1128 4493 1131
rect 4511 1128 4529 1146
rect 8405 1212 8423 1230
rect 8441 1227 8462 1230
rect 8754 1239 8872 1257
rect 8890 1239 8910 1257
rect 8441 1212 8556 1227
rect 8754 1218 8910 1239
rect 8754 1217 8854 1218
rect 8405 1189 8556 1212
rect 4472 1109 4529 1128
rect 4037 1096 4193 1100
rect 7 1049 163 1053
rect 7 1031 125 1049
rect 143 1031 163 1049
rect 7 1010 163 1031
rect 7 1009 107 1010
rect 8 973 50 1009
rect 4037 1080 4098 1096
rect 4466 1066 4527 1082
rect 8514 1153 8556 1189
rect 8755 1181 8797 1217
rect 12784 1288 12845 1304
rect 13213 1274 13274 1290
rect 17261 1361 17303 1397
rect 17204 1360 17304 1361
rect 17148 1339 17304 1360
rect 17148 1321 17168 1339
rect 17186 1321 17304 1339
rect 17148 1317 17304 1321
rect 13118 1270 13274 1274
rect 12782 1242 12839 1261
rect 8755 1158 8906 1181
rect 8457 1152 8557 1153
rect 8401 1131 8557 1152
rect 8755 1143 8870 1158
rect 8401 1113 8421 1131
rect 8439 1113 8557 1131
rect 8849 1140 8870 1143
rect 8888 1140 8906 1158
rect 12782 1224 12800 1242
rect 12818 1239 12839 1242
rect 13118 1252 13236 1270
rect 13254 1252 13274 1270
rect 12818 1224 12933 1239
rect 13118 1231 13274 1252
rect 13118 1230 13218 1231
rect 12782 1201 12933 1224
rect 8849 1121 8906 1140
rect 8401 1109 8557 1113
rect 4371 1062 4527 1066
rect 4371 1044 4489 1062
rect 4507 1044 4527 1062
rect 4371 1023 4527 1044
rect 4371 1022 4471 1023
rect 4372 986 4414 1022
rect 8401 1093 8462 1109
rect 8843 1078 8904 1094
rect 12891 1165 12933 1201
rect 13119 1194 13161 1230
rect 17148 1301 17209 1317
rect 17146 1255 17203 1274
rect 13119 1171 13270 1194
rect 12834 1164 12934 1165
rect 12778 1143 12934 1164
rect 13119 1156 13234 1171
rect 12778 1125 12798 1143
rect 12816 1125 12934 1143
rect 13213 1153 13234 1156
rect 13252 1153 13270 1171
rect 17146 1237 17164 1255
rect 17182 1252 17203 1255
rect 17182 1237 17297 1252
rect 17146 1214 17297 1237
rect 13213 1134 13270 1153
rect 12778 1121 12934 1125
rect 8748 1074 8904 1078
rect 8748 1056 8866 1074
rect 8884 1056 8904 1074
rect 8748 1035 8904 1056
rect 8748 1034 8848 1035
rect 8749 998 8791 1034
rect 12778 1105 12839 1121
rect 13207 1091 13268 1107
rect 17255 1178 17297 1214
rect 17198 1177 17298 1178
rect 17142 1156 17298 1177
rect 17142 1138 17162 1156
rect 17180 1138 17298 1156
rect 17142 1134 17298 1138
rect 13112 1087 13268 1091
rect 13112 1069 13230 1087
rect 13248 1069 13268 1087
rect 13112 1048 13268 1069
rect 13112 1047 13212 1048
rect 13113 1011 13155 1047
rect 17142 1118 17203 1134
rect 8 950 159 973
rect 8 935 123 950
rect 102 932 123 935
rect 141 932 159 950
rect 102 913 159 932
rect 4372 963 4523 986
rect 4372 948 4487 963
rect 4466 945 4487 948
rect 4505 945 4523 963
rect 95 835 156 851
rect 0 831 156 835
rect 0 813 118 831
rect 136 813 156 831
rect 4466 926 4523 945
rect 8749 975 8900 998
rect 8749 960 8864 975
rect 8843 957 8864 960
rect 8882 957 8900 975
rect 4036 893 4093 912
rect 4036 875 4054 893
rect 4072 890 4093 893
rect 4072 875 4187 890
rect 4036 852 4187 875
rect 0 792 156 813
rect 0 791 100 792
rect 1 755 43 791
rect 1 732 152 755
rect 4145 816 4187 852
rect 4459 848 4520 864
rect 4364 844 4520 848
rect 4364 826 4482 844
rect 4500 826 4520 844
rect 8843 938 8900 957
rect 13113 988 13264 1011
rect 13113 973 13228 988
rect 13207 970 13228 973
rect 13246 970 13264 988
rect 8400 906 8457 925
rect 8400 888 8418 906
rect 8436 903 8457 906
rect 8436 888 8551 903
rect 8400 865 8551 888
rect 4088 815 4188 816
rect 4032 794 4188 815
rect 4364 805 4520 826
rect 4364 804 4464 805
rect 4032 776 4052 794
rect 4070 776 4188 794
rect 4032 772 4188 776
rect 4032 756 4093 772
rect 4365 768 4407 804
rect 1 717 116 732
rect 95 714 116 717
rect 134 714 152 732
rect 95 695 152 714
rect 4365 745 4516 768
rect 8509 829 8551 865
rect 8836 860 8897 876
rect 8741 856 8897 860
rect 8741 838 8859 856
rect 8877 838 8897 856
rect 13207 951 13264 970
rect 12777 918 12834 937
rect 12777 900 12795 918
rect 12813 915 12834 918
rect 12813 900 12928 915
rect 12777 877 12928 900
rect 8452 828 8552 829
rect 8396 807 8552 828
rect 8741 817 8897 838
rect 8741 816 8841 817
rect 8396 789 8416 807
rect 8434 789 8552 807
rect 8396 785 8552 789
rect 8396 769 8457 785
rect 8742 780 8784 816
rect 4365 730 4480 745
rect 4459 727 4480 730
rect 4498 727 4516 745
rect 4459 708 4516 727
rect 8742 757 8893 780
rect 12886 841 12928 877
rect 13200 873 13261 889
rect 13105 869 13261 873
rect 13105 851 13223 869
rect 13241 851 13261 869
rect 17141 931 17198 950
rect 17141 913 17159 931
rect 17177 928 17198 931
rect 17177 913 17292 928
rect 17141 890 17292 913
rect 12829 840 12929 841
rect 12773 819 12929 840
rect 13105 830 13261 851
rect 13105 829 13205 830
rect 12773 801 12793 819
rect 12811 801 12929 819
rect 12773 797 12929 801
rect 12773 781 12834 797
rect 13106 793 13148 829
rect 8742 742 8857 757
rect 8836 739 8857 742
rect 8875 739 8893 757
rect 8836 720 8893 739
rect 13106 770 13257 793
rect 17250 854 17292 890
rect 17193 853 17293 854
rect 17137 832 17293 853
rect 17137 814 17157 832
rect 17175 814 17293 832
rect 17137 810 17293 814
rect 17137 794 17198 810
rect 13106 755 13221 770
rect 13200 752 13221 755
rect 13239 752 13257 770
rect 13200 733 13257 752
<< locali >>
rect 8546 8914 8587 8917
rect 2875 8823 2915 8831
rect 2875 8801 2883 8823
rect 2907 8801 2915 8823
rect 3779 8826 4235 8861
rect 8146 8854 9041 8914
rect 8146 8853 8593 8854
rect 7239 8836 7279 8844
rect 253 8682 300 8798
rect 253 8664 263 8682
rect 281 8664 300 8682
rect 253 8660 300 8664
rect 254 8655 291 8660
rect 242 8593 294 8595
rect 240 8589 673 8593
rect 240 8583 679 8589
rect 240 8565 261 8583
rect 279 8565 679 8583
rect 240 8547 679 8565
rect 242 8358 294 8547
rect 640 8522 679 8547
rect 2480 8572 2517 8578
rect 2480 8553 2488 8572
rect 2509 8553 2517 8572
rect 2480 8545 2517 8553
rect 424 8497 611 8521
rect 640 8502 1035 8522
rect 1055 8502 1058 8522
rect 640 8497 1058 8502
rect 424 8426 461 8497
rect 640 8496 983 8497
rect 640 8493 679 8496
rect 945 8495 982 8496
rect 576 8436 607 8437
rect 424 8406 433 8426
rect 453 8406 461 8426
rect 424 8396 461 8406
rect 520 8426 607 8436
rect 520 8406 529 8426
rect 549 8406 607 8426
rect 520 8397 607 8406
rect 520 8396 557 8397
rect 242 8340 258 8358
rect 276 8340 294 8358
rect 576 8346 607 8397
rect 642 8426 679 8493
rect 794 8436 830 8437
rect 642 8406 651 8426
rect 671 8406 679 8426
rect 642 8396 679 8406
rect 738 8426 886 8436
rect 986 8433 1082 8435
rect 738 8406 747 8426
rect 767 8406 857 8426
rect 877 8406 886 8426
rect 738 8397 886 8406
rect 944 8426 1082 8433
rect 944 8406 953 8426
rect 973 8406 1082 8426
rect 944 8397 1082 8406
rect 738 8396 775 8397
rect 468 8343 509 8344
rect 242 8322 294 8340
rect 360 8336 509 8343
rect 360 8316 419 8336
rect 439 8316 478 8336
rect 498 8316 509 8336
rect 360 8308 509 8316
rect 576 8339 733 8346
rect 576 8319 696 8339
rect 716 8319 733 8339
rect 576 8309 733 8319
rect 576 8308 611 8309
rect 576 8287 607 8308
rect 794 8287 830 8397
rect 849 8396 886 8397
rect 945 8396 982 8397
rect 905 8337 995 8343
rect 905 8317 914 8337
rect 934 8335 995 8337
rect 934 8317 959 8335
rect 905 8315 959 8317
rect 979 8315 995 8335
rect 905 8309 995 8315
rect 419 8286 456 8287
rect 418 8277 456 8286
rect 246 8259 286 8269
rect 246 8241 256 8259
rect 274 8241 286 8259
rect 418 8257 427 8277
rect 447 8257 456 8277
rect 418 8249 456 8257
rect 522 8281 607 8287
rect 637 8286 674 8287
rect 522 8261 530 8281
rect 550 8261 607 8281
rect 522 8253 607 8261
rect 636 8277 674 8286
rect 636 8257 645 8277
rect 665 8257 674 8277
rect 522 8252 558 8253
rect 636 8249 674 8257
rect 740 8281 884 8287
rect 740 8261 748 8281
rect 768 8261 801 8281
rect 821 8261 856 8281
rect 876 8261 884 8281
rect 740 8253 884 8261
rect 740 8252 776 8253
rect 848 8252 884 8253
rect 950 8286 987 8287
rect 950 8285 988 8286
rect 950 8277 1014 8285
rect 950 8257 959 8277
rect 979 8263 1014 8277
rect 1034 8263 1037 8283
rect 979 8258 1037 8263
rect 979 8257 1014 8258
rect 246 8185 286 8241
rect 419 8220 456 8249
rect 420 8218 456 8220
rect 420 8196 611 8218
rect 637 8217 674 8249
rect 950 8245 1014 8257
rect 1054 8219 1081 8397
rect 913 8217 1081 8219
rect 637 8207 1081 8217
rect 1222 8313 1409 8337
rect 1440 8318 1833 8338
rect 1853 8318 1856 8338
rect 1440 8313 1856 8318
rect 1222 8242 1259 8313
rect 1440 8312 1781 8313
rect 1374 8252 1405 8253
rect 1222 8222 1231 8242
rect 1251 8222 1259 8242
rect 1222 8212 1259 8222
rect 1318 8242 1405 8252
rect 1318 8222 1327 8242
rect 1347 8222 1405 8242
rect 1318 8213 1405 8222
rect 1318 8212 1355 8213
rect 243 8180 286 8185
rect 634 8191 1081 8207
rect 634 8185 662 8191
rect 913 8190 1081 8191
rect 243 8177 393 8180
rect 634 8177 661 8185
rect 243 8175 661 8177
rect 243 8157 252 8175
rect 270 8157 661 8175
rect 1374 8162 1405 8213
rect 1440 8242 1477 8312
rect 1743 8311 1780 8312
rect 1592 8252 1628 8253
rect 1440 8222 1449 8242
rect 1469 8222 1477 8242
rect 1440 8212 1477 8222
rect 1536 8242 1684 8252
rect 1784 8249 1880 8251
rect 1536 8222 1545 8242
rect 1565 8222 1655 8242
rect 1675 8222 1684 8242
rect 1536 8213 1684 8222
rect 1742 8242 1880 8249
rect 1742 8222 1751 8242
rect 1771 8222 1880 8242
rect 1742 8213 1880 8222
rect 1536 8212 1573 8213
rect 1266 8159 1307 8160
rect 243 8154 661 8157
rect 243 8148 286 8154
rect 246 8145 286 8148
rect 1158 8152 1307 8159
rect 643 8136 683 8137
rect 354 8119 683 8136
rect 1158 8132 1217 8152
rect 1237 8132 1276 8152
rect 1296 8132 1307 8152
rect 1158 8124 1307 8132
rect 1374 8155 1531 8162
rect 1374 8135 1494 8155
rect 1514 8135 1531 8155
rect 1374 8125 1531 8135
rect 1374 8124 1409 8125
rect 238 8076 281 8087
rect 238 8058 250 8076
rect 268 8058 281 8076
rect 238 8032 281 8058
rect 354 8032 381 8119
rect 643 8110 683 8119
rect 238 8011 381 8032
rect 425 8084 459 8100
rect 643 8090 1036 8110
rect 1056 8090 1059 8110
rect 1374 8103 1405 8124
rect 1592 8103 1628 8213
rect 1647 8212 1684 8213
rect 1743 8212 1780 8213
rect 1703 8153 1793 8159
rect 1703 8133 1712 8153
rect 1732 8151 1793 8153
rect 1732 8133 1757 8151
rect 1703 8131 1757 8133
rect 1777 8131 1793 8151
rect 1703 8125 1793 8131
rect 1217 8102 1254 8103
rect 643 8085 1059 8090
rect 1216 8093 1254 8102
rect 643 8084 984 8085
rect 425 8014 462 8084
rect 577 8024 608 8025
rect 238 8009 375 8011
rect 238 7967 281 8009
rect 425 7994 434 8014
rect 454 7994 462 8014
rect 425 7984 462 7994
rect 521 8014 608 8024
rect 521 7994 530 8014
rect 550 7994 608 8014
rect 521 7985 608 7994
rect 521 7984 558 7985
rect 236 7957 281 7967
rect 236 7939 245 7957
rect 263 7939 281 7957
rect 236 7933 281 7939
rect 577 7934 608 7985
rect 643 8014 680 8084
rect 946 8083 983 8084
rect 1216 8073 1225 8093
rect 1245 8073 1254 8093
rect 1216 8065 1254 8073
rect 1320 8097 1405 8103
rect 1435 8102 1472 8103
rect 1320 8077 1328 8097
rect 1348 8077 1405 8097
rect 1320 8069 1405 8077
rect 1434 8093 1472 8102
rect 1434 8073 1443 8093
rect 1463 8073 1472 8093
rect 1320 8068 1356 8069
rect 1434 8065 1472 8073
rect 1538 8097 1682 8103
rect 1538 8077 1546 8097
rect 1566 8078 1598 8097
rect 1619 8078 1654 8097
rect 1566 8077 1654 8078
rect 1674 8077 1682 8097
rect 1538 8069 1682 8077
rect 1538 8068 1574 8069
rect 1646 8068 1682 8069
rect 1748 8102 1785 8103
rect 1748 8101 1786 8102
rect 1748 8093 1812 8101
rect 1748 8073 1757 8093
rect 1777 8079 1812 8093
rect 1832 8079 1835 8099
rect 1777 8074 1835 8079
rect 1777 8073 1812 8074
rect 1217 8036 1254 8065
rect 1218 8034 1254 8036
rect 795 8024 831 8025
rect 643 7994 652 8014
rect 672 7994 680 8014
rect 643 7984 680 7994
rect 739 8014 887 8024
rect 987 8021 1083 8023
rect 739 7994 748 8014
rect 768 7994 858 8014
rect 878 7994 887 8014
rect 739 7985 887 7994
rect 945 8014 1083 8021
rect 945 7994 954 8014
rect 974 7994 1083 8014
rect 1218 8012 1409 8034
rect 1435 8033 1472 8065
rect 1748 8061 1812 8073
rect 1852 8035 1879 8213
rect 2484 8212 2517 8545
rect 2581 8577 2749 8578
rect 2875 8577 2915 8801
rect 3378 8805 3546 8806
rect 3779 8805 3824 8826
rect 3378 8779 3824 8805
rect 3378 8777 3546 8779
rect 3742 8778 3824 8779
rect 3959 8778 4040 8804
rect 4184 8791 4665 8826
rect 7239 8814 7247 8836
rect 7271 8814 7279 8836
rect 3378 8599 3405 8777
rect 3445 8739 3509 8751
rect 3785 8747 3822 8778
rect 4003 8747 4040 8778
rect 4187 8772 4226 8791
rect 4185 8753 4226 8772
rect 3445 8738 3480 8739
rect 3422 8733 3480 8738
rect 3422 8713 3425 8733
rect 3445 8719 3480 8733
rect 3500 8719 3509 8739
rect 3445 8711 3509 8719
rect 3471 8710 3509 8711
rect 3472 8709 3509 8710
rect 3575 8743 3611 8744
rect 3683 8743 3719 8744
rect 3575 8735 3719 8743
rect 3575 8715 3583 8735
rect 3603 8731 3691 8735
rect 3603 8715 3647 8731
rect 3575 8711 3647 8715
rect 3667 8715 3691 8731
rect 3711 8715 3719 8735
rect 3667 8711 3719 8715
rect 3575 8709 3719 8711
rect 3785 8739 3823 8747
rect 3901 8743 3937 8744
rect 3785 8719 3794 8739
rect 3814 8719 3823 8739
rect 3785 8710 3823 8719
rect 3852 8735 3937 8743
rect 3852 8715 3909 8735
rect 3929 8715 3937 8735
rect 3785 8709 3822 8710
rect 3852 8709 3937 8715
rect 4003 8739 4041 8747
rect 4003 8719 4012 8739
rect 4032 8719 4041 8739
rect 4003 8710 4041 8719
rect 4185 8744 4227 8753
rect 4185 8726 4199 8744
rect 4217 8726 4227 8744
rect 4185 8718 4227 8726
rect 4190 8716 4227 8718
rect 4003 8709 4040 8710
rect 3464 8681 3554 8687
rect 3464 8661 3480 8681
rect 3500 8679 3554 8681
rect 3500 8661 3525 8679
rect 3464 8659 3525 8661
rect 3545 8659 3554 8679
rect 3464 8653 3554 8659
rect 3477 8599 3514 8600
rect 3573 8599 3610 8600
rect 3629 8599 3665 8709
rect 3852 8688 3883 8709
rect 4617 8695 4664 8791
rect 3848 8687 3883 8688
rect 3726 8677 3883 8687
rect 3726 8657 3743 8677
rect 3763 8657 3883 8677
rect 3726 8650 3883 8657
rect 3950 8680 4099 8688
rect 3950 8660 3961 8680
rect 3981 8660 4020 8680
rect 4040 8660 4099 8680
rect 4617 8677 4627 8695
rect 4645 8677 4664 8695
rect 4617 8673 4664 8677
rect 4618 8668 4655 8673
rect 3950 8653 4099 8660
rect 3950 8652 3991 8653
rect 4187 8651 4224 8654
rect 3684 8599 3721 8600
rect 3377 8590 3515 8599
rect 2581 8551 3025 8577
rect 2581 8549 2749 8551
rect 2581 8371 2608 8549
rect 2648 8511 2712 8523
rect 2988 8519 3025 8551
rect 3051 8550 3242 8572
rect 3377 8570 3486 8590
rect 3506 8570 3515 8590
rect 3377 8563 3515 8570
rect 3573 8590 3721 8599
rect 3573 8570 3582 8590
rect 3602 8570 3692 8590
rect 3712 8570 3721 8590
rect 3377 8561 3473 8563
rect 3573 8560 3721 8570
rect 3780 8590 3817 8600
rect 3780 8570 3788 8590
rect 3808 8570 3817 8590
rect 3629 8559 3665 8560
rect 3206 8548 3242 8550
rect 3206 8519 3243 8548
rect 2648 8510 2683 8511
rect 2625 8505 2683 8510
rect 2625 8485 2628 8505
rect 2648 8491 2683 8505
rect 2703 8491 2712 8511
rect 2648 8485 2712 8491
rect 2625 8483 2712 8485
rect 2625 8479 2652 8483
rect 2674 8482 2712 8483
rect 2675 8481 2712 8482
rect 2778 8515 2814 8516
rect 2886 8515 2922 8516
rect 2778 8508 2922 8515
rect 2778 8507 2840 8508
rect 2778 8487 2786 8507
rect 2806 8490 2840 8507
rect 2859 8507 2922 8508
rect 2859 8490 2894 8507
rect 2806 8487 2894 8490
rect 2914 8487 2922 8507
rect 2778 8481 2922 8487
rect 2988 8511 3026 8519
rect 3104 8515 3140 8516
rect 2988 8491 2997 8511
rect 3017 8491 3026 8511
rect 2988 8482 3026 8491
rect 3055 8507 3140 8515
rect 3055 8487 3112 8507
rect 3132 8487 3140 8507
rect 2988 8481 3025 8482
rect 3055 8481 3140 8487
rect 3206 8511 3244 8519
rect 3206 8491 3215 8511
rect 3235 8491 3244 8511
rect 3477 8500 3514 8501
rect 3780 8500 3817 8570
rect 3852 8599 3883 8650
rect 4179 8645 4224 8651
rect 4179 8627 4197 8645
rect 4215 8627 4224 8645
rect 4179 8617 4224 8627
rect 3902 8599 3939 8600
rect 3852 8590 3939 8599
rect 3852 8570 3910 8590
rect 3930 8570 3939 8590
rect 3852 8560 3939 8570
rect 3998 8590 4035 8600
rect 3998 8570 4006 8590
rect 4026 8570 4035 8590
rect 4179 8575 4222 8617
rect 4606 8606 4658 8608
rect 4085 8573 4222 8575
rect 3852 8559 3883 8560
rect 3998 8500 4035 8570
rect 3476 8499 3817 8500
rect 3206 8482 3244 8491
rect 3401 8494 3817 8499
rect 3206 8481 3243 8482
rect 2667 8453 2757 8459
rect 2667 8433 2683 8453
rect 2703 8451 2757 8453
rect 2703 8433 2728 8451
rect 2667 8431 2728 8433
rect 2748 8431 2757 8451
rect 2667 8425 2757 8431
rect 2680 8371 2717 8372
rect 2776 8371 2813 8372
rect 2832 8371 2868 8481
rect 3055 8460 3086 8481
rect 3401 8474 3404 8494
rect 3424 8474 3817 8494
rect 4001 8484 4035 8500
rect 4079 8552 4222 8573
rect 4604 8602 5037 8606
rect 4604 8596 5043 8602
rect 4604 8578 4625 8596
rect 4643 8578 5043 8596
rect 4604 8560 5043 8578
rect 3777 8465 3817 8474
rect 4079 8465 4106 8552
rect 4179 8526 4222 8552
rect 4179 8508 4192 8526
rect 4210 8508 4222 8526
rect 4179 8497 4222 8508
rect 3051 8459 3086 8460
rect 2929 8449 3086 8459
rect 2929 8429 2946 8449
rect 2966 8429 3086 8449
rect 2929 8422 3086 8429
rect 3153 8452 3299 8460
rect 3153 8432 3164 8452
rect 3184 8432 3223 8452
rect 3243 8432 3299 8452
rect 3777 8448 4106 8465
rect 3777 8447 3817 8448
rect 3153 8425 3299 8432
rect 4174 8436 4214 8439
rect 4174 8430 4217 8436
rect 3799 8427 4217 8430
rect 3153 8424 3194 8425
rect 2887 8371 2924 8372
rect 2580 8362 2718 8371
rect 2580 8342 2689 8362
rect 2709 8342 2718 8362
rect 2580 8335 2718 8342
rect 2776 8362 2924 8371
rect 2776 8342 2785 8362
rect 2805 8342 2895 8362
rect 2915 8342 2924 8362
rect 2580 8333 2676 8335
rect 2776 8332 2924 8342
rect 2983 8362 3020 8372
rect 2983 8342 2991 8362
rect 3011 8342 3020 8362
rect 2832 8331 2868 8332
rect 2680 8272 2717 8273
rect 2983 8272 3020 8342
rect 3055 8371 3086 8422
rect 3799 8409 4190 8427
rect 4208 8409 4217 8427
rect 3799 8407 4217 8409
rect 3799 8399 3826 8407
rect 4067 8404 4217 8407
rect 3379 8393 3547 8394
rect 3798 8393 3826 8399
rect 3379 8377 3826 8393
rect 4174 8399 4217 8404
rect 3105 8371 3142 8372
rect 3055 8362 3142 8371
rect 3055 8342 3113 8362
rect 3133 8342 3142 8362
rect 3055 8332 3142 8342
rect 3201 8362 3238 8372
rect 3201 8342 3209 8362
rect 3229 8342 3238 8362
rect 3055 8331 3086 8332
rect 2679 8271 3020 8272
rect 3201 8271 3238 8342
rect 2604 8266 3020 8271
rect 2604 8246 2607 8266
rect 2627 8246 3020 8266
rect 3051 8247 3238 8271
rect 3379 8367 3823 8377
rect 3379 8365 3547 8367
rect 2479 8167 2521 8212
rect 3379 8187 3406 8365
rect 3446 8327 3510 8339
rect 3786 8335 3823 8367
rect 3849 8366 4040 8388
rect 4004 8364 4040 8366
rect 4004 8335 4041 8364
rect 4174 8343 4214 8399
rect 3446 8326 3481 8327
rect 3423 8321 3481 8326
rect 3423 8301 3426 8321
rect 3446 8307 3481 8321
rect 3501 8307 3510 8327
rect 3446 8299 3510 8307
rect 3472 8298 3510 8299
rect 3473 8297 3510 8298
rect 3576 8331 3612 8332
rect 3684 8331 3720 8332
rect 3576 8323 3720 8331
rect 3576 8303 3584 8323
rect 3604 8303 3639 8323
rect 3659 8303 3692 8323
rect 3712 8303 3720 8323
rect 3576 8297 3720 8303
rect 3786 8327 3824 8335
rect 3902 8331 3938 8332
rect 3786 8307 3795 8327
rect 3815 8307 3824 8327
rect 3786 8298 3824 8307
rect 3853 8323 3938 8331
rect 3853 8303 3910 8323
rect 3930 8303 3938 8323
rect 3786 8297 3823 8298
rect 3853 8297 3938 8303
rect 4004 8327 4042 8335
rect 4004 8307 4013 8327
rect 4033 8307 4042 8327
rect 4174 8325 4186 8343
rect 4204 8325 4214 8343
rect 4606 8371 4658 8560
rect 5004 8535 5043 8560
rect 6844 8585 6881 8591
rect 6844 8566 6852 8585
rect 6873 8566 6881 8585
rect 6844 8558 6881 8566
rect 4788 8510 4975 8534
rect 5004 8515 5399 8535
rect 5419 8515 5422 8535
rect 5004 8510 5422 8515
rect 4788 8439 4825 8510
rect 5004 8509 5347 8510
rect 5004 8506 5043 8509
rect 5309 8508 5346 8509
rect 4940 8449 4971 8450
rect 4788 8419 4797 8439
rect 4817 8419 4825 8439
rect 4788 8409 4825 8419
rect 4884 8439 4971 8449
rect 4884 8419 4893 8439
rect 4913 8419 4971 8439
rect 4884 8410 4971 8419
rect 4884 8409 4921 8410
rect 4606 8353 4622 8371
rect 4640 8353 4658 8371
rect 4940 8359 4971 8410
rect 5006 8439 5043 8506
rect 5158 8449 5194 8450
rect 5006 8419 5015 8439
rect 5035 8419 5043 8439
rect 5006 8409 5043 8419
rect 5102 8439 5250 8449
rect 5350 8446 5446 8448
rect 5102 8419 5111 8439
rect 5131 8419 5221 8439
rect 5241 8419 5250 8439
rect 5102 8410 5250 8419
rect 5308 8439 5446 8446
rect 5308 8419 5317 8439
rect 5337 8419 5446 8439
rect 5308 8410 5446 8419
rect 5102 8409 5139 8410
rect 4832 8356 4873 8357
rect 4606 8335 4658 8353
rect 4724 8349 4873 8356
rect 4174 8315 4214 8325
rect 4724 8329 4783 8349
rect 4803 8329 4842 8349
rect 4862 8329 4873 8349
rect 4724 8321 4873 8329
rect 4940 8352 5097 8359
rect 4940 8332 5060 8352
rect 5080 8332 5097 8352
rect 4940 8322 5097 8332
rect 4940 8321 4975 8322
rect 4004 8298 4042 8307
rect 4940 8300 4971 8321
rect 5158 8300 5194 8410
rect 5213 8409 5250 8410
rect 5309 8409 5346 8410
rect 5269 8350 5359 8356
rect 5269 8330 5278 8350
rect 5298 8348 5359 8350
rect 5298 8330 5323 8348
rect 5269 8328 5323 8330
rect 5343 8328 5359 8348
rect 5269 8322 5359 8328
rect 4783 8299 4820 8300
rect 4004 8297 4041 8298
rect 3465 8269 3555 8275
rect 3465 8249 3481 8269
rect 3501 8267 3555 8269
rect 3501 8249 3526 8267
rect 3465 8247 3526 8249
rect 3546 8247 3555 8267
rect 3465 8241 3555 8247
rect 3478 8187 3515 8188
rect 3574 8187 3611 8188
rect 3630 8187 3666 8297
rect 3853 8276 3884 8297
rect 4782 8290 4820 8299
rect 3849 8275 3884 8276
rect 3727 8265 3884 8275
rect 3727 8245 3744 8265
rect 3764 8245 3884 8265
rect 3727 8238 3884 8245
rect 3951 8268 4100 8276
rect 3951 8248 3962 8268
rect 3982 8248 4021 8268
rect 4041 8248 4100 8268
rect 4610 8272 4650 8282
rect 3951 8241 4100 8248
rect 4166 8244 4218 8262
rect 3951 8240 3992 8241
rect 3685 8187 3722 8188
rect 3378 8178 3516 8187
rect 2850 8167 2883 8169
rect 2479 8155 2926 8167
rect 1711 8033 1879 8035
rect 1435 8007 1879 8033
rect 945 7985 1083 7994
rect 739 7984 776 7985
rect 236 7930 273 7933
rect 469 7931 510 7932
rect 361 7924 510 7931
rect 361 7904 420 7924
rect 440 7904 479 7924
rect 499 7904 510 7924
rect 361 7896 510 7904
rect 577 7927 734 7934
rect 577 7907 697 7927
rect 717 7907 734 7927
rect 577 7897 734 7907
rect 577 7896 612 7897
rect 577 7875 608 7896
rect 795 7875 831 7985
rect 850 7984 887 7985
rect 946 7984 983 7985
rect 906 7925 996 7931
rect 906 7905 915 7925
rect 935 7923 996 7925
rect 935 7905 960 7923
rect 906 7903 960 7905
rect 980 7903 996 7923
rect 906 7897 996 7903
rect 420 7874 457 7875
rect 233 7866 270 7868
rect 233 7858 275 7866
rect 233 7840 243 7858
rect 261 7840 275 7858
rect 233 7831 275 7840
rect 419 7865 457 7874
rect 419 7845 428 7865
rect 448 7845 457 7865
rect 419 7837 457 7845
rect 523 7869 608 7875
rect 638 7874 675 7875
rect 523 7849 531 7869
rect 551 7849 608 7869
rect 523 7841 608 7849
rect 637 7865 675 7874
rect 637 7845 646 7865
rect 666 7845 675 7865
rect 523 7840 559 7841
rect 637 7837 675 7845
rect 741 7873 885 7875
rect 741 7869 793 7873
rect 741 7849 749 7869
rect 769 7853 793 7869
rect 813 7869 885 7873
rect 813 7853 857 7869
rect 769 7849 857 7853
rect 877 7849 885 7869
rect 741 7841 885 7849
rect 741 7840 777 7841
rect 849 7840 885 7841
rect 951 7874 988 7875
rect 951 7873 989 7874
rect 951 7865 1015 7873
rect 951 7845 960 7865
rect 980 7851 1015 7865
rect 1035 7851 1038 7871
rect 980 7846 1038 7851
rect 980 7845 1015 7846
rect 234 7806 275 7831
rect 420 7806 457 7837
rect 638 7806 675 7837
rect 951 7833 1015 7845
rect 1055 7807 1082 7985
rect 234 7779 283 7806
rect 419 7780 468 7806
rect 637 7805 718 7806
rect 914 7805 1082 7807
rect 637 7780 1082 7805
rect 638 7779 1082 7780
rect 236 7746 283 7779
rect 639 7746 679 7779
rect 914 7778 1082 7779
rect 1545 7783 1585 8007
rect 1711 8006 1879 8007
rect 2482 8141 2926 8155
rect 2482 8139 2650 8141
rect 2482 7961 2509 8139
rect 2549 8101 2613 8113
rect 2889 8109 2926 8141
rect 2952 8140 3143 8162
rect 3378 8158 3487 8178
rect 3507 8158 3516 8178
rect 3378 8151 3516 8158
rect 3574 8178 3722 8187
rect 3574 8158 3583 8178
rect 3603 8158 3693 8178
rect 3713 8158 3722 8178
rect 3378 8149 3474 8151
rect 3574 8148 3722 8158
rect 3781 8178 3818 8188
rect 3781 8158 3789 8178
rect 3809 8158 3818 8178
rect 3630 8147 3666 8148
rect 3107 8138 3143 8140
rect 3107 8109 3144 8138
rect 2549 8100 2584 8101
rect 2526 8095 2584 8100
rect 2526 8075 2529 8095
rect 2549 8081 2584 8095
rect 2604 8081 2613 8101
rect 2549 8073 2613 8081
rect 2575 8072 2613 8073
rect 2576 8071 2613 8072
rect 2679 8105 2715 8106
rect 2787 8105 2823 8106
rect 2679 8099 2823 8105
rect 2679 8097 2740 8099
rect 2679 8077 2687 8097
rect 2707 8082 2740 8097
rect 2759 8097 2823 8099
rect 2759 8082 2795 8097
rect 2707 8077 2795 8082
rect 2815 8077 2823 8097
rect 2679 8071 2823 8077
rect 2889 8101 2927 8109
rect 3005 8105 3041 8106
rect 2889 8081 2898 8101
rect 2918 8081 2927 8101
rect 2889 8072 2927 8081
rect 2956 8097 3041 8105
rect 2956 8077 3013 8097
rect 3033 8077 3041 8097
rect 2889 8071 2926 8072
rect 2956 8071 3041 8077
rect 3107 8101 3145 8109
rect 3107 8081 3116 8101
rect 3136 8081 3145 8101
rect 3781 8091 3818 8158
rect 3853 8187 3884 8238
rect 4166 8226 4184 8244
rect 4202 8226 4218 8244
rect 3903 8187 3940 8188
rect 3853 8178 3940 8187
rect 3853 8158 3911 8178
rect 3931 8158 3940 8178
rect 3853 8148 3940 8158
rect 3999 8178 4036 8188
rect 3999 8158 4007 8178
rect 4027 8158 4036 8178
rect 3853 8147 3884 8148
rect 3478 8088 3515 8089
rect 3781 8088 3820 8091
rect 3477 8087 3820 8088
rect 3999 8087 4036 8158
rect 3107 8072 3145 8081
rect 3402 8082 3820 8087
rect 3107 8071 3144 8072
rect 2568 8043 2658 8049
rect 2568 8023 2584 8043
rect 2604 8041 2658 8043
rect 2604 8023 2629 8041
rect 2568 8021 2629 8023
rect 2649 8021 2658 8041
rect 2568 8015 2658 8021
rect 2581 7961 2618 7962
rect 2677 7961 2714 7962
rect 2733 7961 2769 8071
rect 2956 8050 2987 8071
rect 3402 8062 3405 8082
rect 3425 8062 3820 8082
rect 3849 8063 4036 8087
rect 2952 8049 2987 8050
rect 2830 8039 2987 8049
rect 2830 8019 2847 8039
rect 2867 8019 2987 8039
rect 2830 8012 2987 8019
rect 3054 8042 3203 8050
rect 3054 8022 3065 8042
rect 3085 8022 3124 8042
rect 3144 8022 3203 8042
rect 3054 8015 3203 8022
rect 3781 8037 3820 8062
rect 4166 8037 4218 8226
rect 4610 8254 4620 8272
rect 4638 8254 4650 8272
rect 4782 8270 4791 8290
rect 4811 8270 4820 8290
rect 4782 8262 4820 8270
rect 4886 8294 4971 8300
rect 5001 8299 5038 8300
rect 4886 8274 4894 8294
rect 4914 8274 4971 8294
rect 4886 8266 4971 8274
rect 5000 8290 5038 8299
rect 5000 8270 5009 8290
rect 5029 8270 5038 8290
rect 4886 8265 4922 8266
rect 5000 8262 5038 8270
rect 5104 8294 5248 8300
rect 5104 8274 5112 8294
rect 5132 8274 5165 8294
rect 5185 8274 5220 8294
rect 5240 8274 5248 8294
rect 5104 8266 5248 8274
rect 5104 8265 5140 8266
rect 5212 8265 5248 8266
rect 5314 8299 5351 8300
rect 5314 8298 5352 8299
rect 5314 8290 5378 8298
rect 5314 8270 5323 8290
rect 5343 8276 5378 8290
rect 5398 8276 5401 8296
rect 5343 8271 5401 8276
rect 5343 8270 5378 8271
rect 4610 8198 4650 8254
rect 4783 8233 4820 8262
rect 4784 8231 4820 8233
rect 4784 8209 4975 8231
rect 5001 8230 5038 8262
rect 5314 8258 5378 8270
rect 5418 8232 5445 8410
rect 5277 8230 5445 8232
rect 5001 8220 5445 8230
rect 5586 8326 5773 8350
rect 5804 8331 6197 8351
rect 6217 8331 6220 8351
rect 5804 8326 6220 8331
rect 5586 8255 5623 8326
rect 5804 8325 6145 8326
rect 5738 8265 5769 8266
rect 5586 8235 5595 8255
rect 5615 8235 5623 8255
rect 5586 8225 5623 8235
rect 5682 8255 5769 8265
rect 5682 8235 5691 8255
rect 5711 8235 5769 8255
rect 5682 8226 5769 8235
rect 5682 8225 5719 8226
rect 4607 8193 4650 8198
rect 4998 8204 5445 8220
rect 4998 8198 5026 8204
rect 5277 8203 5445 8204
rect 4607 8190 4757 8193
rect 4998 8190 5025 8198
rect 4607 8188 5025 8190
rect 4607 8170 4616 8188
rect 4634 8170 5025 8188
rect 5738 8175 5769 8226
rect 5804 8255 5841 8325
rect 6107 8324 6144 8325
rect 5956 8265 5992 8266
rect 5804 8235 5813 8255
rect 5833 8235 5841 8255
rect 5804 8225 5841 8235
rect 5900 8255 6048 8265
rect 6148 8262 6244 8264
rect 5900 8235 5909 8255
rect 5929 8235 6019 8255
rect 6039 8235 6048 8255
rect 5900 8226 6048 8235
rect 6106 8255 6244 8262
rect 6106 8235 6115 8255
rect 6135 8235 6244 8255
rect 6106 8226 6244 8235
rect 5900 8225 5937 8226
rect 5630 8172 5671 8173
rect 4607 8167 5025 8170
rect 4607 8161 4650 8167
rect 4610 8158 4650 8161
rect 5522 8165 5671 8172
rect 5007 8149 5047 8150
rect 4718 8132 5047 8149
rect 5522 8145 5581 8165
rect 5601 8145 5640 8165
rect 5660 8145 5671 8165
rect 5522 8137 5671 8145
rect 5738 8168 5895 8175
rect 5738 8148 5858 8168
rect 5878 8148 5895 8168
rect 5738 8138 5895 8148
rect 5738 8137 5773 8138
rect 4602 8089 4645 8100
rect 4602 8071 4614 8089
rect 4632 8071 4645 8089
rect 4602 8045 4645 8071
rect 4718 8045 4745 8132
rect 5007 8123 5047 8132
rect 3781 8019 4220 8037
rect 3054 8014 3095 8015
rect 2788 7961 2825 7962
rect 2481 7952 2619 7961
rect 2481 7932 2590 7952
rect 2610 7932 2619 7952
rect 2481 7925 2619 7932
rect 2677 7952 2825 7961
rect 2677 7932 2686 7952
rect 2706 7932 2796 7952
rect 2816 7932 2825 7952
rect 2481 7923 2577 7925
rect 2677 7922 2825 7932
rect 2884 7952 2921 7962
rect 2884 7932 2892 7952
rect 2912 7932 2921 7952
rect 2733 7921 2769 7922
rect 2581 7862 2618 7863
rect 2884 7862 2921 7932
rect 2956 7961 2987 8012
rect 3781 8001 4181 8019
rect 4199 8001 4220 8019
rect 3781 7995 4220 8001
rect 3787 7991 4220 7995
rect 4602 8024 4745 8045
rect 4789 8097 4823 8113
rect 5007 8103 5400 8123
rect 5420 8103 5423 8123
rect 5738 8116 5769 8137
rect 5956 8116 5992 8226
rect 6011 8225 6048 8226
rect 6107 8225 6144 8226
rect 6067 8166 6157 8172
rect 6067 8146 6076 8166
rect 6096 8164 6157 8166
rect 6096 8146 6121 8164
rect 6067 8144 6121 8146
rect 6141 8144 6157 8164
rect 6067 8138 6157 8144
rect 5581 8115 5618 8116
rect 5007 8098 5423 8103
rect 5580 8106 5618 8115
rect 5007 8097 5348 8098
rect 4789 8027 4826 8097
rect 4941 8037 4972 8038
rect 4602 8022 4739 8024
rect 4166 7989 4218 7991
rect 4602 7980 4645 8022
rect 4789 8007 4798 8027
rect 4818 8007 4826 8027
rect 4789 7997 4826 8007
rect 4885 8027 4972 8037
rect 4885 8007 4894 8027
rect 4914 8007 4972 8027
rect 4885 7998 4972 8007
rect 4885 7997 4922 7998
rect 4600 7970 4645 7980
rect 3006 7961 3043 7962
rect 2956 7952 3043 7961
rect 2956 7932 3014 7952
rect 3034 7932 3043 7952
rect 2956 7922 3043 7932
rect 3102 7952 3139 7962
rect 3102 7932 3110 7952
rect 3130 7932 3139 7952
rect 4600 7952 4609 7970
rect 4627 7952 4645 7970
rect 4600 7946 4645 7952
rect 4941 7947 4972 7998
rect 5007 8027 5044 8097
rect 5310 8096 5347 8097
rect 5580 8086 5589 8106
rect 5609 8086 5618 8106
rect 5580 8078 5618 8086
rect 5684 8110 5769 8116
rect 5799 8115 5836 8116
rect 5684 8090 5692 8110
rect 5712 8090 5769 8110
rect 5684 8082 5769 8090
rect 5798 8106 5836 8115
rect 5798 8086 5807 8106
rect 5827 8086 5836 8106
rect 5684 8081 5720 8082
rect 5798 8078 5836 8086
rect 5902 8110 6046 8116
rect 5902 8090 5910 8110
rect 5930 8091 5962 8110
rect 5983 8091 6018 8110
rect 5930 8090 6018 8091
rect 6038 8090 6046 8110
rect 5902 8082 6046 8090
rect 5902 8081 5938 8082
rect 6010 8081 6046 8082
rect 6112 8115 6149 8116
rect 6112 8114 6150 8115
rect 6112 8106 6176 8114
rect 6112 8086 6121 8106
rect 6141 8092 6176 8106
rect 6196 8092 6199 8112
rect 6141 8087 6199 8092
rect 6141 8086 6176 8087
rect 5581 8049 5618 8078
rect 5582 8047 5618 8049
rect 5159 8037 5195 8038
rect 5007 8007 5016 8027
rect 5036 8007 5044 8027
rect 5007 7997 5044 8007
rect 5103 8027 5251 8037
rect 5351 8034 5447 8036
rect 5103 8007 5112 8027
rect 5132 8007 5222 8027
rect 5242 8007 5251 8027
rect 5103 7998 5251 8007
rect 5309 8027 5447 8034
rect 5309 8007 5318 8027
rect 5338 8007 5447 8027
rect 5582 8025 5773 8047
rect 5799 8046 5836 8078
rect 6112 8074 6176 8086
rect 6216 8048 6243 8226
rect 6848 8225 6881 8558
rect 6945 8590 7113 8591
rect 7239 8590 7279 8814
rect 7742 8818 7910 8819
rect 8146 8818 8195 8853
rect 7742 8792 8195 8818
rect 7742 8790 7910 8792
rect 8106 8791 8188 8792
rect 8328 8791 8406 8817
rect 8546 8795 8593 8853
rect 8994 8849 9041 8854
rect 7742 8612 7769 8790
rect 7809 8752 7873 8764
rect 8149 8760 8186 8791
rect 8367 8760 8404 8791
rect 8546 8782 8594 8795
rect 7809 8751 7844 8752
rect 7786 8746 7844 8751
rect 7786 8726 7789 8746
rect 7809 8732 7844 8746
rect 7864 8732 7873 8752
rect 7809 8724 7873 8732
rect 7835 8723 7873 8724
rect 7836 8722 7873 8723
rect 7939 8756 7975 8757
rect 8047 8756 8083 8757
rect 7939 8748 8083 8756
rect 7939 8728 7947 8748
rect 7967 8744 8055 8748
rect 7967 8728 8011 8744
rect 7939 8724 8011 8728
rect 8031 8728 8055 8744
rect 8075 8728 8083 8748
rect 8031 8724 8083 8728
rect 7939 8722 8083 8724
rect 8149 8752 8187 8760
rect 8265 8756 8301 8757
rect 8149 8732 8158 8752
rect 8178 8732 8187 8752
rect 8149 8723 8187 8732
rect 8216 8748 8301 8756
rect 8216 8728 8273 8748
rect 8293 8728 8301 8748
rect 8149 8722 8186 8723
rect 8216 8722 8301 8728
rect 8367 8752 8405 8760
rect 8367 8732 8376 8752
rect 8396 8732 8405 8752
rect 8367 8723 8405 8732
rect 8549 8757 8594 8782
rect 8549 8739 8563 8757
rect 8581 8739 8594 8757
rect 8549 8731 8594 8739
rect 8554 8729 8594 8731
rect 8994 8787 9042 8849
rect 11616 8848 11656 8856
rect 11616 8826 11624 8848
rect 11648 8826 11656 8848
rect 12520 8851 12976 8886
rect 15980 8861 16020 8869
rect 8367 8722 8404 8723
rect 7828 8694 7918 8700
rect 7828 8674 7844 8694
rect 7864 8692 7918 8694
rect 7864 8674 7889 8692
rect 7828 8672 7889 8674
rect 7909 8672 7918 8692
rect 7828 8666 7918 8672
rect 7841 8612 7878 8613
rect 7937 8612 7974 8613
rect 7993 8612 8029 8722
rect 8216 8701 8247 8722
rect 8994 8707 9041 8787
rect 8212 8700 8247 8701
rect 8090 8690 8247 8700
rect 8090 8670 8107 8690
rect 8127 8670 8247 8690
rect 8090 8663 8247 8670
rect 8314 8693 8463 8701
rect 8314 8673 8325 8693
rect 8345 8673 8384 8693
rect 8404 8673 8463 8693
rect 8994 8689 9004 8707
rect 9022 8689 9041 8707
rect 8994 8685 9041 8689
rect 8995 8680 9032 8685
rect 8314 8666 8463 8673
rect 8314 8665 8355 8666
rect 8551 8664 8588 8667
rect 8048 8612 8085 8613
rect 7741 8603 7879 8612
rect 6945 8564 7389 8590
rect 6945 8562 7113 8564
rect 6945 8384 6972 8562
rect 7012 8524 7076 8536
rect 7352 8532 7389 8564
rect 7415 8563 7606 8585
rect 7741 8583 7850 8603
rect 7870 8583 7879 8603
rect 7741 8576 7879 8583
rect 7937 8603 8085 8612
rect 7937 8583 7946 8603
rect 7966 8583 8056 8603
rect 8076 8583 8085 8603
rect 7741 8574 7837 8576
rect 7937 8573 8085 8583
rect 8144 8603 8181 8613
rect 8144 8583 8152 8603
rect 8172 8583 8181 8603
rect 7993 8572 8029 8573
rect 7570 8561 7606 8563
rect 7570 8532 7607 8561
rect 7012 8523 7047 8524
rect 6989 8518 7047 8523
rect 6989 8498 6992 8518
rect 7012 8504 7047 8518
rect 7067 8504 7076 8524
rect 7012 8498 7076 8504
rect 6989 8496 7076 8498
rect 6989 8492 7016 8496
rect 7038 8495 7076 8496
rect 7039 8494 7076 8495
rect 7142 8528 7178 8529
rect 7250 8528 7286 8529
rect 7142 8521 7286 8528
rect 7142 8520 7204 8521
rect 7142 8500 7150 8520
rect 7170 8503 7204 8520
rect 7223 8520 7286 8521
rect 7223 8503 7258 8520
rect 7170 8500 7258 8503
rect 7278 8500 7286 8520
rect 7142 8494 7286 8500
rect 7352 8524 7390 8532
rect 7468 8528 7504 8529
rect 7352 8504 7361 8524
rect 7381 8504 7390 8524
rect 7352 8495 7390 8504
rect 7419 8520 7504 8528
rect 7419 8500 7476 8520
rect 7496 8500 7504 8520
rect 7352 8494 7389 8495
rect 7419 8494 7504 8500
rect 7570 8524 7608 8532
rect 7570 8504 7579 8524
rect 7599 8504 7608 8524
rect 7841 8513 7878 8514
rect 8144 8513 8181 8583
rect 8216 8612 8247 8663
rect 8543 8658 8588 8664
rect 8543 8640 8561 8658
rect 8579 8640 8588 8658
rect 8543 8630 8588 8640
rect 8266 8612 8303 8613
rect 8216 8603 8303 8612
rect 8216 8583 8274 8603
rect 8294 8583 8303 8603
rect 8216 8573 8303 8583
rect 8362 8603 8399 8613
rect 8362 8583 8370 8603
rect 8390 8583 8399 8603
rect 8543 8588 8586 8630
rect 8983 8618 9035 8620
rect 8449 8586 8586 8588
rect 8216 8572 8247 8573
rect 8362 8513 8399 8583
rect 7840 8512 8181 8513
rect 7570 8495 7608 8504
rect 7765 8507 8181 8512
rect 7570 8494 7607 8495
rect 7031 8466 7121 8472
rect 7031 8446 7047 8466
rect 7067 8464 7121 8466
rect 7067 8446 7092 8464
rect 7031 8444 7092 8446
rect 7112 8444 7121 8464
rect 7031 8438 7121 8444
rect 7044 8384 7081 8385
rect 7140 8384 7177 8385
rect 7196 8384 7232 8494
rect 7419 8473 7450 8494
rect 7765 8487 7768 8507
rect 7788 8487 8181 8507
rect 8365 8497 8399 8513
rect 8443 8565 8586 8586
rect 8981 8614 9414 8618
rect 8981 8608 9420 8614
rect 8981 8590 9002 8608
rect 9020 8590 9420 8608
rect 8981 8572 9420 8590
rect 8141 8478 8181 8487
rect 8443 8478 8470 8565
rect 8543 8539 8586 8565
rect 8543 8521 8556 8539
rect 8574 8521 8586 8539
rect 8543 8510 8586 8521
rect 7415 8472 7450 8473
rect 7293 8462 7450 8472
rect 7293 8442 7310 8462
rect 7330 8442 7450 8462
rect 7293 8435 7450 8442
rect 7517 8465 7663 8473
rect 7517 8445 7528 8465
rect 7548 8445 7587 8465
rect 7607 8445 7663 8465
rect 8141 8461 8470 8478
rect 8141 8460 8181 8461
rect 7517 8438 7663 8445
rect 8538 8449 8578 8452
rect 8538 8443 8581 8449
rect 8163 8440 8581 8443
rect 7517 8437 7558 8438
rect 7251 8384 7288 8385
rect 6944 8375 7082 8384
rect 6944 8355 7053 8375
rect 7073 8355 7082 8375
rect 6944 8348 7082 8355
rect 7140 8375 7288 8384
rect 7140 8355 7149 8375
rect 7169 8355 7259 8375
rect 7279 8355 7288 8375
rect 6944 8346 7040 8348
rect 7140 8345 7288 8355
rect 7347 8375 7384 8385
rect 7347 8355 7355 8375
rect 7375 8355 7384 8375
rect 7196 8344 7232 8345
rect 7044 8285 7081 8286
rect 7347 8285 7384 8355
rect 7419 8384 7450 8435
rect 8163 8422 8554 8440
rect 8572 8422 8581 8440
rect 8163 8420 8581 8422
rect 8163 8412 8190 8420
rect 8431 8417 8581 8420
rect 7743 8406 7911 8407
rect 8162 8406 8190 8412
rect 7743 8390 8190 8406
rect 8538 8412 8581 8417
rect 7469 8384 7506 8385
rect 7419 8375 7506 8384
rect 7419 8355 7477 8375
rect 7497 8355 7506 8375
rect 7419 8345 7506 8355
rect 7565 8375 7602 8385
rect 7565 8355 7573 8375
rect 7593 8355 7602 8375
rect 7419 8344 7450 8345
rect 7043 8284 7384 8285
rect 7565 8284 7602 8355
rect 6968 8279 7384 8284
rect 6968 8259 6971 8279
rect 6991 8259 7384 8279
rect 7415 8260 7602 8284
rect 7743 8380 8187 8390
rect 7743 8378 7911 8380
rect 6843 8180 6885 8225
rect 7743 8200 7770 8378
rect 7810 8340 7874 8352
rect 8150 8348 8187 8380
rect 8213 8379 8404 8401
rect 8368 8377 8404 8379
rect 8368 8348 8405 8377
rect 8538 8356 8578 8412
rect 7810 8339 7845 8340
rect 7787 8334 7845 8339
rect 7787 8314 7790 8334
rect 7810 8320 7845 8334
rect 7865 8320 7874 8340
rect 7810 8312 7874 8320
rect 7836 8311 7874 8312
rect 7837 8310 7874 8311
rect 7940 8344 7976 8345
rect 8048 8344 8084 8345
rect 7940 8336 8084 8344
rect 7940 8316 7948 8336
rect 7968 8316 8003 8336
rect 8023 8316 8056 8336
rect 8076 8316 8084 8336
rect 7940 8310 8084 8316
rect 8150 8340 8188 8348
rect 8266 8344 8302 8345
rect 8150 8320 8159 8340
rect 8179 8320 8188 8340
rect 8150 8311 8188 8320
rect 8217 8336 8302 8344
rect 8217 8316 8274 8336
rect 8294 8316 8302 8336
rect 8150 8310 8187 8311
rect 8217 8310 8302 8316
rect 8368 8340 8406 8348
rect 8368 8320 8377 8340
rect 8397 8320 8406 8340
rect 8538 8338 8550 8356
rect 8568 8338 8578 8356
rect 8983 8383 9035 8572
rect 9381 8547 9420 8572
rect 11221 8597 11258 8603
rect 11221 8578 11229 8597
rect 11250 8578 11258 8597
rect 11221 8570 11258 8578
rect 9165 8522 9352 8546
rect 9381 8527 9776 8547
rect 9796 8527 9799 8547
rect 9381 8522 9799 8527
rect 9165 8451 9202 8522
rect 9381 8521 9724 8522
rect 9381 8518 9420 8521
rect 9686 8520 9723 8521
rect 9317 8461 9348 8462
rect 9165 8431 9174 8451
rect 9194 8431 9202 8451
rect 9165 8421 9202 8431
rect 9261 8451 9348 8461
rect 9261 8431 9270 8451
rect 9290 8431 9348 8451
rect 9261 8422 9348 8431
rect 9261 8421 9298 8422
rect 8983 8365 8999 8383
rect 9017 8365 9035 8383
rect 9317 8371 9348 8422
rect 9383 8451 9420 8518
rect 9535 8461 9571 8462
rect 9383 8431 9392 8451
rect 9412 8431 9420 8451
rect 9383 8421 9420 8431
rect 9479 8451 9627 8461
rect 9727 8458 9823 8460
rect 9479 8431 9488 8451
rect 9508 8431 9598 8451
rect 9618 8431 9627 8451
rect 9479 8422 9627 8431
rect 9685 8451 9823 8458
rect 9685 8431 9694 8451
rect 9714 8431 9823 8451
rect 9685 8422 9823 8431
rect 9479 8421 9516 8422
rect 9209 8368 9250 8369
rect 8983 8347 9035 8365
rect 9101 8361 9250 8368
rect 8538 8328 8578 8338
rect 9101 8341 9160 8361
rect 9180 8341 9219 8361
rect 9239 8341 9250 8361
rect 9101 8333 9250 8341
rect 9317 8364 9474 8371
rect 9317 8344 9437 8364
rect 9457 8344 9474 8364
rect 9317 8334 9474 8344
rect 9317 8333 9352 8334
rect 8368 8311 8406 8320
rect 9317 8312 9348 8333
rect 9535 8312 9571 8422
rect 9590 8421 9627 8422
rect 9686 8421 9723 8422
rect 9646 8362 9736 8368
rect 9646 8342 9655 8362
rect 9675 8360 9736 8362
rect 9675 8342 9700 8360
rect 9646 8340 9700 8342
rect 9720 8340 9736 8360
rect 9646 8334 9736 8340
rect 9160 8311 9197 8312
rect 8368 8310 8405 8311
rect 7829 8282 7919 8288
rect 7829 8262 7845 8282
rect 7865 8280 7919 8282
rect 7865 8262 7890 8280
rect 7829 8260 7890 8262
rect 7910 8260 7919 8280
rect 7829 8254 7919 8260
rect 7842 8200 7879 8201
rect 7938 8200 7975 8201
rect 7994 8200 8030 8310
rect 8217 8289 8248 8310
rect 9159 8302 9197 8311
rect 8213 8288 8248 8289
rect 8091 8278 8248 8288
rect 8091 8258 8108 8278
rect 8128 8258 8248 8278
rect 8091 8251 8248 8258
rect 8315 8281 8464 8289
rect 8315 8261 8326 8281
rect 8346 8261 8385 8281
rect 8405 8261 8464 8281
rect 8987 8284 9027 8294
rect 8315 8254 8464 8261
rect 8530 8257 8582 8275
rect 8315 8253 8356 8254
rect 8049 8200 8086 8201
rect 7742 8191 7880 8200
rect 7214 8180 7247 8182
rect 6843 8168 7290 8180
rect 6075 8046 6243 8048
rect 5799 8020 6243 8046
rect 5309 7998 5447 8007
rect 5103 7997 5140 7998
rect 4600 7943 4637 7946
rect 4833 7944 4874 7945
rect 2956 7921 2987 7922
rect 2580 7861 2921 7862
rect 3102 7861 3139 7932
rect 4725 7937 4874 7944
rect 4169 7924 4206 7929
rect 4160 7920 4207 7924
rect 4160 7902 4179 7920
rect 4197 7902 4207 7920
rect 4725 7917 4784 7937
rect 4804 7917 4843 7937
rect 4863 7917 4874 7937
rect 4725 7909 4874 7917
rect 4941 7940 5098 7947
rect 4941 7920 5061 7940
rect 5081 7920 5098 7940
rect 4941 7910 5098 7920
rect 4941 7909 4976 7910
rect 2505 7856 2921 7861
rect 2505 7836 2508 7856
rect 2528 7836 2921 7856
rect 2952 7837 3139 7861
rect 3764 7859 3804 7864
rect 4160 7859 4207 7902
rect 4941 7888 4972 7909
rect 5159 7888 5195 7998
rect 5214 7997 5251 7998
rect 5310 7997 5347 7998
rect 5270 7938 5360 7944
rect 5270 7918 5279 7938
rect 5299 7936 5360 7938
rect 5299 7918 5324 7936
rect 5270 7916 5324 7918
rect 5344 7916 5360 7936
rect 5270 7910 5360 7916
rect 4784 7887 4821 7888
rect 3764 7820 4207 7859
rect 4597 7879 4634 7881
rect 4597 7871 4639 7879
rect 4597 7853 4607 7871
rect 4625 7853 4639 7871
rect 4597 7844 4639 7853
rect 4783 7878 4821 7887
rect 4783 7858 4792 7878
rect 4812 7858 4821 7878
rect 4783 7850 4821 7858
rect 4887 7882 4972 7888
rect 5002 7887 5039 7888
rect 4887 7862 4895 7882
rect 4915 7862 4972 7882
rect 4887 7854 4972 7862
rect 5001 7878 5039 7887
rect 5001 7858 5010 7878
rect 5030 7858 5039 7878
rect 4887 7853 4923 7854
rect 5001 7850 5039 7858
rect 5105 7886 5249 7888
rect 5105 7882 5157 7886
rect 5105 7862 5113 7882
rect 5133 7866 5157 7882
rect 5177 7882 5249 7886
rect 5177 7866 5221 7882
rect 5133 7862 5221 7866
rect 5241 7862 5249 7882
rect 5105 7854 5249 7862
rect 5105 7853 5141 7854
rect 5213 7853 5249 7854
rect 5315 7887 5352 7888
rect 5315 7886 5353 7887
rect 5315 7878 5379 7886
rect 5315 7858 5324 7878
rect 5344 7864 5379 7878
rect 5399 7864 5402 7884
rect 5344 7859 5402 7864
rect 5344 7858 5379 7859
rect 1545 7761 1553 7783
rect 1577 7761 1585 7783
rect 1545 7753 1585 7761
rect 2858 7805 2898 7813
rect 2858 7783 2866 7805
rect 2890 7783 2898 7805
rect 236 7707 679 7746
rect 236 7664 283 7707
rect 639 7702 679 7707
rect 1304 7705 1491 7729
rect 1522 7710 1915 7730
rect 1935 7710 1938 7730
rect 1522 7705 1938 7710
rect 236 7646 246 7664
rect 264 7646 283 7664
rect 236 7642 283 7646
rect 237 7637 274 7642
rect 1304 7634 1341 7705
rect 1522 7704 1863 7705
rect 1456 7644 1487 7645
rect 1304 7614 1313 7634
rect 1333 7614 1341 7634
rect 1304 7604 1341 7614
rect 1400 7634 1487 7644
rect 1400 7614 1409 7634
rect 1429 7614 1487 7634
rect 1400 7605 1487 7614
rect 1400 7604 1437 7605
rect 225 7575 277 7577
rect 223 7571 656 7575
rect 223 7565 662 7571
rect 223 7547 244 7565
rect 262 7547 662 7565
rect 1456 7554 1487 7605
rect 1522 7634 1559 7704
rect 1825 7703 1862 7704
rect 1674 7644 1710 7645
rect 1522 7614 1531 7634
rect 1551 7614 1559 7634
rect 1522 7604 1559 7614
rect 1618 7634 1766 7644
rect 1866 7641 1962 7643
rect 1618 7614 1627 7634
rect 1647 7614 1737 7634
rect 1757 7614 1766 7634
rect 1618 7605 1766 7614
rect 1824 7634 1962 7641
rect 1824 7614 1833 7634
rect 1853 7614 1962 7634
rect 1824 7605 1962 7614
rect 1618 7604 1655 7605
rect 1348 7551 1389 7552
rect 223 7529 662 7547
rect 225 7340 277 7529
rect 623 7504 662 7529
rect 1240 7544 1389 7551
rect 1240 7524 1299 7544
rect 1319 7524 1358 7544
rect 1378 7524 1389 7544
rect 1240 7516 1389 7524
rect 1456 7547 1613 7554
rect 1456 7527 1576 7547
rect 1596 7527 1613 7547
rect 1456 7517 1613 7527
rect 1456 7516 1491 7517
rect 407 7479 594 7503
rect 623 7484 1018 7504
rect 1038 7484 1041 7504
rect 1456 7495 1487 7516
rect 1674 7495 1710 7605
rect 1729 7604 1766 7605
rect 1825 7604 1862 7605
rect 1785 7545 1875 7551
rect 1785 7525 1794 7545
rect 1814 7543 1875 7545
rect 1814 7525 1839 7543
rect 1785 7523 1839 7525
rect 1859 7523 1875 7543
rect 1785 7517 1875 7523
rect 1299 7494 1336 7495
rect 623 7479 1041 7484
rect 1298 7485 1336 7494
rect 407 7408 444 7479
rect 623 7478 966 7479
rect 623 7475 662 7478
rect 928 7477 965 7478
rect 559 7418 590 7419
rect 407 7388 416 7408
rect 436 7388 444 7408
rect 407 7378 444 7388
rect 503 7408 590 7418
rect 503 7388 512 7408
rect 532 7388 590 7408
rect 503 7379 590 7388
rect 503 7378 540 7379
rect 225 7322 241 7340
rect 259 7322 277 7340
rect 559 7328 590 7379
rect 625 7408 662 7475
rect 1298 7465 1307 7485
rect 1327 7465 1336 7485
rect 1298 7457 1336 7465
rect 1402 7489 1487 7495
rect 1517 7494 1554 7495
rect 1402 7469 1410 7489
rect 1430 7469 1487 7489
rect 1402 7461 1487 7469
rect 1516 7485 1554 7494
rect 1516 7465 1525 7485
rect 1545 7465 1554 7485
rect 1402 7460 1438 7461
rect 1516 7457 1554 7465
rect 1620 7490 1764 7495
rect 1620 7489 1682 7490
rect 1620 7469 1628 7489
rect 1648 7471 1682 7489
rect 1703 7489 1764 7490
rect 1703 7471 1736 7489
rect 1648 7469 1736 7471
rect 1756 7469 1764 7489
rect 1620 7461 1764 7469
rect 1620 7460 1656 7461
rect 1728 7460 1764 7461
rect 1830 7494 1867 7495
rect 1830 7493 1868 7494
rect 1830 7485 1894 7493
rect 1830 7465 1839 7485
rect 1859 7471 1894 7485
rect 1914 7471 1917 7491
rect 1859 7466 1917 7471
rect 1859 7465 1894 7466
rect 1299 7428 1336 7457
rect 1300 7426 1336 7428
rect 777 7418 813 7419
rect 625 7388 634 7408
rect 654 7388 662 7408
rect 625 7378 662 7388
rect 721 7408 869 7418
rect 969 7415 1065 7417
rect 721 7388 730 7408
rect 750 7388 840 7408
rect 860 7388 869 7408
rect 721 7379 869 7388
rect 927 7408 1065 7415
rect 927 7388 936 7408
rect 956 7388 1065 7408
rect 1300 7404 1491 7426
rect 1517 7425 1554 7457
rect 1830 7453 1894 7465
rect 1934 7427 1961 7605
rect 1793 7425 1961 7427
rect 1517 7411 1961 7425
rect 2564 7559 2732 7560
rect 2858 7559 2898 7783
rect 3361 7787 3529 7788
rect 3764 7787 3804 7820
rect 4160 7787 4207 7820
rect 4598 7819 4639 7844
rect 4784 7819 4821 7850
rect 5002 7819 5039 7850
rect 5315 7846 5379 7858
rect 5419 7820 5446 7998
rect 4598 7792 4647 7819
rect 4783 7793 4832 7819
rect 5001 7818 5082 7819
rect 5278 7818 5446 7820
rect 5001 7793 5446 7818
rect 5002 7792 5446 7793
rect 3361 7786 3805 7787
rect 3361 7761 3806 7786
rect 3361 7759 3529 7761
rect 3725 7760 3806 7761
rect 3975 7760 4024 7786
rect 4160 7760 4209 7787
rect 3361 7581 3388 7759
rect 3428 7721 3492 7733
rect 3768 7729 3805 7760
rect 3986 7729 4023 7760
rect 4168 7735 4209 7760
rect 4600 7759 4647 7792
rect 5003 7759 5043 7792
rect 5278 7791 5446 7792
rect 5909 7796 5949 8020
rect 6075 8019 6243 8020
rect 6846 8154 7290 8168
rect 6846 8152 7014 8154
rect 6846 7974 6873 8152
rect 6913 8114 6977 8126
rect 7253 8122 7290 8154
rect 7316 8153 7507 8175
rect 7742 8171 7851 8191
rect 7871 8171 7880 8191
rect 7742 8164 7880 8171
rect 7938 8191 8086 8200
rect 7938 8171 7947 8191
rect 7967 8171 8057 8191
rect 8077 8171 8086 8191
rect 7742 8162 7838 8164
rect 7938 8161 8086 8171
rect 8145 8191 8182 8201
rect 8145 8171 8153 8191
rect 8173 8171 8182 8191
rect 7994 8160 8030 8161
rect 7471 8151 7507 8153
rect 7471 8122 7508 8151
rect 6913 8113 6948 8114
rect 6890 8108 6948 8113
rect 6890 8088 6893 8108
rect 6913 8094 6948 8108
rect 6968 8094 6977 8114
rect 6913 8086 6977 8094
rect 6939 8085 6977 8086
rect 6940 8084 6977 8085
rect 7043 8118 7079 8119
rect 7151 8118 7187 8119
rect 7043 8112 7187 8118
rect 7043 8110 7104 8112
rect 7043 8090 7051 8110
rect 7071 8095 7104 8110
rect 7123 8110 7187 8112
rect 7123 8095 7159 8110
rect 7071 8090 7159 8095
rect 7179 8090 7187 8110
rect 7043 8084 7187 8090
rect 7253 8114 7291 8122
rect 7369 8118 7405 8119
rect 7253 8094 7262 8114
rect 7282 8094 7291 8114
rect 7253 8085 7291 8094
rect 7320 8110 7405 8118
rect 7320 8090 7377 8110
rect 7397 8090 7405 8110
rect 7253 8084 7290 8085
rect 7320 8084 7405 8090
rect 7471 8114 7509 8122
rect 7471 8094 7480 8114
rect 7500 8094 7509 8114
rect 8145 8104 8182 8171
rect 8217 8200 8248 8251
rect 8530 8239 8548 8257
rect 8566 8239 8582 8257
rect 8267 8200 8304 8201
rect 8217 8191 8304 8200
rect 8217 8171 8275 8191
rect 8295 8171 8304 8191
rect 8217 8161 8304 8171
rect 8363 8191 8400 8201
rect 8363 8171 8371 8191
rect 8391 8171 8400 8191
rect 8217 8160 8248 8161
rect 7842 8101 7879 8102
rect 8145 8101 8184 8104
rect 7841 8100 8184 8101
rect 8363 8100 8400 8171
rect 7471 8085 7509 8094
rect 7766 8095 8184 8100
rect 7471 8084 7508 8085
rect 6932 8056 7022 8062
rect 6932 8036 6948 8056
rect 6968 8054 7022 8056
rect 6968 8036 6993 8054
rect 6932 8034 6993 8036
rect 7013 8034 7022 8054
rect 6932 8028 7022 8034
rect 6945 7974 6982 7975
rect 7041 7974 7078 7975
rect 7097 7974 7133 8084
rect 7320 8063 7351 8084
rect 7766 8075 7769 8095
rect 7789 8075 8184 8095
rect 8213 8076 8400 8100
rect 7316 8062 7351 8063
rect 7194 8052 7351 8062
rect 7194 8032 7211 8052
rect 7231 8032 7351 8052
rect 7194 8025 7351 8032
rect 7418 8055 7567 8063
rect 7418 8035 7429 8055
rect 7449 8035 7488 8055
rect 7508 8035 7567 8055
rect 7418 8028 7567 8035
rect 8145 8050 8184 8075
rect 8530 8050 8582 8239
rect 8987 8266 8997 8284
rect 9015 8266 9027 8284
rect 9159 8282 9168 8302
rect 9188 8282 9197 8302
rect 9159 8274 9197 8282
rect 9263 8306 9348 8312
rect 9378 8311 9415 8312
rect 9263 8286 9271 8306
rect 9291 8286 9348 8306
rect 9263 8278 9348 8286
rect 9377 8302 9415 8311
rect 9377 8282 9386 8302
rect 9406 8282 9415 8302
rect 9263 8277 9299 8278
rect 9377 8274 9415 8282
rect 9481 8306 9625 8312
rect 9481 8286 9489 8306
rect 9509 8286 9542 8306
rect 9562 8286 9597 8306
rect 9617 8286 9625 8306
rect 9481 8278 9625 8286
rect 9481 8277 9517 8278
rect 9589 8277 9625 8278
rect 9691 8311 9728 8312
rect 9691 8310 9729 8311
rect 9691 8302 9755 8310
rect 9691 8282 9700 8302
rect 9720 8288 9755 8302
rect 9775 8288 9778 8308
rect 9720 8283 9778 8288
rect 9720 8282 9755 8283
rect 8987 8210 9027 8266
rect 9160 8245 9197 8274
rect 9161 8243 9197 8245
rect 9161 8221 9352 8243
rect 9378 8242 9415 8274
rect 9691 8270 9755 8282
rect 9795 8244 9822 8422
rect 9654 8242 9822 8244
rect 9378 8232 9822 8242
rect 9963 8338 10150 8362
rect 10181 8343 10574 8363
rect 10594 8343 10597 8363
rect 10181 8338 10597 8343
rect 9963 8267 10000 8338
rect 10181 8337 10522 8338
rect 10115 8277 10146 8278
rect 9963 8247 9972 8267
rect 9992 8247 10000 8267
rect 9963 8237 10000 8247
rect 10059 8267 10146 8277
rect 10059 8247 10068 8267
rect 10088 8247 10146 8267
rect 10059 8238 10146 8247
rect 10059 8237 10096 8238
rect 8984 8205 9027 8210
rect 9375 8216 9822 8232
rect 9375 8210 9403 8216
rect 9654 8215 9822 8216
rect 8984 8202 9134 8205
rect 9375 8202 9402 8210
rect 8984 8200 9402 8202
rect 8984 8182 8993 8200
rect 9011 8182 9402 8200
rect 10115 8187 10146 8238
rect 10181 8267 10218 8337
rect 10484 8336 10521 8337
rect 10333 8277 10369 8278
rect 10181 8247 10190 8267
rect 10210 8247 10218 8267
rect 10181 8237 10218 8247
rect 10277 8267 10425 8277
rect 10525 8274 10621 8276
rect 10277 8247 10286 8267
rect 10306 8247 10396 8267
rect 10416 8247 10425 8267
rect 10277 8238 10425 8247
rect 10483 8267 10621 8274
rect 10483 8247 10492 8267
rect 10512 8247 10621 8267
rect 10483 8238 10621 8247
rect 10277 8237 10314 8238
rect 10007 8184 10048 8185
rect 8984 8179 9402 8182
rect 8984 8173 9027 8179
rect 8987 8170 9027 8173
rect 9899 8177 10048 8184
rect 9384 8161 9424 8162
rect 9095 8144 9424 8161
rect 9899 8157 9958 8177
rect 9978 8157 10017 8177
rect 10037 8157 10048 8177
rect 9899 8149 10048 8157
rect 10115 8180 10272 8187
rect 10115 8160 10235 8180
rect 10255 8160 10272 8180
rect 10115 8150 10272 8160
rect 10115 8149 10150 8150
rect 8979 8101 9022 8112
rect 8979 8083 8991 8101
rect 9009 8083 9022 8101
rect 8979 8057 9022 8083
rect 9095 8057 9122 8144
rect 9384 8135 9424 8144
rect 8145 8032 8584 8050
rect 7418 8027 7459 8028
rect 7152 7974 7189 7975
rect 6845 7965 6983 7974
rect 6845 7945 6954 7965
rect 6974 7945 6983 7965
rect 6845 7938 6983 7945
rect 7041 7965 7189 7974
rect 7041 7945 7050 7965
rect 7070 7945 7160 7965
rect 7180 7945 7189 7965
rect 6845 7936 6941 7938
rect 7041 7935 7189 7945
rect 7248 7965 7285 7975
rect 7248 7945 7256 7965
rect 7276 7945 7285 7965
rect 7097 7934 7133 7935
rect 6945 7875 6982 7876
rect 7248 7875 7285 7945
rect 7320 7974 7351 8025
rect 8145 8014 8545 8032
rect 8563 8014 8584 8032
rect 8145 8008 8584 8014
rect 8151 8004 8584 8008
rect 8979 8036 9122 8057
rect 9166 8109 9200 8125
rect 9384 8115 9777 8135
rect 9797 8115 9800 8135
rect 10115 8128 10146 8149
rect 10333 8128 10369 8238
rect 10388 8237 10425 8238
rect 10484 8237 10521 8238
rect 10444 8178 10534 8184
rect 10444 8158 10453 8178
rect 10473 8176 10534 8178
rect 10473 8158 10498 8176
rect 10444 8156 10498 8158
rect 10518 8156 10534 8176
rect 10444 8150 10534 8156
rect 9958 8127 9995 8128
rect 9384 8110 9800 8115
rect 9957 8118 9995 8127
rect 9384 8109 9725 8110
rect 9166 8039 9203 8109
rect 9318 8049 9349 8050
rect 8979 8034 9116 8036
rect 8530 8002 8582 8004
rect 8979 7992 9022 8034
rect 9166 8019 9175 8039
rect 9195 8019 9203 8039
rect 9166 8009 9203 8019
rect 9262 8039 9349 8049
rect 9262 8019 9271 8039
rect 9291 8019 9349 8039
rect 9262 8010 9349 8019
rect 9262 8009 9299 8010
rect 8977 7982 9022 7992
rect 7370 7974 7407 7975
rect 7320 7965 7407 7974
rect 7320 7945 7378 7965
rect 7398 7945 7407 7965
rect 7320 7935 7407 7945
rect 7466 7965 7503 7975
rect 7466 7945 7474 7965
rect 7494 7945 7503 7965
rect 8977 7964 8986 7982
rect 9004 7964 9022 7982
rect 8977 7958 9022 7964
rect 9318 7959 9349 8010
rect 9384 8039 9421 8109
rect 9687 8108 9724 8109
rect 9957 8098 9966 8118
rect 9986 8098 9995 8118
rect 9957 8090 9995 8098
rect 10061 8122 10146 8128
rect 10176 8127 10213 8128
rect 10061 8102 10069 8122
rect 10089 8102 10146 8122
rect 10061 8094 10146 8102
rect 10175 8118 10213 8127
rect 10175 8098 10184 8118
rect 10204 8098 10213 8118
rect 10061 8093 10097 8094
rect 10175 8090 10213 8098
rect 10279 8122 10423 8128
rect 10279 8102 10287 8122
rect 10307 8103 10339 8122
rect 10360 8103 10395 8122
rect 10307 8102 10395 8103
rect 10415 8102 10423 8122
rect 10279 8094 10423 8102
rect 10279 8093 10315 8094
rect 10387 8093 10423 8094
rect 10489 8127 10526 8128
rect 10489 8126 10527 8127
rect 10489 8118 10553 8126
rect 10489 8098 10498 8118
rect 10518 8104 10553 8118
rect 10573 8104 10576 8124
rect 10518 8099 10576 8104
rect 10518 8098 10553 8099
rect 9958 8061 9995 8090
rect 9959 8059 9995 8061
rect 9536 8049 9572 8050
rect 9384 8019 9393 8039
rect 9413 8019 9421 8039
rect 9384 8009 9421 8019
rect 9480 8039 9628 8049
rect 9728 8046 9824 8048
rect 9480 8019 9489 8039
rect 9509 8019 9599 8039
rect 9619 8019 9628 8039
rect 9480 8010 9628 8019
rect 9686 8039 9824 8046
rect 9686 8019 9695 8039
rect 9715 8019 9824 8039
rect 9959 8037 10150 8059
rect 10176 8058 10213 8090
rect 10489 8086 10553 8098
rect 10593 8060 10620 8238
rect 11225 8237 11258 8570
rect 11322 8602 11490 8603
rect 11616 8602 11656 8826
rect 12119 8830 12287 8831
rect 12520 8830 12565 8851
rect 12119 8804 12565 8830
rect 12119 8802 12287 8804
rect 12483 8803 12565 8804
rect 12700 8803 12781 8829
rect 12925 8816 13406 8851
rect 15980 8839 15988 8861
rect 16012 8839 16020 8861
rect 12119 8624 12146 8802
rect 12186 8764 12250 8776
rect 12526 8772 12563 8803
rect 12744 8772 12781 8803
rect 12928 8797 12967 8816
rect 12926 8778 12967 8797
rect 12186 8763 12221 8764
rect 12163 8758 12221 8763
rect 12163 8738 12166 8758
rect 12186 8744 12221 8758
rect 12241 8744 12250 8764
rect 12186 8736 12250 8744
rect 12212 8735 12250 8736
rect 12213 8734 12250 8735
rect 12316 8768 12352 8769
rect 12424 8768 12460 8769
rect 12316 8760 12460 8768
rect 12316 8740 12324 8760
rect 12344 8756 12432 8760
rect 12344 8740 12388 8756
rect 12316 8736 12388 8740
rect 12408 8740 12432 8756
rect 12452 8740 12460 8760
rect 12408 8736 12460 8740
rect 12316 8734 12460 8736
rect 12526 8764 12564 8772
rect 12642 8768 12678 8769
rect 12526 8744 12535 8764
rect 12555 8744 12564 8764
rect 12526 8735 12564 8744
rect 12593 8760 12678 8768
rect 12593 8740 12650 8760
rect 12670 8740 12678 8760
rect 12526 8734 12563 8735
rect 12593 8734 12678 8740
rect 12744 8764 12782 8772
rect 12744 8744 12753 8764
rect 12773 8744 12782 8764
rect 12744 8735 12782 8744
rect 12926 8769 12968 8778
rect 12926 8751 12940 8769
rect 12958 8751 12968 8769
rect 12926 8743 12968 8751
rect 12931 8741 12968 8743
rect 12744 8734 12781 8735
rect 12205 8706 12295 8712
rect 12205 8686 12221 8706
rect 12241 8704 12295 8706
rect 12241 8686 12266 8704
rect 12205 8684 12266 8686
rect 12286 8684 12295 8704
rect 12205 8678 12295 8684
rect 12218 8624 12255 8625
rect 12314 8624 12351 8625
rect 12370 8624 12406 8734
rect 12593 8713 12624 8734
rect 13358 8720 13405 8816
rect 12589 8712 12624 8713
rect 12467 8702 12624 8712
rect 12467 8682 12484 8702
rect 12504 8682 12624 8702
rect 12467 8675 12624 8682
rect 12691 8705 12840 8713
rect 12691 8685 12702 8705
rect 12722 8685 12761 8705
rect 12781 8685 12840 8705
rect 13358 8702 13368 8720
rect 13386 8702 13405 8720
rect 13358 8698 13405 8702
rect 13359 8693 13396 8698
rect 12691 8678 12840 8685
rect 12691 8677 12732 8678
rect 12928 8676 12965 8679
rect 12425 8624 12462 8625
rect 12118 8615 12256 8624
rect 11322 8576 11766 8602
rect 11322 8574 11490 8576
rect 11322 8396 11349 8574
rect 11389 8536 11453 8548
rect 11729 8544 11766 8576
rect 11792 8575 11983 8597
rect 12118 8595 12227 8615
rect 12247 8595 12256 8615
rect 12118 8588 12256 8595
rect 12314 8615 12462 8624
rect 12314 8595 12323 8615
rect 12343 8595 12433 8615
rect 12453 8595 12462 8615
rect 12118 8586 12214 8588
rect 12314 8585 12462 8595
rect 12521 8615 12558 8625
rect 12521 8595 12529 8615
rect 12549 8595 12558 8615
rect 12370 8584 12406 8585
rect 11947 8573 11983 8575
rect 11947 8544 11984 8573
rect 11389 8535 11424 8536
rect 11366 8530 11424 8535
rect 11366 8510 11369 8530
rect 11389 8516 11424 8530
rect 11444 8516 11453 8536
rect 11389 8510 11453 8516
rect 11366 8508 11453 8510
rect 11366 8504 11393 8508
rect 11415 8507 11453 8508
rect 11416 8506 11453 8507
rect 11519 8540 11555 8541
rect 11627 8540 11663 8541
rect 11519 8533 11663 8540
rect 11519 8532 11581 8533
rect 11519 8512 11527 8532
rect 11547 8515 11581 8532
rect 11600 8532 11663 8533
rect 11600 8515 11635 8532
rect 11547 8512 11635 8515
rect 11655 8512 11663 8532
rect 11519 8506 11663 8512
rect 11729 8536 11767 8544
rect 11845 8540 11881 8541
rect 11729 8516 11738 8536
rect 11758 8516 11767 8536
rect 11729 8507 11767 8516
rect 11796 8532 11881 8540
rect 11796 8512 11853 8532
rect 11873 8512 11881 8532
rect 11729 8506 11766 8507
rect 11796 8506 11881 8512
rect 11947 8536 11985 8544
rect 11947 8516 11956 8536
rect 11976 8516 11985 8536
rect 12218 8525 12255 8526
rect 12521 8525 12558 8595
rect 12593 8624 12624 8675
rect 12920 8670 12965 8676
rect 12920 8652 12938 8670
rect 12956 8652 12965 8670
rect 12920 8642 12965 8652
rect 12643 8624 12680 8625
rect 12593 8615 12680 8624
rect 12593 8595 12651 8615
rect 12671 8595 12680 8615
rect 12593 8585 12680 8595
rect 12739 8615 12776 8625
rect 12739 8595 12747 8615
rect 12767 8595 12776 8615
rect 12920 8600 12963 8642
rect 13347 8631 13399 8633
rect 12826 8598 12963 8600
rect 12593 8584 12624 8585
rect 12739 8525 12776 8595
rect 12217 8524 12558 8525
rect 11947 8507 11985 8516
rect 12142 8519 12558 8524
rect 11947 8506 11984 8507
rect 11408 8478 11498 8484
rect 11408 8458 11424 8478
rect 11444 8476 11498 8478
rect 11444 8458 11469 8476
rect 11408 8456 11469 8458
rect 11489 8456 11498 8476
rect 11408 8450 11498 8456
rect 11421 8396 11458 8397
rect 11517 8396 11554 8397
rect 11573 8396 11609 8506
rect 11796 8485 11827 8506
rect 12142 8499 12145 8519
rect 12165 8499 12558 8519
rect 12742 8509 12776 8525
rect 12820 8577 12963 8598
rect 13345 8627 13778 8631
rect 13345 8621 13784 8627
rect 13345 8603 13366 8621
rect 13384 8603 13784 8621
rect 13345 8585 13784 8603
rect 12518 8490 12558 8499
rect 12820 8490 12847 8577
rect 12920 8551 12963 8577
rect 12920 8533 12933 8551
rect 12951 8533 12963 8551
rect 12920 8522 12963 8533
rect 11792 8484 11827 8485
rect 11670 8474 11827 8484
rect 11670 8454 11687 8474
rect 11707 8454 11827 8474
rect 11670 8447 11827 8454
rect 11894 8477 12040 8485
rect 11894 8457 11905 8477
rect 11925 8457 11964 8477
rect 11984 8457 12040 8477
rect 12518 8473 12847 8490
rect 12518 8472 12558 8473
rect 11894 8450 12040 8457
rect 12915 8461 12955 8464
rect 12915 8455 12958 8461
rect 12540 8452 12958 8455
rect 11894 8449 11935 8450
rect 11628 8396 11665 8397
rect 11321 8387 11459 8396
rect 11321 8367 11430 8387
rect 11450 8367 11459 8387
rect 11321 8360 11459 8367
rect 11517 8387 11665 8396
rect 11517 8367 11526 8387
rect 11546 8367 11636 8387
rect 11656 8367 11665 8387
rect 11321 8358 11417 8360
rect 11517 8357 11665 8367
rect 11724 8387 11761 8397
rect 11724 8367 11732 8387
rect 11752 8367 11761 8387
rect 11573 8356 11609 8357
rect 11421 8297 11458 8298
rect 11724 8297 11761 8367
rect 11796 8396 11827 8447
rect 12540 8434 12931 8452
rect 12949 8434 12958 8452
rect 12540 8432 12958 8434
rect 12540 8424 12567 8432
rect 12808 8429 12958 8432
rect 12120 8418 12288 8419
rect 12539 8418 12567 8424
rect 12120 8402 12567 8418
rect 12915 8424 12958 8429
rect 11846 8396 11883 8397
rect 11796 8387 11883 8396
rect 11796 8367 11854 8387
rect 11874 8367 11883 8387
rect 11796 8357 11883 8367
rect 11942 8387 11979 8397
rect 11942 8367 11950 8387
rect 11970 8367 11979 8387
rect 11796 8356 11827 8357
rect 11420 8296 11761 8297
rect 11942 8296 11979 8367
rect 11345 8291 11761 8296
rect 11345 8271 11348 8291
rect 11368 8271 11761 8291
rect 11792 8272 11979 8296
rect 12120 8392 12564 8402
rect 12120 8390 12288 8392
rect 11220 8192 11262 8237
rect 12120 8212 12147 8390
rect 12187 8352 12251 8364
rect 12527 8360 12564 8392
rect 12590 8391 12781 8413
rect 12745 8389 12781 8391
rect 12745 8360 12782 8389
rect 12915 8368 12955 8424
rect 12187 8351 12222 8352
rect 12164 8346 12222 8351
rect 12164 8326 12167 8346
rect 12187 8332 12222 8346
rect 12242 8332 12251 8352
rect 12187 8324 12251 8332
rect 12213 8323 12251 8324
rect 12214 8322 12251 8323
rect 12317 8356 12353 8357
rect 12425 8356 12461 8357
rect 12317 8348 12461 8356
rect 12317 8328 12325 8348
rect 12345 8328 12380 8348
rect 12400 8328 12433 8348
rect 12453 8328 12461 8348
rect 12317 8322 12461 8328
rect 12527 8352 12565 8360
rect 12643 8356 12679 8357
rect 12527 8332 12536 8352
rect 12556 8332 12565 8352
rect 12527 8323 12565 8332
rect 12594 8348 12679 8356
rect 12594 8328 12651 8348
rect 12671 8328 12679 8348
rect 12527 8322 12564 8323
rect 12594 8322 12679 8328
rect 12745 8352 12783 8360
rect 12745 8332 12754 8352
rect 12774 8332 12783 8352
rect 12915 8350 12927 8368
rect 12945 8350 12955 8368
rect 13347 8396 13399 8585
rect 13745 8560 13784 8585
rect 15585 8610 15622 8616
rect 15585 8591 15593 8610
rect 15614 8591 15622 8610
rect 15585 8583 15622 8591
rect 13529 8535 13716 8559
rect 13745 8540 14140 8560
rect 14160 8540 14163 8560
rect 13745 8535 14163 8540
rect 13529 8464 13566 8535
rect 13745 8534 14088 8535
rect 13745 8531 13784 8534
rect 14050 8533 14087 8534
rect 13681 8474 13712 8475
rect 13529 8444 13538 8464
rect 13558 8444 13566 8464
rect 13529 8434 13566 8444
rect 13625 8464 13712 8474
rect 13625 8444 13634 8464
rect 13654 8444 13712 8464
rect 13625 8435 13712 8444
rect 13625 8434 13662 8435
rect 13347 8378 13363 8396
rect 13381 8378 13399 8396
rect 13681 8384 13712 8435
rect 13747 8464 13784 8531
rect 13899 8474 13935 8475
rect 13747 8444 13756 8464
rect 13776 8444 13784 8464
rect 13747 8434 13784 8444
rect 13843 8464 13991 8474
rect 14091 8471 14187 8473
rect 13843 8444 13852 8464
rect 13872 8444 13962 8464
rect 13982 8444 13991 8464
rect 13843 8435 13991 8444
rect 14049 8464 14187 8471
rect 14049 8444 14058 8464
rect 14078 8444 14187 8464
rect 14049 8435 14187 8444
rect 13843 8434 13880 8435
rect 13573 8381 13614 8382
rect 13347 8360 13399 8378
rect 13465 8374 13614 8381
rect 12915 8340 12955 8350
rect 13465 8354 13524 8374
rect 13544 8354 13583 8374
rect 13603 8354 13614 8374
rect 13465 8346 13614 8354
rect 13681 8377 13838 8384
rect 13681 8357 13801 8377
rect 13821 8357 13838 8377
rect 13681 8347 13838 8357
rect 13681 8346 13716 8347
rect 12745 8323 12783 8332
rect 13681 8325 13712 8346
rect 13899 8325 13935 8435
rect 13954 8434 13991 8435
rect 14050 8434 14087 8435
rect 14010 8375 14100 8381
rect 14010 8355 14019 8375
rect 14039 8373 14100 8375
rect 14039 8355 14064 8373
rect 14010 8353 14064 8355
rect 14084 8353 14100 8373
rect 14010 8347 14100 8353
rect 13524 8324 13561 8325
rect 12745 8322 12782 8323
rect 12206 8294 12296 8300
rect 12206 8274 12222 8294
rect 12242 8292 12296 8294
rect 12242 8274 12267 8292
rect 12206 8272 12267 8274
rect 12287 8272 12296 8292
rect 12206 8266 12296 8272
rect 12219 8212 12256 8213
rect 12315 8212 12352 8213
rect 12371 8212 12407 8322
rect 12594 8301 12625 8322
rect 13523 8315 13561 8324
rect 12590 8300 12625 8301
rect 12468 8290 12625 8300
rect 12468 8270 12485 8290
rect 12505 8270 12625 8290
rect 12468 8263 12625 8270
rect 12692 8293 12841 8301
rect 12692 8273 12703 8293
rect 12723 8273 12762 8293
rect 12782 8273 12841 8293
rect 13351 8297 13391 8307
rect 12692 8266 12841 8273
rect 12907 8269 12959 8287
rect 12692 8265 12733 8266
rect 12426 8212 12463 8213
rect 12119 8203 12257 8212
rect 11591 8192 11624 8194
rect 11220 8180 11667 8192
rect 10452 8058 10620 8060
rect 10176 8032 10620 8058
rect 9686 8010 9824 8019
rect 9480 8009 9517 8010
rect 8977 7955 9014 7958
rect 9210 7956 9251 7957
rect 7320 7934 7351 7935
rect 6944 7874 7285 7875
rect 7466 7874 7503 7945
rect 9102 7949 9251 7956
rect 8533 7937 8570 7942
rect 8524 7933 8571 7937
rect 8524 7915 8543 7933
rect 8561 7915 8571 7933
rect 9102 7929 9161 7949
rect 9181 7929 9220 7949
rect 9240 7929 9251 7949
rect 9102 7921 9251 7929
rect 9318 7952 9475 7959
rect 9318 7932 9438 7952
rect 9458 7932 9475 7952
rect 9318 7922 9475 7932
rect 9318 7921 9353 7922
rect 6869 7869 7285 7874
rect 6869 7849 6872 7869
rect 6892 7849 7285 7869
rect 7316 7850 7503 7874
rect 8128 7872 8168 7877
rect 8524 7872 8571 7915
rect 9318 7900 9349 7921
rect 9536 7900 9572 8010
rect 9591 8009 9628 8010
rect 9687 8009 9724 8010
rect 9647 7950 9737 7956
rect 9647 7930 9656 7950
rect 9676 7948 9737 7950
rect 9676 7930 9701 7948
rect 9647 7928 9701 7930
rect 9721 7928 9737 7948
rect 9647 7922 9737 7928
rect 9161 7899 9198 7900
rect 8128 7833 8571 7872
rect 8974 7891 9011 7893
rect 8974 7883 9016 7891
rect 8974 7865 8984 7883
rect 9002 7865 9016 7883
rect 8974 7856 9016 7865
rect 9160 7890 9198 7899
rect 9160 7870 9169 7890
rect 9189 7870 9198 7890
rect 9160 7862 9198 7870
rect 9264 7894 9349 7900
rect 9379 7899 9416 7900
rect 9264 7874 9272 7894
rect 9292 7874 9349 7894
rect 9264 7866 9349 7874
rect 9378 7890 9416 7899
rect 9378 7870 9387 7890
rect 9407 7870 9416 7890
rect 9264 7865 9300 7866
rect 9378 7862 9416 7870
rect 9482 7898 9626 7900
rect 9482 7894 9534 7898
rect 9482 7874 9490 7894
rect 9510 7878 9534 7894
rect 9554 7894 9626 7898
rect 9554 7878 9598 7894
rect 9510 7874 9598 7878
rect 9618 7874 9626 7894
rect 9482 7866 9626 7874
rect 9482 7865 9518 7866
rect 9590 7865 9626 7866
rect 9692 7899 9729 7900
rect 9692 7898 9730 7899
rect 9692 7890 9756 7898
rect 9692 7870 9701 7890
rect 9721 7876 9756 7890
rect 9776 7876 9779 7896
rect 9721 7871 9779 7876
rect 9721 7870 9756 7871
rect 5909 7774 5917 7796
rect 5941 7774 5949 7796
rect 5909 7766 5949 7774
rect 7222 7818 7262 7826
rect 7222 7796 7230 7818
rect 7254 7796 7262 7818
rect 3428 7720 3463 7721
rect 3405 7715 3463 7720
rect 3405 7695 3408 7715
rect 3428 7701 3463 7715
rect 3483 7701 3492 7721
rect 3428 7693 3492 7701
rect 3454 7692 3492 7693
rect 3455 7691 3492 7692
rect 3558 7725 3594 7726
rect 3666 7725 3702 7726
rect 3558 7717 3702 7725
rect 3558 7697 3566 7717
rect 3586 7713 3674 7717
rect 3586 7697 3630 7713
rect 3558 7693 3630 7697
rect 3650 7697 3674 7713
rect 3694 7697 3702 7717
rect 3650 7693 3702 7697
rect 3558 7691 3702 7693
rect 3768 7721 3806 7729
rect 3884 7725 3920 7726
rect 3768 7701 3777 7721
rect 3797 7701 3806 7721
rect 3768 7692 3806 7701
rect 3835 7717 3920 7725
rect 3835 7697 3892 7717
rect 3912 7697 3920 7717
rect 3768 7691 3805 7692
rect 3835 7691 3920 7697
rect 3986 7721 4024 7729
rect 3986 7701 3995 7721
rect 4015 7701 4024 7721
rect 3986 7692 4024 7701
rect 4168 7726 4210 7735
rect 4168 7708 4182 7726
rect 4200 7708 4210 7726
rect 4168 7700 4210 7708
rect 4173 7698 4210 7700
rect 4600 7720 5043 7759
rect 3986 7691 4023 7692
rect 3447 7663 3537 7669
rect 3447 7643 3463 7663
rect 3483 7661 3537 7663
rect 3483 7643 3508 7661
rect 3447 7641 3508 7643
rect 3528 7641 3537 7661
rect 3447 7635 3537 7641
rect 3460 7581 3497 7582
rect 3556 7581 3593 7582
rect 3612 7581 3648 7691
rect 3835 7670 3866 7691
rect 4600 7677 4647 7720
rect 5003 7715 5043 7720
rect 5668 7718 5855 7742
rect 5886 7723 6279 7743
rect 6299 7723 6302 7743
rect 5886 7718 6302 7723
rect 3831 7669 3866 7670
rect 3709 7659 3866 7669
rect 3709 7639 3726 7659
rect 3746 7639 3866 7659
rect 3709 7632 3866 7639
rect 3933 7662 4082 7670
rect 3933 7642 3944 7662
rect 3964 7642 4003 7662
rect 4023 7642 4082 7662
rect 4600 7659 4610 7677
rect 4628 7659 4647 7677
rect 4600 7655 4647 7659
rect 4601 7650 4638 7655
rect 3933 7635 4082 7642
rect 5668 7647 5705 7718
rect 5886 7717 6227 7718
rect 5820 7657 5851 7658
rect 3933 7634 3974 7635
rect 4170 7633 4207 7636
rect 3667 7581 3704 7582
rect 3360 7572 3498 7581
rect 2564 7533 3008 7559
rect 2564 7531 2732 7533
rect 1517 7399 1964 7411
rect 1560 7397 1593 7399
rect 927 7379 1065 7388
rect 721 7378 758 7379
rect 451 7325 492 7326
rect 225 7304 277 7322
rect 343 7318 492 7325
rect 343 7298 402 7318
rect 422 7298 461 7318
rect 481 7298 492 7318
rect 343 7290 492 7298
rect 559 7321 716 7328
rect 559 7301 679 7321
rect 699 7301 716 7321
rect 559 7291 716 7301
rect 559 7290 594 7291
rect 559 7269 590 7290
rect 777 7269 813 7379
rect 832 7378 869 7379
rect 928 7378 965 7379
rect 888 7319 978 7325
rect 888 7299 897 7319
rect 917 7317 978 7319
rect 917 7299 942 7317
rect 888 7297 942 7299
rect 962 7297 978 7317
rect 888 7291 978 7297
rect 402 7268 439 7269
rect 401 7259 439 7268
rect 229 7241 269 7251
rect 229 7223 239 7241
rect 257 7223 269 7241
rect 401 7239 410 7259
rect 430 7239 439 7259
rect 401 7231 439 7239
rect 505 7263 590 7269
rect 620 7268 657 7269
rect 505 7243 513 7263
rect 533 7243 590 7263
rect 505 7235 590 7243
rect 619 7259 657 7268
rect 619 7239 628 7259
rect 648 7239 657 7259
rect 505 7234 541 7235
rect 619 7231 657 7239
rect 723 7263 867 7269
rect 723 7243 731 7263
rect 751 7243 784 7263
rect 804 7243 839 7263
rect 859 7243 867 7263
rect 723 7235 867 7243
rect 723 7234 759 7235
rect 831 7234 867 7235
rect 933 7268 970 7269
rect 933 7267 971 7268
rect 933 7259 997 7267
rect 933 7239 942 7259
rect 962 7245 997 7259
rect 1017 7245 1020 7265
rect 962 7240 1020 7245
rect 962 7239 997 7240
rect 229 7167 269 7223
rect 402 7202 439 7231
rect 403 7200 439 7202
rect 403 7178 594 7200
rect 620 7199 657 7231
rect 933 7227 997 7239
rect 1037 7201 1064 7379
rect 1922 7354 1964 7399
rect 896 7199 1064 7201
rect 620 7189 1064 7199
rect 1205 7295 1392 7319
rect 1423 7300 1816 7320
rect 1836 7300 1839 7320
rect 1423 7295 1839 7300
rect 1205 7224 1242 7295
rect 1423 7294 1764 7295
rect 1357 7234 1388 7235
rect 1205 7204 1214 7224
rect 1234 7204 1242 7224
rect 1205 7194 1242 7204
rect 1301 7224 1388 7234
rect 1301 7204 1310 7224
rect 1330 7204 1388 7224
rect 1301 7195 1388 7204
rect 1301 7194 1338 7195
rect 226 7162 269 7167
rect 617 7173 1064 7189
rect 617 7167 645 7173
rect 896 7172 1064 7173
rect 226 7159 376 7162
rect 617 7159 644 7167
rect 226 7157 644 7159
rect 226 7139 235 7157
rect 253 7139 644 7157
rect 1357 7144 1388 7195
rect 1423 7224 1460 7294
rect 1726 7293 1763 7294
rect 1575 7234 1611 7235
rect 1423 7204 1432 7224
rect 1452 7204 1460 7224
rect 1423 7194 1460 7204
rect 1519 7224 1667 7234
rect 1767 7231 1863 7233
rect 1519 7204 1528 7224
rect 1548 7204 1638 7224
rect 1658 7204 1667 7224
rect 1519 7195 1667 7204
rect 1725 7224 1863 7231
rect 1725 7204 1734 7224
rect 1754 7204 1863 7224
rect 1725 7195 1863 7204
rect 1519 7194 1556 7195
rect 1249 7141 1290 7142
rect 226 7136 644 7139
rect 226 7130 269 7136
rect 229 7127 269 7130
rect 1144 7134 1290 7141
rect 626 7118 666 7119
rect 337 7101 666 7118
rect 1144 7114 1200 7134
rect 1220 7114 1259 7134
rect 1279 7114 1290 7134
rect 1144 7106 1290 7114
rect 1357 7137 1514 7144
rect 1357 7117 1477 7137
rect 1497 7117 1514 7137
rect 1357 7107 1514 7117
rect 1357 7106 1392 7107
rect 221 7058 264 7069
rect 221 7040 233 7058
rect 251 7040 264 7058
rect 221 7014 264 7040
rect 337 7014 364 7101
rect 626 7092 666 7101
rect 221 6993 364 7014
rect 408 7066 442 7082
rect 626 7072 1019 7092
rect 1039 7072 1042 7092
rect 1357 7085 1388 7106
rect 1575 7085 1611 7195
rect 1630 7194 1667 7195
rect 1726 7194 1763 7195
rect 1686 7135 1776 7141
rect 1686 7115 1695 7135
rect 1715 7133 1776 7135
rect 1715 7115 1740 7133
rect 1686 7113 1740 7115
rect 1760 7113 1776 7133
rect 1686 7107 1776 7113
rect 1200 7084 1237 7085
rect 626 7067 1042 7072
rect 1199 7075 1237 7084
rect 626 7066 967 7067
rect 408 6996 445 7066
rect 560 7006 591 7007
rect 221 6991 358 6993
rect 221 6949 264 6991
rect 408 6976 417 6996
rect 437 6976 445 6996
rect 408 6966 445 6976
rect 504 6996 591 7006
rect 504 6976 513 6996
rect 533 6976 591 6996
rect 504 6967 591 6976
rect 504 6966 541 6967
rect 219 6939 264 6949
rect 219 6921 228 6939
rect 246 6921 264 6939
rect 219 6915 264 6921
rect 560 6916 591 6967
rect 626 6996 663 7066
rect 929 7065 966 7066
rect 1199 7055 1208 7075
rect 1228 7055 1237 7075
rect 1199 7047 1237 7055
rect 1303 7079 1388 7085
rect 1418 7084 1455 7085
rect 1303 7059 1311 7079
rect 1331 7059 1388 7079
rect 1303 7051 1388 7059
rect 1417 7075 1455 7084
rect 1417 7055 1426 7075
rect 1446 7055 1455 7075
rect 1303 7050 1339 7051
rect 1417 7047 1455 7055
rect 1521 7079 1665 7085
rect 1521 7059 1529 7079
rect 1549 7076 1637 7079
rect 1549 7059 1584 7076
rect 1521 7058 1584 7059
rect 1603 7059 1637 7076
rect 1657 7059 1665 7079
rect 1603 7058 1665 7059
rect 1521 7051 1665 7058
rect 1521 7050 1557 7051
rect 1629 7050 1665 7051
rect 1731 7084 1768 7085
rect 1731 7083 1769 7084
rect 1791 7083 1818 7087
rect 1731 7081 1818 7083
rect 1731 7075 1795 7081
rect 1731 7055 1740 7075
rect 1760 7061 1795 7075
rect 1815 7061 1818 7081
rect 1760 7056 1818 7061
rect 1760 7055 1795 7056
rect 1200 7018 1237 7047
rect 1201 7016 1237 7018
rect 778 7006 814 7007
rect 626 6976 635 6996
rect 655 6976 663 6996
rect 626 6966 663 6976
rect 722 6996 870 7006
rect 970 7003 1066 7005
rect 722 6976 731 6996
rect 751 6976 841 6996
rect 861 6976 870 6996
rect 722 6967 870 6976
rect 928 6996 1066 7003
rect 928 6976 937 6996
rect 957 6976 1066 6996
rect 1201 6994 1392 7016
rect 1418 7015 1455 7047
rect 1731 7043 1795 7055
rect 1835 7017 1862 7195
rect 1694 7015 1862 7017
rect 1418 6989 1862 7015
rect 928 6967 1066 6976
rect 722 6966 759 6967
rect 219 6912 256 6915
rect 452 6913 493 6914
rect 344 6906 493 6913
rect 344 6886 403 6906
rect 423 6886 462 6906
rect 482 6886 493 6906
rect 344 6878 493 6886
rect 560 6909 717 6916
rect 560 6889 680 6909
rect 700 6889 717 6909
rect 560 6879 717 6889
rect 560 6878 595 6879
rect 560 6857 591 6878
rect 778 6857 814 6967
rect 833 6966 870 6967
rect 929 6966 966 6967
rect 889 6907 979 6913
rect 889 6887 898 6907
rect 918 6905 979 6907
rect 918 6887 943 6905
rect 889 6885 943 6887
rect 963 6885 979 6905
rect 889 6879 979 6885
rect 403 6856 440 6857
rect 215 6848 253 6850
rect 215 6840 258 6848
rect 215 6822 226 6840
rect 244 6822 258 6840
rect 215 6795 258 6822
rect 402 6847 440 6856
rect 402 6827 411 6847
rect 431 6827 440 6847
rect 402 6819 440 6827
rect 506 6851 591 6857
rect 621 6856 658 6857
rect 506 6831 514 6851
rect 534 6831 591 6851
rect 506 6823 591 6831
rect 620 6847 658 6856
rect 620 6827 629 6847
rect 649 6827 658 6847
rect 506 6822 542 6823
rect 620 6819 658 6827
rect 724 6855 868 6857
rect 724 6851 776 6855
rect 724 6831 732 6851
rect 752 6835 776 6851
rect 796 6851 868 6855
rect 796 6835 840 6851
rect 752 6831 840 6835
rect 860 6831 868 6851
rect 724 6823 868 6831
rect 724 6822 760 6823
rect 832 6822 868 6823
rect 934 6856 971 6857
rect 934 6855 972 6856
rect 934 6847 998 6855
rect 934 6827 943 6847
rect 963 6833 998 6847
rect 1018 6833 1021 6853
rect 963 6828 1021 6833
rect 963 6827 998 6828
rect 216 6788 258 6795
rect 403 6788 440 6819
rect 621 6788 658 6819
rect 934 6815 998 6827
rect 1038 6789 1065 6967
rect 216 6748 261 6788
rect 403 6763 548 6788
rect 621 6787 701 6788
rect 897 6787 1065 6789
rect 621 6771 1065 6787
rect 405 6762 548 6763
rect 620 6761 1065 6771
rect 216 6727 263 6748
rect 620 6727 661 6761
rect 897 6760 1065 6761
rect 1528 6765 1568 6989
rect 1694 6988 1862 6989
rect 1926 7021 1959 7354
rect 2564 7353 2591 7531
rect 2631 7493 2695 7505
rect 2971 7501 3008 7533
rect 3034 7532 3225 7554
rect 3360 7552 3469 7572
rect 3489 7552 3498 7572
rect 3360 7545 3498 7552
rect 3556 7572 3704 7581
rect 3556 7552 3565 7572
rect 3585 7552 3675 7572
rect 3695 7552 3704 7572
rect 3360 7543 3456 7545
rect 3556 7542 3704 7552
rect 3763 7572 3800 7582
rect 3763 7552 3771 7572
rect 3791 7552 3800 7572
rect 3612 7541 3648 7542
rect 3189 7530 3225 7532
rect 3189 7501 3226 7530
rect 2631 7492 2666 7493
rect 2608 7487 2666 7492
rect 2608 7467 2611 7487
rect 2631 7473 2666 7487
rect 2686 7473 2695 7493
rect 2631 7465 2695 7473
rect 2657 7464 2695 7465
rect 2658 7463 2695 7464
rect 2761 7497 2797 7498
rect 2869 7497 2905 7498
rect 2761 7489 2905 7497
rect 2761 7469 2769 7489
rect 2789 7488 2877 7489
rect 2789 7469 2824 7488
rect 2845 7469 2877 7488
rect 2897 7469 2905 7489
rect 2761 7463 2905 7469
rect 2971 7493 3009 7501
rect 3087 7497 3123 7498
rect 2971 7473 2980 7493
rect 3000 7473 3009 7493
rect 2971 7464 3009 7473
rect 3038 7489 3123 7497
rect 3038 7469 3095 7489
rect 3115 7469 3123 7489
rect 2971 7463 3008 7464
rect 3038 7463 3123 7469
rect 3189 7493 3227 7501
rect 3189 7473 3198 7493
rect 3218 7473 3227 7493
rect 3460 7482 3497 7483
rect 3763 7482 3800 7552
rect 3835 7581 3866 7632
rect 4162 7627 4207 7633
rect 4162 7609 4180 7627
rect 4198 7609 4207 7627
rect 5668 7627 5677 7647
rect 5697 7627 5705 7647
rect 5668 7617 5705 7627
rect 5764 7647 5851 7657
rect 5764 7627 5773 7647
rect 5793 7627 5851 7647
rect 5764 7618 5851 7627
rect 5764 7617 5801 7618
rect 4162 7599 4207 7609
rect 3885 7581 3922 7582
rect 3835 7572 3922 7581
rect 3835 7552 3893 7572
rect 3913 7552 3922 7572
rect 3835 7542 3922 7552
rect 3981 7572 4018 7582
rect 3981 7552 3989 7572
rect 4009 7552 4018 7572
rect 4162 7557 4205 7599
rect 4589 7588 4641 7590
rect 4068 7555 4205 7557
rect 3835 7541 3866 7542
rect 3981 7482 4018 7552
rect 3459 7481 3800 7482
rect 3189 7464 3227 7473
rect 3384 7476 3800 7481
rect 3189 7463 3226 7464
rect 2650 7435 2740 7441
rect 2650 7415 2666 7435
rect 2686 7433 2740 7435
rect 2686 7415 2711 7433
rect 2650 7413 2711 7415
rect 2731 7413 2740 7433
rect 2650 7407 2740 7413
rect 2663 7353 2700 7354
rect 2759 7353 2796 7354
rect 2815 7353 2851 7463
rect 3038 7442 3069 7463
rect 3384 7456 3387 7476
rect 3407 7456 3800 7476
rect 3984 7466 4018 7482
rect 4062 7534 4205 7555
rect 4587 7584 5020 7588
rect 4587 7578 5026 7584
rect 4587 7560 4608 7578
rect 4626 7560 5026 7578
rect 5820 7567 5851 7618
rect 5886 7647 5923 7717
rect 6189 7716 6226 7717
rect 6038 7657 6074 7658
rect 5886 7627 5895 7647
rect 5915 7627 5923 7647
rect 5886 7617 5923 7627
rect 5982 7647 6130 7657
rect 6230 7654 6326 7656
rect 5982 7627 5991 7647
rect 6011 7627 6101 7647
rect 6121 7627 6130 7647
rect 5982 7618 6130 7627
rect 6188 7647 6326 7654
rect 6188 7627 6197 7647
rect 6217 7627 6326 7647
rect 6188 7618 6326 7627
rect 5982 7617 6019 7618
rect 5712 7564 5753 7565
rect 4587 7542 5026 7560
rect 3760 7447 3800 7456
rect 4062 7447 4089 7534
rect 4162 7508 4205 7534
rect 4162 7490 4175 7508
rect 4193 7490 4205 7508
rect 4162 7479 4205 7490
rect 3034 7441 3069 7442
rect 2912 7431 3069 7441
rect 2912 7411 2929 7431
rect 2949 7411 3069 7431
rect 2912 7404 3069 7411
rect 3136 7434 3285 7442
rect 3136 7414 3147 7434
rect 3167 7414 3206 7434
rect 3226 7414 3285 7434
rect 3760 7430 4089 7447
rect 3760 7429 3800 7430
rect 3136 7407 3285 7414
rect 4157 7418 4197 7421
rect 4157 7412 4200 7418
rect 3782 7409 4200 7412
rect 3136 7406 3177 7407
rect 2870 7353 2907 7354
rect 2563 7344 2701 7353
rect 2426 7334 2462 7340
rect 2426 7316 2431 7334
rect 2453 7316 2462 7334
rect 2426 7312 2462 7316
rect 2563 7324 2672 7344
rect 2692 7324 2701 7344
rect 2563 7317 2701 7324
rect 2759 7344 2907 7353
rect 2759 7324 2768 7344
rect 2788 7324 2878 7344
rect 2898 7324 2907 7344
rect 2563 7315 2659 7317
rect 2759 7314 2907 7324
rect 2966 7344 3003 7354
rect 2966 7324 2974 7344
rect 2994 7324 3003 7344
rect 2815 7313 2851 7314
rect 2429 7153 2462 7312
rect 2663 7254 2700 7255
rect 2966 7254 3003 7324
rect 3038 7353 3069 7404
rect 3782 7391 4173 7409
rect 4191 7391 4200 7409
rect 3782 7389 4200 7391
rect 3782 7381 3809 7389
rect 4050 7386 4200 7389
rect 3362 7375 3530 7376
rect 3781 7375 3809 7381
rect 3362 7359 3809 7375
rect 4157 7381 4200 7386
rect 3088 7353 3125 7354
rect 3038 7344 3125 7353
rect 3038 7324 3096 7344
rect 3116 7324 3125 7344
rect 3038 7314 3125 7324
rect 3184 7344 3221 7354
rect 3184 7324 3192 7344
rect 3212 7324 3221 7344
rect 3038 7313 3069 7314
rect 2662 7253 3003 7254
rect 3184 7253 3221 7324
rect 2587 7248 3003 7253
rect 2587 7228 2590 7248
rect 2610 7228 3003 7248
rect 3034 7229 3221 7253
rect 3362 7349 3806 7359
rect 3362 7347 3530 7349
rect 3362 7169 3389 7347
rect 3429 7309 3493 7321
rect 3769 7317 3806 7349
rect 3832 7348 4023 7370
rect 3987 7346 4023 7348
rect 3987 7317 4024 7346
rect 4157 7325 4197 7381
rect 3429 7308 3464 7309
rect 3406 7303 3464 7308
rect 3406 7283 3409 7303
rect 3429 7289 3464 7303
rect 3484 7289 3493 7309
rect 3429 7281 3493 7289
rect 3455 7280 3493 7281
rect 3456 7279 3493 7280
rect 3559 7313 3595 7314
rect 3667 7313 3703 7314
rect 3559 7305 3703 7313
rect 3559 7285 3567 7305
rect 3587 7285 3622 7305
rect 3642 7285 3675 7305
rect 3695 7285 3703 7305
rect 3559 7279 3703 7285
rect 3769 7309 3807 7317
rect 3885 7313 3921 7314
rect 3769 7289 3778 7309
rect 3798 7289 3807 7309
rect 3769 7280 3807 7289
rect 3836 7305 3921 7313
rect 3836 7285 3893 7305
rect 3913 7285 3921 7305
rect 3769 7279 3806 7280
rect 3836 7279 3921 7285
rect 3987 7309 4025 7317
rect 3987 7289 3996 7309
rect 4016 7289 4025 7309
rect 4157 7307 4169 7325
rect 4187 7307 4197 7325
rect 4589 7353 4641 7542
rect 4987 7517 5026 7542
rect 5604 7557 5753 7564
rect 5604 7537 5663 7557
rect 5683 7537 5722 7557
rect 5742 7537 5753 7557
rect 5604 7529 5753 7537
rect 5820 7560 5977 7567
rect 5820 7540 5940 7560
rect 5960 7540 5977 7560
rect 5820 7530 5977 7540
rect 5820 7529 5855 7530
rect 4771 7492 4958 7516
rect 4987 7497 5382 7517
rect 5402 7497 5405 7517
rect 5820 7508 5851 7529
rect 6038 7508 6074 7618
rect 6093 7617 6130 7618
rect 6189 7617 6226 7618
rect 6149 7558 6239 7564
rect 6149 7538 6158 7558
rect 6178 7556 6239 7558
rect 6178 7538 6203 7556
rect 6149 7536 6203 7538
rect 6223 7536 6239 7556
rect 6149 7530 6239 7536
rect 5663 7507 5700 7508
rect 4987 7492 5405 7497
rect 5662 7498 5700 7507
rect 4771 7421 4808 7492
rect 4987 7491 5330 7492
rect 4987 7488 5026 7491
rect 5292 7490 5329 7491
rect 4923 7431 4954 7432
rect 4771 7401 4780 7421
rect 4800 7401 4808 7421
rect 4771 7391 4808 7401
rect 4867 7421 4954 7431
rect 4867 7401 4876 7421
rect 4896 7401 4954 7421
rect 4867 7392 4954 7401
rect 4867 7391 4904 7392
rect 4589 7335 4605 7353
rect 4623 7335 4641 7353
rect 4923 7341 4954 7392
rect 4989 7421 5026 7488
rect 5662 7478 5671 7498
rect 5691 7478 5700 7498
rect 5662 7470 5700 7478
rect 5766 7502 5851 7508
rect 5881 7507 5918 7508
rect 5766 7482 5774 7502
rect 5794 7482 5851 7502
rect 5766 7474 5851 7482
rect 5880 7498 5918 7507
rect 5880 7478 5889 7498
rect 5909 7478 5918 7498
rect 5766 7473 5802 7474
rect 5880 7470 5918 7478
rect 5984 7503 6128 7508
rect 5984 7502 6046 7503
rect 5984 7482 5992 7502
rect 6012 7484 6046 7502
rect 6067 7502 6128 7503
rect 6067 7484 6100 7502
rect 6012 7482 6100 7484
rect 6120 7482 6128 7502
rect 5984 7474 6128 7482
rect 5984 7473 6020 7474
rect 6092 7473 6128 7474
rect 6194 7507 6231 7508
rect 6194 7506 6232 7507
rect 6194 7498 6258 7506
rect 6194 7478 6203 7498
rect 6223 7484 6258 7498
rect 6278 7484 6281 7504
rect 6223 7479 6281 7484
rect 6223 7478 6258 7479
rect 5663 7441 5700 7470
rect 5664 7439 5700 7441
rect 5141 7431 5177 7432
rect 4989 7401 4998 7421
rect 5018 7401 5026 7421
rect 4989 7391 5026 7401
rect 5085 7421 5233 7431
rect 5333 7428 5429 7430
rect 5085 7401 5094 7421
rect 5114 7401 5204 7421
rect 5224 7401 5233 7421
rect 5085 7392 5233 7401
rect 5291 7421 5429 7428
rect 5291 7401 5300 7421
rect 5320 7401 5429 7421
rect 5664 7417 5855 7439
rect 5881 7438 5918 7470
rect 6194 7466 6258 7478
rect 6298 7440 6325 7618
rect 6157 7438 6325 7440
rect 5881 7424 6325 7438
rect 6928 7572 7096 7573
rect 7222 7572 7262 7796
rect 7725 7800 7893 7801
rect 8128 7800 8168 7833
rect 8524 7800 8571 7833
rect 8975 7831 9016 7856
rect 9161 7831 9198 7862
rect 9379 7831 9416 7862
rect 9692 7858 9756 7870
rect 9796 7832 9823 8010
rect 8975 7804 9024 7831
rect 9160 7805 9209 7831
rect 9378 7830 9459 7831
rect 9655 7830 9823 7832
rect 9378 7805 9823 7830
rect 9379 7804 9823 7805
rect 7725 7799 8169 7800
rect 7725 7774 8170 7799
rect 7725 7772 7893 7774
rect 8089 7773 8170 7774
rect 8339 7773 8388 7799
rect 8524 7773 8573 7800
rect 7725 7594 7752 7772
rect 7792 7734 7856 7746
rect 8132 7742 8169 7773
rect 8350 7742 8387 7773
rect 8532 7748 8573 7773
rect 8977 7771 9024 7804
rect 9380 7771 9420 7804
rect 9655 7803 9823 7804
rect 10286 7808 10326 8032
rect 10452 8031 10620 8032
rect 11223 8166 11667 8180
rect 11223 8164 11391 8166
rect 11223 7986 11250 8164
rect 11290 8126 11354 8138
rect 11630 8134 11667 8166
rect 11693 8165 11884 8187
rect 12119 8183 12228 8203
rect 12248 8183 12257 8203
rect 12119 8176 12257 8183
rect 12315 8203 12463 8212
rect 12315 8183 12324 8203
rect 12344 8183 12434 8203
rect 12454 8183 12463 8203
rect 12119 8174 12215 8176
rect 12315 8173 12463 8183
rect 12522 8203 12559 8213
rect 12522 8183 12530 8203
rect 12550 8183 12559 8203
rect 12371 8172 12407 8173
rect 11848 8163 11884 8165
rect 11848 8134 11885 8163
rect 11290 8125 11325 8126
rect 11267 8120 11325 8125
rect 11267 8100 11270 8120
rect 11290 8106 11325 8120
rect 11345 8106 11354 8126
rect 11290 8098 11354 8106
rect 11316 8097 11354 8098
rect 11317 8096 11354 8097
rect 11420 8130 11456 8131
rect 11528 8130 11564 8131
rect 11420 8124 11564 8130
rect 11420 8122 11481 8124
rect 11420 8102 11428 8122
rect 11448 8107 11481 8122
rect 11500 8122 11564 8124
rect 11500 8107 11536 8122
rect 11448 8102 11536 8107
rect 11556 8102 11564 8122
rect 11420 8096 11564 8102
rect 11630 8126 11668 8134
rect 11746 8130 11782 8131
rect 11630 8106 11639 8126
rect 11659 8106 11668 8126
rect 11630 8097 11668 8106
rect 11697 8122 11782 8130
rect 11697 8102 11754 8122
rect 11774 8102 11782 8122
rect 11630 8096 11667 8097
rect 11697 8096 11782 8102
rect 11848 8126 11886 8134
rect 11848 8106 11857 8126
rect 11877 8106 11886 8126
rect 12522 8116 12559 8183
rect 12594 8212 12625 8263
rect 12907 8251 12925 8269
rect 12943 8251 12959 8269
rect 12644 8212 12681 8213
rect 12594 8203 12681 8212
rect 12594 8183 12652 8203
rect 12672 8183 12681 8203
rect 12594 8173 12681 8183
rect 12740 8203 12777 8213
rect 12740 8183 12748 8203
rect 12768 8183 12777 8203
rect 12594 8172 12625 8173
rect 12219 8113 12256 8114
rect 12522 8113 12561 8116
rect 12218 8112 12561 8113
rect 12740 8112 12777 8183
rect 11848 8097 11886 8106
rect 12143 8107 12561 8112
rect 11848 8096 11885 8097
rect 11309 8068 11399 8074
rect 11309 8048 11325 8068
rect 11345 8066 11399 8068
rect 11345 8048 11370 8066
rect 11309 8046 11370 8048
rect 11390 8046 11399 8066
rect 11309 8040 11399 8046
rect 11322 7986 11359 7987
rect 11418 7986 11455 7987
rect 11474 7986 11510 8096
rect 11697 8075 11728 8096
rect 12143 8087 12146 8107
rect 12166 8087 12561 8107
rect 12590 8088 12777 8112
rect 11693 8074 11728 8075
rect 11571 8064 11728 8074
rect 11571 8044 11588 8064
rect 11608 8044 11728 8064
rect 11571 8037 11728 8044
rect 11795 8067 11944 8075
rect 11795 8047 11806 8067
rect 11826 8047 11865 8067
rect 11885 8047 11944 8067
rect 11795 8040 11944 8047
rect 12522 8062 12561 8087
rect 12907 8062 12959 8251
rect 13351 8279 13361 8297
rect 13379 8279 13391 8297
rect 13523 8295 13532 8315
rect 13552 8295 13561 8315
rect 13523 8287 13561 8295
rect 13627 8319 13712 8325
rect 13742 8324 13779 8325
rect 13627 8299 13635 8319
rect 13655 8299 13712 8319
rect 13627 8291 13712 8299
rect 13741 8315 13779 8324
rect 13741 8295 13750 8315
rect 13770 8295 13779 8315
rect 13627 8290 13663 8291
rect 13741 8287 13779 8295
rect 13845 8319 13989 8325
rect 13845 8299 13853 8319
rect 13873 8299 13906 8319
rect 13926 8299 13961 8319
rect 13981 8299 13989 8319
rect 13845 8291 13989 8299
rect 13845 8290 13881 8291
rect 13953 8290 13989 8291
rect 14055 8324 14092 8325
rect 14055 8323 14093 8324
rect 14055 8315 14119 8323
rect 14055 8295 14064 8315
rect 14084 8301 14119 8315
rect 14139 8301 14142 8321
rect 14084 8296 14142 8301
rect 14084 8295 14119 8296
rect 13351 8223 13391 8279
rect 13524 8258 13561 8287
rect 13525 8256 13561 8258
rect 13525 8234 13716 8256
rect 13742 8255 13779 8287
rect 14055 8283 14119 8295
rect 14159 8257 14186 8435
rect 14018 8255 14186 8257
rect 13742 8245 14186 8255
rect 14327 8351 14514 8375
rect 14545 8356 14938 8376
rect 14958 8356 14961 8376
rect 14545 8351 14961 8356
rect 14327 8280 14364 8351
rect 14545 8350 14886 8351
rect 14479 8290 14510 8291
rect 14327 8260 14336 8280
rect 14356 8260 14364 8280
rect 14327 8250 14364 8260
rect 14423 8280 14510 8290
rect 14423 8260 14432 8280
rect 14452 8260 14510 8280
rect 14423 8251 14510 8260
rect 14423 8250 14460 8251
rect 13348 8218 13391 8223
rect 13739 8229 14186 8245
rect 13739 8223 13767 8229
rect 14018 8228 14186 8229
rect 13348 8215 13498 8218
rect 13739 8215 13766 8223
rect 13348 8213 13766 8215
rect 13348 8195 13357 8213
rect 13375 8195 13766 8213
rect 14479 8200 14510 8251
rect 14545 8280 14582 8350
rect 14848 8349 14885 8350
rect 14697 8290 14733 8291
rect 14545 8260 14554 8280
rect 14574 8260 14582 8280
rect 14545 8250 14582 8260
rect 14641 8280 14789 8290
rect 14889 8287 14985 8289
rect 14641 8260 14650 8280
rect 14670 8260 14760 8280
rect 14780 8260 14789 8280
rect 14641 8251 14789 8260
rect 14847 8280 14985 8287
rect 14847 8260 14856 8280
rect 14876 8260 14985 8280
rect 14847 8251 14985 8260
rect 14641 8250 14678 8251
rect 14371 8197 14412 8198
rect 13348 8192 13766 8195
rect 13348 8186 13391 8192
rect 13351 8183 13391 8186
rect 14263 8190 14412 8197
rect 13748 8174 13788 8175
rect 13459 8157 13788 8174
rect 14263 8170 14322 8190
rect 14342 8170 14381 8190
rect 14401 8170 14412 8190
rect 14263 8162 14412 8170
rect 14479 8193 14636 8200
rect 14479 8173 14599 8193
rect 14619 8173 14636 8193
rect 14479 8163 14636 8173
rect 14479 8162 14514 8163
rect 13343 8114 13386 8125
rect 13343 8096 13355 8114
rect 13373 8096 13386 8114
rect 13343 8070 13386 8096
rect 13459 8070 13486 8157
rect 13748 8148 13788 8157
rect 12522 8044 12961 8062
rect 11795 8039 11836 8040
rect 11529 7986 11566 7987
rect 11222 7977 11360 7986
rect 11222 7957 11331 7977
rect 11351 7957 11360 7977
rect 11222 7950 11360 7957
rect 11418 7977 11566 7986
rect 11418 7957 11427 7977
rect 11447 7957 11537 7977
rect 11557 7957 11566 7977
rect 11222 7948 11318 7950
rect 11418 7947 11566 7957
rect 11625 7977 11662 7987
rect 11625 7957 11633 7977
rect 11653 7957 11662 7977
rect 11474 7946 11510 7947
rect 11322 7887 11359 7888
rect 11625 7887 11662 7957
rect 11697 7986 11728 8037
rect 12522 8026 12922 8044
rect 12940 8026 12961 8044
rect 12522 8020 12961 8026
rect 12528 8016 12961 8020
rect 13343 8049 13486 8070
rect 13530 8122 13564 8138
rect 13748 8128 14141 8148
rect 14161 8128 14164 8148
rect 14479 8141 14510 8162
rect 14697 8141 14733 8251
rect 14752 8250 14789 8251
rect 14848 8250 14885 8251
rect 14808 8191 14898 8197
rect 14808 8171 14817 8191
rect 14837 8189 14898 8191
rect 14837 8171 14862 8189
rect 14808 8169 14862 8171
rect 14882 8169 14898 8189
rect 14808 8163 14898 8169
rect 14322 8140 14359 8141
rect 13748 8123 14164 8128
rect 14321 8131 14359 8140
rect 13748 8122 14089 8123
rect 13530 8052 13567 8122
rect 13682 8062 13713 8063
rect 13343 8047 13480 8049
rect 12907 8014 12959 8016
rect 13343 8005 13386 8047
rect 13530 8032 13539 8052
rect 13559 8032 13567 8052
rect 13530 8022 13567 8032
rect 13626 8052 13713 8062
rect 13626 8032 13635 8052
rect 13655 8032 13713 8052
rect 13626 8023 13713 8032
rect 13626 8022 13663 8023
rect 13341 7995 13386 8005
rect 11747 7986 11784 7987
rect 11697 7977 11784 7986
rect 11697 7957 11755 7977
rect 11775 7957 11784 7977
rect 11697 7947 11784 7957
rect 11843 7977 11880 7987
rect 11843 7957 11851 7977
rect 11871 7957 11880 7977
rect 13341 7977 13350 7995
rect 13368 7977 13386 7995
rect 13341 7971 13386 7977
rect 13682 7972 13713 8023
rect 13748 8052 13785 8122
rect 14051 8121 14088 8122
rect 14321 8111 14330 8131
rect 14350 8111 14359 8131
rect 14321 8103 14359 8111
rect 14425 8135 14510 8141
rect 14540 8140 14577 8141
rect 14425 8115 14433 8135
rect 14453 8115 14510 8135
rect 14425 8107 14510 8115
rect 14539 8131 14577 8140
rect 14539 8111 14548 8131
rect 14568 8111 14577 8131
rect 14425 8106 14461 8107
rect 14539 8103 14577 8111
rect 14643 8135 14787 8141
rect 14643 8115 14651 8135
rect 14671 8116 14703 8135
rect 14724 8116 14759 8135
rect 14671 8115 14759 8116
rect 14779 8115 14787 8135
rect 14643 8107 14787 8115
rect 14643 8106 14679 8107
rect 14751 8106 14787 8107
rect 14853 8140 14890 8141
rect 14853 8139 14891 8140
rect 14853 8131 14917 8139
rect 14853 8111 14862 8131
rect 14882 8117 14917 8131
rect 14937 8117 14940 8137
rect 14882 8112 14940 8117
rect 14882 8111 14917 8112
rect 14322 8074 14359 8103
rect 14323 8072 14359 8074
rect 13900 8062 13936 8063
rect 13748 8032 13757 8052
rect 13777 8032 13785 8052
rect 13748 8022 13785 8032
rect 13844 8052 13992 8062
rect 14092 8059 14188 8061
rect 13844 8032 13853 8052
rect 13873 8032 13963 8052
rect 13983 8032 13992 8052
rect 13844 8023 13992 8032
rect 14050 8052 14188 8059
rect 14050 8032 14059 8052
rect 14079 8032 14188 8052
rect 14323 8050 14514 8072
rect 14540 8071 14577 8103
rect 14853 8099 14917 8111
rect 14957 8073 14984 8251
rect 15589 8250 15622 8583
rect 15686 8615 15854 8616
rect 15980 8615 16020 8839
rect 16483 8843 16651 8844
rect 16483 8842 16927 8843
rect 17290 8842 17331 8843
rect 16483 8817 17331 8842
rect 16483 8815 16651 8817
rect 16847 8816 17331 8817
rect 16483 8637 16510 8815
rect 16550 8777 16614 8789
rect 16890 8785 16927 8816
rect 17108 8785 17145 8816
rect 17290 8791 17331 8816
rect 16550 8776 16585 8777
rect 16527 8771 16585 8776
rect 16527 8751 16530 8771
rect 16550 8757 16585 8771
rect 16605 8757 16614 8777
rect 16550 8749 16614 8757
rect 16576 8748 16614 8749
rect 16577 8747 16614 8748
rect 16680 8781 16716 8782
rect 16788 8781 16824 8782
rect 16680 8773 16824 8781
rect 16680 8753 16688 8773
rect 16708 8769 16796 8773
rect 16708 8753 16752 8769
rect 16680 8749 16752 8753
rect 16772 8753 16796 8769
rect 16816 8753 16824 8773
rect 16772 8749 16824 8753
rect 16680 8747 16824 8749
rect 16890 8777 16928 8785
rect 17006 8781 17042 8782
rect 16890 8757 16899 8777
rect 16919 8757 16928 8777
rect 16890 8748 16928 8757
rect 16957 8773 17042 8781
rect 16957 8753 17014 8773
rect 17034 8753 17042 8773
rect 16890 8747 16927 8748
rect 16957 8747 17042 8753
rect 17108 8777 17146 8785
rect 17108 8757 17117 8777
rect 17137 8757 17146 8777
rect 17108 8748 17146 8757
rect 17290 8782 17332 8791
rect 17290 8764 17304 8782
rect 17322 8764 17332 8782
rect 17290 8756 17332 8764
rect 17295 8754 17332 8756
rect 17108 8747 17145 8748
rect 16569 8719 16659 8725
rect 16569 8699 16585 8719
rect 16605 8717 16659 8719
rect 16605 8699 16630 8717
rect 16569 8697 16630 8699
rect 16650 8697 16659 8717
rect 16569 8691 16659 8697
rect 16582 8637 16619 8638
rect 16678 8637 16715 8638
rect 16734 8637 16770 8747
rect 16957 8726 16988 8747
rect 16953 8725 16988 8726
rect 16831 8715 16988 8725
rect 16831 8695 16848 8715
rect 16868 8695 16988 8715
rect 16831 8688 16988 8695
rect 17055 8718 17204 8726
rect 17055 8698 17066 8718
rect 17086 8698 17125 8718
rect 17145 8698 17204 8718
rect 17055 8691 17204 8698
rect 17055 8690 17096 8691
rect 17292 8689 17329 8692
rect 16789 8637 16826 8638
rect 16482 8628 16620 8637
rect 15686 8589 16130 8615
rect 15686 8587 15854 8589
rect 15686 8409 15713 8587
rect 15753 8549 15817 8561
rect 16093 8557 16130 8589
rect 16156 8588 16347 8610
rect 16482 8608 16591 8628
rect 16611 8608 16620 8628
rect 16482 8601 16620 8608
rect 16678 8628 16826 8637
rect 16678 8608 16687 8628
rect 16707 8608 16797 8628
rect 16817 8608 16826 8628
rect 16482 8599 16578 8601
rect 16678 8598 16826 8608
rect 16885 8628 16922 8638
rect 16885 8608 16893 8628
rect 16913 8608 16922 8628
rect 16734 8597 16770 8598
rect 16311 8586 16347 8588
rect 16311 8557 16348 8586
rect 15753 8548 15788 8549
rect 15730 8543 15788 8548
rect 15730 8523 15733 8543
rect 15753 8529 15788 8543
rect 15808 8529 15817 8549
rect 15753 8523 15817 8529
rect 15730 8521 15817 8523
rect 15730 8517 15757 8521
rect 15779 8520 15817 8521
rect 15780 8519 15817 8520
rect 15883 8553 15919 8554
rect 15991 8553 16027 8554
rect 15883 8546 16027 8553
rect 15883 8545 15945 8546
rect 15883 8525 15891 8545
rect 15911 8528 15945 8545
rect 15964 8545 16027 8546
rect 15964 8528 15999 8545
rect 15911 8525 15999 8528
rect 16019 8525 16027 8545
rect 15883 8519 16027 8525
rect 16093 8549 16131 8557
rect 16209 8553 16245 8554
rect 16093 8529 16102 8549
rect 16122 8529 16131 8549
rect 16093 8520 16131 8529
rect 16160 8545 16245 8553
rect 16160 8525 16217 8545
rect 16237 8525 16245 8545
rect 16093 8519 16130 8520
rect 16160 8519 16245 8525
rect 16311 8549 16349 8557
rect 16311 8529 16320 8549
rect 16340 8529 16349 8549
rect 16582 8538 16619 8539
rect 16885 8538 16922 8608
rect 16957 8637 16988 8688
rect 17284 8683 17329 8689
rect 17284 8665 17302 8683
rect 17320 8665 17329 8683
rect 17284 8655 17329 8665
rect 17007 8637 17044 8638
rect 16957 8628 17044 8637
rect 16957 8608 17015 8628
rect 17035 8608 17044 8628
rect 16957 8598 17044 8608
rect 17103 8628 17140 8638
rect 17103 8608 17111 8628
rect 17131 8608 17140 8628
rect 17284 8613 17327 8655
rect 17190 8611 17327 8613
rect 16957 8597 16988 8598
rect 17103 8538 17140 8608
rect 16581 8537 16922 8538
rect 16311 8520 16349 8529
rect 16506 8532 16922 8537
rect 16311 8519 16348 8520
rect 15772 8491 15862 8497
rect 15772 8471 15788 8491
rect 15808 8489 15862 8491
rect 15808 8471 15833 8489
rect 15772 8469 15833 8471
rect 15853 8469 15862 8489
rect 15772 8463 15862 8469
rect 15785 8409 15822 8410
rect 15881 8409 15918 8410
rect 15937 8409 15973 8519
rect 16160 8498 16191 8519
rect 16506 8512 16509 8532
rect 16529 8512 16922 8532
rect 17106 8522 17140 8538
rect 17184 8590 17327 8611
rect 16882 8503 16922 8512
rect 17184 8503 17211 8590
rect 17284 8564 17327 8590
rect 17284 8546 17297 8564
rect 17315 8546 17327 8564
rect 17284 8535 17327 8546
rect 16156 8497 16191 8498
rect 16034 8487 16191 8497
rect 16034 8467 16051 8487
rect 16071 8467 16191 8487
rect 16034 8460 16191 8467
rect 16258 8490 16404 8498
rect 16258 8470 16269 8490
rect 16289 8470 16328 8490
rect 16348 8470 16404 8490
rect 16882 8486 17211 8503
rect 16882 8485 16922 8486
rect 16258 8463 16404 8470
rect 17279 8474 17319 8477
rect 17279 8468 17322 8474
rect 16904 8465 17322 8468
rect 16258 8462 16299 8463
rect 15992 8409 16029 8410
rect 15685 8400 15823 8409
rect 15685 8380 15794 8400
rect 15814 8380 15823 8400
rect 15685 8373 15823 8380
rect 15881 8400 16029 8409
rect 15881 8380 15890 8400
rect 15910 8380 16000 8400
rect 16020 8380 16029 8400
rect 15685 8371 15781 8373
rect 15881 8370 16029 8380
rect 16088 8400 16125 8410
rect 16088 8380 16096 8400
rect 16116 8380 16125 8400
rect 15937 8369 15973 8370
rect 15785 8310 15822 8311
rect 16088 8310 16125 8380
rect 16160 8409 16191 8460
rect 16904 8447 17295 8465
rect 17313 8447 17322 8465
rect 16904 8445 17322 8447
rect 16904 8437 16931 8445
rect 17172 8442 17322 8445
rect 16484 8431 16652 8432
rect 16903 8431 16931 8437
rect 16484 8415 16931 8431
rect 17279 8437 17322 8442
rect 16210 8409 16247 8410
rect 16160 8400 16247 8409
rect 16160 8380 16218 8400
rect 16238 8380 16247 8400
rect 16160 8370 16247 8380
rect 16306 8400 16343 8410
rect 16306 8380 16314 8400
rect 16334 8380 16343 8400
rect 16160 8369 16191 8370
rect 15784 8309 16125 8310
rect 16306 8309 16343 8380
rect 15709 8304 16125 8309
rect 15709 8284 15712 8304
rect 15732 8284 16125 8304
rect 16156 8285 16343 8309
rect 16484 8405 16928 8415
rect 16484 8403 16652 8405
rect 15584 8205 15626 8250
rect 16484 8225 16511 8403
rect 16551 8365 16615 8377
rect 16891 8373 16928 8405
rect 16954 8404 17145 8426
rect 17109 8402 17145 8404
rect 17109 8373 17146 8402
rect 17279 8381 17319 8437
rect 16551 8364 16586 8365
rect 16528 8359 16586 8364
rect 16528 8339 16531 8359
rect 16551 8345 16586 8359
rect 16606 8345 16615 8365
rect 16551 8337 16615 8345
rect 16577 8336 16615 8337
rect 16578 8335 16615 8336
rect 16681 8369 16717 8370
rect 16789 8369 16825 8370
rect 16681 8361 16825 8369
rect 16681 8341 16689 8361
rect 16709 8341 16744 8361
rect 16764 8341 16797 8361
rect 16817 8341 16825 8361
rect 16681 8335 16825 8341
rect 16891 8365 16929 8373
rect 17007 8369 17043 8370
rect 16891 8345 16900 8365
rect 16920 8345 16929 8365
rect 16891 8336 16929 8345
rect 16958 8361 17043 8369
rect 16958 8341 17015 8361
rect 17035 8341 17043 8361
rect 16891 8335 16928 8336
rect 16958 8335 17043 8341
rect 17109 8365 17147 8373
rect 17109 8345 17118 8365
rect 17138 8345 17147 8365
rect 17279 8363 17291 8381
rect 17309 8363 17319 8381
rect 17279 8353 17319 8363
rect 17109 8336 17147 8345
rect 17109 8335 17146 8336
rect 16570 8307 16660 8313
rect 16570 8287 16586 8307
rect 16606 8305 16660 8307
rect 16606 8287 16631 8305
rect 16570 8285 16631 8287
rect 16651 8285 16660 8305
rect 16570 8279 16660 8285
rect 16583 8225 16620 8226
rect 16679 8225 16716 8226
rect 16735 8225 16771 8335
rect 16958 8314 16989 8335
rect 16954 8313 16989 8314
rect 16832 8303 16989 8313
rect 16832 8283 16849 8303
rect 16869 8283 16989 8303
rect 16832 8276 16989 8283
rect 17056 8306 17205 8314
rect 17056 8286 17067 8306
rect 17087 8286 17126 8306
rect 17146 8286 17205 8306
rect 17056 8279 17205 8286
rect 17271 8282 17323 8300
rect 17056 8278 17097 8279
rect 16790 8225 16827 8226
rect 16483 8216 16621 8225
rect 15955 8205 15988 8207
rect 15584 8193 16031 8205
rect 14816 8071 14984 8073
rect 14540 8045 14984 8071
rect 14050 8023 14188 8032
rect 13844 8022 13881 8023
rect 13341 7968 13378 7971
rect 13574 7969 13615 7970
rect 11697 7946 11728 7947
rect 11321 7886 11662 7887
rect 11843 7886 11880 7957
rect 13466 7962 13615 7969
rect 12910 7949 12947 7954
rect 12901 7945 12948 7949
rect 12901 7927 12920 7945
rect 12938 7927 12948 7945
rect 13466 7942 13525 7962
rect 13545 7942 13584 7962
rect 13604 7942 13615 7962
rect 13466 7934 13615 7942
rect 13682 7965 13839 7972
rect 13682 7945 13802 7965
rect 13822 7945 13839 7965
rect 13682 7935 13839 7945
rect 13682 7934 13717 7935
rect 11246 7881 11662 7886
rect 11246 7861 11249 7881
rect 11269 7861 11662 7881
rect 11693 7862 11880 7886
rect 12505 7884 12545 7889
rect 12901 7884 12948 7927
rect 13682 7913 13713 7934
rect 13900 7913 13936 8023
rect 13955 8022 13992 8023
rect 14051 8022 14088 8023
rect 14011 7963 14101 7969
rect 14011 7943 14020 7963
rect 14040 7961 14101 7963
rect 14040 7943 14065 7961
rect 14011 7941 14065 7943
rect 14085 7941 14101 7961
rect 14011 7935 14101 7941
rect 13525 7912 13562 7913
rect 12505 7845 12948 7884
rect 13338 7904 13375 7906
rect 13338 7896 13380 7904
rect 13338 7878 13348 7896
rect 13366 7878 13380 7896
rect 13338 7869 13380 7878
rect 13524 7903 13562 7912
rect 13524 7883 13533 7903
rect 13553 7883 13562 7903
rect 13524 7875 13562 7883
rect 13628 7907 13713 7913
rect 13743 7912 13780 7913
rect 13628 7887 13636 7907
rect 13656 7887 13713 7907
rect 13628 7879 13713 7887
rect 13742 7903 13780 7912
rect 13742 7883 13751 7903
rect 13771 7883 13780 7903
rect 13628 7878 13664 7879
rect 13742 7875 13780 7883
rect 13846 7911 13990 7913
rect 13846 7907 13898 7911
rect 13846 7887 13854 7907
rect 13874 7891 13898 7907
rect 13918 7907 13990 7911
rect 13918 7891 13962 7907
rect 13874 7887 13962 7891
rect 13982 7887 13990 7907
rect 13846 7879 13990 7887
rect 13846 7878 13882 7879
rect 13954 7878 13990 7879
rect 14056 7912 14093 7913
rect 14056 7911 14094 7912
rect 14056 7903 14120 7911
rect 14056 7883 14065 7903
rect 14085 7889 14120 7903
rect 14140 7889 14143 7909
rect 14085 7884 14143 7889
rect 14085 7883 14120 7884
rect 10286 7786 10294 7808
rect 10318 7786 10326 7808
rect 10286 7778 10326 7786
rect 11599 7830 11639 7838
rect 11599 7808 11607 7830
rect 11631 7808 11639 7830
rect 7792 7733 7827 7734
rect 7769 7728 7827 7733
rect 7769 7708 7772 7728
rect 7792 7714 7827 7728
rect 7847 7714 7856 7734
rect 7792 7706 7856 7714
rect 7818 7705 7856 7706
rect 7819 7704 7856 7705
rect 7922 7738 7958 7739
rect 8030 7738 8066 7739
rect 7922 7730 8066 7738
rect 7922 7710 7930 7730
rect 7950 7726 8038 7730
rect 7950 7710 7994 7726
rect 7922 7706 7994 7710
rect 8014 7710 8038 7726
rect 8058 7710 8066 7730
rect 8014 7706 8066 7710
rect 7922 7704 8066 7706
rect 8132 7734 8170 7742
rect 8248 7738 8284 7739
rect 8132 7714 8141 7734
rect 8161 7714 8170 7734
rect 8132 7705 8170 7714
rect 8199 7730 8284 7738
rect 8199 7710 8256 7730
rect 8276 7710 8284 7730
rect 8132 7704 8169 7705
rect 8199 7704 8284 7710
rect 8350 7734 8388 7742
rect 8350 7714 8359 7734
rect 8379 7714 8388 7734
rect 8350 7705 8388 7714
rect 8532 7739 8574 7748
rect 8532 7721 8546 7739
rect 8564 7721 8574 7739
rect 8532 7713 8574 7721
rect 8537 7711 8574 7713
rect 8977 7732 9420 7771
rect 8350 7704 8387 7705
rect 7811 7676 7901 7682
rect 7811 7656 7827 7676
rect 7847 7674 7901 7676
rect 7847 7656 7872 7674
rect 7811 7654 7872 7656
rect 7892 7654 7901 7674
rect 7811 7648 7901 7654
rect 7824 7594 7861 7595
rect 7920 7594 7957 7595
rect 7976 7594 8012 7704
rect 8199 7683 8230 7704
rect 8977 7689 9024 7732
rect 9380 7727 9420 7732
rect 10045 7730 10232 7754
rect 10263 7735 10656 7755
rect 10676 7735 10679 7755
rect 10263 7730 10679 7735
rect 8195 7682 8230 7683
rect 8073 7672 8230 7682
rect 8073 7652 8090 7672
rect 8110 7652 8230 7672
rect 8073 7645 8230 7652
rect 8297 7675 8446 7683
rect 8297 7655 8308 7675
rect 8328 7655 8367 7675
rect 8387 7655 8446 7675
rect 8977 7671 8987 7689
rect 9005 7671 9024 7689
rect 8977 7667 9024 7671
rect 8978 7662 9015 7667
rect 8297 7648 8446 7655
rect 10045 7659 10082 7730
rect 10263 7729 10604 7730
rect 10197 7669 10228 7670
rect 8297 7647 8338 7648
rect 8534 7646 8571 7649
rect 8031 7594 8068 7595
rect 7724 7585 7862 7594
rect 6928 7546 7372 7572
rect 6928 7544 7096 7546
rect 5881 7412 6328 7424
rect 5924 7410 5957 7412
rect 5291 7392 5429 7401
rect 5085 7391 5122 7392
rect 4815 7338 4856 7339
rect 4589 7317 4641 7335
rect 4707 7331 4856 7338
rect 4157 7297 4197 7307
rect 4707 7311 4766 7331
rect 4786 7311 4825 7331
rect 4845 7311 4856 7331
rect 4707 7303 4856 7311
rect 4923 7334 5080 7341
rect 4923 7314 5043 7334
rect 5063 7314 5080 7334
rect 4923 7304 5080 7314
rect 4923 7303 4958 7304
rect 3987 7280 4025 7289
rect 4923 7282 4954 7303
rect 5141 7282 5177 7392
rect 5196 7391 5233 7392
rect 5292 7391 5329 7392
rect 5252 7332 5342 7338
rect 5252 7312 5261 7332
rect 5281 7330 5342 7332
rect 5281 7312 5306 7330
rect 5252 7310 5306 7312
rect 5326 7310 5342 7330
rect 5252 7304 5342 7310
rect 4766 7281 4803 7282
rect 3987 7279 4024 7280
rect 3448 7251 3538 7257
rect 3448 7231 3464 7251
rect 3484 7249 3538 7251
rect 3484 7231 3509 7249
rect 3448 7229 3509 7231
rect 3529 7229 3538 7249
rect 3448 7223 3538 7229
rect 3461 7169 3498 7170
rect 3557 7169 3594 7170
rect 3613 7169 3649 7279
rect 3836 7258 3867 7279
rect 4765 7272 4803 7281
rect 3832 7257 3867 7258
rect 3710 7247 3867 7257
rect 3710 7227 3727 7247
rect 3747 7227 3867 7247
rect 3710 7220 3867 7227
rect 3934 7250 4083 7258
rect 3934 7230 3945 7250
rect 3965 7230 4004 7250
rect 4024 7230 4083 7250
rect 4593 7254 4633 7264
rect 3934 7223 4083 7230
rect 4149 7226 4201 7244
rect 3934 7222 3975 7223
rect 3668 7169 3705 7170
rect 3361 7160 3499 7169
rect 2428 7152 2465 7153
rect 2399 7151 2567 7152
rect 2693 7151 2733 7153
rect 2224 7142 2263 7148
rect 2224 7120 2232 7142
rect 2256 7120 2263 7142
rect 1926 7013 1963 7021
rect 1926 6994 1934 7013
rect 1955 6994 1963 7013
rect 1926 6988 1963 6994
rect 1528 6743 1536 6765
rect 1560 6743 1568 6765
rect 1528 6735 1568 6743
rect 216 6697 661 6727
rect 1699 6710 1764 6711
rect 216 6694 639 6697
rect 216 6646 263 6694
rect 216 6628 226 6646
rect 244 6628 263 6646
rect 216 6624 263 6628
rect 1350 6685 1537 6709
rect 1568 6690 1961 6710
rect 1981 6690 1984 6710
rect 1568 6685 1984 6690
rect 217 6619 254 6624
rect 1350 6614 1387 6685
rect 1568 6684 1909 6685
rect 1502 6624 1533 6625
rect 1350 6594 1359 6614
rect 1379 6594 1387 6614
rect 1350 6584 1387 6594
rect 1446 6614 1533 6624
rect 1446 6594 1455 6614
rect 1475 6594 1533 6614
rect 1446 6585 1533 6594
rect 1446 6584 1483 6585
rect 205 6557 257 6559
rect 203 6553 636 6557
rect 203 6547 642 6553
rect 203 6529 224 6547
rect 242 6529 642 6547
rect 1502 6534 1533 6585
rect 1568 6614 1605 6684
rect 1871 6683 1908 6684
rect 1720 6624 1756 6625
rect 1568 6594 1577 6614
rect 1597 6594 1605 6614
rect 1568 6584 1605 6594
rect 1664 6614 1812 6624
rect 1912 6621 2008 6623
rect 1664 6594 1673 6614
rect 1693 6594 1783 6614
rect 1803 6594 1812 6614
rect 1664 6585 1812 6594
rect 1870 6614 2008 6621
rect 1870 6594 1879 6614
rect 1899 6594 2008 6614
rect 1870 6585 2008 6594
rect 1664 6584 1701 6585
rect 1394 6531 1435 6532
rect 203 6511 642 6529
rect 205 6322 257 6511
rect 603 6486 642 6511
rect 1286 6524 1435 6531
rect 1286 6504 1345 6524
rect 1365 6504 1404 6524
rect 1424 6504 1435 6524
rect 1286 6496 1435 6504
rect 1502 6527 1659 6534
rect 1502 6507 1622 6527
rect 1642 6507 1659 6527
rect 1502 6497 1659 6507
rect 1502 6496 1537 6497
rect 387 6461 574 6485
rect 603 6466 998 6486
rect 1018 6466 1021 6486
rect 1502 6475 1533 6496
rect 1720 6475 1756 6585
rect 1775 6584 1812 6585
rect 1871 6584 1908 6585
rect 1831 6525 1921 6531
rect 1831 6505 1840 6525
rect 1860 6523 1921 6525
rect 1860 6505 1885 6523
rect 1831 6503 1885 6505
rect 1905 6503 1921 6523
rect 1831 6497 1921 6503
rect 1345 6474 1382 6475
rect 603 6461 1021 6466
rect 1344 6465 1382 6474
rect 387 6390 424 6461
rect 603 6460 946 6461
rect 603 6457 642 6460
rect 908 6459 945 6460
rect 539 6400 570 6401
rect 387 6370 396 6390
rect 416 6370 424 6390
rect 387 6360 424 6370
rect 483 6390 570 6400
rect 483 6370 492 6390
rect 512 6370 570 6390
rect 483 6361 570 6370
rect 483 6360 520 6361
rect 205 6304 221 6322
rect 239 6304 257 6322
rect 539 6310 570 6361
rect 605 6390 642 6457
rect 1344 6445 1353 6465
rect 1373 6445 1382 6465
rect 1344 6437 1382 6445
rect 1448 6469 1533 6475
rect 1563 6474 1600 6475
rect 1448 6449 1456 6469
rect 1476 6449 1533 6469
rect 1448 6441 1533 6449
rect 1562 6465 1600 6474
rect 1562 6445 1571 6465
rect 1591 6445 1600 6465
rect 1448 6440 1484 6441
rect 1562 6437 1600 6445
rect 1666 6469 1810 6475
rect 1666 6449 1674 6469
rect 1694 6468 1782 6469
rect 1694 6450 1729 6468
rect 1747 6450 1782 6468
rect 1694 6449 1782 6450
rect 1802 6449 1810 6469
rect 1666 6441 1810 6449
rect 1666 6440 1702 6441
rect 1774 6440 1810 6441
rect 1876 6474 1913 6475
rect 1876 6473 1914 6474
rect 1876 6465 1940 6473
rect 1876 6445 1885 6465
rect 1905 6451 1940 6465
rect 1960 6451 1963 6471
rect 1905 6446 1963 6451
rect 1905 6445 1940 6446
rect 1345 6408 1382 6437
rect 1346 6406 1382 6408
rect 757 6400 793 6401
rect 605 6370 614 6390
rect 634 6370 642 6390
rect 605 6360 642 6370
rect 701 6390 849 6400
rect 949 6397 1045 6399
rect 701 6370 710 6390
rect 730 6370 820 6390
rect 840 6370 849 6390
rect 701 6361 849 6370
rect 907 6390 1045 6397
rect 907 6370 916 6390
rect 936 6370 1045 6390
rect 1346 6384 1537 6406
rect 1563 6405 1600 6437
rect 1876 6433 1940 6445
rect 1980 6409 2007 6585
rect 1926 6407 2007 6409
rect 1839 6405 2007 6407
rect 1563 6379 2007 6405
rect 1673 6377 1713 6379
rect 1839 6378 2007 6379
rect 907 6361 1045 6370
rect 1948 6376 2007 6378
rect 701 6360 738 6361
rect 431 6307 472 6308
rect 205 6286 257 6304
rect 323 6300 472 6307
rect 323 6280 382 6300
rect 402 6280 441 6300
rect 461 6280 472 6300
rect 323 6272 472 6280
rect 539 6303 696 6310
rect 539 6283 659 6303
rect 679 6283 696 6303
rect 539 6273 696 6283
rect 539 6272 574 6273
rect 539 6251 570 6272
rect 757 6251 793 6361
rect 812 6360 849 6361
rect 908 6360 945 6361
rect 868 6301 958 6307
rect 868 6281 877 6301
rect 897 6299 958 6301
rect 897 6281 922 6299
rect 868 6279 922 6281
rect 942 6279 958 6299
rect 868 6273 958 6279
rect 382 6250 419 6251
rect 381 6241 419 6250
rect 209 6223 249 6233
rect 209 6205 219 6223
rect 237 6205 249 6223
rect 381 6221 390 6241
rect 410 6221 419 6241
rect 381 6213 419 6221
rect 485 6245 570 6251
rect 600 6250 637 6251
rect 485 6225 493 6245
rect 513 6225 570 6245
rect 485 6217 570 6225
rect 599 6241 637 6250
rect 599 6221 608 6241
rect 628 6221 637 6241
rect 485 6216 521 6217
rect 599 6213 637 6221
rect 703 6245 847 6251
rect 703 6225 711 6245
rect 731 6225 764 6245
rect 784 6225 819 6245
rect 839 6225 847 6245
rect 703 6217 847 6225
rect 703 6216 739 6217
rect 811 6216 847 6217
rect 913 6250 950 6251
rect 913 6249 951 6250
rect 913 6241 977 6249
rect 913 6221 922 6241
rect 942 6227 977 6241
rect 997 6227 1000 6247
rect 942 6222 1000 6227
rect 942 6221 977 6222
rect 209 6149 249 6205
rect 382 6184 419 6213
rect 383 6182 419 6184
rect 383 6160 574 6182
rect 600 6181 637 6213
rect 913 6209 977 6221
rect 1017 6183 1044 6361
rect 1948 6358 1977 6376
rect 876 6181 1044 6183
rect 600 6171 1044 6181
rect 1185 6277 1372 6301
rect 1403 6282 1796 6302
rect 1816 6282 1819 6302
rect 1403 6277 1819 6282
rect 1185 6206 1222 6277
rect 1403 6276 1744 6277
rect 1337 6216 1368 6217
rect 1185 6186 1194 6206
rect 1214 6186 1222 6206
rect 1185 6176 1222 6186
rect 1281 6206 1368 6216
rect 1281 6186 1290 6206
rect 1310 6186 1368 6206
rect 1281 6177 1368 6186
rect 1281 6176 1318 6177
rect 206 6144 249 6149
rect 597 6155 1044 6171
rect 597 6149 625 6155
rect 876 6154 1044 6155
rect 206 6141 356 6144
rect 597 6141 624 6149
rect 206 6139 624 6141
rect 206 6121 215 6139
rect 233 6121 624 6139
rect 1337 6126 1368 6177
rect 1403 6206 1440 6276
rect 1706 6275 1743 6276
rect 1555 6216 1591 6217
rect 1403 6186 1412 6206
rect 1432 6186 1440 6206
rect 1403 6176 1440 6186
rect 1499 6206 1647 6216
rect 1747 6213 1843 6215
rect 1499 6186 1508 6206
rect 1528 6186 1618 6206
rect 1638 6186 1647 6206
rect 1499 6177 1647 6186
rect 1705 6206 1843 6213
rect 1705 6186 1714 6206
rect 1734 6186 1843 6206
rect 1705 6177 1843 6186
rect 1499 6176 1536 6177
rect 1229 6123 1270 6124
rect 206 6118 624 6121
rect 206 6112 249 6118
rect 209 6109 249 6112
rect 1121 6116 1270 6123
rect 606 6100 646 6101
rect 317 6083 646 6100
rect 1121 6096 1180 6116
rect 1200 6096 1239 6116
rect 1259 6096 1270 6116
rect 1121 6088 1270 6096
rect 1337 6119 1494 6126
rect 1337 6099 1457 6119
rect 1477 6099 1494 6119
rect 1337 6089 1494 6099
rect 1337 6088 1372 6089
rect 201 6040 244 6051
rect 201 6022 213 6040
rect 231 6022 244 6040
rect 201 5996 244 6022
rect 317 5996 344 6083
rect 606 6074 646 6083
rect 201 5975 344 5996
rect 388 6048 422 6064
rect 606 6054 999 6074
rect 1019 6054 1022 6074
rect 1337 6067 1368 6088
rect 1555 6067 1591 6177
rect 1610 6176 1647 6177
rect 1706 6176 1743 6177
rect 1666 6117 1756 6123
rect 1666 6097 1675 6117
rect 1695 6115 1756 6117
rect 1695 6097 1720 6115
rect 1666 6095 1720 6097
rect 1740 6095 1756 6115
rect 1666 6089 1756 6095
rect 1180 6066 1217 6067
rect 606 6049 1022 6054
rect 1179 6057 1217 6066
rect 606 6048 947 6049
rect 388 5978 425 6048
rect 540 5988 571 5989
rect 201 5973 338 5975
rect 201 5931 244 5973
rect 388 5958 397 5978
rect 417 5958 425 5978
rect 388 5948 425 5958
rect 484 5978 571 5988
rect 484 5958 493 5978
rect 513 5958 571 5978
rect 484 5949 571 5958
rect 484 5948 521 5949
rect 199 5921 244 5931
rect 199 5903 208 5921
rect 226 5903 244 5921
rect 199 5897 244 5903
rect 540 5898 571 5949
rect 606 5978 643 6048
rect 909 6047 946 6048
rect 1179 6037 1188 6057
rect 1208 6037 1217 6057
rect 1179 6029 1217 6037
rect 1283 6061 1368 6067
rect 1398 6066 1435 6067
rect 1283 6041 1291 6061
rect 1311 6041 1368 6061
rect 1283 6033 1368 6041
rect 1397 6057 1435 6066
rect 1397 6037 1406 6057
rect 1426 6037 1435 6057
rect 1283 6032 1319 6033
rect 1397 6029 1435 6037
rect 1501 6061 1645 6067
rect 1501 6041 1509 6061
rect 1529 6042 1561 6061
rect 1582 6042 1617 6061
rect 1529 6041 1617 6042
rect 1637 6041 1645 6061
rect 1501 6033 1645 6041
rect 1501 6032 1537 6033
rect 1609 6032 1645 6033
rect 1711 6066 1748 6067
rect 1711 6065 1749 6066
rect 1711 6057 1775 6065
rect 1711 6037 1720 6057
rect 1740 6043 1775 6057
rect 1795 6043 1798 6063
rect 1740 6038 1798 6043
rect 1740 6037 1775 6038
rect 1180 6000 1217 6029
rect 1181 5998 1217 6000
rect 758 5988 794 5989
rect 606 5958 615 5978
rect 635 5958 643 5978
rect 606 5948 643 5958
rect 702 5978 850 5988
rect 950 5985 1046 5987
rect 702 5958 711 5978
rect 731 5958 821 5978
rect 841 5958 850 5978
rect 702 5949 850 5958
rect 908 5978 1046 5985
rect 908 5958 917 5978
rect 937 5958 1046 5978
rect 1181 5976 1372 5998
rect 1398 5997 1435 6029
rect 1711 6025 1775 6037
rect 1815 5999 1842 6177
rect 1674 5997 1842 5999
rect 1398 5971 1842 5997
rect 908 5949 1046 5958
rect 702 5948 739 5949
rect 199 5894 236 5897
rect 432 5895 473 5896
rect 324 5888 473 5895
rect 324 5868 383 5888
rect 403 5868 442 5888
rect 462 5868 473 5888
rect 324 5860 473 5868
rect 540 5891 697 5898
rect 540 5871 660 5891
rect 680 5871 697 5891
rect 540 5861 697 5871
rect 540 5860 575 5861
rect 540 5839 571 5860
rect 758 5839 794 5949
rect 813 5948 850 5949
rect 909 5948 946 5949
rect 869 5889 959 5895
rect 869 5869 878 5889
rect 898 5887 959 5889
rect 898 5869 923 5887
rect 869 5867 923 5869
rect 943 5867 959 5887
rect 869 5861 959 5867
rect 383 5838 420 5839
rect 196 5830 233 5832
rect 196 5822 238 5830
rect 196 5804 206 5822
rect 224 5804 238 5822
rect 196 5795 238 5804
rect 382 5829 420 5838
rect 382 5809 391 5829
rect 411 5809 420 5829
rect 382 5801 420 5809
rect 486 5833 571 5839
rect 601 5838 638 5839
rect 486 5813 494 5833
rect 514 5813 571 5833
rect 486 5805 571 5813
rect 600 5829 638 5838
rect 600 5809 609 5829
rect 629 5809 638 5829
rect 486 5804 522 5805
rect 600 5801 638 5809
rect 704 5837 848 5839
rect 704 5833 756 5837
rect 704 5813 712 5833
rect 732 5817 756 5833
rect 776 5833 848 5837
rect 776 5817 820 5833
rect 732 5813 820 5817
rect 840 5813 848 5833
rect 704 5805 848 5813
rect 704 5804 740 5805
rect 812 5804 848 5805
rect 914 5838 951 5839
rect 914 5837 952 5838
rect 914 5829 978 5837
rect 914 5809 923 5829
rect 943 5815 978 5829
rect 998 5815 1001 5835
rect 943 5810 1001 5815
rect 943 5809 978 5810
rect 197 5770 238 5795
rect 383 5770 420 5801
rect 601 5770 638 5801
rect 914 5797 978 5809
rect 1018 5771 1045 5949
rect 197 5743 246 5770
rect 382 5744 431 5770
rect 600 5769 681 5770
rect 877 5769 1045 5771
rect 600 5744 1045 5769
rect 601 5743 1045 5744
rect 199 5710 246 5743
rect 602 5710 642 5743
rect 877 5742 1045 5743
rect 1508 5747 1548 5971
rect 1674 5970 1842 5971
rect 1508 5725 1516 5747
rect 1540 5725 1548 5747
rect 1508 5717 1548 5725
rect 199 5671 642 5710
rect 199 5628 246 5671
rect 602 5666 642 5671
rect 1267 5669 1454 5693
rect 1485 5674 1878 5694
rect 1898 5674 1901 5694
rect 1485 5669 1901 5674
rect 199 5610 209 5628
rect 227 5610 246 5628
rect 199 5606 246 5610
rect 200 5601 237 5606
rect 1267 5598 1304 5669
rect 1485 5668 1826 5669
rect 1419 5608 1450 5609
rect 1267 5578 1276 5598
rect 1296 5578 1304 5598
rect 1267 5568 1304 5578
rect 1363 5598 1450 5608
rect 1363 5578 1372 5598
rect 1392 5578 1450 5598
rect 1363 5569 1450 5578
rect 1363 5568 1400 5569
rect 188 5539 240 5541
rect 186 5535 619 5539
rect 186 5529 625 5535
rect 186 5511 207 5529
rect 225 5511 625 5529
rect 1419 5518 1450 5569
rect 1485 5598 1522 5668
rect 1788 5667 1825 5668
rect 1637 5608 1673 5609
rect 1485 5578 1494 5598
rect 1514 5578 1522 5598
rect 1485 5568 1522 5578
rect 1581 5598 1729 5608
rect 1829 5605 1925 5607
rect 1581 5578 1590 5598
rect 1610 5578 1700 5598
rect 1720 5578 1729 5598
rect 1581 5569 1729 5578
rect 1787 5598 1925 5605
rect 1787 5578 1796 5598
rect 1816 5578 1925 5598
rect 1787 5569 1925 5578
rect 1581 5568 1618 5569
rect 1311 5515 1352 5516
rect 186 5493 625 5511
rect 188 5304 240 5493
rect 586 5468 625 5493
rect 1203 5508 1352 5515
rect 1203 5488 1262 5508
rect 1282 5488 1321 5508
rect 1341 5488 1352 5508
rect 1203 5480 1352 5488
rect 1419 5511 1576 5518
rect 1419 5491 1539 5511
rect 1559 5491 1576 5511
rect 1419 5481 1576 5491
rect 1419 5480 1454 5481
rect 370 5443 557 5467
rect 586 5448 981 5468
rect 1001 5448 1004 5468
rect 1419 5459 1450 5480
rect 1637 5459 1673 5569
rect 1692 5568 1729 5569
rect 1788 5568 1825 5569
rect 1748 5509 1838 5515
rect 1748 5489 1757 5509
rect 1777 5507 1838 5509
rect 1777 5489 1802 5507
rect 1748 5487 1802 5489
rect 1822 5487 1838 5507
rect 1748 5481 1838 5487
rect 1262 5458 1299 5459
rect 586 5443 1004 5448
rect 1261 5449 1299 5458
rect 370 5372 407 5443
rect 586 5442 929 5443
rect 586 5439 625 5442
rect 891 5441 928 5442
rect 522 5382 553 5383
rect 370 5352 379 5372
rect 399 5352 407 5372
rect 370 5342 407 5352
rect 466 5372 553 5382
rect 466 5352 475 5372
rect 495 5352 553 5372
rect 466 5343 553 5352
rect 466 5342 503 5343
rect 188 5286 204 5304
rect 222 5286 240 5304
rect 522 5292 553 5343
rect 588 5372 625 5439
rect 1261 5429 1270 5449
rect 1290 5429 1299 5449
rect 1261 5421 1299 5429
rect 1365 5453 1450 5459
rect 1480 5458 1517 5459
rect 1365 5433 1373 5453
rect 1393 5433 1450 5453
rect 1365 5425 1450 5433
rect 1479 5449 1517 5458
rect 1479 5429 1488 5449
rect 1508 5429 1517 5449
rect 1365 5424 1401 5425
rect 1479 5421 1517 5429
rect 1583 5453 1727 5459
rect 1583 5433 1591 5453
rect 1611 5448 1699 5453
rect 1611 5433 1647 5448
rect 1583 5431 1647 5433
rect 1666 5433 1699 5448
rect 1719 5433 1727 5453
rect 1666 5431 1727 5433
rect 1583 5425 1727 5431
rect 1583 5424 1619 5425
rect 1691 5424 1727 5425
rect 1793 5458 1830 5459
rect 1793 5457 1831 5458
rect 1793 5449 1857 5457
rect 1793 5429 1802 5449
rect 1822 5435 1857 5449
rect 1877 5435 1880 5455
rect 1822 5430 1880 5435
rect 1822 5429 1857 5430
rect 1262 5392 1299 5421
rect 1263 5390 1299 5392
rect 740 5382 776 5383
rect 588 5352 597 5372
rect 617 5352 625 5372
rect 588 5342 625 5352
rect 684 5372 832 5382
rect 932 5379 1028 5381
rect 684 5352 693 5372
rect 713 5352 803 5372
rect 823 5352 832 5372
rect 684 5343 832 5352
rect 890 5372 1028 5379
rect 890 5352 899 5372
rect 919 5352 1028 5372
rect 1263 5368 1454 5390
rect 1480 5389 1517 5421
rect 1793 5417 1857 5429
rect 1897 5391 1924 5569
rect 1756 5389 1924 5391
rect 1480 5375 1924 5389
rect 1948 5412 1976 6358
rect 1948 5382 1993 5412
rect 1480 5363 1927 5375
rect 1523 5361 1556 5363
rect 890 5343 1028 5352
rect 684 5342 721 5343
rect 414 5289 455 5290
rect 188 5268 240 5286
rect 306 5282 455 5289
rect 306 5262 365 5282
rect 385 5262 424 5282
rect 444 5262 455 5282
rect 306 5254 455 5262
rect 522 5285 679 5292
rect 522 5265 642 5285
rect 662 5265 679 5285
rect 522 5255 679 5265
rect 522 5254 557 5255
rect 522 5233 553 5254
rect 740 5233 776 5343
rect 795 5342 832 5343
rect 891 5342 928 5343
rect 851 5283 941 5289
rect 851 5263 860 5283
rect 880 5281 941 5283
rect 880 5263 905 5281
rect 851 5261 905 5263
rect 925 5261 941 5281
rect 851 5255 941 5261
rect 365 5232 402 5233
rect 364 5223 402 5232
rect 192 5205 232 5215
rect 192 5187 202 5205
rect 220 5187 232 5205
rect 364 5203 373 5223
rect 393 5203 402 5223
rect 364 5195 402 5203
rect 468 5227 553 5233
rect 583 5232 620 5233
rect 468 5207 476 5227
rect 496 5207 553 5227
rect 468 5199 553 5207
rect 582 5223 620 5232
rect 582 5203 591 5223
rect 611 5203 620 5223
rect 468 5198 504 5199
rect 582 5195 620 5203
rect 686 5227 830 5233
rect 686 5207 694 5227
rect 714 5207 747 5227
rect 767 5207 802 5227
rect 822 5207 830 5227
rect 686 5199 830 5207
rect 686 5198 722 5199
rect 794 5198 830 5199
rect 896 5232 933 5233
rect 896 5231 934 5232
rect 896 5223 960 5231
rect 896 5203 905 5223
rect 925 5209 960 5223
rect 980 5209 983 5229
rect 925 5204 983 5209
rect 925 5203 960 5204
rect 192 5131 232 5187
rect 365 5166 402 5195
rect 366 5164 402 5166
rect 366 5142 557 5164
rect 583 5163 620 5195
rect 896 5191 960 5203
rect 1000 5165 1027 5343
rect 1885 5318 1927 5363
rect 1948 5364 1959 5382
rect 1981 5364 1993 5382
rect 1948 5358 1993 5364
rect 1949 5357 1993 5358
rect 859 5163 1027 5165
rect 583 5153 1027 5163
rect 1168 5259 1355 5283
rect 1386 5264 1779 5284
rect 1799 5264 1802 5284
rect 1386 5259 1802 5264
rect 1168 5188 1205 5259
rect 1386 5258 1727 5259
rect 1320 5198 1351 5199
rect 1168 5168 1177 5188
rect 1197 5168 1205 5188
rect 1168 5158 1205 5168
rect 1264 5188 1351 5198
rect 1264 5168 1273 5188
rect 1293 5168 1351 5188
rect 1264 5159 1351 5168
rect 1264 5158 1301 5159
rect 189 5126 232 5131
rect 580 5137 1027 5153
rect 580 5131 608 5137
rect 859 5136 1027 5137
rect 189 5123 339 5126
rect 580 5123 607 5131
rect 189 5121 607 5123
rect 189 5103 198 5121
rect 216 5103 607 5121
rect 1320 5108 1351 5159
rect 1386 5188 1423 5258
rect 1689 5257 1726 5258
rect 1538 5198 1574 5199
rect 1386 5168 1395 5188
rect 1415 5168 1423 5188
rect 1386 5158 1423 5168
rect 1482 5188 1630 5198
rect 1730 5195 1826 5197
rect 1482 5168 1491 5188
rect 1511 5168 1601 5188
rect 1621 5168 1630 5188
rect 1482 5159 1630 5168
rect 1688 5188 1826 5195
rect 1688 5168 1697 5188
rect 1717 5168 1826 5188
rect 1688 5159 1826 5168
rect 1482 5158 1519 5159
rect 1212 5105 1253 5106
rect 189 5100 607 5103
rect 189 5094 232 5100
rect 192 5091 232 5094
rect 1107 5098 1253 5105
rect 589 5082 629 5083
rect 300 5065 629 5082
rect 1107 5078 1163 5098
rect 1183 5078 1222 5098
rect 1242 5078 1253 5098
rect 1107 5070 1253 5078
rect 1320 5101 1477 5108
rect 1320 5081 1440 5101
rect 1460 5081 1477 5101
rect 1320 5071 1477 5081
rect 1320 5070 1355 5071
rect 184 5022 227 5033
rect 184 5004 196 5022
rect 214 5004 227 5022
rect 184 4978 227 5004
rect 300 4978 327 5065
rect 589 5056 629 5065
rect 184 4957 327 4978
rect 371 5030 405 5046
rect 589 5036 982 5056
rect 1002 5036 1005 5056
rect 1320 5049 1351 5070
rect 1538 5049 1574 5159
rect 1593 5158 1630 5159
rect 1689 5158 1726 5159
rect 1649 5099 1739 5105
rect 1649 5079 1658 5099
rect 1678 5097 1739 5099
rect 1678 5079 1703 5097
rect 1649 5077 1703 5079
rect 1723 5077 1739 5097
rect 1649 5071 1739 5077
rect 1163 5048 1200 5049
rect 589 5031 1005 5036
rect 1162 5039 1200 5048
rect 589 5030 930 5031
rect 371 4960 408 5030
rect 523 4970 554 4971
rect 184 4955 321 4957
rect 184 4913 227 4955
rect 371 4940 380 4960
rect 400 4940 408 4960
rect 371 4930 408 4940
rect 467 4960 554 4970
rect 467 4940 476 4960
rect 496 4940 554 4960
rect 467 4931 554 4940
rect 467 4930 504 4931
rect 182 4903 227 4913
rect 182 4885 191 4903
rect 209 4885 227 4903
rect 182 4879 227 4885
rect 523 4880 554 4931
rect 589 4960 626 5030
rect 892 5029 929 5030
rect 1162 5019 1171 5039
rect 1191 5019 1200 5039
rect 1162 5011 1200 5019
rect 1266 5043 1351 5049
rect 1381 5048 1418 5049
rect 1266 5023 1274 5043
rect 1294 5023 1351 5043
rect 1266 5015 1351 5023
rect 1380 5039 1418 5048
rect 1380 5019 1389 5039
rect 1409 5019 1418 5039
rect 1266 5014 1302 5015
rect 1380 5011 1418 5019
rect 1484 5043 1628 5049
rect 1484 5023 1492 5043
rect 1512 5040 1600 5043
rect 1512 5023 1547 5040
rect 1484 5022 1547 5023
rect 1566 5023 1600 5040
rect 1620 5023 1628 5043
rect 1566 5022 1628 5023
rect 1484 5015 1628 5022
rect 1484 5014 1520 5015
rect 1592 5014 1628 5015
rect 1694 5048 1731 5049
rect 1694 5047 1732 5048
rect 1754 5047 1781 5051
rect 1694 5045 1781 5047
rect 1694 5039 1758 5045
rect 1694 5019 1703 5039
rect 1723 5025 1758 5039
rect 1778 5025 1781 5045
rect 1723 5020 1781 5025
rect 1723 5019 1758 5020
rect 1163 4982 1200 5011
rect 1164 4980 1200 4982
rect 741 4970 777 4971
rect 589 4940 598 4960
rect 618 4940 626 4960
rect 589 4930 626 4940
rect 685 4960 833 4970
rect 933 4967 1029 4969
rect 685 4940 694 4960
rect 714 4940 804 4960
rect 824 4940 833 4960
rect 685 4931 833 4940
rect 891 4960 1029 4967
rect 891 4940 900 4960
rect 920 4940 1029 4960
rect 1164 4958 1355 4980
rect 1381 4979 1418 5011
rect 1694 5007 1758 5019
rect 1798 4981 1825 5159
rect 1657 4979 1825 4981
rect 1381 4953 1825 4979
rect 891 4931 1029 4940
rect 685 4930 722 4931
rect 182 4876 219 4879
rect 415 4877 456 4878
rect 307 4870 456 4877
rect 307 4850 366 4870
rect 386 4850 425 4870
rect 445 4850 456 4870
rect 307 4842 456 4850
rect 523 4873 680 4880
rect 523 4853 643 4873
rect 663 4853 680 4873
rect 523 4843 680 4853
rect 523 4842 558 4843
rect 523 4821 554 4842
rect 741 4821 777 4931
rect 796 4930 833 4931
rect 892 4930 929 4931
rect 852 4871 942 4877
rect 852 4851 861 4871
rect 881 4869 942 4871
rect 881 4851 906 4869
rect 852 4849 906 4851
rect 926 4849 942 4869
rect 852 4843 942 4849
rect 366 4820 403 4821
rect 179 4812 216 4814
rect 179 4804 221 4812
rect 179 4786 189 4804
rect 207 4786 221 4804
rect 179 4777 221 4786
rect 365 4811 403 4820
rect 365 4791 374 4811
rect 394 4791 403 4811
rect 365 4783 403 4791
rect 469 4815 554 4821
rect 584 4820 621 4821
rect 469 4795 477 4815
rect 497 4795 554 4815
rect 469 4787 554 4795
rect 583 4811 621 4820
rect 583 4791 592 4811
rect 612 4791 621 4811
rect 469 4786 505 4787
rect 583 4783 621 4791
rect 687 4819 831 4821
rect 687 4815 739 4819
rect 687 4795 695 4815
rect 715 4799 739 4815
rect 759 4815 831 4819
rect 759 4799 803 4815
rect 715 4795 803 4799
rect 823 4795 831 4815
rect 687 4787 831 4795
rect 687 4786 723 4787
rect 795 4786 831 4787
rect 897 4820 934 4821
rect 897 4819 935 4820
rect 897 4811 961 4819
rect 897 4791 906 4811
rect 926 4797 961 4811
rect 981 4797 984 4817
rect 926 4792 984 4797
rect 926 4791 961 4792
rect 180 4752 221 4777
rect 366 4752 403 4783
rect 584 4752 621 4783
rect 897 4779 961 4791
rect 1001 4753 1028 4931
rect 180 4718 223 4752
rect 362 4726 429 4752
rect 584 4751 664 4752
rect 860 4751 1028 4753
rect 584 4725 1028 4751
rect 180 4707 227 4718
rect 584 4708 619 4725
rect 860 4724 1028 4725
rect 1491 4729 1531 4953
rect 1657 4952 1825 4953
rect 1889 4985 1922 5318
rect 2224 5305 2263 7120
rect 2399 7126 2843 7151
rect 2399 6945 2426 7126
rect 2568 7125 2843 7126
rect 2466 7085 2530 7097
rect 2806 7093 2843 7125
rect 2869 7124 3060 7146
rect 3361 7140 3470 7160
rect 3490 7140 3499 7160
rect 3361 7133 3499 7140
rect 3557 7160 3705 7169
rect 3557 7140 3566 7160
rect 3586 7140 3676 7160
rect 3696 7140 3705 7160
rect 3361 7131 3457 7133
rect 3557 7130 3705 7140
rect 3764 7160 3801 7170
rect 3764 7140 3772 7160
rect 3792 7140 3801 7160
rect 3613 7129 3649 7130
rect 3024 7122 3060 7124
rect 3024 7093 3061 7122
rect 2466 7084 2501 7085
rect 2443 7079 2501 7084
rect 2443 7059 2446 7079
rect 2466 7065 2501 7079
rect 2521 7065 2530 7085
rect 2466 7057 2530 7065
rect 2492 7056 2530 7057
rect 2493 7055 2530 7056
rect 2596 7089 2632 7090
rect 2704 7089 2740 7090
rect 2596 7081 2740 7089
rect 2596 7061 2604 7081
rect 2624 7079 2712 7081
rect 2624 7061 2657 7079
rect 2596 7057 2657 7061
rect 2680 7061 2712 7079
rect 2732 7061 2740 7081
rect 2680 7057 2740 7061
rect 2596 7055 2740 7057
rect 2806 7085 2844 7093
rect 2922 7089 2958 7090
rect 2806 7065 2815 7085
rect 2835 7065 2844 7085
rect 2806 7056 2844 7065
rect 2873 7081 2958 7089
rect 2873 7061 2930 7081
rect 2950 7061 2958 7081
rect 2806 7055 2843 7056
rect 2873 7055 2958 7061
rect 3024 7085 3062 7093
rect 3024 7065 3033 7085
rect 3053 7065 3062 7085
rect 3764 7073 3801 7140
rect 3836 7169 3867 7220
rect 4149 7208 4167 7226
rect 4185 7208 4201 7226
rect 3886 7169 3923 7170
rect 3836 7160 3923 7169
rect 3836 7140 3894 7160
rect 3914 7140 3923 7160
rect 3836 7130 3923 7140
rect 3982 7160 4019 7170
rect 3982 7140 3990 7160
rect 4010 7140 4019 7160
rect 3836 7129 3867 7130
rect 3461 7070 3498 7071
rect 3764 7070 3803 7073
rect 3460 7069 3803 7070
rect 3982 7069 4019 7140
rect 3024 7056 3062 7065
rect 3385 7064 3803 7069
rect 3024 7055 3061 7056
rect 2485 7027 2575 7033
rect 2485 7007 2501 7027
rect 2521 7025 2575 7027
rect 2521 7007 2546 7025
rect 2485 7005 2546 7007
rect 2566 7005 2575 7025
rect 2485 6999 2575 7005
rect 2498 6945 2535 6946
rect 2594 6945 2631 6946
rect 2650 6945 2686 7055
rect 2873 7034 2904 7055
rect 3385 7044 3388 7064
rect 3408 7044 3803 7064
rect 3832 7045 4019 7069
rect 2869 7033 2904 7034
rect 2747 7023 2904 7033
rect 2747 7003 2764 7023
rect 2784 7003 2904 7023
rect 2747 6996 2904 7003
rect 2971 7026 3120 7034
rect 2971 7006 2982 7026
rect 3002 7006 3041 7026
rect 3061 7006 3120 7026
rect 2971 6999 3120 7006
rect 3764 7019 3803 7044
rect 4149 7019 4201 7208
rect 4593 7236 4603 7254
rect 4621 7236 4633 7254
rect 4765 7252 4774 7272
rect 4794 7252 4803 7272
rect 4765 7244 4803 7252
rect 4869 7276 4954 7282
rect 4984 7281 5021 7282
rect 4869 7256 4877 7276
rect 4897 7256 4954 7276
rect 4869 7248 4954 7256
rect 4983 7272 5021 7281
rect 4983 7252 4992 7272
rect 5012 7252 5021 7272
rect 4869 7247 4905 7248
rect 4983 7244 5021 7252
rect 5087 7276 5231 7282
rect 5087 7256 5095 7276
rect 5115 7256 5148 7276
rect 5168 7256 5203 7276
rect 5223 7256 5231 7276
rect 5087 7248 5231 7256
rect 5087 7247 5123 7248
rect 5195 7247 5231 7248
rect 5297 7281 5334 7282
rect 5297 7280 5335 7281
rect 5297 7272 5361 7280
rect 5297 7252 5306 7272
rect 5326 7258 5361 7272
rect 5381 7258 5384 7278
rect 5326 7253 5384 7258
rect 5326 7252 5361 7253
rect 4593 7180 4633 7236
rect 4766 7215 4803 7244
rect 4767 7213 4803 7215
rect 4767 7191 4958 7213
rect 4984 7212 5021 7244
rect 5297 7240 5361 7252
rect 5401 7214 5428 7392
rect 6286 7367 6328 7412
rect 5260 7212 5428 7214
rect 4984 7202 5428 7212
rect 5569 7308 5756 7332
rect 5787 7313 6180 7333
rect 6200 7313 6203 7333
rect 5787 7308 6203 7313
rect 5569 7237 5606 7308
rect 5787 7307 6128 7308
rect 5721 7247 5752 7248
rect 5569 7217 5578 7237
rect 5598 7217 5606 7237
rect 5569 7207 5606 7217
rect 5665 7237 5752 7247
rect 5665 7217 5674 7237
rect 5694 7217 5752 7237
rect 5665 7208 5752 7217
rect 5665 7207 5702 7208
rect 4590 7175 4633 7180
rect 4981 7186 5428 7202
rect 4981 7180 5009 7186
rect 5260 7185 5428 7186
rect 4590 7172 4740 7175
rect 4981 7172 5008 7180
rect 4590 7170 5008 7172
rect 4590 7152 4599 7170
rect 4617 7152 5008 7170
rect 5721 7157 5752 7208
rect 5787 7237 5824 7307
rect 6090 7306 6127 7307
rect 5939 7247 5975 7248
rect 5787 7217 5796 7237
rect 5816 7217 5824 7237
rect 5787 7207 5824 7217
rect 5883 7237 6031 7247
rect 6131 7244 6227 7246
rect 5883 7217 5892 7237
rect 5912 7217 6002 7237
rect 6022 7217 6031 7237
rect 5883 7208 6031 7217
rect 6089 7237 6227 7244
rect 6089 7217 6098 7237
rect 6118 7217 6227 7237
rect 6089 7208 6227 7217
rect 5883 7207 5920 7208
rect 5613 7154 5654 7155
rect 4590 7149 5008 7152
rect 4590 7143 4633 7149
rect 4593 7140 4633 7143
rect 5508 7147 5654 7154
rect 4990 7131 5030 7132
rect 4701 7114 5030 7131
rect 5508 7127 5564 7147
rect 5584 7127 5623 7147
rect 5643 7127 5654 7147
rect 5508 7119 5654 7127
rect 5721 7150 5878 7157
rect 5721 7130 5841 7150
rect 5861 7130 5878 7150
rect 5721 7120 5878 7130
rect 5721 7119 5756 7120
rect 4585 7071 4628 7082
rect 4585 7053 4597 7071
rect 4615 7053 4628 7071
rect 4585 7027 4628 7053
rect 4701 7027 4728 7114
rect 4990 7105 5030 7114
rect 3764 7001 4203 7019
rect 2971 6998 3012 6999
rect 2705 6945 2742 6946
rect 2398 6936 2536 6945
rect 2398 6916 2507 6936
rect 2527 6916 2536 6936
rect 2398 6909 2536 6916
rect 2594 6936 2742 6945
rect 2594 6916 2603 6936
rect 2623 6916 2713 6936
rect 2733 6916 2742 6936
rect 2398 6907 2494 6909
rect 2594 6906 2742 6916
rect 2801 6936 2838 6946
rect 2801 6916 2809 6936
rect 2829 6916 2838 6936
rect 2650 6905 2686 6906
rect 2498 6846 2535 6847
rect 2801 6846 2838 6916
rect 2873 6945 2904 6996
rect 3764 6983 4164 7001
rect 4182 6983 4203 7001
rect 3764 6977 4203 6983
rect 3770 6973 4203 6977
rect 4585 7006 4728 7027
rect 4772 7079 4806 7095
rect 4990 7085 5383 7105
rect 5403 7085 5406 7105
rect 5721 7098 5752 7119
rect 5939 7098 5975 7208
rect 5994 7207 6031 7208
rect 6090 7207 6127 7208
rect 6050 7148 6140 7154
rect 6050 7128 6059 7148
rect 6079 7146 6140 7148
rect 6079 7128 6104 7146
rect 6050 7126 6104 7128
rect 6124 7126 6140 7146
rect 6050 7120 6140 7126
rect 5564 7097 5601 7098
rect 4990 7080 5406 7085
rect 5563 7088 5601 7097
rect 4990 7079 5331 7080
rect 4772 7009 4809 7079
rect 4924 7019 4955 7020
rect 4585 7004 4722 7006
rect 4149 6971 4201 6973
rect 4585 6962 4628 7004
rect 4772 6989 4781 7009
rect 4801 6989 4809 7009
rect 4772 6979 4809 6989
rect 4868 7009 4955 7019
rect 4868 6989 4877 7009
rect 4897 6989 4955 7009
rect 4868 6980 4955 6989
rect 4868 6979 4905 6980
rect 4583 6952 4628 6962
rect 2923 6945 2960 6946
rect 2873 6936 2960 6945
rect 2873 6916 2931 6936
rect 2951 6916 2960 6936
rect 2873 6906 2960 6916
rect 3019 6936 3056 6946
rect 3019 6916 3027 6936
rect 3047 6916 3056 6936
rect 4583 6934 4592 6952
rect 4610 6934 4628 6952
rect 4583 6928 4628 6934
rect 4924 6929 4955 6980
rect 4990 7009 5027 7079
rect 5293 7078 5330 7079
rect 5563 7068 5572 7088
rect 5592 7068 5601 7088
rect 5563 7060 5601 7068
rect 5667 7092 5752 7098
rect 5782 7097 5819 7098
rect 5667 7072 5675 7092
rect 5695 7072 5752 7092
rect 5667 7064 5752 7072
rect 5781 7088 5819 7097
rect 5781 7068 5790 7088
rect 5810 7068 5819 7088
rect 5667 7063 5703 7064
rect 5781 7060 5819 7068
rect 5885 7092 6029 7098
rect 5885 7072 5893 7092
rect 5913 7089 6001 7092
rect 5913 7072 5948 7089
rect 5885 7071 5948 7072
rect 5967 7072 6001 7089
rect 6021 7072 6029 7092
rect 5967 7071 6029 7072
rect 5885 7064 6029 7071
rect 5885 7063 5921 7064
rect 5993 7063 6029 7064
rect 6095 7097 6132 7098
rect 6095 7096 6133 7097
rect 6155 7096 6182 7100
rect 6095 7094 6182 7096
rect 6095 7088 6159 7094
rect 6095 7068 6104 7088
rect 6124 7074 6159 7088
rect 6179 7074 6182 7094
rect 6124 7069 6182 7074
rect 6124 7068 6159 7069
rect 5564 7031 5601 7060
rect 5565 7029 5601 7031
rect 5142 7019 5178 7020
rect 4990 6989 4999 7009
rect 5019 6989 5027 7009
rect 4990 6979 5027 6989
rect 5086 7009 5234 7019
rect 5334 7016 5430 7018
rect 5086 6989 5095 7009
rect 5115 6989 5205 7009
rect 5225 6989 5234 7009
rect 5086 6980 5234 6989
rect 5292 7009 5430 7016
rect 5292 6989 5301 7009
rect 5321 6989 5430 7009
rect 5565 7007 5756 7029
rect 5782 7028 5819 7060
rect 6095 7056 6159 7068
rect 6199 7030 6226 7208
rect 6058 7028 6226 7030
rect 5782 7002 6226 7028
rect 5292 6980 5430 6989
rect 5086 6979 5123 6980
rect 4583 6925 4620 6928
rect 4816 6926 4857 6927
rect 2873 6905 2904 6906
rect 2497 6845 2838 6846
rect 3019 6845 3056 6916
rect 4708 6919 4857 6926
rect 4152 6906 4189 6911
rect 2422 6840 2838 6845
rect 2422 6820 2425 6840
rect 2445 6820 2838 6840
rect 2869 6821 3056 6845
rect 4143 6902 4190 6906
rect 4143 6884 4162 6902
rect 4180 6884 4190 6902
rect 4708 6899 4767 6919
rect 4787 6899 4826 6919
rect 4846 6899 4857 6919
rect 4708 6891 4857 6899
rect 4924 6922 5081 6929
rect 4924 6902 5044 6922
rect 5064 6902 5081 6922
rect 4924 6892 5081 6902
rect 4924 6891 4959 6892
rect 4143 6836 4190 6884
rect 4924 6870 4955 6891
rect 5142 6870 5178 6980
rect 5197 6979 5234 6980
rect 5293 6979 5330 6980
rect 5253 6920 5343 6926
rect 5253 6900 5262 6920
rect 5282 6918 5343 6920
rect 5282 6900 5307 6918
rect 5253 6898 5307 6900
rect 5327 6898 5343 6918
rect 5253 6892 5343 6898
rect 4767 6869 4804 6870
rect 3767 6833 4190 6836
rect 2642 6819 2707 6820
rect 3745 6803 4190 6833
rect 4579 6861 4617 6863
rect 4579 6853 4622 6861
rect 4579 6835 4590 6853
rect 4608 6835 4622 6853
rect 4579 6808 4622 6835
rect 4766 6860 4804 6869
rect 4766 6840 4775 6860
rect 4795 6840 4804 6860
rect 4766 6832 4804 6840
rect 4870 6864 4955 6870
rect 4985 6869 5022 6870
rect 4870 6844 4878 6864
rect 4898 6844 4955 6864
rect 4870 6836 4955 6844
rect 4984 6860 5022 6869
rect 4984 6840 4993 6860
rect 5013 6840 5022 6860
rect 4870 6835 4906 6836
rect 4984 6832 5022 6840
rect 5088 6868 5232 6870
rect 5088 6864 5140 6868
rect 5088 6844 5096 6864
rect 5116 6848 5140 6864
rect 5160 6864 5232 6868
rect 5160 6848 5204 6864
rect 5116 6844 5204 6848
rect 5224 6844 5232 6864
rect 5088 6836 5232 6844
rect 5088 6835 5124 6836
rect 5196 6835 5232 6836
rect 5298 6869 5335 6870
rect 5298 6868 5336 6869
rect 5298 6860 5362 6868
rect 5298 6840 5307 6860
rect 5327 6846 5362 6860
rect 5382 6846 5385 6866
rect 5327 6841 5385 6846
rect 5327 6840 5362 6841
rect 2838 6787 2878 6795
rect 2838 6765 2846 6787
rect 2870 6765 2878 6787
rect 2443 6536 2480 6542
rect 2443 6517 2451 6536
rect 2472 6517 2480 6536
rect 2443 6509 2480 6517
rect 2447 6176 2480 6509
rect 2544 6541 2712 6542
rect 2838 6541 2878 6765
rect 3341 6769 3509 6770
rect 3745 6769 3786 6803
rect 4143 6782 4190 6803
rect 3341 6759 3786 6769
rect 3858 6767 4001 6768
rect 3341 6743 3785 6759
rect 3341 6741 3509 6743
rect 3705 6742 3785 6743
rect 3858 6742 4003 6767
rect 4145 6742 4190 6782
rect 3341 6563 3368 6741
rect 3408 6703 3472 6715
rect 3748 6711 3785 6742
rect 3966 6711 4003 6742
rect 4148 6735 4190 6742
rect 4580 6801 4622 6808
rect 4767 6801 4804 6832
rect 4985 6801 5022 6832
rect 5298 6828 5362 6840
rect 5402 6802 5429 6980
rect 4580 6761 4625 6801
rect 4767 6776 4912 6801
rect 4985 6800 5065 6801
rect 5261 6800 5429 6802
rect 4985 6784 5429 6800
rect 4769 6775 4912 6776
rect 4984 6774 5429 6784
rect 4580 6740 4627 6761
rect 4984 6740 5025 6774
rect 5261 6773 5429 6774
rect 5892 6778 5932 7002
rect 6058 7001 6226 7002
rect 6290 7034 6323 7367
rect 6928 7366 6955 7544
rect 6995 7506 7059 7518
rect 7335 7514 7372 7546
rect 7398 7545 7589 7567
rect 7724 7565 7833 7585
rect 7853 7565 7862 7585
rect 7724 7558 7862 7565
rect 7920 7585 8068 7594
rect 7920 7565 7929 7585
rect 7949 7565 8039 7585
rect 8059 7565 8068 7585
rect 7724 7556 7820 7558
rect 7920 7555 8068 7565
rect 8127 7585 8164 7595
rect 8127 7565 8135 7585
rect 8155 7565 8164 7585
rect 7976 7554 8012 7555
rect 7553 7543 7589 7545
rect 7553 7514 7590 7543
rect 6995 7505 7030 7506
rect 6972 7500 7030 7505
rect 6972 7480 6975 7500
rect 6995 7486 7030 7500
rect 7050 7486 7059 7506
rect 6995 7478 7059 7486
rect 7021 7477 7059 7478
rect 7022 7476 7059 7477
rect 7125 7510 7161 7511
rect 7233 7510 7269 7511
rect 7125 7502 7269 7510
rect 7125 7482 7133 7502
rect 7153 7501 7241 7502
rect 7153 7482 7188 7501
rect 7209 7482 7241 7501
rect 7261 7482 7269 7502
rect 7125 7476 7269 7482
rect 7335 7506 7373 7514
rect 7451 7510 7487 7511
rect 7335 7486 7344 7506
rect 7364 7486 7373 7506
rect 7335 7477 7373 7486
rect 7402 7502 7487 7510
rect 7402 7482 7459 7502
rect 7479 7482 7487 7502
rect 7335 7476 7372 7477
rect 7402 7476 7487 7482
rect 7553 7506 7591 7514
rect 7553 7486 7562 7506
rect 7582 7486 7591 7506
rect 7824 7495 7861 7496
rect 8127 7495 8164 7565
rect 8199 7594 8230 7645
rect 8526 7640 8571 7646
rect 8526 7622 8544 7640
rect 8562 7622 8571 7640
rect 10045 7639 10054 7659
rect 10074 7639 10082 7659
rect 10045 7629 10082 7639
rect 10141 7659 10228 7669
rect 10141 7639 10150 7659
rect 10170 7639 10228 7659
rect 10141 7630 10228 7639
rect 10141 7629 10178 7630
rect 8526 7612 8571 7622
rect 8249 7594 8286 7595
rect 8199 7585 8286 7594
rect 8199 7565 8257 7585
rect 8277 7565 8286 7585
rect 8199 7555 8286 7565
rect 8345 7585 8382 7595
rect 8345 7565 8353 7585
rect 8373 7565 8382 7585
rect 8526 7570 8569 7612
rect 8966 7600 9018 7602
rect 8432 7568 8569 7570
rect 8199 7554 8230 7555
rect 8345 7495 8382 7565
rect 7823 7494 8164 7495
rect 7553 7477 7591 7486
rect 7748 7489 8164 7494
rect 7553 7476 7590 7477
rect 7014 7448 7104 7454
rect 7014 7428 7030 7448
rect 7050 7446 7104 7448
rect 7050 7428 7075 7446
rect 7014 7426 7075 7428
rect 7095 7426 7104 7446
rect 7014 7420 7104 7426
rect 7027 7366 7064 7367
rect 7123 7366 7160 7367
rect 7179 7366 7215 7476
rect 7402 7455 7433 7476
rect 7748 7469 7751 7489
rect 7771 7469 8164 7489
rect 8348 7479 8382 7495
rect 8426 7547 8569 7568
rect 8964 7596 9397 7600
rect 8964 7590 9403 7596
rect 8964 7572 8985 7590
rect 9003 7572 9403 7590
rect 10197 7579 10228 7630
rect 10263 7659 10300 7729
rect 10566 7728 10603 7729
rect 10415 7669 10451 7670
rect 10263 7639 10272 7659
rect 10292 7639 10300 7659
rect 10263 7629 10300 7639
rect 10359 7659 10507 7669
rect 10607 7666 10703 7668
rect 10359 7639 10368 7659
rect 10388 7639 10478 7659
rect 10498 7639 10507 7659
rect 10359 7630 10507 7639
rect 10565 7659 10703 7666
rect 10565 7639 10574 7659
rect 10594 7639 10703 7659
rect 10565 7630 10703 7639
rect 10359 7629 10396 7630
rect 10089 7576 10130 7577
rect 8964 7554 9403 7572
rect 8124 7460 8164 7469
rect 8426 7460 8453 7547
rect 8526 7521 8569 7547
rect 8526 7503 8539 7521
rect 8557 7503 8569 7521
rect 8526 7492 8569 7503
rect 7398 7454 7433 7455
rect 7276 7444 7433 7454
rect 7276 7424 7293 7444
rect 7313 7424 7433 7444
rect 7276 7417 7433 7424
rect 7500 7447 7649 7455
rect 7500 7427 7511 7447
rect 7531 7427 7570 7447
rect 7590 7427 7649 7447
rect 8124 7443 8453 7460
rect 8124 7442 8164 7443
rect 7500 7420 7649 7427
rect 8521 7431 8561 7434
rect 8521 7425 8564 7431
rect 8146 7422 8564 7425
rect 7500 7419 7541 7420
rect 7234 7366 7271 7367
rect 6927 7357 7065 7366
rect 6790 7347 6826 7353
rect 6790 7329 6795 7347
rect 6817 7329 6826 7347
rect 6790 7325 6826 7329
rect 6927 7337 7036 7357
rect 7056 7337 7065 7357
rect 6927 7330 7065 7337
rect 7123 7357 7271 7366
rect 7123 7337 7132 7357
rect 7152 7337 7242 7357
rect 7262 7337 7271 7357
rect 6927 7328 7023 7330
rect 7123 7327 7271 7337
rect 7330 7357 7367 7367
rect 7330 7337 7338 7357
rect 7358 7337 7367 7357
rect 7179 7326 7215 7327
rect 6793 7166 6826 7325
rect 7027 7267 7064 7268
rect 7330 7267 7367 7337
rect 7402 7366 7433 7417
rect 8146 7404 8537 7422
rect 8555 7404 8564 7422
rect 8146 7402 8564 7404
rect 8146 7394 8173 7402
rect 8414 7399 8564 7402
rect 7726 7388 7894 7389
rect 8145 7388 8173 7394
rect 7726 7372 8173 7388
rect 8521 7394 8564 7399
rect 7452 7366 7489 7367
rect 7402 7357 7489 7366
rect 7402 7337 7460 7357
rect 7480 7337 7489 7357
rect 7402 7327 7489 7337
rect 7548 7357 7585 7367
rect 7548 7337 7556 7357
rect 7576 7337 7585 7357
rect 7402 7326 7433 7327
rect 7026 7266 7367 7267
rect 7548 7266 7585 7337
rect 6951 7261 7367 7266
rect 6951 7241 6954 7261
rect 6974 7241 7367 7261
rect 7398 7242 7585 7266
rect 7726 7362 8170 7372
rect 7726 7360 7894 7362
rect 7726 7182 7753 7360
rect 7793 7322 7857 7334
rect 8133 7330 8170 7362
rect 8196 7361 8387 7383
rect 8351 7359 8387 7361
rect 8351 7330 8388 7359
rect 8521 7338 8561 7394
rect 7793 7321 7828 7322
rect 7770 7316 7828 7321
rect 7770 7296 7773 7316
rect 7793 7302 7828 7316
rect 7848 7302 7857 7322
rect 7793 7294 7857 7302
rect 7819 7293 7857 7294
rect 7820 7292 7857 7293
rect 7923 7326 7959 7327
rect 8031 7326 8067 7327
rect 7923 7318 8067 7326
rect 7923 7298 7931 7318
rect 7951 7298 7986 7318
rect 8006 7298 8039 7318
rect 8059 7298 8067 7318
rect 7923 7292 8067 7298
rect 8133 7322 8171 7330
rect 8249 7326 8285 7327
rect 8133 7302 8142 7322
rect 8162 7302 8171 7322
rect 8133 7293 8171 7302
rect 8200 7318 8285 7326
rect 8200 7298 8257 7318
rect 8277 7298 8285 7318
rect 8133 7292 8170 7293
rect 8200 7292 8285 7298
rect 8351 7322 8389 7330
rect 8351 7302 8360 7322
rect 8380 7302 8389 7322
rect 8521 7320 8533 7338
rect 8551 7320 8561 7338
rect 8966 7365 9018 7554
rect 9364 7529 9403 7554
rect 9981 7569 10130 7576
rect 9981 7549 10040 7569
rect 10060 7549 10099 7569
rect 10119 7549 10130 7569
rect 9981 7541 10130 7549
rect 10197 7572 10354 7579
rect 10197 7552 10317 7572
rect 10337 7552 10354 7572
rect 10197 7542 10354 7552
rect 10197 7541 10232 7542
rect 9148 7504 9335 7528
rect 9364 7509 9759 7529
rect 9779 7509 9782 7529
rect 10197 7520 10228 7541
rect 10415 7520 10451 7630
rect 10470 7629 10507 7630
rect 10566 7629 10603 7630
rect 10526 7570 10616 7576
rect 10526 7550 10535 7570
rect 10555 7568 10616 7570
rect 10555 7550 10580 7568
rect 10526 7548 10580 7550
rect 10600 7548 10616 7568
rect 10526 7542 10616 7548
rect 10040 7519 10077 7520
rect 9364 7504 9782 7509
rect 10039 7510 10077 7519
rect 9148 7433 9185 7504
rect 9364 7503 9707 7504
rect 9364 7500 9403 7503
rect 9669 7502 9706 7503
rect 9300 7443 9331 7444
rect 9148 7413 9157 7433
rect 9177 7413 9185 7433
rect 9148 7403 9185 7413
rect 9244 7433 9331 7443
rect 9244 7413 9253 7433
rect 9273 7413 9331 7433
rect 9244 7404 9331 7413
rect 9244 7403 9281 7404
rect 8966 7347 8982 7365
rect 9000 7347 9018 7365
rect 9300 7353 9331 7404
rect 9366 7433 9403 7500
rect 10039 7490 10048 7510
rect 10068 7490 10077 7510
rect 10039 7482 10077 7490
rect 10143 7514 10228 7520
rect 10258 7519 10295 7520
rect 10143 7494 10151 7514
rect 10171 7494 10228 7514
rect 10143 7486 10228 7494
rect 10257 7510 10295 7519
rect 10257 7490 10266 7510
rect 10286 7490 10295 7510
rect 10143 7485 10179 7486
rect 10257 7482 10295 7490
rect 10361 7515 10505 7520
rect 10361 7514 10423 7515
rect 10361 7494 10369 7514
rect 10389 7496 10423 7514
rect 10444 7514 10505 7515
rect 10444 7496 10477 7514
rect 10389 7494 10477 7496
rect 10497 7494 10505 7514
rect 10361 7486 10505 7494
rect 10361 7485 10397 7486
rect 10469 7485 10505 7486
rect 10571 7519 10608 7520
rect 10571 7518 10609 7519
rect 10571 7510 10635 7518
rect 10571 7490 10580 7510
rect 10600 7496 10635 7510
rect 10655 7496 10658 7516
rect 10600 7491 10658 7496
rect 10600 7490 10635 7491
rect 10040 7453 10077 7482
rect 10041 7451 10077 7453
rect 9518 7443 9554 7444
rect 9366 7413 9375 7433
rect 9395 7413 9403 7433
rect 9366 7403 9403 7413
rect 9462 7433 9610 7443
rect 9710 7440 9806 7442
rect 9462 7413 9471 7433
rect 9491 7413 9581 7433
rect 9601 7413 9610 7433
rect 9462 7404 9610 7413
rect 9668 7433 9806 7440
rect 9668 7413 9677 7433
rect 9697 7413 9806 7433
rect 10041 7429 10232 7451
rect 10258 7450 10295 7482
rect 10571 7478 10635 7490
rect 10675 7452 10702 7630
rect 10534 7450 10702 7452
rect 10258 7436 10702 7450
rect 11305 7584 11473 7585
rect 11599 7584 11639 7808
rect 12102 7812 12270 7813
rect 12505 7812 12545 7845
rect 12901 7812 12948 7845
rect 13339 7844 13380 7869
rect 13525 7844 13562 7875
rect 13743 7844 13780 7875
rect 14056 7871 14120 7883
rect 14160 7845 14187 8023
rect 13339 7817 13388 7844
rect 13524 7818 13573 7844
rect 13742 7843 13823 7844
rect 14019 7843 14187 7845
rect 13742 7818 14187 7843
rect 13743 7817 14187 7818
rect 12102 7811 12546 7812
rect 12102 7786 12547 7811
rect 12102 7784 12270 7786
rect 12466 7785 12547 7786
rect 12716 7785 12765 7811
rect 12901 7785 12950 7812
rect 12102 7606 12129 7784
rect 12169 7746 12233 7758
rect 12509 7754 12546 7785
rect 12727 7754 12764 7785
rect 12909 7760 12950 7785
rect 13341 7784 13388 7817
rect 13744 7784 13784 7817
rect 14019 7816 14187 7817
rect 14650 7821 14690 8045
rect 14816 8044 14984 8045
rect 15587 8179 16031 8193
rect 15587 8177 15755 8179
rect 15587 7999 15614 8177
rect 15654 8139 15718 8151
rect 15994 8147 16031 8179
rect 16057 8178 16248 8200
rect 16483 8196 16592 8216
rect 16612 8196 16621 8216
rect 16483 8189 16621 8196
rect 16679 8216 16827 8225
rect 16679 8196 16688 8216
rect 16708 8196 16798 8216
rect 16818 8196 16827 8216
rect 16483 8187 16579 8189
rect 16679 8186 16827 8196
rect 16886 8216 16923 8226
rect 16886 8196 16894 8216
rect 16914 8196 16923 8216
rect 16735 8185 16771 8186
rect 16212 8176 16248 8178
rect 16212 8147 16249 8176
rect 15654 8138 15689 8139
rect 15631 8133 15689 8138
rect 15631 8113 15634 8133
rect 15654 8119 15689 8133
rect 15709 8119 15718 8139
rect 15654 8111 15718 8119
rect 15680 8110 15718 8111
rect 15681 8109 15718 8110
rect 15784 8143 15820 8144
rect 15892 8143 15928 8144
rect 15784 8137 15928 8143
rect 15784 8135 15845 8137
rect 15784 8115 15792 8135
rect 15812 8120 15845 8135
rect 15864 8135 15928 8137
rect 15864 8120 15900 8135
rect 15812 8115 15900 8120
rect 15920 8115 15928 8135
rect 15784 8109 15928 8115
rect 15994 8139 16032 8147
rect 16110 8143 16146 8144
rect 15994 8119 16003 8139
rect 16023 8119 16032 8139
rect 15994 8110 16032 8119
rect 16061 8135 16146 8143
rect 16061 8115 16118 8135
rect 16138 8115 16146 8135
rect 15994 8109 16031 8110
rect 16061 8109 16146 8115
rect 16212 8139 16250 8147
rect 16212 8119 16221 8139
rect 16241 8119 16250 8139
rect 16886 8129 16923 8196
rect 16958 8225 16989 8276
rect 17271 8264 17289 8282
rect 17307 8264 17323 8282
rect 17008 8225 17045 8226
rect 16958 8216 17045 8225
rect 16958 8196 17016 8216
rect 17036 8196 17045 8216
rect 16958 8186 17045 8196
rect 17104 8216 17141 8226
rect 17104 8196 17112 8216
rect 17132 8196 17141 8216
rect 16958 8185 16989 8186
rect 16583 8126 16620 8127
rect 16886 8126 16925 8129
rect 16582 8125 16925 8126
rect 17104 8125 17141 8196
rect 16212 8110 16250 8119
rect 16507 8120 16925 8125
rect 16212 8109 16249 8110
rect 15673 8081 15763 8087
rect 15673 8061 15689 8081
rect 15709 8079 15763 8081
rect 15709 8061 15734 8079
rect 15673 8059 15734 8061
rect 15754 8059 15763 8079
rect 15673 8053 15763 8059
rect 15686 7999 15723 8000
rect 15782 7999 15819 8000
rect 15838 7999 15874 8109
rect 16061 8088 16092 8109
rect 16507 8100 16510 8120
rect 16530 8100 16925 8120
rect 16954 8101 17141 8125
rect 16057 8087 16092 8088
rect 15935 8077 16092 8087
rect 15935 8057 15952 8077
rect 15972 8057 16092 8077
rect 15935 8050 16092 8057
rect 16159 8080 16308 8088
rect 16159 8060 16170 8080
rect 16190 8060 16229 8080
rect 16249 8060 16308 8080
rect 16159 8053 16308 8060
rect 16886 8075 16925 8100
rect 17271 8075 17323 8264
rect 16886 8057 17325 8075
rect 16159 8052 16200 8053
rect 15893 7999 15930 8000
rect 15586 7990 15724 7999
rect 15586 7970 15695 7990
rect 15715 7970 15724 7990
rect 15586 7963 15724 7970
rect 15782 7990 15930 7999
rect 15782 7970 15791 7990
rect 15811 7970 15901 7990
rect 15921 7970 15930 7990
rect 15586 7961 15682 7963
rect 15782 7960 15930 7970
rect 15989 7990 16026 8000
rect 15989 7970 15997 7990
rect 16017 7970 16026 7990
rect 15838 7959 15874 7960
rect 15686 7900 15723 7901
rect 15989 7900 16026 7970
rect 16061 7999 16092 8050
rect 16886 8039 17286 8057
rect 17304 8039 17325 8057
rect 16886 8033 17325 8039
rect 16892 8029 17325 8033
rect 17271 8027 17323 8029
rect 16111 7999 16148 8000
rect 16061 7990 16148 7999
rect 16061 7970 16119 7990
rect 16139 7970 16148 7990
rect 16061 7960 16148 7970
rect 16207 7990 16244 8000
rect 16207 7970 16215 7990
rect 16235 7970 16244 7990
rect 16061 7959 16092 7960
rect 15685 7899 16026 7900
rect 16207 7899 16244 7970
rect 17274 7962 17311 7967
rect 17265 7958 17312 7962
rect 17265 7940 17284 7958
rect 17302 7940 17312 7958
rect 15610 7894 16026 7899
rect 15610 7874 15613 7894
rect 15633 7874 16026 7894
rect 16057 7875 16244 7899
rect 16869 7897 16909 7902
rect 17265 7897 17312 7940
rect 16869 7858 17312 7897
rect 14650 7799 14658 7821
rect 14682 7799 14690 7821
rect 14650 7791 14690 7799
rect 15963 7843 16003 7851
rect 15963 7821 15971 7843
rect 15995 7821 16003 7843
rect 12169 7745 12204 7746
rect 12146 7740 12204 7745
rect 12146 7720 12149 7740
rect 12169 7726 12204 7740
rect 12224 7726 12233 7746
rect 12169 7718 12233 7726
rect 12195 7717 12233 7718
rect 12196 7716 12233 7717
rect 12299 7750 12335 7751
rect 12407 7750 12443 7751
rect 12299 7742 12443 7750
rect 12299 7722 12307 7742
rect 12327 7738 12415 7742
rect 12327 7722 12371 7738
rect 12299 7718 12371 7722
rect 12391 7722 12415 7738
rect 12435 7722 12443 7742
rect 12391 7718 12443 7722
rect 12299 7716 12443 7718
rect 12509 7746 12547 7754
rect 12625 7750 12661 7751
rect 12509 7726 12518 7746
rect 12538 7726 12547 7746
rect 12509 7717 12547 7726
rect 12576 7742 12661 7750
rect 12576 7722 12633 7742
rect 12653 7722 12661 7742
rect 12509 7716 12546 7717
rect 12576 7716 12661 7722
rect 12727 7746 12765 7754
rect 12727 7726 12736 7746
rect 12756 7726 12765 7746
rect 12727 7717 12765 7726
rect 12909 7751 12951 7760
rect 12909 7733 12923 7751
rect 12941 7733 12951 7751
rect 12909 7725 12951 7733
rect 12914 7723 12951 7725
rect 13341 7745 13784 7784
rect 12727 7716 12764 7717
rect 12188 7688 12278 7694
rect 12188 7668 12204 7688
rect 12224 7686 12278 7688
rect 12224 7668 12249 7686
rect 12188 7666 12249 7668
rect 12269 7666 12278 7686
rect 12188 7660 12278 7666
rect 12201 7606 12238 7607
rect 12297 7606 12334 7607
rect 12353 7606 12389 7716
rect 12576 7695 12607 7716
rect 13341 7702 13388 7745
rect 13744 7740 13784 7745
rect 14409 7743 14596 7767
rect 14627 7748 15020 7768
rect 15040 7748 15043 7768
rect 14627 7743 15043 7748
rect 12572 7694 12607 7695
rect 12450 7684 12607 7694
rect 12450 7664 12467 7684
rect 12487 7664 12607 7684
rect 12450 7657 12607 7664
rect 12674 7687 12823 7695
rect 12674 7667 12685 7687
rect 12705 7667 12744 7687
rect 12764 7667 12823 7687
rect 13341 7684 13351 7702
rect 13369 7684 13388 7702
rect 13341 7680 13388 7684
rect 13342 7675 13379 7680
rect 12674 7660 12823 7667
rect 14409 7672 14446 7743
rect 14627 7742 14968 7743
rect 14561 7682 14592 7683
rect 12674 7659 12715 7660
rect 12911 7658 12948 7661
rect 12408 7606 12445 7607
rect 12101 7597 12239 7606
rect 11305 7558 11749 7584
rect 11305 7556 11473 7558
rect 10258 7424 10705 7436
rect 10301 7422 10334 7424
rect 9668 7404 9806 7413
rect 9462 7403 9499 7404
rect 9192 7350 9233 7351
rect 8966 7329 9018 7347
rect 9084 7343 9233 7350
rect 8521 7310 8561 7320
rect 9084 7323 9143 7343
rect 9163 7323 9202 7343
rect 9222 7323 9233 7343
rect 9084 7315 9233 7323
rect 9300 7346 9457 7353
rect 9300 7326 9420 7346
rect 9440 7326 9457 7346
rect 9300 7316 9457 7326
rect 9300 7315 9335 7316
rect 8351 7293 8389 7302
rect 9300 7294 9331 7315
rect 9518 7294 9554 7404
rect 9573 7403 9610 7404
rect 9669 7403 9706 7404
rect 9629 7344 9719 7350
rect 9629 7324 9638 7344
rect 9658 7342 9719 7344
rect 9658 7324 9683 7342
rect 9629 7322 9683 7324
rect 9703 7322 9719 7342
rect 9629 7316 9719 7322
rect 9143 7293 9180 7294
rect 8351 7292 8388 7293
rect 7812 7264 7902 7270
rect 7812 7244 7828 7264
rect 7848 7262 7902 7264
rect 7848 7244 7873 7262
rect 7812 7242 7873 7244
rect 7893 7242 7902 7262
rect 7812 7236 7902 7242
rect 7825 7182 7862 7183
rect 7921 7182 7958 7183
rect 7977 7182 8013 7292
rect 8200 7271 8231 7292
rect 9142 7284 9180 7293
rect 8196 7270 8231 7271
rect 8074 7260 8231 7270
rect 8074 7240 8091 7260
rect 8111 7240 8231 7260
rect 8074 7233 8231 7240
rect 8298 7263 8447 7271
rect 8298 7243 8309 7263
rect 8329 7243 8368 7263
rect 8388 7243 8447 7263
rect 8970 7266 9010 7276
rect 8298 7236 8447 7243
rect 8513 7239 8565 7257
rect 8298 7235 8339 7236
rect 8032 7182 8069 7183
rect 7725 7173 7863 7182
rect 6792 7165 6829 7166
rect 6763 7164 6931 7165
rect 7057 7164 7097 7166
rect 6588 7155 6627 7161
rect 6588 7133 6596 7155
rect 6620 7133 6627 7155
rect 6290 7026 6327 7034
rect 6290 7007 6298 7026
rect 6319 7007 6327 7026
rect 6290 7001 6327 7007
rect 5892 6756 5900 6778
rect 5924 6756 5932 6778
rect 5892 6748 5932 6756
rect 3408 6702 3443 6703
rect 3385 6697 3443 6702
rect 3385 6677 3388 6697
rect 3408 6683 3443 6697
rect 3463 6683 3472 6703
rect 3408 6675 3472 6683
rect 3434 6674 3472 6675
rect 3435 6673 3472 6674
rect 3538 6707 3574 6708
rect 3646 6707 3682 6708
rect 3538 6699 3682 6707
rect 3538 6679 3546 6699
rect 3566 6695 3654 6699
rect 3566 6679 3610 6695
rect 3538 6675 3610 6679
rect 3630 6679 3654 6695
rect 3674 6679 3682 6699
rect 3630 6675 3682 6679
rect 3538 6673 3682 6675
rect 3748 6703 3786 6711
rect 3864 6707 3900 6708
rect 3748 6683 3757 6703
rect 3777 6683 3786 6703
rect 3748 6674 3786 6683
rect 3815 6699 3900 6707
rect 3815 6679 3872 6699
rect 3892 6679 3900 6699
rect 3748 6673 3785 6674
rect 3815 6673 3900 6679
rect 3966 6703 4004 6711
rect 3966 6683 3975 6703
rect 3995 6683 4004 6703
rect 3966 6674 4004 6683
rect 4148 6708 4191 6735
rect 4148 6690 4162 6708
rect 4180 6690 4191 6708
rect 4148 6682 4191 6690
rect 4153 6680 4191 6682
rect 4580 6710 5025 6740
rect 6063 6723 6128 6724
rect 4580 6707 5003 6710
rect 3966 6673 4003 6674
rect 3427 6645 3517 6651
rect 3427 6625 3443 6645
rect 3463 6643 3517 6645
rect 3463 6625 3488 6643
rect 3427 6623 3488 6625
rect 3508 6623 3517 6643
rect 3427 6617 3517 6623
rect 3440 6563 3477 6564
rect 3536 6563 3573 6564
rect 3592 6563 3628 6673
rect 3815 6652 3846 6673
rect 4580 6659 4627 6707
rect 3811 6651 3846 6652
rect 3689 6641 3846 6651
rect 3689 6621 3706 6641
rect 3726 6621 3846 6641
rect 3689 6614 3846 6621
rect 3913 6644 4062 6652
rect 3913 6624 3924 6644
rect 3944 6624 3983 6644
rect 4003 6624 4062 6644
rect 4580 6641 4590 6659
rect 4608 6641 4627 6659
rect 4580 6637 4627 6641
rect 5714 6698 5901 6722
rect 5932 6703 6325 6723
rect 6345 6703 6348 6723
rect 5932 6698 6348 6703
rect 4581 6632 4618 6637
rect 3913 6617 4062 6624
rect 5714 6627 5751 6698
rect 5932 6697 6273 6698
rect 5866 6637 5897 6638
rect 3913 6616 3954 6617
rect 4150 6615 4187 6618
rect 3647 6563 3684 6564
rect 3340 6554 3478 6563
rect 2544 6515 2988 6541
rect 2544 6513 2712 6515
rect 2544 6335 2571 6513
rect 2611 6475 2675 6487
rect 2951 6483 2988 6515
rect 3014 6514 3205 6536
rect 3340 6534 3449 6554
rect 3469 6534 3478 6554
rect 3340 6527 3478 6534
rect 3536 6554 3684 6563
rect 3536 6534 3545 6554
rect 3565 6534 3655 6554
rect 3675 6534 3684 6554
rect 3340 6525 3436 6527
rect 3536 6524 3684 6534
rect 3743 6554 3780 6564
rect 3743 6534 3751 6554
rect 3771 6534 3780 6554
rect 3592 6523 3628 6524
rect 3169 6512 3205 6514
rect 3169 6483 3206 6512
rect 2611 6474 2646 6475
rect 2588 6469 2646 6474
rect 2588 6449 2591 6469
rect 2611 6455 2646 6469
rect 2666 6455 2675 6475
rect 2611 6449 2675 6455
rect 2588 6447 2675 6449
rect 2588 6443 2615 6447
rect 2637 6446 2675 6447
rect 2638 6445 2675 6446
rect 2741 6479 2777 6480
rect 2849 6479 2885 6480
rect 2741 6472 2885 6479
rect 2741 6471 2803 6472
rect 2741 6451 2749 6471
rect 2769 6454 2803 6471
rect 2822 6471 2885 6472
rect 2822 6454 2857 6471
rect 2769 6451 2857 6454
rect 2877 6451 2885 6471
rect 2741 6445 2885 6451
rect 2951 6475 2989 6483
rect 3067 6479 3103 6480
rect 2951 6455 2960 6475
rect 2980 6455 2989 6475
rect 2951 6446 2989 6455
rect 3018 6471 3103 6479
rect 3018 6451 3075 6471
rect 3095 6451 3103 6471
rect 2951 6445 2988 6446
rect 3018 6445 3103 6451
rect 3169 6475 3207 6483
rect 3169 6455 3178 6475
rect 3198 6455 3207 6475
rect 3440 6464 3477 6465
rect 3743 6464 3780 6534
rect 3815 6563 3846 6614
rect 4142 6609 4187 6615
rect 4142 6591 4160 6609
rect 4178 6591 4187 6609
rect 5714 6607 5723 6627
rect 5743 6607 5751 6627
rect 5714 6597 5751 6607
rect 5810 6627 5897 6637
rect 5810 6607 5819 6627
rect 5839 6607 5897 6627
rect 5810 6598 5897 6607
rect 5810 6597 5847 6598
rect 4142 6581 4187 6591
rect 3865 6563 3902 6564
rect 3815 6554 3902 6563
rect 3815 6534 3873 6554
rect 3893 6534 3902 6554
rect 3815 6524 3902 6534
rect 3961 6554 3998 6564
rect 3961 6534 3969 6554
rect 3989 6534 3998 6554
rect 4142 6539 4185 6581
rect 4569 6570 4621 6572
rect 4048 6537 4185 6539
rect 3815 6523 3846 6524
rect 3961 6464 3998 6534
rect 3439 6463 3780 6464
rect 3169 6446 3207 6455
rect 3364 6458 3780 6463
rect 3169 6445 3206 6446
rect 2630 6417 2720 6423
rect 2630 6397 2646 6417
rect 2666 6415 2720 6417
rect 2666 6397 2691 6415
rect 2630 6395 2691 6397
rect 2711 6395 2720 6415
rect 2630 6389 2720 6395
rect 2643 6335 2680 6336
rect 2739 6335 2776 6336
rect 2795 6335 2831 6445
rect 3018 6424 3049 6445
rect 3364 6438 3367 6458
rect 3387 6438 3780 6458
rect 3964 6448 3998 6464
rect 4042 6516 4185 6537
rect 4567 6566 5000 6570
rect 4567 6560 5006 6566
rect 4567 6542 4588 6560
rect 4606 6542 5006 6560
rect 5866 6547 5897 6598
rect 5932 6627 5969 6697
rect 6235 6696 6272 6697
rect 6084 6637 6120 6638
rect 5932 6607 5941 6627
rect 5961 6607 5969 6627
rect 5932 6597 5969 6607
rect 6028 6627 6176 6637
rect 6276 6634 6372 6636
rect 6028 6607 6037 6627
rect 6057 6607 6147 6627
rect 6167 6607 6176 6627
rect 6028 6598 6176 6607
rect 6234 6627 6372 6634
rect 6234 6607 6243 6627
rect 6263 6607 6372 6627
rect 6234 6598 6372 6607
rect 6028 6597 6065 6598
rect 5758 6544 5799 6545
rect 4567 6524 5006 6542
rect 3740 6429 3780 6438
rect 4042 6429 4069 6516
rect 4142 6490 4185 6516
rect 4142 6472 4155 6490
rect 4173 6472 4185 6490
rect 4142 6461 4185 6472
rect 3014 6423 3049 6424
rect 2892 6413 3049 6423
rect 2892 6393 2909 6413
rect 2929 6393 3049 6413
rect 2892 6386 3049 6393
rect 3116 6416 3262 6424
rect 3116 6396 3127 6416
rect 3147 6396 3186 6416
rect 3206 6396 3262 6416
rect 3740 6412 4069 6429
rect 3740 6411 3780 6412
rect 3116 6389 3262 6396
rect 4137 6400 4177 6403
rect 4137 6394 4180 6400
rect 3762 6391 4180 6394
rect 3116 6388 3157 6389
rect 2850 6335 2887 6336
rect 2543 6326 2681 6335
rect 2543 6306 2652 6326
rect 2672 6306 2681 6326
rect 2543 6299 2681 6306
rect 2739 6326 2887 6335
rect 2739 6306 2748 6326
rect 2768 6306 2858 6326
rect 2878 6306 2887 6326
rect 2543 6297 2639 6299
rect 2739 6296 2887 6306
rect 2946 6326 2983 6336
rect 2946 6306 2954 6326
rect 2974 6306 2983 6326
rect 2795 6295 2831 6296
rect 2643 6236 2680 6237
rect 2946 6236 2983 6306
rect 3018 6335 3049 6386
rect 3762 6373 4153 6391
rect 4171 6373 4180 6391
rect 3762 6371 4180 6373
rect 3762 6363 3789 6371
rect 4030 6368 4180 6371
rect 3342 6357 3510 6358
rect 3761 6357 3789 6363
rect 3342 6341 3789 6357
rect 4137 6363 4180 6368
rect 3068 6335 3105 6336
rect 3018 6326 3105 6335
rect 3018 6306 3076 6326
rect 3096 6306 3105 6326
rect 3018 6296 3105 6306
rect 3164 6326 3201 6336
rect 3164 6306 3172 6326
rect 3192 6306 3201 6326
rect 3018 6295 3049 6296
rect 2642 6235 2983 6236
rect 3164 6235 3201 6306
rect 2567 6230 2983 6235
rect 2567 6210 2570 6230
rect 2590 6210 2983 6230
rect 3014 6211 3201 6235
rect 3342 6331 3786 6341
rect 3342 6329 3510 6331
rect 2442 6131 2484 6176
rect 3342 6151 3369 6329
rect 3409 6291 3473 6303
rect 3749 6299 3786 6331
rect 3812 6330 4003 6352
rect 3967 6328 4003 6330
rect 3967 6299 4004 6328
rect 4137 6307 4177 6363
rect 3409 6290 3444 6291
rect 3386 6285 3444 6290
rect 3386 6265 3389 6285
rect 3409 6271 3444 6285
rect 3464 6271 3473 6291
rect 3409 6263 3473 6271
rect 3435 6262 3473 6263
rect 3436 6261 3473 6262
rect 3539 6295 3575 6296
rect 3647 6295 3683 6296
rect 3539 6287 3683 6295
rect 3539 6267 3547 6287
rect 3567 6267 3602 6287
rect 3622 6267 3655 6287
rect 3675 6267 3683 6287
rect 3539 6261 3683 6267
rect 3749 6291 3787 6299
rect 3865 6295 3901 6296
rect 3749 6271 3758 6291
rect 3778 6271 3787 6291
rect 3749 6262 3787 6271
rect 3816 6287 3901 6295
rect 3816 6267 3873 6287
rect 3893 6267 3901 6287
rect 3749 6261 3786 6262
rect 3816 6261 3901 6267
rect 3967 6291 4005 6299
rect 3967 6271 3976 6291
rect 3996 6271 4005 6291
rect 4137 6289 4149 6307
rect 4167 6289 4177 6307
rect 4569 6335 4621 6524
rect 4967 6499 5006 6524
rect 5650 6537 5799 6544
rect 5650 6517 5709 6537
rect 5729 6517 5768 6537
rect 5788 6517 5799 6537
rect 5650 6509 5799 6517
rect 5866 6540 6023 6547
rect 5866 6520 5986 6540
rect 6006 6520 6023 6540
rect 5866 6510 6023 6520
rect 5866 6509 5901 6510
rect 4751 6474 4938 6498
rect 4967 6479 5362 6499
rect 5382 6479 5385 6499
rect 5866 6488 5897 6509
rect 6084 6488 6120 6598
rect 6139 6597 6176 6598
rect 6235 6597 6272 6598
rect 6195 6538 6285 6544
rect 6195 6518 6204 6538
rect 6224 6536 6285 6538
rect 6224 6518 6249 6536
rect 6195 6516 6249 6518
rect 6269 6516 6285 6536
rect 6195 6510 6285 6516
rect 5709 6487 5746 6488
rect 4967 6474 5385 6479
rect 5708 6478 5746 6487
rect 4751 6403 4788 6474
rect 4967 6473 5310 6474
rect 4967 6470 5006 6473
rect 5272 6472 5309 6473
rect 4903 6413 4934 6414
rect 4751 6383 4760 6403
rect 4780 6383 4788 6403
rect 4751 6373 4788 6383
rect 4847 6403 4934 6413
rect 4847 6383 4856 6403
rect 4876 6383 4934 6403
rect 4847 6374 4934 6383
rect 4847 6373 4884 6374
rect 4569 6317 4585 6335
rect 4603 6317 4621 6335
rect 4903 6323 4934 6374
rect 4969 6403 5006 6470
rect 5708 6458 5717 6478
rect 5737 6458 5746 6478
rect 5708 6450 5746 6458
rect 5812 6482 5897 6488
rect 5927 6487 5964 6488
rect 5812 6462 5820 6482
rect 5840 6462 5897 6482
rect 5812 6454 5897 6462
rect 5926 6478 5964 6487
rect 5926 6458 5935 6478
rect 5955 6458 5964 6478
rect 5812 6453 5848 6454
rect 5926 6450 5964 6458
rect 6030 6482 6174 6488
rect 6030 6462 6038 6482
rect 6058 6481 6146 6482
rect 6058 6463 6093 6481
rect 6111 6463 6146 6481
rect 6058 6462 6146 6463
rect 6166 6462 6174 6482
rect 6030 6454 6174 6462
rect 6030 6453 6066 6454
rect 6138 6453 6174 6454
rect 6240 6487 6277 6488
rect 6240 6486 6278 6487
rect 6240 6478 6304 6486
rect 6240 6458 6249 6478
rect 6269 6464 6304 6478
rect 6324 6464 6327 6484
rect 6269 6459 6327 6464
rect 6269 6458 6304 6459
rect 5709 6421 5746 6450
rect 5710 6419 5746 6421
rect 5121 6413 5157 6414
rect 4969 6383 4978 6403
rect 4998 6383 5006 6403
rect 4969 6373 5006 6383
rect 5065 6403 5213 6413
rect 5313 6410 5409 6412
rect 5065 6383 5074 6403
rect 5094 6383 5184 6403
rect 5204 6383 5213 6403
rect 5065 6374 5213 6383
rect 5271 6403 5409 6410
rect 5271 6383 5280 6403
rect 5300 6383 5409 6403
rect 5710 6397 5901 6419
rect 5927 6418 5964 6450
rect 6240 6446 6304 6458
rect 6344 6422 6371 6598
rect 6290 6420 6371 6422
rect 6203 6418 6371 6420
rect 5927 6392 6371 6418
rect 6037 6390 6077 6392
rect 6203 6391 6371 6392
rect 5271 6374 5409 6383
rect 6312 6389 6371 6391
rect 5065 6373 5102 6374
rect 4795 6320 4836 6321
rect 4569 6299 4621 6317
rect 4687 6313 4836 6320
rect 4137 6279 4177 6289
rect 4687 6293 4746 6313
rect 4766 6293 4805 6313
rect 4825 6293 4836 6313
rect 4687 6285 4836 6293
rect 4903 6316 5060 6323
rect 4903 6296 5023 6316
rect 5043 6296 5060 6316
rect 4903 6286 5060 6296
rect 4903 6285 4938 6286
rect 3967 6262 4005 6271
rect 4903 6264 4934 6285
rect 5121 6264 5157 6374
rect 5176 6373 5213 6374
rect 5272 6373 5309 6374
rect 5232 6314 5322 6320
rect 5232 6294 5241 6314
rect 5261 6312 5322 6314
rect 5261 6294 5286 6312
rect 5232 6292 5286 6294
rect 5306 6292 5322 6312
rect 5232 6286 5322 6292
rect 4746 6263 4783 6264
rect 3967 6261 4004 6262
rect 3428 6233 3518 6239
rect 3428 6213 3444 6233
rect 3464 6231 3518 6233
rect 3464 6213 3489 6231
rect 3428 6211 3489 6213
rect 3509 6211 3518 6231
rect 3428 6205 3518 6211
rect 3441 6151 3478 6152
rect 3537 6151 3574 6152
rect 3593 6151 3629 6261
rect 3816 6240 3847 6261
rect 4745 6254 4783 6263
rect 3812 6239 3847 6240
rect 3690 6229 3847 6239
rect 3690 6209 3707 6229
rect 3727 6209 3847 6229
rect 3690 6202 3847 6209
rect 3914 6232 4063 6240
rect 3914 6212 3925 6232
rect 3945 6212 3984 6232
rect 4004 6212 4063 6232
rect 4573 6236 4613 6246
rect 3914 6205 4063 6212
rect 4129 6208 4181 6226
rect 3914 6204 3955 6205
rect 3648 6151 3685 6152
rect 3341 6142 3479 6151
rect 2813 6131 2846 6133
rect 2442 6119 2889 6131
rect 2445 6105 2889 6119
rect 2445 6103 2613 6105
rect 2445 5925 2472 6103
rect 2512 6065 2576 6077
rect 2852 6073 2889 6105
rect 2915 6104 3106 6126
rect 3341 6122 3450 6142
rect 3470 6122 3479 6142
rect 3341 6115 3479 6122
rect 3537 6142 3685 6151
rect 3537 6122 3546 6142
rect 3566 6122 3656 6142
rect 3676 6122 3685 6142
rect 3341 6113 3437 6115
rect 3537 6112 3685 6122
rect 3744 6142 3781 6152
rect 3744 6122 3752 6142
rect 3772 6122 3781 6142
rect 3593 6111 3629 6112
rect 3070 6102 3106 6104
rect 3070 6073 3107 6102
rect 2512 6064 2547 6065
rect 2489 6059 2547 6064
rect 2489 6039 2492 6059
rect 2512 6045 2547 6059
rect 2567 6045 2576 6065
rect 2512 6037 2576 6045
rect 2538 6036 2576 6037
rect 2539 6035 2576 6036
rect 2642 6069 2678 6070
rect 2750 6069 2786 6070
rect 2642 6061 2786 6069
rect 2642 6041 2650 6061
rect 2670 6059 2758 6061
rect 2670 6041 2703 6059
rect 2642 6040 2703 6041
rect 2724 6041 2758 6059
rect 2778 6041 2786 6061
rect 2724 6040 2786 6041
rect 2642 6035 2786 6040
rect 2852 6065 2890 6073
rect 2968 6069 3004 6070
rect 2852 6045 2861 6065
rect 2881 6045 2890 6065
rect 2852 6036 2890 6045
rect 2919 6061 3004 6069
rect 2919 6041 2976 6061
rect 2996 6041 3004 6061
rect 2852 6035 2889 6036
rect 2919 6035 3004 6041
rect 3070 6065 3108 6073
rect 3070 6045 3079 6065
rect 3099 6045 3108 6065
rect 3744 6055 3781 6122
rect 3816 6151 3847 6202
rect 4129 6190 4147 6208
rect 4165 6190 4181 6208
rect 3866 6151 3903 6152
rect 3816 6142 3903 6151
rect 3816 6122 3874 6142
rect 3894 6122 3903 6142
rect 3816 6112 3903 6122
rect 3962 6142 3999 6152
rect 3962 6122 3970 6142
rect 3990 6122 3999 6142
rect 3816 6111 3847 6112
rect 3441 6052 3478 6053
rect 3744 6052 3783 6055
rect 3440 6051 3783 6052
rect 3962 6051 3999 6122
rect 3070 6036 3108 6045
rect 3365 6046 3783 6051
rect 3070 6035 3107 6036
rect 2531 6007 2621 6013
rect 2531 5987 2547 6007
rect 2567 6005 2621 6007
rect 2567 5987 2592 6005
rect 2531 5985 2592 5987
rect 2612 5985 2621 6005
rect 2531 5979 2621 5985
rect 2544 5925 2581 5926
rect 2640 5925 2677 5926
rect 2696 5925 2732 6035
rect 2919 6014 2950 6035
rect 3365 6026 3368 6046
rect 3388 6026 3783 6046
rect 3812 6027 3999 6051
rect 2915 6013 2950 6014
rect 2793 6003 2950 6013
rect 2793 5983 2810 6003
rect 2830 5983 2950 6003
rect 2793 5976 2950 5983
rect 3017 6006 3166 6014
rect 3017 5986 3028 6006
rect 3048 5986 3087 6006
rect 3107 5986 3166 6006
rect 3017 5979 3166 5986
rect 3744 6001 3783 6026
rect 4129 6001 4181 6190
rect 4573 6218 4583 6236
rect 4601 6218 4613 6236
rect 4745 6234 4754 6254
rect 4774 6234 4783 6254
rect 4745 6226 4783 6234
rect 4849 6258 4934 6264
rect 4964 6263 5001 6264
rect 4849 6238 4857 6258
rect 4877 6238 4934 6258
rect 4849 6230 4934 6238
rect 4963 6254 5001 6263
rect 4963 6234 4972 6254
rect 4992 6234 5001 6254
rect 4849 6229 4885 6230
rect 4963 6226 5001 6234
rect 5067 6258 5211 6264
rect 5067 6238 5075 6258
rect 5095 6238 5128 6258
rect 5148 6238 5183 6258
rect 5203 6238 5211 6258
rect 5067 6230 5211 6238
rect 5067 6229 5103 6230
rect 5175 6229 5211 6230
rect 5277 6263 5314 6264
rect 5277 6262 5315 6263
rect 5277 6254 5341 6262
rect 5277 6234 5286 6254
rect 5306 6240 5341 6254
rect 5361 6240 5364 6260
rect 5306 6235 5364 6240
rect 5306 6234 5341 6235
rect 4573 6162 4613 6218
rect 4746 6197 4783 6226
rect 4747 6195 4783 6197
rect 4747 6173 4938 6195
rect 4964 6194 5001 6226
rect 5277 6222 5341 6234
rect 5381 6196 5408 6374
rect 6312 6371 6341 6389
rect 5240 6194 5408 6196
rect 4964 6184 5408 6194
rect 5549 6290 5736 6314
rect 5767 6295 6160 6315
rect 6180 6295 6183 6315
rect 5767 6290 6183 6295
rect 5549 6219 5586 6290
rect 5767 6289 6108 6290
rect 5701 6229 5732 6230
rect 5549 6199 5558 6219
rect 5578 6199 5586 6219
rect 5549 6189 5586 6199
rect 5645 6219 5732 6229
rect 5645 6199 5654 6219
rect 5674 6199 5732 6219
rect 5645 6190 5732 6199
rect 5645 6189 5682 6190
rect 4570 6157 4613 6162
rect 4961 6168 5408 6184
rect 4961 6162 4989 6168
rect 5240 6167 5408 6168
rect 4570 6154 4720 6157
rect 4961 6154 4988 6162
rect 4570 6152 4988 6154
rect 4570 6134 4579 6152
rect 4597 6134 4988 6152
rect 5701 6139 5732 6190
rect 5767 6219 5804 6289
rect 6070 6288 6107 6289
rect 5919 6229 5955 6230
rect 5767 6199 5776 6219
rect 5796 6199 5804 6219
rect 5767 6189 5804 6199
rect 5863 6219 6011 6229
rect 6111 6226 6207 6228
rect 5863 6199 5872 6219
rect 5892 6199 5982 6219
rect 6002 6199 6011 6219
rect 5863 6190 6011 6199
rect 6069 6219 6207 6226
rect 6069 6199 6078 6219
rect 6098 6199 6207 6219
rect 6069 6190 6207 6199
rect 5863 6189 5900 6190
rect 5593 6136 5634 6137
rect 4570 6131 4988 6134
rect 4570 6125 4613 6131
rect 4573 6122 4613 6125
rect 5485 6129 5634 6136
rect 4970 6113 5010 6114
rect 4681 6096 5010 6113
rect 5485 6109 5544 6129
rect 5564 6109 5603 6129
rect 5623 6109 5634 6129
rect 5485 6101 5634 6109
rect 5701 6132 5858 6139
rect 5701 6112 5821 6132
rect 5841 6112 5858 6132
rect 5701 6102 5858 6112
rect 5701 6101 5736 6102
rect 4565 6053 4608 6064
rect 4565 6035 4577 6053
rect 4595 6035 4608 6053
rect 4565 6009 4608 6035
rect 4681 6009 4708 6096
rect 4970 6087 5010 6096
rect 3744 5983 4183 6001
rect 3017 5978 3058 5979
rect 2751 5925 2788 5926
rect 2444 5916 2582 5925
rect 2444 5896 2553 5916
rect 2573 5896 2582 5916
rect 2444 5889 2582 5896
rect 2640 5916 2788 5925
rect 2640 5896 2649 5916
rect 2669 5896 2759 5916
rect 2779 5896 2788 5916
rect 2444 5887 2540 5889
rect 2640 5886 2788 5896
rect 2847 5916 2884 5926
rect 2847 5896 2855 5916
rect 2875 5896 2884 5916
rect 2696 5885 2732 5886
rect 2544 5826 2581 5827
rect 2847 5826 2884 5896
rect 2919 5925 2950 5976
rect 3744 5965 4144 5983
rect 4162 5965 4183 5983
rect 3744 5959 4183 5965
rect 3750 5955 4183 5959
rect 4565 5988 4708 6009
rect 4752 6061 4786 6077
rect 4970 6067 5363 6087
rect 5383 6067 5386 6087
rect 5701 6080 5732 6101
rect 5919 6080 5955 6190
rect 5974 6189 6011 6190
rect 6070 6189 6107 6190
rect 6030 6130 6120 6136
rect 6030 6110 6039 6130
rect 6059 6128 6120 6130
rect 6059 6110 6084 6128
rect 6030 6108 6084 6110
rect 6104 6108 6120 6128
rect 6030 6102 6120 6108
rect 5544 6079 5581 6080
rect 4970 6062 5386 6067
rect 5543 6070 5581 6079
rect 4970 6061 5311 6062
rect 4752 5991 4789 6061
rect 4904 6001 4935 6002
rect 4565 5986 4702 5988
rect 4129 5953 4181 5955
rect 4565 5944 4608 5986
rect 4752 5971 4761 5991
rect 4781 5971 4789 5991
rect 4752 5961 4789 5971
rect 4848 5991 4935 6001
rect 4848 5971 4857 5991
rect 4877 5971 4935 5991
rect 4848 5962 4935 5971
rect 4848 5961 4885 5962
rect 4563 5934 4608 5944
rect 2969 5925 3006 5926
rect 2919 5916 3006 5925
rect 2919 5896 2977 5916
rect 2997 5896 3006 5916
rect 2919 5886 3006 5896
rect 3065 5916 3102 5926
rect 3065 5896 3073 5916
rect 3093 5896 3102 5916
rect 4563 5916 4572 5934
rect 4590 5916 4608 5934
rect 4563 5910 4608 5916
rect 4904 5911 4935 5962
rect 4970 5991 5007 6061
rect 5273 6060 5310 6061
rect 5543 6050 5552 6070
rect 5572 6050 5581 6070
rect 5543 6042 5581 6050
rect 5647 6074 5732 6080
rect 5762 6079 5799 6080
rect 5647 6054 5655 6074
rect 5675 6054 5732 6074
rect 5647 6046 5732 6054
rect 5761 6070 5799 6079
rect 5761 6050 5770 6070
rect 5790 6050 5799 6070
rect 5647 6045 5683 6046
rect 5761 6042 5799 6050
rect 5865 6074 6009 6080
rect 5865 6054 5873 6074
rect 5893 6055 5925 6074
rect 5946 6055 5981 6074
rect 5893 6054 5981 6055
rect 6001 6054 6009 6074
rect 5865 6046 6009 6054
rect 5865 6045 5901 6046
rect 5973 6045 6009 6046
rect 6075 6079 6112 6080
rect 6075 6078 6113 6079
rect 6075 6070 6139 6078
rect 6075 6050 6084 6070
rect 6104 6056 6139 6070
rect 6159 6056 6162 6076
rect 6104 6051 6162 6056
rect 6104 6050 6139 6051
rect 5544 6013 5581 6042
rect 5545 6011 5581 6013
rect 5122 6001 5158 6002
rect 4970 5971 4979 5991
rect 4999 5971 5007 5991
rect 4970 5961 5007 5971
rect 5066 5991 5214 6001
rect 5314 5998 5410 6000
rect 5066 5971 5075 5991
rect 5095 5971 5185 5991
rect 5205 5971 5214 5991
rect 5066 5962 5214 5971
rect 5272 5991 5410 5998
rect 5272 5971 5281 5991
rect 5301 5971 5410 5991
rect 5545 5989 5736 6011
rect 5762 6010 5799 6042
rect 6075 6038 6139 6050
rect 6179 6012 6206 6190
rect 6038 6010 6206 6012
rect 5762 5984 6206 6010
rect 5272 5962 5410 5971
rect 5066 5961 5103 5962
rect 4563 5907 4600 5910
rect 4796 5908 4837 5909
rect 2919 5885 2950 5886
rect 2543 5825 2884 5826
rect 3065 5825 3102 5896
rect 4688 5901 4837 5908
rect 4132 5888 4169 5893
rect 4123 5884 4170 5888
rect 4123 5866 4142 5884
rect 4160 5866 4170 5884
rect 4688 5881 4747 5901
rect 4767 5881 4806 5901
rect 4826 5881 4837 5901
rect 4688 5873 4837 5881
rect 4904 5904 5061 5911
rect 4904 5884 5024 5904
rect 5044 5884 5061 5904
rect 4904 5874 5061 5884
rect 4904 5873 4939 5874
rect 2468 5820 2884 5825
rect 2468 5800 2471 5820
rect 2491 5800 2884 5820
rect 2915 5801 3102 5825
rect 3727 5823 3767 5828
rect 4123 5823 4170 5866
rect 4904 5852 4935 5873
rect 5122 5852 5158 5962
rect 5177 5961 5214 5962
rect 5273 5961 5310 5962
rect 5233 5902 5323 5908
rect 5233 5882 5242 5902
rect 5262 5900 5323 5902
rect 5262 5882 5287 5900
rect 5233 5880 5287 5882
rect 5307 5880 5323 5900
rect 5233 5874 5323 5880
rect 4747 5851 4784 5852
rect 3727 5784 4170 5823
rect 4560 5843 4597 5845
rect 4560 5835 4602 5843
rect 4560 5817 4570 5835
rect 4588 5817 4602 5835
rect 4560 5808 4602 5817
rect 4746 5842 4784 5851
rect 4746 5822 4755 5842
rect 4775 5822 4784 5842
rect 4746 5814 4784 5822
rect 4850 5846 4935 5852
rect 4965 5851 5002 5852
rect 4850 5826 4858 5846
rect 4878 5826 4935 5846
rect 4850 5818 4935 5826
rect 4964 5842 5002 5851
rect 4964 5822 4973 5842
rect 4993 5822 5002 5842
rect 4850 5817 4886 5818
rect 4964 5814 5002 5822
rect 5068 5850 5212 5852
rect 5068 5846 5120 5850
rect 5068 5826 5076 5846
rect 5096 5830 5120 5846
rect 5140 5846 5212 5850
rect 5140 5830 5184 5846
rect 5096 5826 5184 5830
rect 5204 5826 5212 5846
rect 5068 5818 5212 5826
rect 5068 5817 5104 5818
rect 5176 5817 5212 5818
rect 5278 5851 5315 5852
rect 5278 5850 5316 5851
rect 5278 5842 5342 5850
rect 5278 5822 5287 5842
rect 5307 5828 5342 5842
rect 5362 5828 5365 5848
rect 5307 5823 5365 5828
rect 5307 5822 5342 5823
rect 2821 5769 2861 5777
rect 2821 5747 2829 5769
rect 2853 5747 2861 5769
rect 2527 5523 2695 5524
rect 2821 5523 2861 5747
rect 3324 5751 3492 5752
rect 3727 5751 3767 5784
rect 4123 5751 4170 5784
rect 4561 5783 4602 5808
rect 4747 5783 4784 5814
rect 4965 5783 5002 5814
rect 5278 5810 5342 5822
rect 5382 5784 5409 5962
rect 4561 5756 4610 5783
rect 4746 5757 4795 5783
rect 4964 5782 5045 5783
rect 5241 5782 5409 5784
rect 4964 5757 5409 5782
rect 4965 5756 5409 5757
rect 3324 5750 3768 5751
rect 3324 5725 3769 5750
rect 3324 5723 3492 5725
rect 3688 5724 3769 5725
rect 3938 5724 3987 5750
rect 4123 5724 4172 5751
rect 3324 5545 3351 5723
rect 3391 5685 3455 5697
rect 3731 5693 3768 5724
rect 3949 5693 3986 5724
rect 4131 5699 4172 5724
rect 4563 5723 4610 5756
rect 4966 5723 5006 5756
rect 5241 5755 5409 5756
rect 5872 5760 5912 5984
rect 6038 5983 6206 5984
rect 5872 5738 5880 5760
rect 5904 5738 5912 5760
rect 5872 5730 5912 5738
rect 3391 5684 3426 5685
rect 3368 5679 3426 5684
rect 3368 5659 3371 5679
rect 3391 5665 3426 5679
rect 3446 5665 3455 5685
rect 3391 5657 3455 5665
rect 3417 5656 3455 5657
rect 3418 5655 3455 5656
rect 3521 5689 3557 5690
rect 3629 5689 3665 5690
rect 3521 5681 3665 5689
rect 3521 5661 3529 5681
rect 3549 5677 3637 5681
rect 3549 5661 3593 5677
rect 3521 5657 3593 5661
rect 3613 5661 3637 5677
rect 3657 5661 3665 5681
rect 3613 5657 3665 5661
rect 3521 5655 3665 5657
rect 3731 5685 3769 5693
rect 3847 5689 3883 5690
rect 3731 5665 3740 5685
rect 3760 5665 3769 5685
rect 3731 5656 3769 5665
rect 3798 5681 3883 5689
rect 3798 5661 3855 5681
rect 3875 5661 3883 5681
rect 3731 5655 3768 5656
rect 3798 5655 3883 5661
rect 3949 5685 3987 5693
rect 3949 5665 3958 5685
rect 3978 5665 3987 5685
rect 3949 5656 3987 5665
rect 4131 5690 4173 5699
rect 4131 5672 4145 5690
rect 4163 5672 4173 5690
rect 4131 5664 4173 5672
rect 4136 5662 4173 5664
rect 4563 5684 5006 5723
rect 3949 5655 3986 5656
rect 3410 5627 3500 5633
rect 3410 5607 3426 5627
rect 3446 5625 3500 5627
rect 3446 5607 3471 5625
rect 3410 5605 3471 5607
rect 3491 5605 3500 5625
rect 3410 5599 3500 5605
rect 3423 5545 3460 5546
rect 3519 5545 3556 5546
rect 3575 5545 3611 5655
rect 3798 5634 3829 5655
rect 4563 5641 4610 5684
rect 4966 5679 5006 5684
rect 5631 5682 5818 5706
rect 5849 5687 6242 5707
rect 6262 5687 6265 5707
rect 5849 5682 6265 5687
rect 3794 5633 3829 5634
rect 3672 5623 3829 5633
rect 3672 5603 3689 5623
rect 3709 5603 3829 5623
rect 3672 5596 3829 5603
rect 3896 5626 4045 5634
rect 3896 5606 3907 5626
rect 3927 5606 3966 5626
rect 3986 5606 4045 5626
rect 4563 5623 4573 5641
rect 4591 5623 4610 5641
rect 4563 5619 4610 5623
rect 4564 5614 4601 5619
rect 3896 5599 4045 5606
rect 5631 5611 5668 5682
rect 5849 5681 6190 5682
rect 5783 5621 5814 5622
rect 3896 5598 3937 5599
rect 4133 5597 4170 5600
rect 3630 5545 3667 5546
rect 3323 5536 3461 5545
rect 2527 5497 2971 5523
rect 2527 5495 2695 5497
rect 2527 5317 2554 5495
rect 2594 5457 2658 5469
rect 2934 5465 2971 5497
rect 2997 5496 3188 5518
rect 3323 5516 3432 5536
rect 3452 5516 3461 5536
rect 3323 5509 3461 5516
rect 3519 5536 3667 5545
rect 3519 5516 3528 5536
rect 3548 5516 3638 5536
rect 3658 5516 3667 5536
rect 3323 5507 3419 5509
rect 3519 5506 3667 5516
rect 3726 5536 3763 5546
rect 3726 5516 3734 5536
rect 3754 5516 3763 5536
rect 3575 5505 3611 5506
rect 3152 5494 3188 5496
rect 3152 5465 3189 5494
rect 2594 5456 2629 5457
rect 2571 5451 2629 5456
rect 2571 5431 2574 5451
rect 2594 5437 2629 5451
rect 2649 5437 2658 5457
rect 2594 5429 2658 5437
rect 2620 5428 2658 5429
rect 2621 5427 2658 5428
rect 2724 5461 2760 5462
rect 2832 5461 2868 5462
rect 2724 5453 2868 5461
rect 2724 5433 2732 5453
rect 2752 5452 2840 5453
rect 2752 5433 2787 5452
rect 2808 5433 2840 5452
rect 2860 5433 2868 5453
rect 2724 5427 2868 5433
rect 2934 5457 2972 5465
rect 3050 5461 3086 5462
rect 2934 5437 2943 5457
rect 2963 5437 2972 5457
rect 2934 5428 2972 5437
rect 3001 5453 3086 5461
rect 3001 5433 3058 5453
rect 3078 5433 3086 5453
rect 2934 5427 2971 5428
rect 3001 5427 3086 5433
rect 3152 5457 3190 5465
rect 3152 5437 3161 5457
rect 3181 5437 3190 5457
rect 3423 5446 3460 5447
rect 3726 5446 3763 5516
rect 3798 5545 3829 5596
rect 4125 5591 4170 5597
rect 4125 5573 4143 5591
rect 4161 5573 4170 5591
rect 5631 5591 5640 5611
rect 5660 5591 5668 5611
rect 5631 5581 5668 5591
rect 5727 5611 5814 5621
rect 5727 5591 5736 5611
rect 5756 5591 5814 5611
rect 5727 5582 5814 5591
rect 5727 5581 5764 5582
rect 4125 5563 4170 5573
rect 3848 5545 3885 5546
rect 3798 5536 3885 5545
rect 3798 5516 3856 5536
rect 3876 5516 3885 5536
rect 3798 5506 3885 5516
rect 3944 5536 3981 5546
rect 3944 5516 3952 5536
rect 3972 5516 3981 5536
rect 4125 5521 4168 5563
rect 4552 5552 4604 5554
rect 4031 5519 4168 5521
rect 3798 5505 3829 5506
rect 3944 5446 3981 5516
rect 3422 5445 3763 5446
rect 3152 5428 3190 5437
rect 3347 5440 3763 5445
rect 3152 5427 3189 5428
rect 2613 5399 2703 5405
rect 2613 5379 2629 5399
rect 2649 5397 2703 5399
rect 2649 5379 2674 5397
rect 2613 5377 2674 5379
rect 2694 5377 2703 5397
rect 2613 5371 2703 5377
rect 2626 5317 2663 5318
rect 2722 5317 2759 5318
rect 2778 5317 2814 5427
rect 3001 5406 3032 5427
rect 3347 5420 3350 5440
rect 3370 5420 3763 5440
rect 3947 5430 3981 5446
rect 4025 5498 4168 5519
rect 4550 5548 4983 5552
rect 4550 5542 4989 5548
rect 4550 5524 4571 5542
rect 4589 5524 4989 5542
rect 5783 5531 5814 5582
rect 5849 5611 5886 5681
rect 6152 5680 6189 5681
rect 6001 5621 6037 5622
rect 5849 5591 5858 5611
rect 5878 5591 5886 5611
rect 5849 5581 5886 5591
rect 5945 5611 6093 5621
rect 6193 5618 6289 5620
rect 5945 5591 5954 5611
rect 5974 5591 6064 5611
rect 6084 5591 6093 5611
rect 5945 5582 6093 5591
rect 6151 5611 6289 5618
rect 6151 5591 6160 5611
rect 6180 5591 6289 5611
rect 6151 5582 6289 5591
rect 5945 5581 5982 5582
rect 5675 5528 5716 5529
rect 4550 5506 4989 5524
rect 3723 5411 3763 5420
rect 4025 5411 4052 5498
rect 4125 5472 4168 5498
rect 4125 5454 4138 5472
rect 4156 5454 4168 5472
rect 4125 5443 4168 5454
rect 2997 5405 3032 5406
rect 2875 5395 3032 5405
rect 2875 5375 2892 5395
rect 2912 5375 3032 5395
rect 2875 5368 3032 5375
rect 3099 5398 3248 5406
rect 3099 5378 3110 5398
rect 3130 5378 3169 5398
rect 3189 5378 3248 5398
rect 3723 5394 4052 5411
rect 3723 5393 3763 5394
rect 3099 5371 3248 5378
rect 4120 5382 4160 5385
rect 4120 5376 4163 5382
rect 3745 5373 4163 5376
rect 3099 5370 3140 5371
rect 2833 5317 2870 5318
rect 2526 5308 2664 5317
rect 2224 5133 2264 5305
rect 2526 5288 2635 5308
rect 2655 5288 2664 5308
rect 2526 5281 2664 5288
rect 2722 5308 2870 5317
rect 2722 5288 2731 5308
rect 2751 5288 2841 5308
rect 2861 5288 2870 5308
rect 2526 5279 2622 5281
rect 2722 5278 2870 5288
rect 2929 5308 2966 5318
rect 2929 5288 2937 5308
rect 2957 5288 2966 5308
rect 2778 5277 2814 5278
rect 2626 5218 2663 5219
rect 2929 5218 2966 5288
rect 3001 5317 3032 5368
rect 3745 5355 4136 5373
rect 4154 5355 4163 5373
rect 3745 5353 4163 5355
rect 3745 5345 3772 5353
rect 4013 5350 4163 5353
rect 3325 5339 3493 5340
rect 3744 5339 3772 5345
rect 3325 5323 3772 5339
rect 4120 5345 4163 5350
rect 3051 5317 3088 5318
rect 3001 5308 3088 5317
rect 3001 5288 3059 5308
rect 3079 5288 3088 5308
rect 3001 5278 3088 5288
rect 3147 5308 3184 5318
rect 3147 5288 3155 5308
rect 3175 5288 3184 5308
rect 3001 5277 3032 5278
rect 2625 5217 2966 5218
rect 3147 5217 3184 5288
rect 2550 5212 2966 5217
rect 2550 5192 2553 5212
rect 2573 5192 2966 5212
rect 2997 5193 3184 5217
rect 3325 5313 3769 5323
rect 3325 5311 3493 5313
rect 3325 5133 3352 5311
rect 3392 5273 3456 5285
rect 3732 5281 3769 5313
rect 3795 5312 3986 5334
rect 3950 5310 3986 5312
rect 3950 5281 3987 5310
rect 4120 5289 4160 5345
rect 3392 5272 3427 5273
rect 3369 5267 3427 5272
rect 3369 5247 3372 5267
rect 3392 5253 3427 5267
rect 3447 5253 3456 5273
rect 3392 5245 3456 5253
rect 3418 5244 3456 5245
rect 3419 5243 3456 5244
rect 3522 5277 3558 5278
rect 3630 5277 3666 5278
rect 3522 5269 3666 5277
rect 3522 5249 3530 5269
rect 3550 5249 3585 5269
rect 3605 5249 3638 5269
rect 3658 5249 3666 5269
rect 3522 5243 3666 5249
rect 3732 5273 3770 5281
rect 3848 5277 3884 5278
rect 3732 5253 3741 5273
rect 3761 5253 3770 5273
rect 3732 5244 3770 5253
rect 3799 5269 3884 5277
rect 3799 5249 3856 5269
rect 3876 5249 3884 5269
rect 3732 5243 3769 5244
rect 3799 5243 3884 5249
rect 3950 5273 3988 5281
rect 3950 5253 3959 5273
rect 3979 5253 3988 5273
rect 4120 5271 4132 5289
rect 4150 5271 4160 5289
rect 4552 5317 4604 5506
rect 4950 5481 4989 5506
rect 5567 5521 5716 5528
rect 5567 5501 5626 5521
rect 5646 5501 5685 5521
rect 5705 5501 5716 5521
rect 5567 5493 5716 5501
rect 5783 5524 5940 5531
rect 5783 5504 5903 5524
rect 5923 5504 5940 5524
rect 5783 5494 5940 5504
rect 5783 5493 5818 5494
rect 4734 5456 4921 5480
rect 4950 5461 5345 5481
rect 5365 5461 5368 5481
rect 5783 5472 5814 5493
rect 6001 5472 6037 5582
rect 6056 5581 6093 5582
rect 6152 5581 6189 5582
rect 6112 5522 6202 5528
rect 6112 5502 6121 5522
rect 6141 5520 6202 5522
rect 6141 5502 6166 5520
rect 6112 5500 6166 5502
rect 6186 5500 6202 5520
rect 6112 5494 6202 5500
rect 5626 5471 5663 5472
rect 4950 5456 5368 5461
rect 5625 5462 5663 5471
rect 4734 5385 4771 5456
rect 4950 5455 5293 5456
rect 4950 5452 4989 5455
rect 5255 5454 5292 5455
rect 4886 5395 4917 5396
rect 4734 5365 4743 5385
rect 4763 5365 4771 5385
rect 4734 5355 4771 5365
rect 4830 5385 4917 5395
rect 4830 5365 4839 5385
rect 4859 5365 4917 5385
rect 4830 5356 4917 5365
rect 4830 5355 4867 5356
rect 4552 5299 4568 5317
rect 4586 5299 4604 5317
rect 4886 5305 4917 5356
rect 4952 5385 4989 5452
rect 5625 5442 5634 5462
rect 5654 5442 5663 5462
rect 5625 5434 5663 5442
rect 5729 5466 5814 5472
rect 5844 5471 5881 5472
rect 5729 5446 5737 5466
rect 5757 5446 5814 5466
rect 5729 5438 5814 5446
rect 5843 5462 5881 5471
rect 5843 5442 5852 5462
rect 5872 5442 5881 5462
rect 5729 5437 5765 5438
rect 5843 5434 5881 5442
rect 5947 5466 6091 5472
rect 5947 5446 5955 5466
rect 5975 5461 6063 5466
rect 5975 5446 6011 5461
rect 5947 5444 6011 5446
rect 6030 5446 6063 5461
rect 6083 5446 6091 5466
rect 6030 5444 6091 5446
rect 5947 5438 6091 5444
rect 5947 5437 5983 5438
rect 6055 5437 6091 5438
rect 6157 5471 6194 5472
rect 6157 5470 6195 5471
rect 6157 5462 6221 5470
rect 6157 5442 6166 5462
rect 6186 5448 6221 5462
rect 6241 5448 6244 5468
rect 6186 5443 6244 5448
rect 6186 5442 6221 5443
rect 5626 5405 5663 5434
rect 5627 5403 5663 5405
rect 5104 5395 5140 5396
rect 4952 5365 4961 5385
rect 4981 5365 4989 5385
rect 4952 5355 4989 5365
rect 5048 5385 5196 5395
rect 5296 5392 5392 5394
rect 5048 5365 5057 5385
rect 5077 5365 5167 5385
rect 5187 5365 5196 5385
rect 5048 5356 5196 5365
rect 5254 5385 5392 5392
rect 5254 5365 5263 5385
rect 5283 5365 5392 5385
rect 5627 5381 5818 5403
rect 5844 5402 5881 5434
rect 6157 5430 6221 5442
rect 6261 5404 6288 5582
rect 6120 5402 6288 5404
rect 5844 5388 6288 5402
rect 6312 5425 6340 6371
rect 6312 5395 6357 5425
rect 5844 5376 6291 5388
rect 5887 5374 5920 5376
rect 5254 5356 5392 5365
rect 5048 5355 5085 5356
rect 4778 5302 4819 5303
rect 4552 5281 4604 5299
rect 4670 5295 4819 5302
rect 4120 5261 4160 5271
rect 4670 5275 4729 5295
rect 4749 5275 4788 5295
rect 4808 5275 4819 5295
rect 4670 5267 4819 5275
rect 4886 5298 5043 5305
rect 4886 5278 5006 5298
rect 5026 5278 5043 5298
rect 4886 5268 5043 5278
rect 4886 5267 4921 5268
rect 3950 5244 3988 5253
rect 4886 5246 4917 5267
rect 5104 5246 5140 5356
rect 5159 5355 5196 5356
rect 5255 5355 5292 5356
rect 5215 5296 5305 5302
rect 5215 5276 5224 5296
rect 5244 5294 5305 5296
rect 5244 5276 5269 5294
rect 5215 5274 5269 5276
rect 5289 5274 5305 5294
rect 5215 5268 5305 5274
rect 4729 5245 4766 5246
rect 3950 5243 3987 5244
rect 3411 5215 3501 5221
rect 3411 5195 3427 5215
rect 3447 5213 3501 5215
rect 3447 5195 3472 5213
rect 3411 5193 3472 5195
rect 3492 5193 3501 5213
rect 3411 5187 3501 5193
rect 3424 5133 3461 5134
rect 3520 5133 3557 5134
rect 3576 5133 3612 5243
rect 3799 5222 3830 5243
rect 4728 5236 4766 5245
rect 3795 5221 3830 5222
rect 3673 5211 3830 5221
rect 3673 5191 3690 5211
rect 3710 5191 3830 5211
rect 3673 5184 3830 5191
rect 3897 5214 4046 5222
rect 3897 5194 3908 5214
rect 3928 5194 3967 5214
rect 3987 5194 4046 5214
rect 4556 5218 4596 5228
rect 3897 5187 4046 5194
rect 4112 5190 4164 5208
rect 3897 5186 3938 5187
rect 3631 5133 3668 5134
rect 2225 5118 2264 5133
rect 3324 5124 3462 5133
rect 2225 5117 2391 5118
rect 2517 5117 2557 5119
rect 2225 5091 2667 5117
rect 2225 5089 2391 5091
rect 1889 4977 1926 4985
rect 1889 4958 1897 4977
rect 1918 4958 1926 4977
rect 1889 4952 1926 4958
rect 2225 4911 2250 5089
rect 2290 5051 2354 5063
rect 2630 5059 2667 5091
rect 2693 5090 2884 5112
rect 3324 5104 3433 5124
rect 3453 5104 3462 5124
rect 3324 5097 3462 5104
rect 3520 5124 3668 5133
rect 3520 5104 3529 5124
rect 3549 5104 3639 5124
rect 3659 5104 3668 5124
rect 3324 5095 3420 5097
rect 3520 5094 3668 5104
rect 3727 5124 3764 5134
rect 3727 5104 3735 5124
rect 3755 5104 3764 5124
rect 3576 5093 3612 5094
rect 2848 5088 2884 5090
rect 2848 5059 2885 5088
rect 2290 5050 2325 5051
rect 2267 5045 2325 5050
rect 2267 5025 2270 5045
rect 2290 5031 2325 5045
rect 2345 5031 2354 5051
rect 2290 5023 2354 5031
rect 2316 5022 2354 5023
rect 2317 5021 2354 5022
rect 2420 5055 2456 5056
rect 2528 5055 2564 5056
rect 2420 5050 2564 5055
rect 2420 5047 2482 5050
rect 2420 5027 2428 5047
rect 2448 5027 2482 5047
rect 2420 5024 2482 5027
rect 2508 5047 2564 5050
rect 2508 5027 2536 5047
rect 2556 5027 2564 5047
rect 2508 5024 2564 5027
rect 2420 5021 2564 5024
rect 2630 5051 2668 5059
rect 2746 5055 2782 5056
rect 2630 5031 2639 5051
rect 2659 5031 2668 5051
rect 2630 5022 2668 5031
rect 2697 5047 2782 5055
rect 2697 5027 2754 5047
rect 2774 5027 2782 5047
rect 2630 5021 2667 5022
rect 2697 5021 2782 5027
rect 2848 5051 2886 5059
rect 2848 5031 2857 5051
rect 2877 5031 2886 5051
rect 3727 5037 3764 5104
rect 3799 5133 3830 5184
rect 4112 5172 4130 5190
rect 4148 5172 4164 5190
rect 3849 5133 3886 5134
rect 3799 5124 3886 5133
rect 3799 5104 3857 5124
rect 3877 5104 3886 5124
rect 3799 5094 3886 5104
rect 3945 5124 3982 5134
rect 3945 5104 3953 5124
rect 3973 5104 3982 5124
rect 3799 5093 3830 5094
rect 3424 5034 3461 5035
rect 3727 5034 3766 5037
rect 3423 5033 3766 5034
rect 3945 5033 3982 5104
rect 2848 5022 2886 5031
rect 3348 5028 3766 5033
rect 2848 5021 2885 5022
rect 2309 4993 2399 4999
rect 2309 4973 2325 4993
rect 2345 4991 2399 4993
rect 2345 4973 2370 4991
rect 2309 4971 2370 4973
rect 2390 4971 2399 4991
rect 2309 4965 2399 4971
rect 2322 4911 2359 4912
rect 2418 4911 2455 4912
rect 2474 4911 2510 5021
rect 2697 5000 2728 5021
rect 3348 5008 3351 5028
rect 3371 5008 3766 5028
rect 3795 5009 3982 5033
rect 2693 4999 2728 5000
rect 2571 4989 2728 4999
rect 2571 4969 2588 4989
rect 2608 4969 2728 4989
rect 2571 4962 2728 4969
rect 2795 4992 2944 5000
rect 2795 4972 2806 4992
rect 2826 4972 2865 4992
rect 2885 4972 2944 4992
rect 2795 4965 2944 4972
rect 3727 4983 3766 5008
rect 4112 4983 4164 5172
rect 4556 5200 4566 5218
rect 4584 5200 4596 5218
rect 4728 5216 4737 5236
rect 4757 5216 4766 5236
rect 4728 5208 4766 5216
rect 4832 5240 4917 5246
rect 4947 5245 4984 5246
rect 4832 5220 4840 5240
rect 4860 5220 4917 5240
rect 4832 5212 4917 5220
rect 4946 5236 4984 5245
rect 4946 5216 4955 5236
rect 4975 5216 4984 5236
rect 4832 5211 4868 5212
rect 4946 5208 4984 5216
rect 5050 5240 5194 5246
rect 5050 5220 5058 5240
rect 5078 5220 5111 5240
rect 5131 5220 5166 5240
rect 5186 5220 5194 5240
rect 5050 5212 5194 5220
rect 5050 5211 5086 5212
rect 5158 5211 5194 5212
rect 5260 5245 5297 5246
rect 5260 5244 5298 5245
rect 5260 5236 5324 5244
rect 5260 5216 5269 5236
rect 5289 5222 5324 5236
rect 5344 5222 5347 5242
rect 5289 5217 5347 5222
rect 5289 5216 5324 5217
rect 4556 5144 4596 5200
rect 4729 5179 4766 5208
rect 4730 5177 4766 5179
rect 4730 5155 4921 5177
rect 4947 5176 4984 5208
rect 5260 5204 5324 5216
rect 5364 5178 5391 5356
rect 6249 5331 6291 5376
rect 6312 5377 6323 5395
rect 6345 5377 6357 5395
rect 6312 5371 6357 5377
rect 6313 5370 6357 5371
rect 5223 5176 5391 5178
rect 4947 5166 5391 5176
rect 5532 5272 5719 5296
rect 5750 5277 6143 5297
rect 6163 5277 6166 5297
rect 5750 5272 6166 5277
rect 5532 5201 5569 5272
rect 5750 5271 6091 5272
rect 5684 5211 5715 5212
rect 5532 5181 5541 5201
rect 5561 5181 5569 5201
rect 5532 5171 5569 5181
rect 5628 5201 5715 5211
rect 5628 5181 5637 5201
rect 5657 5181 5715 5201
rect 5628 5172 5715 5181
rect 5628 5171 5665 5172
rect 4553 5139 4596 5144
rect 4944 5150 5391 5166
rect 4944 5144 4972 5150
rect 5223 5149 5391 5150
rect 4553 5136 4703 5139
rect 4944 5136 4971 5144
rect 4553 5134 4971 5136
rect 4553 5116 4562 5134
rect 4580 5116 4971 5134
rect 5684 5121 5715 5172
rect 5750 5201 5787 5271
rect 6053 5270 6090 5271
rect 5902 5211 5938 5212
rect 5750 5181 5759 5201
rect 5779 5181 5787 5201
rect 5750 5171 5787 5181
rect 5846 5201 5994 5211
rect 6094 5208 6190 5210
rect 5846 5181 5855 5201
rect 5875 5181 5965 5201
rect 5985 5181 5994 5201
rect 5846 5172 5994 5181
rect 6052 5201 6190 5208
rect 6052 5181 6061 5201
rect 6081 5181 6190 5201
rect 6052 5172 6190 5181
rect 5846 5171 5883 5172
rect 5576 5118 5617 5119
rect 4553 5113 4971 5116
rect 4553 5107 4596 5113
rect 4556 5104 4596 5107
rect 5471 5111 5617 5118
rect 4953 5095 4993 5096
rect 4664 5078 4993 5095
rect 5471 5091 5527 5111
rect 5547 5091 5586 5111
rect 5606 5091 5617 5111
rect 5471 5083 5617 5091
rect 5684 5114 5841 5121
rect 5684 5094 5804 5114
rect 5824 5094 5841 5114
rect 5684 5084 5841 5094
rect 5684 5083 5719 5084
rect 4548 5035 4591 5046
rect 4548 5017 4560 5035
rect 4578 5017 4591 5035
rect 4548 4991 4591 5017
rect 4664 4991 4691 5078
rect 4953 5069 4993 5078
rect 3727 4965 4166 4983
rect 2795 4964 2836 4965
rect 2529 4911 2566 4912
rect 2225 4902 2360 4911
rect 2225 4882 2331 4902
rect 2351 4882 2360 4902
rect 2225 4875 2360 4882
rect 2418 4902 2566 4911
rect 2418 4882 2427 4902
rect 2447 4882 2537 4902
rect 2557 4882 2566 4902
rect 2225 4873 2318 4875
rect 2418 4872 2566 4882
rect 2625 4902 2662 4912
rect 2625 4882 2633 4902
rect 2653 4882 2662 4902
rect 2474 4871 2510 4872
rect 2322 4812 2359 4813
rect 2625 4812 2662 4882
rect 2697 4911 2728 4962
rect 3727 4947 4127 4965
rect 4145 4947 4166 4965
rect 3727 4941 4166 4947
rect 3733 4937 4166 4941
rect 4548 4970 4691 4991
rect 4735 5043 4769 5059
rect 4953 5049 5346 5069
rect 5366 5049 5369 5069
rect 5684 5062 5715 5083
rect 5902 5062 5938 5172
rect 5957 5171 5994 5172
rect 6053 5171 6090 5172
rect 6013 5112 6103 5118
rect 6013 5092 6022 5112
rect 6042 5110 6103 5112
rect 6042 5092 6067 5110
rect 6013 5090 6067 5092
rect 6087 5090 6103 5110
rect 6013 5084 6103 5090
rect 5527 5061 5564 5062
rect 4953 5044 5369 5049
rect 5526 5052 5564 5061
rect 4953 5043 5294 5044
rect 4735 4973 4772 5043
rect 4887 4983 4918 4984
rect 4548 4968 4685 4970
rect 4112 4935 4164 4937
rect 4548 4926 4591 4968
rect 4735 4953 4744 4973
rect 4764 4953 4772 4973
rect 4735 4943 4772 4953
rect 4831 4973 4918 4983
rect 4831 4953 4840 4973
rect 4860 4953 4918 4973
rect 4831 4944 4918 4953
rect 4831 4943 4868 4944
rect 4546 4916 4591 4926
rect 2747 4911 2784 4912
rect 2697 4902 2784 4911
rect 2697 4882 2755 4902
rect 2775 4882 2784 4902
rect 2697 4872 2784 4882
rect 2843 4902 2880 4912
rect 2843 4882 2851 4902
rect 2871 4882 2880 4902
rect 4546 4898 4555 4916
rect 4573 4898 4591 4916
rect 4546 4892 4591 4898
rect 4887 4893 4918 4944
rect 4953 4973 4990 5043
rect 5256 5042 5293 5043
rect 5526 5032 5535 5052
rect 5555 5032 5564 5052
rect 5526 5024 5564 5032
rect 5630 5056 5715 5062
rect 5745 5061 5782 5062
rect 5630 5036 5638 5056
rect 5658 5036 5715 5056
rect 5630 5028 5715 5036
rect 5744 5052 5782 5061
rect 5744 5032 5753 5052
rect 5773 5032 5782 5052
rect 5630 5027 5666 5028
rect 5744 5024 5782 5032
rect 5848 5056 5992 5062
rect 5848 5036 5856 5056
rect 5876 5053 5964 5056
rect 5876 5036 5911 5053
rect 5848 5035 5911 5036
rect 5930 5036 5964 5053
rect 5984 5036 5992 5056
rect 5930 5035 5992 5036
rect 5848 5028 5992 5035
rect 5848 5027 5884 5028
rect 5956 5027 5992 5028
rect 6058 5061 6095 5062
rect 6058 5060 6096 5061
rect 6118 5060 6145 5064
rect 6058 5058 6145 5060
rect 6058 5052 6122 5058
rect 6058 5032 6067 5052
rect 6087 5038 6122 5052
rect 6142 5038 6145 5058
rect 6087 5033 6145 5038
rect 6087 5032 6122 5033
rect 5527 4995 5564 5024
rect 5528 4993 5564 4995
rect 5105 4983 5141 4984
rect 4953 4953 4962 4973
rect 4982 4953 4990 4973
rect 4953 4943 4990 4953
rect 5049 4973 5197 4983
rect 5297 4980 5393 4982
rect 5049 4953 5058 4973
rect 5078 4953 5168 4973
rect 5188 4953 5197 4973
rect 5049 4944 5197 4953
rect 5255 4973 5393 4980
rect 5255 4953 5264 4973
rect 5284 4953 5393 4973
rect 5528 4971 5719 4993
rect 5745 4992 5782 5024
rect 6058 5020 6122 5032
rect 6162 4994 6189 5172
rect 6021 4992 6189 4994
rect 5745 4966 6189 4992
rect 5255 4944 5393 4953
rect 5049 4943 5086 4944
rect 4546 4889 4583 4892
rect 4779 4890 4820 4891
rect 2697 4871 2728 4872
rect 2321 4811 2662 4812
rect 2843 4811 2880 4882
rect 4671 4883 4820 4890
rect 4115 4870 4152 4875
rect 2246 4806 2662 4811
rect 2246 4786 2249 4806
rect 2269 4786 2662 4806
rect 2693 4787 2880 4811
rect 4106 4866 4153 4870
rect 4106 4848 4125 4866
rect 4143 4848 4153 4866
rect 4671 4863 4730 4883
rect 4750 4863 4789 4883
rect 4809 4863 4820 4883
rect 4671 4855 4820 4863
rect 4887 4886 5044 4893
rect 4887 4866 5007 4886
rect 5027 4866 5044 4886
rect 4887 4856 5044 4866
rect 4887 4855 4922 4856
rect 3714 4789 3752 4790
rect 4106 4789 4153 4848
rect 4887 4834 4918 4855
rect 5105 4834 5141 4944
rect 5160 4943 5197 4944
rect 5256 4943 5293 4944
rect 5216 4884 5306 4890
rect 5216 4864 5225 4884
rect 5245 4882 5306 4884
rect 5245 4864 5270 4882
rect 5216 4862 5270 4864
rect 5290 4862 5306 4882
rect 5216 4856 5306 4862
rect 4730 4833 4767 4834
rect 4543 4825 4580 4827
rect 4543 4817 4585 4825
rect 4543 4799 4553 4817
rect 4571 4799 4585 4817
rect 4543 4790 4585 4799
rect 4729 4824 4767 4833
rect 4729 4804 4738 4824
rect 4758 4804 4767 4824
rect 4729 4796 4767 4804
rect 4833 4828 4918 4834
rect 4948 4833 4985 4834
rect 4833 4808 4841 4828
rect 4861 4808 4918 4828
rect 4833 4800 4918 4808
rect 4947 4824 4985 4833
rect 4947 4804 4956 4824
rect 4976 4804 4985 4824
rect 4833 4799 4869 4800
rect 4947 4796 4985 4804
rect 5051 4832 5195 4834
rect 5051 4828 5103 4832
rect 5051 4808 5059 4828
rect 5079 4812 5103 4828
rect 5123 4828 5195 4832
rect 5123 4812 5167 4828
rect 5079 4808 5167 4812
rect 5187 4808 5195 4828
rect 5051 4800 5195 4808
rect 5051 4799 5087 4800
rect 5159 4799 5195 4800
rect 5261 4833 5298 4834
rect 5261 4832 5299 4833
rect 5261 4824 5325 4832
rect 5261 4804 5270 4824
rect 5290 4810 5325 4824
rect 5345 4810 5348 4830
rect 5290 4805 5348 4810
rect 5290 4804 5325 4805
rect 2466 4785 2531 4786
rect 581 4707 619 4708
rect 180 4669 619 4707
rect 1491 4707 1499 4729
rect 1523 4707 1531 4729
rect 1491 4699 1531 4707
rect 2802 4751 2842 4759
rect 2802 4729 2810 4751
rect 2834 4729 2842 4751
rect 3714 4751 4153 4789
rect 3714 4750 3752 4751
rect 1802 4672 1867 4673
rect 180 4610 227 4669
rect 581 4668 619 4669
rect 180 4592 190 4610
rect 208 4592 227 4610
rect 180 4588 227 4592
rect 1453 4647 1640 4671
rect 1671 4652 2064 4672
rect 2084 4652 2087 4672
rect 1671 4647 2087 4652
rect 181 4583 218 4588
rect 1453 4576 1490 4647
rect 1671 4646 2012 4647
rect 1605 4586 1636 4587
rect 1453 4556 1462 4576
rect 1482 4556 1490 4576
rect 1453 4546 1490 4556
rect 1549 4576 1636 4586
rect 1549 4556 1558 4576
rect 1578 4556 1636 4576
rect 1549 4547 1636 4556
rect 1549 4546 1586 4547
rect 169 4521 221 4523
rect 167 4517 600 4521
rect 167 4511 606 4517
rect 167 4493 188 4511
rect 206 4493 606 4511
rect 1605 4496 1636 4547
rect 1671 4576 1708 4646
rect 1974 4645 2011 4646
rect 1823 4586 1859 4587
rect 1671 4556 1680 4576
rect 1700 4556 1708 4576
rect 1671 4546 1708 4556
rect 1767 4576 1915 4586
rect 2015 4583 2111 4585
rect 1767 4556 1776 4576
rect 1796 4556 1886 4576
rect 1906 4556 1915 4576
rect 1767 4547 1915 4556
rect 1973 4576 2111 4583
rect 1973 4556 1982 4576
rect 2002 4556 2111 4576
rect 1973 4547 2111 4556
rect 1767 4546 1804 4547
rect 1497 4493 1538 4494
rect 167 4475 606 4493
rect 169 4286 221 4475
rect 567 4450 606 4475
rect 1389 4486 1538 4493
rect 1389 4466 1448 4486
rect 1468 4466 1507 4486
rect 1527 4466 1538 4486
rect 1389 4458 1538 4466
rect 1605 4489 1762 4496
rect 1605 4469 1725 4489
rect 1745 4469 1762 4489
rect 1605 4459 1762 4469
rect 1605 4458 1640 4459
rect 351 4425 538 4449
rect 567 4430 962 4450
rect 982 4430 985 4450
rect 1605 4437 1636 4458
rect 1823 4437 1859 4547
rect 1878 4546 1915 4547
rect 1974 4546 2011 4547
rect 1934 4487 2024 4493
rect 1934 4467 1943 4487
rect 1963 4485 2024 4487
rect 1963 4467 1988 4485
rect 1934 4465 1988 4467
rect 2008 4465 2024 4485
rect 1934 4459 2024 4465
rect 1448 4436 1485 4437
rect 567 4425 985 4430
rect 1447 4427 1485 4436
rect 351 4354 388 4425
rect 567 4424 910 4425
rect 567 4421 606 4424
rect 872 4423 909 4424
rect 503 4364 534 4365
rect 351 4334 360 4354
rect 380 4334 388 4354
rect 351 4324 388 4334
rect 447 4354 534 4364
rect 447 4334 456 4354
rect 476 4334 534 4354
rect 447 4325 534 4334
rect 447 4324 484 4325
rect 169 4268 185 4286
rect 203 4268 221 4286
rect 503 4274 534 4325
rect 569 4354 606 4421
rect 1447 4407 1456 4427
rect 1476 4407 1485 4427
rect 1447 4399 1485 4407
rect 1551 4431 1636 4437
rect 1666 4436 1703 4437
rect 1551 4411 1559 4431
rect 1579 4411 1636 4431
rect 1551 4403 1636 4411
rect 1665 4427 1703 4436
rect 1665 4407 1674 4427
rect 1694 4407 1703 4427
rect 1551 4402 1587 4403
rect 1665 4399 1703 4407
rect 1769 4431 1913 4437
rect 1769 4411 1777 4431
rect 1797 4425 1885 4431
rect 1797 4411 1826 4425
rect 1769 4403 1826 4411
rect 1769 4402 1805 4403
rect 1849 4411 1885 4425
rect 1905 4411 1913 4431
rect 1849 4403 1913 4411
rect 1877 4402 1913 4403
rect 1979 4436 2016 4437
rect 1979 4435 2017 4436
rect 1979 4427 2043 4435
rect 1979 4407 1988 4427
rect 2008 4413 2043 4427
rect 2063 4413 2066 4433
rect 2008 4408 2066 4413
rect 2008 4407 2043 4408
rect 1448 4370 1485 4399
rect 1449 4368 1485 4370
rect 721 4364 757 4365
rect 569 4334 578 4354
rect 598 4334 606 4354
rect 569 4324 606 4334
rect 665 4354 813 4364
rect 913 4361 1009 4363
rect 665 4334 674 4354
rect 694 4334 784 4354
rect 804 4334 813 4354
rect 665 4325 813 4334
rect 871 4354 1009 4361
rect 871 4334 880 4354
rect 900 4334 1009 4354
rect 1449 4346 1640 4368
rect 1666 4367 1703 4399
rect 1979 4395 2043 4407
rect 2083 4369 2110 4547
rect 2407 4500 2444 4506
rect 2407 4481 2415 4500
rect 2436 4481 2444 4500
rect 2407 4473 2444 4481
rect 1942 4367 2110 4369
rect 1666 4341 2110 4367
rect 1776 4339 1816 4341
rect 1942 4340 2110 4341
rect 871 4325 1009 4334
rect 2069 4335 2110 4340
rect 665 4324 702 4325
rect 395 4271 436 4272
rect 169 4250 221 4268
rect 287 4264 436 4271
rect 287 4244 346 4264
rect 366 4244 405 4264
rect 425 4244 436 4264
rect 287 4236 436 4244
rect 503 4267 660 4274
rect 503 4247 623 4267
rect 643 4247 660 4267
rect 503 4237 660 4247
rect 503 4236 538 4237
rect 503 4215 534 4236
rect 721 4215 757 4325
rect 776 4324 813 4325
rect 872 4324 909 4325
rect 832 4265 922 4271
rect 832 4245 841 4265
rect 861 4263 922 4265
rect 861 4245 886 4263
rect 832 4243 886 4245
rect 906 4243 922 4263
rect 832 4237 922 4243
rect 346 4214 383 4215
rect 345 4205 383 4214
rect 173 4187 213 4197
rect 173 4169 183 4187
rect 201 4169 213 4187
rect 345 4185 354 4205
rect 374 4185 383 4205
rect 345 4177 383 4185
rect 449 4209 534 4215
rect 564 4214 601 4215
rect 449 4189 457 4209
rect 477 4189 534 4209
rect 449 4181 534 4189
rect 563 4205 601 4214
rect 563 4185 572 4205
rect 592 4185 601 4205
rect 449 4180 485 4181
rect 563 4177 601 4185
rect 667 4209 811 4215
rect 667 4189 675 4209
rect 695 4189 728 4209
rect 748 4189 783 4209
rect 803 4189 811 4209
rect 667 4181 811 4189
rect 667 4180 703 4181
rect 775 4180 811 4181
rect 877 4214 914 4215
rect 877 4213 915 4214
rect 877 4205 941 4213
rect 877 4185 886 4205
rect 906 4191 941 4205
rect 961 4191 964 4211
rect 906 4186 964 4191
rect 906 4185 941 4186
rect 173 4113 213 4169
rect 346 4148 383 4177
rect 347 4146 383 4148
rect 347 4124 538 4146
rect 564 4145 601 4177
rect 877 4173 941 4185
rect 981 4147 1008 4325
rect 840 4145 1008 4147
rect 564 4135 1008 4145
rect 1149 4241 1336 4265
rect 1367 4246 1760 4266
rect 1780 4246 1783 4266
rect 1367 4241 1783 4246
rect 1149 4170 1186 4241
rect 1367 4240 1708 4241
rect 1301 4180 1332 4181
rect 1149 4150 1158 4170
rect 1178 4150 1186 4170
rect 1149 4140 1186 4150
rect 1245 4170 1332 4180
rect 1245 4150 1254 4170
rect 1274 4150 1332 4170
rect 1245 4141 1332 4150
rect 1245 4140 1282 4141
rect 170 4108 213 4113
rect 561 4119 1008 4135
rect 561 4113 589 4119
rect 840 4118 1008 4119
rect 170 4105 320 4108
rect 561 4105 588 4113
rect 170 4103 588 4105
rect 170 4085 179 4103
rect 197 4085 588 4103
rect 1301 4090 1332 4141
rect 1367 4170 1404 4240
rect 1670 4239 1707 4240
rect 1519 4180 1555 4181
rect 1367 4150 1376 4170
rect 1396 4150 1404 4170
rect 1367 4140 1404 4150
rect 1463 4170 1611 4180
rect 1711 4177 1807 4179
rect 1463 4150 1472 4170
rect 1492 4150 1582 4170
rect 1602 4150 1611 4170
rect 1463 4141 1611 4150
rect 1669 4170 1807 4177
rect 1669 4150 1678 4170
rect 1698 4150 1807 4170
rect 2069 4153 2109 4335
rect 1669 4141 1807 4150
rect 1463 4140 1500 4141
rect 1193 4087 1234 4088
rect 170 4082 588 4085
rect 170 4076 213 4082
rect 173 4073 213 4076
rect 1085 4080 1234 4087
rect 570 4064 610 4065
rect 281 4047 610 4064
rect 1085 4060 1144 4080
rect 1164 4060 1203 4080
rect 1223 4060 1234 4080
rect 1085 4052 1234 4060
rect 1301 4083 1458 4090
rect 1301 4063 1421 4083
rect 1441 4063 1458 4083
rect 1301 4053 1458 4063
rect 1301 4052 1336 4053
rect 165 4004 208 4015
rect 165 3986 177 4004
rect 195 3986 208 4004
rect 165 3960 208 3986
rect 281 3960 308 4047
rect 570 4038 610 4047
rect 165 3939 308 3960
rect 352 4012 386 4028
rect 570 4018 963 4038
rect 983 4018 986 4038
rect 1301 4031 1332 4052
rect 1519 4031 1555 4141
rect 1574 4140 1611 4141
rect 1670 4140 1707 4141
rect 1630 4081 1720 4087
rect 1630 4061 1639 4081
rect 1659 4079 1720 4081
rect 1659 4061 1684 4079
rect 1630 4059 1684 4061
rect 1704 4059 1720 4079
rect 1630 4053 1720 4059
rect 1144 4030 1181 4031
rect 570 4013 986 4018
rect 1143 4021 1181 4030
rect 570 4012 911 4013
rect 352 3942 389 4012
rect 504 3952 535 3953
rect 165 3937 302 3939
rect 165 3895 208 3937
rect 352 3922 361 3942
rect 381 3922 389 3942
rect 352 3912 389 3922
rect 448 3942 535 3952
rect 448 3922 457 3942
rect 477 3922 535 3942
rect 448 3913 535 3922
rect 448 3912 485 3913
rect 163 3885 208 3895
rect 163 3867 172 3885
rect 190 3867 208 3885
rect 163 3861 208 3867
rect 504 3862 535 3913
rect 570 3942 607 4012
rect 873 4011 910 4012
rect 1143 4001 1152 4021
rect 1172 4001 1181 4021
rect 1143 3993 1181 4001
rect 1247 4025 1332 4031
rect 1362 4030 1399 4031
rect 1247 4005 1255 4025
rect 1275 4005 1332 4025
rect 1247 3997 1332 4005
rect 1361 4021 1399 4030
rect 1361 4001 1370 4021
rect 1390 4001 1399 4021
rect 1247 3996 1283 3997
rect 1361 3993 1399 4001
rect 1465 4025 1609 4031
rect 1465 4005 1473 4025
rect 1493 4006 1525 4025
rect 1546 4006 1581 4025
rect 1493 4005 1581 4006
rect 1601 4005 1609 4025
rect 1465 3997 1609 4005
rect 1465 3996 1501 3997
rect 1573 3996 1609 3997
rect 1675 4030 1712 4031
rect 1675 4029 1713 4030
rect 1675 4021 1739 4029
rect 1675 4001 1684 4021
rect 1704 4007 1739 4021
rect 1759 4007 1762 4027
rect 1704 4002 1762 4007
rect 1704 4001 1739 4002
rect 1144 3964 1181 3993
rect 1145 3962 1181 3964
rect 722 3952 758 3953
rect 570 3922 579 3942
rect 599 3922 607 3942
rect 570 3912 607 3922
rect 666 3942 814 3952
rect 914 3949 1010 3951
rect 666 3922 675 3942
rect 695 3922 785 3942
rect 805 3922 814 3942
rect 666 3913 814 3922
rect 872 3942 1010 3949
rect 872 3922 881 3942
rect 901 3922 1010 3942
rect 1145 3940 1336 3962
rect 1362 3961 1399 3993
rect 1675 3989 1739 4001
rect 1779 3963 1806 4141
rect 1638 3961 1806 3963
rect 1362 3935 1806 3961
rect 872 3913 1010 3922
rect 666 3912 703 3913
rect 163 3858 200 3861
rect 396 3859 437 3860
rect 288 3852 437 3859
rect 288 3832 347 3852
rect 367 3832 406 3852
rect 426 3832 437 3852
rect 288 3824 437 3832
rect 504 3855 661 3862
rect 504 3835 624 3855
rect 644 3835 661 3855
rect 504 3825 661 3835
rect 504 3824 539 3825
rect 504 3803 535 3824
rect 722 3803 758 3913
rect 777 3912 814 3913
rect 873 3912 910 3913
rect 833 3853 923 3859
rect 833 3833 842 3853
rect 862 3851 923 3853
rect 862 3833 887 3851
rect 833 3831 887 3833
rect 907 3831 923 3851
rect 833 3825 923 3831
rect 347 3802 384 3803
rect 160 3794 197 3796
rect 160 3786 202 3794
rect 160 3768 170 3786
rect 188 3768 202 3786
rect 160 3759 202 3768
rect 346 3793 384 3802
rect 346 3773 355 3793
rect 375 3773 384 3793
rect 346 3765 384 3773
rect 450 3797 535 3803
rect 565 3802 602 3803
rect 450 3777 458 3797
rect 478 3777 535 3797
rect 450 3769 535 3777
rect 564 3793 602 3802
rect 564 3773 573 3793
rect 593 3773 602 3793
rect 450 3768 486 3769
rect 564 3765 602 3773
rect 668 3801 812 3803
rect 668 3797 720 3801
rect 668 3777 676 3797
rect 696 3781 720 3797
rect 740 3797 812 3801
rect 740 3781 784 3797
rect 696 3777 784 3781
rect 804 3777 812 3797
rect 668 3769 812 3777
rect 668 3768 704 3769
rect 776 3768 812 3769
rect 878 3802 915 3803
rect 878 3801 916 3802
rect 878 3793 942 3801
rect 878 3773 887 3793
rect 907 3779 942 3793
rect 962 3779 965 3799
rect 907 3774 965 3779
rect 907 3773 942 3774
rect 161 3734 202 3759
rect 347 3734 384 3765
rect 565 3734 602 3765
rect 878 3761 942 3773
rect 982 3735 1009 3913
rect 161 3707 210 3734
rect 346 3708 395 3734
rect 564 3733 645 3734
rect 841 3733 1009 3735
rect 564 3708 1009 3733
rect 565 3707 1009 3708
rect 163 3674 210 3707
rect 566 3674 606 3707
rect 841 3706 1009 3707
rect 1472 3711 1512 3935
rect 1638 3934 1806 3935
rect 1472 3689 1480 3711
rect 1504 3689 1512 3711
rect 1472 3681 1512 3689
rect 163 3635 606 3674
rect 163 3592 210 3635
rect 566 3630 606 3635
rect 1231 3633 1418 3657
rect 1449 3638 1842 3658
rect 1862 3638 1865 3658
rect 1449 3633 1865 3638
rect 163 3574 173 3592
rect 191 3574 210 3592
rect 163 3570 210 3574
rect 164 3565 201 3570
rect 1231 3562 1268 3633
rect 1449 3632 1790 3633
rect 1383 3572 1414 3573
rect 1231 3542 1240 3562
rect 1260 3542 1268 3562
rect 1231 3532 1268 3542
rect 1327 3562 1414 3572
rect 1327 3542 1336 3562
rect 1356 3542 1414 3562
rect 1327 3533 1414 3542
rect 1327 3532 1364 3533
rect 152 3503 204 3505
rect 150 3499 583 3503
rect 150 3493 589 3499
rect 150 3475 171 3493
rect 189 3475 589 3493
rect 1383 3482 1414 3533
rect 1449 3562 1486 3632
rect 1752 3631 1789 3632
rect 1601 3572 1637 3573
rect 1449 3542 1458 3562
rect 1478 3542 1486 3562
rect 1449 3532 1486 3542
rect 1545 3562 1693 3572
rect 1793 3569 1889 3571
rect 1545 3542 1554 3562
rect 1574 3542 1664 3562
rect 1684 3542 1693 3562
rect 1545 3533 1693 3542
rect 1751 3562 1889 3569
rect 1751 3542 1760 3562
rect 1780 3542 1889 3562
rect 1751 3533 1889 3542
rect 1545 3532 1582 3533
rect 1275 3479 1316 3480
rect 150 3457 589 3475
rect 152 3268 204 3457
rect 550 3432 589 3457
rect 1167 3472 1316 3479
rect 1167 3452 1226 3472
rect 1246 3452 1285 3472
rect 1305 3452 1316 3472
rect 1167 3444 1316 3452
rect 1383 3475 1540 3482
rect 1383 3455 1503 3475
rect 1523 3455 1540 3475
rect 1383 3445 1540 3455
rect 1383 3444 1418 3445
rect 334 3407 521 3431
rect 550 3412 945 3432
rect 965 3412 968 3432
rect 1383 3423 1414 3444
rect 1601 3423 1637 3533
rect 1656 3532 1693 3533
rect 1752 3532 1789 3533
rect 1712 3473 1802 3479
rect 1712 3453 1721 3473
rect 1741 3471 1802 3473
rect 1741 3453 1766 3471
rect 1712 3451 1766 3453
rect 1786 3451 1802 3471
rect 1712 3445 1802 3451
rect 1226 3422 1263 3423
rect 550 3407 968 3412
rect 1225 3413 1263 3422
rect 334 3336 371 3407
rect 550 3406 893 3407
rect 550 3403 589 3406
rect 855 3405 892 3406
rect 486 3346 517 3347
rect 334 3316 343 3336
rect 363 3316 371 3336
rect 334 3306 371 3316
rect 430 3336 517 3346
rect 430 3316 439 3336
rect 459 3316 517 3336
rect 430 3307 517 3316
rect 430 3306 467 3307
rect 152 3250 168 3268
rect 186 3250 204 3268
rect 486 3256 517 3307
rect 552 3336 589 3403
rect 1225 3393 1234 3413
rect 1254 3393 1263 3413
rect 1225 3385 1263 3393
rect 1329 3417 1414 3423
rect 1444 3422 1481 3423
rect 1329 3397 1337 3417
rect 1357 3397 1414 3417
rect 1329 3389 1414 3397
rect 1443 3413 1481 3422
rect 1443 3393 1452 3413
rect 1472 3393 1481 3413
rect 1329 3388 1365 3389
rect 1443 3385 1481 3393
rect 1547 3418 1691 3423
rect 1547 3417 1609 3418
rect 1547 3397 1555 3417
rect 1575 3399 1609 3417
rect 1630 3417 1691 3418
rect 1630 3399 1663 3417
rect 1575 3397 1663 3399
rect 1683 3397 1691 3417
rect 1547 3389 1691 3397
rect 1547 3388 1583 3389
rect 1655 3388 1691 3389
rect 1757 3422 1794 3423
rect 1757 3421 1795 3422
rect 1757 3413 1821 3421
rect 1757 3393 1766 3413
rect 1786 3399 1821 3413
rect 1841 3399 1844 3419
rect 1786 3394 1844 3399
rect 1786 3393 1821 3394
rect 1226 3356 1263 3385
rect 1227 3354 1263 3356
rect 704 3346 740 3347
rect 552 3316 561 3336
rect 581 3316 589 3336
rect 552 3306 589 3316
rect 648 3336 796 3346
rect 896 3343 992 3345
rect 648 3316 657 3336
rect 677 3316 767 3336
rect 787 3316 796 3336
rect 648 3307 796 3316
rect 854 3336 992 3343
rect 854 3316 863 3336
rect 883 3316 992 3336
rect 1227 3332 1418 3354
rect 1444 3353 1481 3385
rect 1757 3381 1821 3393
rect 1861 3355 1888 3533
rect 1720 3353 1888 3355
rect 1444 3339 1888 3353
rect 1444 3327 1891 3339
rect 1487 3325 1520 3327
rect 854 3307 992 3316
rect 648 3306 685 3307
rect 378 3253 419 3254
rect 152 3232 204 3250
rect 270 3246 419 3253
rect 270 3226 329 3246
rect 349 3226 388 3246
rect 408 3226 419 3246
rect 270 3218 419 3226
rect 486 3249 643 3256
rect 486 3229 606 3249
rect 626 3229 643 3249
rect 486 3219 643 3229
rect 486 3218 521 3219
rect 486 3197 517 3218
rect 704 3197 740 3307
rect 759 3306 796 3307
rect 855 3306 892 3307
rect 815 3247 905 3253
rect 815 3227 824 3247
rect 844 3245 905 3247
rect 844 3227 869 3245
rect 815 3225 869 3227
rect 889 3225 905 3245
rect 815 3219 905 3225
rect 329 3196 366 3197
rect 328 3187 366 3196
rect 156 3169 196 3179
rect 156 3151 166 3169
rect 184 3151 196 3169
rect 328 3167 337 3187
rect 357 3167 366 3187
rect 328 3159 366 3167
rect 432 3191 517 3197
rect 547 3196 584 3197
rect 432 3171 440 3191
rect 460 3171 517 3191
rect 432 3163 517 3171
rect 546 3187 584 3196
rect 546 3167 555 3187
rect 575 3167 584 3187
rect 432 3162 468 3163
rect 546 3159 584 3167
rect 650 3191 794 3197
rect 650 3171 658 3191
rect 678 3171 711 3191
rect 731 3171 766 3191
rect 786 3171 794 3191
rect 650 3163 794 3171
rect 650 3162 686 3163
rect 758 3162 794 3163
rect 860 3196 897 3197
rect 860 3195 898 3196
rect 860 3187 924 3195
rect 860 3167 869 3187
rect 889 3173 924 3187
rect 944 3173 947 3193
rect 889 3168 947 3173
rect 889 3167 924 3168
rect 156 3095 196 3151
rect 329 3130 366 3159
rect 330 3128 366 3130
rect 330 3106 521 3128
rect 547 3127 584 3159
rect 860 3155 924 3167
rect 964 3129 991 3307
rect 1849 3282 1891 3327
rect 823 3127 991 3129
rect 547 3117 991 3127
rect 1132 3223 1319 3247
rect 1350 3228 1743 3248
rect 1763 3228 1766 3248
rect 1350 3223 1766 3228
rect 1132 3152 1169 3223
rect 1350 3222 1691 3223
rect 1284 3162 1315 3163
rect 1132 3132 1141 3152
rect 1161 3132 1169 3152
rect 1132 3122 1169 3132
rect 1228 3152 1315 3162
rect 1228 3132 1237 3152
rect 1257 3132 1315 3152
rect 1228 3123 1315 3132
rect 1228 3122 1265 3123
rect 153 3090 196 3095
rect 544 3101 991 3117
rect 544 3095 572 3101
rect 823 3100 991 3101
rect 153 3087 303 3090
rect 544 3087 571 3095
rect 153 3085 571 3087
rect 153 3067 162 3085
rect 180 3067 571 3085
rect 1284 3072 1315 3123
rect 1350 3152 1387 3222
rect 1653 3221 1690 3222
rect 1502 3162 1538 3163
rect 1350 3132 1359 3152
rect 1379 3132 1387 3152
rect 1350 3122 1387 3132
rect 1446 3152 1594 3162
rect 1694 3159 1790 3161
rect 1446 3132 1455 3152
rect 1475 3132 1565 3152
rect 1585 3132 1594 3152
rect 1446 3123 1594 3132
rect 1652 3152 1790 3159
rect 1652 3132 1661 3152
rect 1681 3132 1790 3152
rect 1652 3123 1790 3132
rect 1446 3122 1483 3123
rect 1176 3069 1217 3070
rect 153 3064 571 3067
rect 153 3058 196 3064
rect 156 3055 196 3058
rect 1071 3062 1217 3069
rect 553 3046 593 3047
rect 264 3029 593 3046
rect 1071 3042 1127 3062
rect 1147 3042 1186 3062
rect 1206 3042 1217 3062
rect 1071 3034 1217 3042
rect 1284 3065 1441 3072
rect 1284 3045 1404 3065
rect 1424 3045 1441 3065
rect 1284 3035 1441 3045
rect 1284 3034 1319 3035
rect 148 2986 191 2997
rect 148 2968 160 2986
rect 178 2968 191 2986
rect 148 2942 191 2968
rect 264 2942 291 3029
rect 553 3020 593 3029
rect 148 2921 291 2942
rect 335 2994 369 3010
rect 553 3000 946 3020
rect 966 3000 969 3020
rect 1284 3013 1315 3034
rect 1502 3013 1538 3123
rect 1557 3122 1594 3123
rect 1653 3122 1690 3123
rect 1613 3063 1703 3069
rect 1613 3043 1622 3063
rect 1642 3061 1703 3063
rect 1642 3043 1667 3061
rect 1613 3041 1667 3043
rect 1687 3041 1703 3061
rect 1613 3035 1703 3041
rect 1127 3012 1164 3013
rect 553 2995 969 3000
rect 1126 3003 1164 3012
rect 553 2994 894 2995
rect 335 2924 372 2994
rect 487 2934 518 2935
rect 148 2919 285 2921
rect 148 2877 191 2919
rect 335 2904 344 2924
rect 364 2904 372 2924
rect 335 2894 372 2904
rect 431 2924 518 2934
rect 431 2904 440 2924
rect 460 2904 518 2924
rect 431 2895 518 2904
rect 431 2894 468 2895
rect 146 2867 191 2877
rect 146 2849 155 2867
rect 173 2849 191 2867
rect 146 2843 191 2849
rect 487 2844 518 2895
rect 553 2924 590 2994
rect 856 2993 893 2994
rect 1126 2983 1135 3003
rect 1155 2983 1164 3003
rect 1126 2975 1164 2983
rect 1230 3007 1315 3013
rect 1345 3012 1382 3013
rect 1230 2987 1238 3007
rect 1258 2987 1315 3007
rect 1230 2979 1315 2987
rect 1344 3003 1382 3012
rect 1344 2983 1353 3003
rect 1373 2983 1382 3003
rect 1230 2978 1266 2979
rect 1344 2975 1382 2983
rect 1448 3007 1592 3013
rect 1448 2987 1456 3007
rect 1476 3004 1564 3007
rect 1476 2987 1511 3004
rect 1448 2986 1511 2987
rect 1530 2987 1564 3004
rect 1584 2987 1592 3007
rect 1530 2986 1592 2987
rect 1448 2979 1592 2986
rect 1448 2978 1484 2979
rect 1556 2978 1592 2979
rect 1658 3012 1695 3013
rect 1658 3011 1696 3012
rect 1718 3011 1745 3015
rect 1658 3009 1745 3011
rect 1658 3003 1722 3009
rect 1658 2983 1667 3003
rect 1687 2989 1722 3003
rect 1742 2989 1745 3009
rect 1687 2984 1745 2989
rect 1687 2983 1722 2984
rect 1127 2946 1164 2975
rect 1128 2944 1164 2946
rect 705 2934 741 2935
rect 553 2904 562 2924
rect 582 2904 590 2924
rect 553 2894 590 2904
rect 649 2924 797 2934
rect 897 2931 993 2933
rect 649 2904 658 2924
rect 678 2904 768 2924
rect 788 2904 797 2924
rect 649 2895 797 2904
rect 855 2924 993 2931
rect 855 2904 864 2924
rect 884 2904 993 2924
rect 1128 2922 1319 2944
rect 1345 2943 1382 2975
rect 1658 2971 1722 2983
rect 1762 2945 1789 3123
rect 1621 2943 1789 2945
rect 1345 2917 1789 2943
rect 855 2895 993 2904
rect 649 2894 686 2895
rect 146 2840 183 2843
rect 379 2841 420 2842
rect 271 2834 420 2841
rect 271 2814 330 2834
rect 350 2814 389 2834
rect 409 2814 420 2834
rect 271 2806 420 2814
rect 487 2837 644 2844
rect 487 2817 607 2837
rect 627 2817 644 2837
rect 487 2807 644 2817
rect 487 2806 522 2807
rect 487 2785 518 2806
rect 705 2785 741 2895
rect 760 2894 797 2895
rect 856 2894 893 2895
rect 816 2835 906 2841
rect 816 2815 825 2835
rect 845 2833 906 2835
rect 845 2815 870 2833
rect 816 2813 870 2815
rect 890 2813 906 2833
rect 816 2807 906 2813
rect 330 2784 367 2785
rect 142 2776 180 2778
rect 142 2768 185 2776
rect 142 2750 153 2768
rect 171 2750 185 2768
rect 142 2723 185 2750
rect 329 2775 367 2784
rect 329 2755 338 2775
rect 358 2755 367 2775
rect 329 2747 367 2755
rect 433 2779 518 2785
rect 548 2784 585 2785
rect 433 2759 441 2779
rect 461 2759 518 2779
rect 433 2751 518 2759
rect 547 2775 585 2784
rect 547 2755 556 2775
rect 576 2755 585 2775
rect 433 2750 469 2751
rect 547 2747 585 2755
rect 651 2783 795 2785
rect 651 2779 703 2783
rect 651 2759 659 2779
rect 679 2763 703 2779
rect 723 2779 795 2783
rect 723 2763 767 2779
rect 679 2759 767 2763
rect 787 2759 795 2779
rect 651 2751 795 2759
rect 651 2750 687 2751
rect 759 2750 795 2751
rect 861 2784 898 2785
rect 861 2783 899 2784
rect 861 2775 925 2783
rect 861 2755 870 2775
rect 890 2761 925 2775
rect 945 2761 948 2781
rect 890 2756 948 2761
rect 890 2755 925 2756
rect 143 2716 185 2723
rect 330 2716 367 2747
rect 548 2716 585 2747
rect 861 2743 925 2755
rect 965 2717 992 2895
rect 143 2676 188 2716
rect 330 2691 475 2716
rect 548 2715 628 2716
rect 824 2715 992 2717
rect 548 2699 992 2715
rect 332 2690 475 2691
rect 547 2689 992 2699
rect 143 2655 190 2676
rect 547 2655 588 2689
rect 824 2688 992 2689
rect 1455 2693 1495 2917
rect 1621 2916 1789 2917
rect 1853 2949 1886 3282
rect 1853 2941 1890 2949
rect 1853 2922 1861 2941
rect 1882 2922 1890 2941
rect 1853 2916 1890 2922
rect 1455 2671 1463 2693
rect 1487 2671 1495 2693
rect 1455 2663 1495 2671
rect 143 2625 588 2655
rect 1626 2638 1691 2639
rect 143 2622 566 2625
rect 143 2574 190 2622
rect 143 2556 153 2574
rect 171 2556 190 2574
rect 143 2552 190 2556
rect 1277 2613 1464 2637
rect 1495 2618 1888 2638
rect 1908 2618 1911 2638
rect 1495 2613 1911 2618
rect 144 2547 181 2552
rect 1277 2542 1314 2613
rect 1495 2612 1836 2613
rect 1429 2552 1460 2553
rect 1277 2522 1286 2542
rect 1306 2522 1314 2542
rect 1277 2512 1314 2522
rect 1373 2542 1460 2552
rect 1373 2522 1382 2542
rect 1402 2522 1460 2542
rect 1373 2513 1460 2522
rect 1373 2512 1410 2513
rect 132 2485 184 2487
rect 130 2481 563 2485
rect 130 2475 569 2481
rect 130 2457 151 2475
rect 169 2457 569 2475
rect 1429 2462 1460 2513
rect 1495 2542 1532 2612
rect 1798 2611 1835 2612
rect 1647 2552 1683 2553
rect 1495 2522 1504 2542
rect 1524 2522 1532 2542
rect 1495 2512 1532 2522
rect 1591 2542 1739 2552
rect 1839 2549 1935 2551
rect 1591 2522 1600 2542
rect 1620 2522 1710 2542
rect 1730 2522 1739 2542
rect 1591 2513 1739 2522
rect 1797 2542 1935 2549
rect 1797 2522 1806 2542
rect 1826 2522 1935 2542
rect 1797 2513 1935 2522
rect 1591 2512 1628 2513
rect 1321 2459 1362 2460
rect 130 2439 569 2457
rect 132 2250 184 2439
rect 530 2414 569 2439
rect 1213 2452 1362 2459
rect 1213 2432 1272 2452
rect 1292 2432 1331 2452
rect 1351 2432 1362 2452
rect 1213 2424 1362 2432
rect 1429 2455 1586 2462
rect 1429 2435 1549 2455
rect 1569 2435 1586 2455
rect 1429 2425 1586 2435
rect 1429 2424 1464 2425
rect 314 2389 501 2413
rect 530 2394 925 2414
rect 945 2394 948 2414
rect 1429 2403 1460 2424
rect 1647 2403 1683 2513
rect 1702 2512 1739 2513
rect 1798 2512 1835 2513
rect 1758 2453 1848 2459
rect 1758 2433 1767 2453
rect 1787 2451 1848 2453
rect 1787 2433 1812 2451
rect 1758 2431 1812 2433
rect 1832 2431 1848 2451
rect 1758 2425 1848 2431
rect 1272 2402 1309 2403
rect 530 2389 948 2394
rect 1271 2393 1309 2402
rect 314 2318 351 2389
rect 530 2388 873 2389
rect 530 2385 569 2388
rect 835 2387 872 2388
rect 466 2328 497 2329
rect 314 2298 323 2318
rect 343 2298 351 2318
rect 314 2288 351 2298
rect 410 2318 497 2328
rect 410 2298 419 2318
rect 439 2298 497 2318
rect 410 2289 497 2298
rect 410 2288 447 2289
rect 132 2232 148 2250
rect 166 2232 184 2250
rect 466 2238 497 2289
rect 532 2318 569 2385
rect 1271 2373 1280 2393
rect 1300 2373 1309 2393
rect 1271 2365 1309 2373
rect 1375 2397 1460 2403
rect 1490 2402 1527 2403
rect 1375 2377 1383 2397
rect 1403 2377 1460 2397
rect 1375 2369 1460 2377
rect 1489 2393 1527 2402
rect 1489 2373 1498 2393
rect 1518 2373 1527 2393
rect 1375 2368 1411 2369
rect 1489 2365 1527 2373
rect 1593 2401 1737 2403
rect 1593 2397 1653 2401
rect 1593 2377 1601 2397
rect 1621 2379 1653 2397
rect 1676 2397 1737 2401
rect 1676 2379 1709 2397
rect 1621 2377 1709 2379
rect 1729 2377 1737 2397
rect 1593 2369 1737 2377
rect 1593 2368 1629 2369
rect 1701 2368 1737 2369
rect 1803 2402 1840 2403
rect 1803 2401 1841 2402
rect 1803 2393 1867 2401
rect 1803 2373 1812 2393
rect 1832 2379 1867 2393
rect 1887 2379 1890 2399
rect 1832 2374 1890 2379
rect 1832 2373 1867 2374
rect 1272 2336 1309 2365
rect 1273 2334 1309 2336
rect 684 2328 720 2329
rect 532 2298 541 2318
rect 561 2298 569 2318
rect 532 2288 569 2298
rect 628 2318 776 2328
rect 876 2325 972 2327
rect 628 2298 637 2318
rect 657 2298 747 2318
rect 767 2298 776 2318
rect 628 2289 776 2298
rect 834 2318 972 2325
rect 834 2298 843 2318
rect 863 2298 972 2318
rect 1273 2312 1464 2334
rect 1490 2333 1527 2365
rect 1803 2361 1867 2373
rect 1490 2332 1765 2333
rect 1907 2332 1934 2513
rect 1490 2307 1934 2332
rect 2070 2338 2109 4153
rect 2411 4140 2444 4473
rect 2508 4505 2676 4506
rect 2802 4505 2842 4729
rect 3305 4733 3473 4734
rect 3714 4733 3749 4750
rect 4106 4740 4153 4751
rect 3305 4707 3749 4733
rect 3305 4705 3473 4707
rect 3669 4706 3749 4707
rect 3904 4706 3971 4732
rect 4110 4706 4153 4740
rect 3305 4527 3332 4705
rect 3372 4667 3436 4679
rect 3712 4675 3749 4706
rect 3930 4675 3967 4706
rect 4112 4681 4153 4706
rect 4544 4765 4585 4790
rect 4730 4765 4767 4796
rect 4948 4765 4985 4796
rect 5261 4792 5325 4804
rect 5365 4766 5392 4944
rect 4544 4731 4587 4765
rect 4726 4739 4793 4765
rect 4948 4764 5028 4765
rect 5224 4764 5392 4766
rect 4948 4738 5392 4764
rect 4544 4720 4591 4731
rect 4948 4721 4983 4738
rect 5224 4737 5392 4738
rect 5855 4742 5895 4966
rect 6021 4965 6189 4966
rect 6253 4998 6286 5331
rect 6588 5318 6627 7133
rect 6763 7139 7207 7164
rect 6763 6958 6790 7139
rect 6932 7138 7207 7139
rect 6830 7098 6894 7110
rect 7170 7106 7207 7138
rect 7233 7137 7424 7159
rect 7725 7153 7834 7173
rect 7854 7153 7863 7173
rect 7725 7146 7863 7153
rect 7921 7173 8069 7182
rect 7921 7153 7930 7173
rect 7950 7153 8040 7173
rect 8060 7153 8069 7173
rect 7725 7144 7821 7146
rect 7921 7143 8069 7153
rect 8128 7173 8165 7183
rect 8128 7153 8136 7173
rect 8156 7153 8165 7173
rect 7977 7142 8013 7143
rect 7388 7135 7424 7137
rect 7388 7106 7425 7135
rect 6830 7097 6865 7098
rect 6807 7092 6865 7097
rect 6807 7072 6810 7092
rect 6830 7078 6865 7092
rect 6885 7078 6894 7098
rect 6830 7070 6894 7078
rect 6856 7069 6894 7070
rect 6857 7068 6894 7069
rect 6960 7102 6996 7103
rect 7068 7102 7104 7103
rect 6960 7094 7104 7102
rect 6960 7074 6968 7094
rect 6988 7092 7076 7094
rect 6988 7074 7021 7092
rect 6960 7070 7021 7074
rect 7044 7074 7076 7092
rect 7096 7074 7104 7094
rect 7044 7070 7104 7074
rect 6960 7068 7104 7070
rect 7170 7098 7208 7106
rect 7286 7102 7322 7103
rect 7170 7078 7179 7098
rect 7199 7078 7208 7098
rect 7170 7069 7208 7078
rect 7237 7094 7322 7102
rect 7237 7074 7294 7094
rect 7314 7074 7322 7094
rect 7170 7068 7207 7069
rect 7237 7068 7322 7074
rect 7388 7098 7426 7106
rect 7388 7078 7397 7098
rect 7417 7078 7426 7098
rect 8128 7086 8165 7153
rect 8200 7182 8231 7233
rect 8513 7221 8531 7239
rect 8549 7221 8565 7239
rect 8250 7182 8287 7183
rect 8200 7173 8287 7182
rect 8200 7153 8258 7173
rect 8278 7153 8287 7173
rect 8200 7143 8287 7153
rect 8346 7173 8383 7183
rect 8346 7153 8354 7173
rect 8374 7153 8383 7173
rect 8200 7142 8231 7143
rect 7825 7083 7862 7084
rect 8128 7083 8167 7086
rect 7824 7082 8167 7083
rect 8346 7082 8383 7153
rect 7388 7069 7426 7078
rect 7749 7077 8167 7082
rect 7388 7068 7425 7069
rect 6849 7040 6939 7046
rect 6849 7020 6865 7040
rect 6885 7038 6939 7040
rect 6885 7020 6910 7038
rect 6849 7018 6910 7020
rect 6930 7018 6939 7038
rect 6849 7012 6939 7018
rect 6862 6958 6899 6959
rect 6958 6958 6995 6959
rect 7014 6958 7050 7068
rect 7237 7047 7268 7068
rect 7749 7057 7752 7077
rect 7772 7057 8167 7077
rect 8196 7058 8383 7082
rect 7233 7046 7268 7047
rect 7111 7036 7268 7046
rect 7111 7016 7128 7036
rect 7148 7016 7268 7036
rect 7111 7009 7268 7016
rect 7335 7039 7484 7047
rect 7335 7019 7346 7039
rect 7366 7019 7405 7039
rect 7425 7019 7484 7039
rect 7335 7012 7484 7019
rect 8128 7032 8167 7057
rect 8513 7032 8565 7221
rect 8970 7248 8980 7266
rect 8998 7248 9010 7266
rect 9142 7264 9151 7284
rect 9171 7264 9180 7284
rect 9142 7256 9180 7264
rect 9246 7288 9331 7294
rect 9361 7293 9398 7294
rect 9246 7268 9254 7288
rect 9274 7268 9331 7288
rect 9246 7260 9331 7268
rect 9360 7284 9398 7293
rect 9360 7264 9369 7284
rect 9389 7264 9398 7284
rect 9246 7259 9282 7260
rect 9360 7256 9398 7264
rect 9464 7288 9608 7294
rect 9464 7268 9472 7288
rect 9492 7268 9525 7288
rect 9545 7268 9580 7288
rect 9600 7268 9608 7288
rect 9464 7260 9608 7268
rect 9464 7259 9500 7260
rect 9572 7259 9608 7260
rect 9674 7293 9711 7294
rect 9674 7292 9712 7293
rect 9674 7284 9738 7292
rect 9674 7264 9683 7284
rect 9703 7270 9738 7284
rect 9758 7270 9761 7290
rect 9703 7265 9761 7270
rect 9703 7264 9738 7265
rect 8970 7192 9010 7248
rect 9143 7227 9180 7256
rect 9144 7225 9180 7227
rect 9144 7203 9335 7225
rect 9361 7224 9398 7256
rect 9674 7252 9738 7264
rect 9778 7226 9805 7404
rect 10663 7379 10705 7424
rect 9637 7224 9805 7226
rect 9361 7214 9805 7224
rect 9946 7320 10133 7344
rect 10164 7325 10557 7345
rect 10577 7325 10580 7345
rect 10164 7320 10580 7325
rect 9946 7249 9983 7320
rect 10164 7319 10505 7320
rect 10098 7259 10129 7260
rect 9946 7229 9955 7249
rect 9975 7229 9983 7249
rect 9946 7219 9983 7229
rect 10042 7249 10129 7259
rect 10042 7229 10051 7249
rect 10071 7229 10129 7249
rect 10042 7220 10129 7229
rect 10042 7219 10079 7220
rect 8967 7187 9010 7192
rect 9358 7198 9805 7214
rect 9358 7192 9386 7198
rect 9637 7197 9805 7198
rect 8967 7184 9117 7187
rect 9358 7184 9385 7192
rect 8967 7182 9385 7184
rect 8967 7164 8976 7182
rect 8994 7164 9385 7182
rect 10098 7169 10129 7220
rect 10164 7249 10201 7319
rect 10467 7318 10504 7319
rect 10316 7259 10352 7260
rect 10164 7229 10173 7249
rect 10193 7229 10201 7249
rect 10164 7219 10201 7229
rect 10260 7249 10408 7259
rect 10508 7256 10604 7258
rect 10260 7229 10269 7249
rect 10289 7229 10379 7249
rect 10399 7229 10408 7249
rect 10260 7220 10408 7229
rect 10466 7249 10604 7256
rect 10466 7229 10475 7249
rect 10495 7229 10604 7249
rect 10466 7220 10604 7229
rect 10260 7219 10297 7220
rect 9990 7166 10031 7167
rect 8967 7161 9385 7164
rect 8967 7155 9010 7161
rect 8970 7152 9010 7155
rect 9885 7159 10031 7166
rect 9367 7143 9407 7144
rect 9078 7126 9407 7143
rect 9885 7139 9941 7159
rect 9961 7139 10000 7159
rect 10020 7139 10031 7159
rect 9885 7131 10031 7139
rect 10098 7162 10255 7169
rect 10098 7142 10218 7162
rect 10238 7142 10255 7162
rect 10098 7132 10255 7142
rect 10098 7131 10133 7132
rect 8962 7083 9005 7094
rect 8962 7065 8974 7083
rect 8992 7065 9005 7083
rect 8962 7039 9005 7065
rect 9078 7039 9105 7126
rect 9367 7117 9407 7126
rect 8128 7014 8567 7032
rect 7335 7011 7376 7012
rect 7069 6958 7106 6959
rect 6762 6949 6900 6958
rect 6762 6929 6871 6949
rect 6891 6929 6900 6949
rect 6762 6922 6900 6929
rect 6958 6949 7106 6958
rect 6958 6929 6967 6949
rect 6987 6929 7077 6949
rect 7097 6929 7106 6949
rect 6762 6920 6858 6922
rect 6958 6919 7106 6929
rect 7165 6949 7202 6959
rect 7165 6929 7173 6949
rect 7193 6929 7202 6949
rect 7014 6918 7050 6919
rect 6862 6859 6899 6860
rect 7165 6859 7202 6929
rect 7237 6958 7268 7009
rect 8128 6996 8528 7014
rect 8546 6996 8567 7014
rect 8128 6990 8567 6996
rect 8134 6986 8567 6990
rect 8962 7018 9105 7039
rect 9149 7091 9183 7107
rect 9367 7097 9760 7117
rect 9780 7097 9783 7117
rect 10098 7110 10129 7131
rect 10316 7110 10352 7220
rect 10371 7219 10408 7220
rect 10467 7219 10504 7220
rect 10427 7160 10517 7166
rect 10427 7140 10436 7160
rect 10456 7158 10517 7160
rect 10456 7140 10481 7158
rect 10427 7138 10481 7140
rect 10501 7138 10517 7158
rect 10427 7132 10517 7138
rect 9941 7109 9978 7110
rect 9367 7092 9783 7097
rect 9940 7100 9978 7109
rect 9367 7091 9708 7092
rect 9149 7021 9186 7091
rect 9301 7031 9332 7032
rect 8962 7016 9099 7018
rect 8513 6984 8565 6986
rect 8962 6974 9005 7016
rect 9149 7001 9158 7021
rect 9178 7001 9186 7021
rect 9149 6991 9186 7001
rect 9245 7021 9332 7031
rect 9245 7001 9254 7021
rect 9274 7001 9332 7021
rect 9245 6992 9332 7001
rect 9245 6991 9282 6992
rect 8960 6964 9005 6974
rect 7287 6958 7324 6959
rect 7237 6949 7324 6958
rect 7237 6929 7295 6949
rect 7315 6929 7324 6949
rect 7237 6919 7324 6929
rect 7383 6949 7420 6959
rect 7383 6929 7391 6949
rect 7411 6929 7420 6949
rect 8960 6946 8969 6964
rect 8987 6946 9005 6964
rect 8960 6940 9005 6946
rect 9301 6941 9332 6992
rect 9367 7021 9404 7091
rect 9670 7090 9707 7091
rect 9940 7080 9949 7100
rect 9969 7080 9978 7100
rect 9940 7072 9978 7080
rect 10044 7104 10129 7110
rect 10159 7109 10196 7110
rect 10044 7084 10052 7104
rect 10072 7084 10129 7104
rect 10044 7076 10129 7084
rect 10158 7100 10196 7109
rect 10158 7080 10167 7100
rect 10187 7080 10196 7100
rect 10044 7075 10080 7076
rect 10158 7072 10196 7080
rect 10262 7104 10406 7110
rect 10262 7084 10270 7104
rect 10290 7101 10378 7104
rect 10290 7084 10325 7101
rect 10262 7083 10325 7084
rect 10344 7084 10378 7101
rect 10398 7084 10406 7104
rect 10344 7083 10406 7084
rect 10262 7076 10406 7083
rect 10262 7075 10298 7076
rect 10370 7075 10406 7076
rect 10472 7109 10509 7110
rect 10472 7108 10510 7109
rect 10532 7108 10559 7112
rect 10472 7106 10559 7108
rect 10472 7100 10536 7106
rect 10472 7080 10481 7100
rect 10501 7086 10536 7100
rect 10556 7086 10559 7106
rect 10501 7081 10559 7086
rect 10501 7080 10536 7081
rect 9941 7043 9978 7072
rect 9942 7041 9978 7043
rect 9519 7031 9555 7032
rect 9367 7001 9376 7021
rect 9396 7001 9404 7021
rect 9367 6991 9404 7001
rect 9463 7021 9611 7031
rect 9711 7028 9807 7030
rect 9463 7001 9472 7021
rect 9492 7001 9582 7021
rect 9602 7001 9611 7021
rect 9463 6992 9611 7001
rect 9669 7021 9807 7028
rect 9669 7001 9678 7021
rect 9698 7001 9807 7021
rect 9942 7019 10133 7041
rect 10159 7040 10196 7072
rect 10472 7068 10536 7080
rect 10576 7042 10603 7220
rect 10435 7040 10603 7042
rect 10159 7014 10603 7040
rect 9669 6992 9807 7001
rect 9463 6991 9500 6992
rect 8960 6937 8997 6940
rect 9193 6938 9234 6939
rect 7237 6918 7268 6919
rect 6861 6858 7202 6859
rect 7383 6858 7420 6929
rect 9085 6931 9234 6938
rect 8516 6919 8553 6924
rect 6786 6853 7202 6858
rect 6786 6833 6789 6853
rect 6809 6833 7202 6853
rect 7233 6834 7420 6858
rect 8507 6915 8554 6919
rect 8507 6897 8526 6915
rect 8544 6897 8554 6915
rect 9085 6911 9144 6931
rect 9164 6911 9203 6931
rect 9223 6911 9234 6931
rect 9085 6903 9234 6911
rect 9301 6934 9458 6941
rect 9301 6914 9421 6934
rect 9441 6914 9458 6934
rect 9301 6904 9458 6914
rect 9301 6903 9336 6904
rect 8507 6849 8554 6897
rect 9301 6882 9332 6903
rect 9519 6882 9555 6992
rect 9574 6991 9611 6992
rect 9670 6991 9707 6992
rect 9630 6932 9720 6938
rect 9630 6912 9639 6932
rect 9659 6930 9720 6932
rect 9659 6912 9684 6930
rect 9630 6910 9684 6912
rect 9704 6910 9720 6930
rect 9630 6904 9720 6910
rect 9144 6881 9181 6882
rect 8131 6846 8554 6849
rect 7006 6832 7071 6833
rect 8109 6816 8554 6846
rect 8956 6873 8994 6875
rect 8956 6865 8999 6873
rect 8956 6847 8967 6865
rect 8985 6847 8999 6865
rect 8956 6820 8999 6847
rect 9143 6872 9181 6881
rect 9143 6852 9152 6872
rect 9172 6852 9181 6872
rect 9143 6844 9181 6852
rect 9247 6876 9332 6882
rect 9362 6881 9399 6882
rect 9247 6856 9255 6876
rect 9275 6856 9332 6876
rect 9247 6848 9332 6856
rect 9361 6872 9399 6881
rect 9361 6852 9370 6872
rect 9390 6852 9399 6872
rect 9247 6847 9283 6848
rect 9361 6844 9399 6852
rect 9465 6880 9609 6882
rect 9465 6876 9517 6880
rect 9465 6856 9473 6876
rect 9493 6860 9517 6876
rect 9537 6876 9609 6880
rect 9537 6860 9581 6876
rect 9493 6856 9581 6860
rect 9601 6856 9609 6876
rect 9465 6848 9609 6856
rect 9465 6847 9501 6848
rect 9573 6847 9609 6848
rect 9675 6881 9712 6882
rect 9675 6880 9713 6881
rect 9675 6872 9739 6880
rect 9675 6852 9684 6872
rect 9704 6858 9739 6872
rect 9759 6858 9762 6878
rect 9704 6853 9762 6858
rect 9704 6852 9739 6853
rect 7202 6800 7242 6808
rect 7202 6778 7210 6800
rect 7234 6778 7242 6800
rect 6807 6549 6844 6555
rect 6807 6530 6815 6549
rect 6836 6530 6844 6549
rect 6807 6522 6844 6530
rect 6811 6189 6844 6522
rect 6908 6554 7076 6555
rect 7202 6554 7242 6778
rect 7705 6782 7873 6783
rect 8109 6782 8150 6816
rect 8507 6795 8554 6816
rect 7705 6772 8150 6782
rect 8222 6780 8365 6781
rect 7705 6756 8149 6772
rect 7705 6754 7873 6756
rect 8069 6755 8149 6756
rect 8222 6755 8367 6780
rect 8509 6755 8554 6795
rect 7705 6576 7732 6754
rect 7772 6716 7836 6728
rect 8112 6724 8149 6755
rect 8330 6724 8367 6755
rect 8512 6748 8554 6755
rect 8957 6813 8999 6820
rect 9144 6813 9181 6844
rect 9362 6813 9399 6844
rect 9675 6840 9739 6852
rect 9779 6814 9806 6992
rect 8957 6773 9002 6813
rect 9144 6788 9289 6813
rect 9362 6812 9442 6813
rect 9638 6812 9806 6814
rect 9362 6796 9806 6812
rect 9146 6787 9289 6788
rect 9361 6786 9806 6796
rect 8957 6752 9004 6773
rect 9361 6752 9402 6786
rect 9638 6785 9806 6786
rect 10269 6790 10309 7014
rect 10435 7013 10603 7014
rect 10667 7046 10700 7379
rect 11305 7378 11332 7556
rect 11372 7518 11436 7530
rect 11712 7526 11749 7558
rect 11775 7557 11966 7579
rect 12101 7577 12210 7597
rect 12230 7577 12239 7597
rect 12101 7570 12239 7577
rect 12297 7597 12445 7606
rect 12297 7577 12306 7597
rect 12326 7577 12416 7597
rect 12436 7577 12445 7597
rect 12101 7568 12197 7570
rect 12297 7567 12445 7577
rect 12504 7597 12541 7607
rect 12504 7577 12512 7597
rect 12532 7577 12541 7597
rect 12353 7566 12389 7567
rect 11930 7555 11966 7557
rect 11930 7526 11967 7555
rect 11372 7517 11407 7518
rect 11349 7512 11407 7517
rect 11349 7492 11352 7512
rect 11372 7498 11407 7512
rect 11427 7498 11436 7518
rect 11372 7490 11436 7498
rect 11398 7489 11436 7490
rect 11399 7488 11436 7489
rect 11502 7522 11538 7523
rect 11610 7522 11646 7523
rect 11502 7514 11646 7522
rect 11502 7494 11510 7514
rect 11530 7513 11618 7514
rect 11530 7494 11565 7513
rect 11586 7494 11618 7513
rect 11638 7494 11646 7514
rect 11502 7488 11646 7494
rect 11712 7518 11750 7526
rect 11828 7522 11864 7523
rect 11712 7498 11721 7518
rect 11741 7498 11750 7518
rect 11712 7489 11750 7498
rect 11779 7514 11864 7522
rect 11779 7494 11836 7514
rect 11856 7494 11864 7514
rect 11712 7488 11749 7489
rect 11779 7488 11864 7494
rect 11930 7518 11968 7526
rect 11930 7498 11939 7518
rect 11959 7498 11968 7518
rect 12201 7507 12238 7508
rect 12504 7507 12541 7577
rect 12576 7606 12607 7657
rect 12903 7652 12948 7658
rect 12903 7634 12921 7652
rect 12939 7634 12948 7652
rect 14409 7652 14418 7672
rect 14438 7652 14446 7672
rect 14409 7642 14446 7652
rect 14505 7672 14592 7682
rect 14505 7652 14514 7672
rect 14534 7652 14592 7672
rect 14505 7643 14592 7652
rect 14505 7642 14542 7643
rect 12903 7624 12948 7634
rect 12626 7606 12663 7607
rect 12576 7597 12663 7606
rect 12576 7577 12634 7597
rect 12654 7577 12663 7597
rect 12576 7567 12663 7577
rect 12722 7597 12759 7607
rect 12722 7577 12730 7597
rect 12750 7577 12759 7597
rect 12903 7582 12946 7624
rect 13330 7613 13382 7615
rect 12809 7580 12946 7582
rect 12576 7566 12607 7567
rect 12722 7507 12759 7577
rect 12200 7506 12541 7507
rect 11930 7489 11968 7498
rect 12125 7501 12541 7506
rect 11930 7488 11967 7489
rect 11391 7460 11481 7466
rect 11391 7440 11407 7460
rect 11427 7458 11481 7460
rect 11427 7440 11452 7458
rect 11391 7438 11452 7440
rect 11472 7438 11481 7458
rect 11391 7432 11481 7438
rect 11404 7378 11441 7379
rect 11500 7378 11537 7379
rect 11556 7378 11592 7488
rect 11779 7467 11810 7488
rect 12125 7481 12128 7501
rect 12148 7481 12541 7501
rect 12725 7491 12759 7507
rect 12803 7559 12946 7580
rect 13328 7609 13761 7613
rect 13328 7603 13767 7609
rect 13328 7585 13349 7603
rect 13367 7585 13767 7603
rect 14561 7592 14592 7643
rect 14627 7672 14664 7742
rect 14930 7741 14967 7742
rect 14779 7682 14815 7683
rect 14627 7652 14636 7672
rect 14656 7652 14664 7672
rect 14627 7642 14664 7652
rect 14723 7672 14871 7682
rect 14971 7679 15067 7681
rect 14723 7652 14732 7672
rect 14752 7652 14842 7672
rect 14862 7652 14871 7672
rect 14723 7643 14871 7652
rect 14929 7672 15067 7679
rect 14929 7652 14938 7672
rect 14958 7652 15067 7672
rect 14929 7643 15067 7652
rect 14723 7642 14760 7643
rect 14453 7589 14494 7590
rect 13328 7567 13767 7585
rect 12501 7472 12541 7481
rect 12803 7472 12830 7559
rect 12903 7533 12946 7559
rect 12903 7515 12916 7533
rect 12934 7515 12946 7533
rect 12903 7504 12946 7515
rect 11775 7466 11810 7467
rect 11653 7456 11810 7466
rect 11653 7436 11670 7456
rect 11690 7436 11810 7456
rect 11653 7429 11810 7436
rect 11877 7459 12026 7467
rect 11877 7439 11888 7459
rect 11908 7439 11947 7459
rect 11967 7439 12026 7459
rect 12501 7455 12830 7472
rect 12501 7454 12541 7455
rect 11877 7432 12026 7439
rect 12898 7443 12938 7446
rect 12898 7437 12941 7443
rect 12523 7434 12941 7437
rect 11877 7431 11918 7432
rect 11611 7378 11648 7379
rect 11304 7369 11442 7378
rect 11167 7359 11203 7365
rect 11167 7341 11172 7359
rect 11194 7341 11203 7359
rect 11167 7337 11203 7341
rect 11304 7349 11413 7369
rect 11433 7349 11442 7369
rect 11304 7342 11442 7349
rect 11500 7369 11648 7378
rect 11500 7349 11509 7369
rect 11529 7349 11619 7369
rect 11639 7349 11648 7369
rect 11304 7340 11400 7342
rect 11500 7339 11648 7349
rect 11707 7369 11744 7379
rect 11707 7349 11715 7369
rect 11735 7349 11744 7369
rect 11556 7338 11592 7339
rect 11170 7178 11203 7337
rect 11404 7279 11441 7280
rect 11707 7279 11744 7349
rect 11779 7378 11810 7429
rect 12523 7416 12914 7434
rect 12932 7416 12941 7434
rect 12523 7414 12941 7416
rect 12523 7406 12550 7414
rect 12791 7411 12941 7414
rect 12103 7400 12271 7401
rect 12522 7400 12550 7406
rect 12103 7384 12550 7400
rect 12898 7406 12941 7411
rect 11829 7378 11866 7379
rect 11779 7369 11866 7378
rect 11779 7349 11837 7369
rect 11857 7349 11866 7369
rect 11779 7339 11866 7349
rect 11925 7369 11962 7379
rect 11925 7349 11933 7369
rect 11953 7349 11962 7369
rect 11779 7338 11810 7339
rect 11403 7278 11744 7279
rect 11925 7278 11962 7349
rect 11328 7273 11744 7278
rect 11328 7253 11331 7273
rect 11351 7253 11744 7273
rect 11775 7254 11962 7278
rect 12103 7374 12547 7384
rect 12103 7372 12271 7374
rect 12103 7194 12130 7372
rect 12170 7334 12234 7346
rect 12510 7342 12547 7374
rect 12573 7373 12764 7395
rect 12728 7371 12764 7373
rect 12728 7342 12765 7371
rect 12898 7350 12938 7406
rect 12170 7333 12205 7334
rect 12147 7328 12205 7333
rect 12147 7308 12150 7328
rect 12170 7314 12205 7328
rect 12225 7314 12234 7334
rect 12170 7306 12234 7314
rect 12196 7305 12234 7306
rect 12197 7304 12234 7305
rect 12300 7338 12336 7339
rect 12408 7338 12444 7339
rect 12300 7330 12444 7338
rect 12300 7310 12308 7330
rect 12328 7310 12363 7330
rect 12383 7310 12416 7330
rect 12436 7310 12444 7330
rect 12300 7304 12444 7310
rect 12510 7334 12548 7342
rect 12626 7338 12662 7339
rect 12510 7314 12519 7334
rect 12539 7314 12548 7334
rect 12510 7305 12548 7314
rect 12577 7330 12662 7338
rect 12577 7310 12634 7330
rect 12654 7310 12662 7330
rect 12510 7304 12547 7305
rect 12577 7304 12662 7310
rect 12728 7334 12766 7342
rect 12728 7314 12737 7334
rect 12757 7314 12766 7334
rect 12898 7332 12910 7350
rect 12928 7332 12938 7350
rect 13330 7378 13382 7567
rect 13728 7542 13767 7567
rect 14345 7582 14494 7589
rect 14345 7562 14404 7582
rect 14424 7562 14463 7582
rect 14483 7562 14494 7582
rect 14345 7554 14494 7562
rect 14561 7585 14718 7592
rect 14561 7565 14681 7585
rect 14701 7565 14718 7585
rect 14561 7555 14718 7565
rect 14561 7554 14596 7555
rect 13512 7517 13699 7541
rect 13728 7522 14123 7542
rect 14143 7522 14146 7542
rect 14561 7533 14592 7554
rect 14779 7533 14815 7643
rect 14834 7642 14871 7643
rect 14930 7642 14967 7643
rect 14890 7583 14980 7589
rect 14890 7563 14899 7583
rect 14919 7581 14980 7583
rect 14919 7563 14944 7581
rect 14890 7561 14944 7563
rect 14964 7561 14980 7581
rect 14890 7555 14980 7561
rect 14404 7532 14441 7533
rect 13728 7517 14146 7522
rect 14403 7523 14441 7532
rect 13512 7446 13549 7517
rect 13728 7516 14071 7517
rect 13728 7513 13767 7516
rect 14033 7515 14070 7516
rect 13664 7456 13695 7457
rect 13512 7426 13521 7446
rect 13541 7426 13549 7446
rect 13512 7416 13549 7426
rect 13608 7446 13695 7456
rect 13608 7426 13617 7446
rect 13637 7426 13695 7446
rect 13608 7417 13695 7426
rect 13608 7416 13645 7417
rect 13330 7360 13346 7378
rect 13364 7360 13382 7378
rect 13664 7366 13695 7417
rect 13730 7446 13767 7513
rect 14403 7503 14412 7523
rect 14432 7503 14441 7523
rect 14403 7495 14441 7503
rect 14507 7527 14592 7533
rect 14622 7532 14659 7533
rect 14507 7507 14515 7527
rect 14535 7507 14592 7527
rect 14507 7499 14592 7507
rect 14621 7523 14659 7532
rect 14621 7503 14630 7523
rect 14650 7503 14659 7523
rect 14507 7498 14543 7499
rect 14621 7495 14659 7503
rect 14725 7528 14869 7533
rect 14725 7527 14787 7528
rect 14725 7507 14733 7527
rect 14753 7509 14787 7527
rect 14808 7527 14869 7528
rect 14808 7509 14841 7527
rect 14753 7507 14841 7509
rect 14861 7507 14869 7527
rect 14725 7499 14869 7507
rect 14725 7498 14761 7499
rect 14833 7498 14869 7499
rect 14935 7532 14972 7533
rect 14935 7531 14973 7532
rect 14935 7523 14999 7531
rect 14935 7503 14944 7523
rect 14964 7509 14999 7523
rect 15019 7509 15022 7529
rect 14964 7504 15022 7509
rect 14964 7503 14999 7504
rect 14404 7466 14441 7495
rect 14405 7464 14441 7466
rect 13882 7456 13918 7457
rect 13730 7426 13739 7446
rect 13759 7426 13767 7446
rect 13730 7416 13767 7426
rect 13826 7446 13974 7456
rect 14074 7453 14170 7455
rect 13826 7426 13835 7446
rect 13855 7426 13945 7446
rect 13965 7426 13974 7446
rect 13826 7417 13974 7426
rect 14032 7446 14170 7453
rect 14032 7426 14041 7446
rect 14061 7426 14170 7446
rect 14405 7442 14596 7464
rect 14622 7463 14659 7495
rect 14935 7491 14999 7503
rect 15039 7465 15066 7643
rect 14898 7463 15066 7465
rect 14622 7449 15066 7463
rect 15669 7597 15837 7598
rect 15963 7597 16003 7821
rect 16466 7825 16634 7826
rect 16869 7825 16909 7858
rect 17265 7825 17312 7858
rect 16466 7824 16910 7825
rect 16466 7799 16911 7824
rect 16466 7797 16634 7799
rect 16830 7798 16911 7799
rect 17080 7798 17129 7824
rect 17265 7798 17314 7825
rect 16466 7619 16493 7797
rect 16533 7759 16597 7771
rect 16873 7767 16910 7798
rect 17091 7767 17128 7798
rect 17273 7773 17314 7798
rect 16533 7758 16568 7759
rect 16510 7753 16568 7758
rect 16510 7733 16513 7753
rect 16533 7739 16568 7753
rect 16588 7739 16597 7759
rect 16533 7731 16597 7739
rect 16559 7730 16597 7731
rect 16560 7729 16597 7730
rect 16663 7763 16699 7764
rect 16771 7763 16807 7764
rect 16663 7755 16807 7763
rect 16663 7735 16671 7755
rect 16691 7751 16779 7755
rect 16691 7735 16735 7751
rect 16663 7731 16735 7735
rect 16755 7735 16779 7751
rect 16799 7735 16807 7755
rect 16755 7731 16807 7735
rect 16663 7729 16807 7731
rect 16873 7759 16911 7767
rect 16989 7763 17025 7764
rect 16873 7739 16882 7759
rect 16902 7739 16911 7759
rect 16873 7730 16911 7739
rect 16940 7755 17025 7763
rect 16940 7735 16997 7755
rect 17017 7735 17025 7755
rect 16873 7729 16910 7730
rect 16940 7729 17025 7735
rect 17091 7759 17129 7767
rect 17091 7739 17100 7759
rect 17120 7739 17129 7759
rect 17091 7730 17129 7739
rect 17273 7764 17315 7773
rect 17273 7746 17287 7764
rect 17305 7746 17315 7764
rect 17273 7738 17315 7746
rect 17278 7736 17315 7738
rect 17091 7729 17128 7730
rect 16552 7701 16642 7707
rect 16552 7681 16568 7701
rect 16588 7699 16642 7701
rect 16588 7681 16613 7699
rect 16552 7679 16613 7681
rect 16633 7679 16642 7699
rect 16552 7673 16642 7679
rect 16565 7619 16602 7620
rect 16661 7619 16698 7620
rect 16717 7619 16753 7729
rect 16940 7708 16971 7729
rect 16936 7707 16971 7708
rect 16814 7697 16971 7707
rect 16814 7677 16831 7697
rect 16851 7677 16971 7697
rect 16814 7670 16971 7677
rect 17038 7700 17187 7708
rect 17038 7680 17049 7700
rect 17069 7680 17108 7700
rect 17128 7680 17187 7700
rect 17038 7673 17187 7680
rect 17038 7672 17079 7673
rect 17275 7671 17312 7674
rect 16772 7619 16809 7620
rect 16465 7610 16603 7619
rect 15669 7571 16113 7597
rect 15669 7569 15837 7571
rect 14622 7437 15069 7449
rect 14665 7435 14698 7437
rect 14032 7417 14170 7426
rect 13826 7416 13863 7417
rect 13556 7363 13597 7364
rect 13330 7342 13382 7360
rect 13448 7356 13597 7363
rect 12898 7322 12938 7332
rect 13448 7336 13507 7356
rect 13527 7336 13566 7356
rect 13586 7336 13597 7356
rect 13448 7328 13597 7336
rect 13664 7359 13821 7366
rect 13664 7339 13784 7359
rect 13804 7339 13821 7359
rect 13664 7329 13821 7339
rect 13664 7328 13699 7329
rect 12728 7305 12766 7314
rect 13664 7307 13695 7328
rect 13882 7307 13918 7417
rect 13937 7416 13974 7417
rect 14033 7416 14070 7417
rect 13993 7357 14083 7363
rect 13993 7337 14002 7357
rect 14022 7355 14083 7357
rect 14022 7337 14047 7355
rect 13993 7335 14047 7337
rect 14067 7335 14083 7355
rect 13993 7329 14083 7335
rect 13507 7306 13544 7307
rect 12728 7304 12765 7305
rect 12189 7276 12279 7282
rect 12189 7256 12205 7276
rect 12225 7274 12279 7276
rect 12225 7256 12250 7274
rect 12189 7254 12250 7256
rect 12270 7254 12279 7274
rect 12189 7248 12279 7254
rect 12202 7194 12239 7195
rect 12298 7194 12335 7195
rect 12354 7194 12390 7304
rect 12577 7283 12608 7304
rect 13506 7297 13544 7306
rect 12573 7282 12608 7283
rect 12451 7272 12608 7282
rect 12451 7252 12468 7272
rect 12488 7252 12608 7272
rect 12451 7245 12608 7252
rect 12675 7275 12824 7283
rect 12675 7255 12686 7275
rect 12706 7255 12745 7275
rect 12765 7255 12824 7275
rect 13334 7279 13374 7289
rect 12675 7248 12824 7255
rect 12890 7251 12942 7269
rect 12675 7247 12716 7248
rect 12409 7194 12446 7195
rect 12102 7185 12240 7194
rect 11169 7177 11206 7178
rect 11140 7176 11308 7177
rect 11434 7176 11474 7178
rect 10965 7167 11004 7173
rect 10965 7145 10973 7167
rect 10997 7145 11004 7167
rect 10667 7038 10704 7046
rect 10667 7019 10675 7038
rect 10696 7019 10704 7038
rect 10667 7013 10704 7019
rect 10269 6768 10277 6790
rect 10301 6768 10309 6790
rect 10269 6760 10309 6768
rect 7772 6715 7807 6716
rect 7749 6710 7807 6715
rect 7749 6690 7752 6710
rect 7772 6696 7807 6710
rect 7827 6696 7836 6716
rect 7772 6688 7836 6696
rect 7798 6687 7836 6688
rect 7799 6686 7836 6687
rect 7902 6720 7938 6721
rect 8010 6720 8046 6721
rect 7902 6712 8046 6720
rect 7902 6692 7910 6712
rect 7930 6708 8018 6712
rect 7930 6692 7974 6708
rect 7902 6688 7974 6692
rect 7994 6692 8018 6708
rect 8038 6692 8046 6712
rect 7994 6688 8046 6692
rect 7902 6686 8046 6688
rect 8112 6716 8150 6724
rect 8228 6720 8264 6721
rect 8112 6696 8121 6716
rect 8141 6696 8150 6716
rect 8112 6687 8150 6696
rect 8179 6712 8264 6720
rect 8179 6692 8236 6712
rect 8256 6692 8264 6712
rect 8112 6686 8149 6687
rect 8179 6686 8264 6692
rect 8330 6716 8368 6724
rect 8330 6696 8339 6716
rect 8359 6696 8368 6716
rect 8330 6687 8368 6696
rect 8512 6721 8555 6748
rect 8512 6703 8526 6721
rect 8544 6703 8555 6721
rect 8512 6695 8555 6703
rect 8517 6693 8555 6695
rect 8957 6722 9402 6752
rect 10440 6735 10505 6736
rect 8957 6719 9380 6722
rect 8330 6686 8367 6687
rect 7791 6658 7881 6664
rect 7791 6638 7807 6658
rect 7827 6656 7881 6658
rect 7827 6638 7852 6656
rect 7791 6636 7852 6638
rect 7872 6636 7881 6656
rect 7791 6630 7881 6636
rect 7804 6576 7841 6577
rect 7900 6576 7937 6577
rect 7956 6576 7992 6686
rect 8179 6665 8210 6686
rect 8957 6671 9004 6719
rect 8175 6664 8210 6665
rect 8053 6654 8210 6664
rect 8053 6634 8070 6654
rect 8090 6634 8210 6654
rect 8053 6627 8210 6634
rect 8277 6657 8426 6665
rect 8277 6637 8288 6657
rect 8308 6637 8347 6657
rect 8367 6637 8426 6657
rect 8957 6653 8967 6671
rect 8985 6653 9004 6671
rect 8957 6649 9004 6653
rect 10091 6710 10278 6734
rect 10309 6715 10702 6735
rect 10722 6715 10725 6735
rect 10309 6710 10725 6715
rect 8958 6644 8995 6649
rect 8277 6630 8426 6637
rect 10091 6639 10128 6710
rect 10309 6709 10650 6710
rect 10243 6649 10274 6650
rect 8277 6629 8318 6630
rect 8514 6628 8551 6631
rect 8011 6576 8048 6577
rect 7704 6567 7842 6576
rect 6908 6528 7352 6554
rect 6908 6526 7076 6528
rect 6908 6348 6935 6526
rect 6975 6488 7039 6500
rect 7315 6496 7352 6528
rect 7378 6527 7569 6549
rect 7704 6547 7813 6567
rect 7833 6547 7842 6567
rect 7704 6540 7842 6547
rect 7900 6567 8048 6576
rect 7900 6547 7909 6567
rect 7929 6547 8019 6567
rect 8039 6547 8048 6567
rect 7704 6538 7800 6540
rect 7900 6537 8048 6547
rect 8107 6567 8144 6577
rect 8107 6547 8115 6567
rect 8135 6547 8144 6567
rect 7956 6536 7992 6537
rect 7533 6525 7569 6527
rect 7533 6496 7570 6525
rect 6975 6487 7010 6488
rect 6952 6482 7010 6487
rect 6952 6462 6955 6482
rect 6975 6468 7010 6482
rect 7030 6468 7039 6488
rect 6975 6462 7039 6468
rect 6952 6460 7039 6462
rect 6952 6456 6979 6460
rect 7001 6459 7039 6460
rect 7002 6458 7039 6459
rect 7105 6492 7141 6493
rect 7213 6492 7249 6493
rect 7105 6485 7249 6492
rect 7105 6484 7167 6485
rect 7105 6464 7113 6484
rect 7133 6467 7167 6484
rect 7186 6484 7249 6485
rect 7186 6467 7221 6484
rect 7133 6464 7221 6467
rect 7241 6464 7249 6484
rect 7105 6458 7249 6464
rect 7315 6488 7353 6496
rect 7431 6492 7467 6493
rect 7315 6468 7324 6488
rect 7344 6468 7353 6488
rect 7315 6459 7353 6468
rect 7382 6484 7467 6492
rect 7382 6464 7439 6484
rect 7459 6464 7467 6484
rect 7315 6458 7352 6459
rect 7382 6458 7467 6464
rect 7533 6488 7571 6496
rect 7533 6468 7542 6488
rect 7562 6468 7571 6488
rect 7804 6477 7841 6478
rect 8107 6477 8144 6547
rect 8179 6576 8210 6627
rect 8506 6622 8551 6628
rect 8506 6604 8524 6622
rect 8542 6604 8551 6622
rect 10091 6619 10100 6639
rect 10120 6619 10128 6639
rect 10091 6609 10128 6619
rect 10187 6639 10274 6649
rect 10187 6619 10196 6639
rect 10216 6619 10274 6639
rect 10187 6610 10274 6619
rect 10187 6609 10224 6610
rect 8506 6594 8551 6604
rect 8229 6576 8266 6577
rect 8179 6567 8266 6576
rect 8179 6547 8237 6567
rect 8257 6547 8266 6567
rect 8179 6537 8266 6547
rect 8325 6567 8362 6577
rect 8325 6547 8333 6567
rect 8353 6547 8362 6567
rect 8506 6552 8549 6594
rect 8946 6582 8998 6584
rect 8412 6550 8549 6552
rect 8179 6536 8210 6537
rect 8325 6477 8362 6547
rect 7803 6476 8144 6477
rect 7533 6459 7571 6468
rect 7728 6471 8144 6476
rect 7533 6458 7570 6459
rect 6994 6430 7084 6436
rect 6994 6410 7010 6430
rect 7030 6428 7084 6430
rect 7030 6410 7055 6428
rect 6994 6408 7055 6410
rect 7075 6408 7084 6428
rect 6994 6402 7084 6408
rect 7007 6348 7044 6349
rect 7103 6348 7140 6349
rect 7159 6348 7195 6458
rect 7382 6437 7413 6458
rect 7728 6451 7731 6471
rect 7751 6451 8144 6471
rect 8328 6461 8362 6477
rect 8406 6529 8549 6550
rect 8944 6578 9377 6582
rect 8944 6572 9383 6578
rect 8944 6554 8965 6572
rect 8983 6554 9383 6572
rect 10243 6559 10274 6610
rect 10309 6639 10346 6709
rect 10612 6708 10649 6709
rect 10461 6649 10497 6650
rect 10309 6619 10318 6639
rect 10338 6619 10346 6639
rect 10309 6609 10346 6619
rect 10405 6639 10553 6649
rect 10653 6646 10749 6648
rect 10405 6619 10414 6639
rect 10434 6619 10524 6639
rect 10544 6619 10553 6639
rect 10405 6610 10553 6619
rect 10611 6639 10749 6646
rect 10611 6619 10620 6639
rect 10640 6619 10749 6639
rect 10611 6610 10749 6619
rect 10405 6609 10442 6610
rect 10135 6556 10176 6557
rect 8944 6536 9383 6554
rect 8104 6442 8144 6451
rect 8406 6442 8433 6529
rect 8506 6503 8549 6529
rect 8506 6485 8519 6503
rect 8537 6485 8549 6503
rect 8506 6474 8549 6485
rect 7378 6436 7413 6437
rect 7256 6426 7413 6436
rect 7256 6406 7273 6426
rect 7293 6406 7413 6426
rect 7256 6399 7413 6406
rect 7480 6429 7626 6437
rect 7480 6409 7491 6429
rect 7511 6409 7550 6429
rect 7570 6409 7626 6429
rect 8104 6425 8433 6442
rect 8104 6424 8144 6425
rect 7480 6402 7626 6409
rect 8501 6413 8541 6416
rect 8501 6407 8544 6413
rect 8126 6404 8544 6407
rect 7480 6401 7521 6402
rect 7214 6348 7251 6349
rect 6907 6339 7045 6348
rect 6907 6319 7016 6339
rect 7036 6319 7045 6339
rect 6907 6312 7045 6319
rect 7103 6339 7251 6348
rect 7103 6319 7112 6339
rect 7132 6319 7222 6339
rect 7242 6319 7251 6339
rect 6907 6310 7003 6312
rect 7103 6309 7251 6319
rect 7310 6339 7347 6349
rect 7310 6319 7318 6339
rect 7338 6319 7347 6339
rect 7159 6308 7195 6309
rect 7007 6249 7044 6250
rect 7310 6249 7347 6319
rect 7382 6348 7413 6399
rect 8126 6386 8517 6404
rect 8535 6386 8544 6404
rect 8126 6384 8544 6386
rect 8126 6376 8153 6384
rect 8394 6381 8544 6384
rect 7706 6370 7874 6371
rect 8125 6370 8153 6376
rect 7706 6354 8153 6370
rect 8501 6376 8544 6381
rect 7432 6348 7469 6349
rect 7382 6339 7469 6348
rect 7382 6319 7440 6339
rect 7460 6319 7469 6339
rect 7382 6309 7469 6319
rect 7528 6339 7565 6349
rect 7528 6319 7536 6339
rect 7556 6319 7565 6339
rect 7382 6308 7413 6309
rect 7006 6248 7347 6249
rect 7528 6248 7565 6319
rect 6931 6243 7347 6248
rect 6931 6223 6934 6243
rect 6954 6223 7347 6243
rect 7378 6224 7565 6248
rect 7706 6344 8150 6354
rect 7706 6342 7874 6344
rect 6806 6144 6848 6189
rect 7706 6164 7733 6342
rect 7773 6304 7837 6316
rect 8113 6312 8150 6344
rect 8176 6343 8367 6365
rect 8331 6341 8367 6343
rect 8331 6312 8368 6341
rect 8501 6320 8541 6376
rect 7773 6303 7808 6304
rect 7750 6298 7808 6303
rect 7750 6278 7753 6298
rect 7773 6284 7808 6298
rect 7828 6284 7837 6304
rect 7773 6276 7837 6284
rect 7799 6275 7837 6276
rect 7800 6274 7837 6275
rect 7903 6308 7939 6309
rect 8011 6308 8047 6309
rect 7903 6300 8047 6308
rect 7903 6280 7911 6300
rect 7931 6280 7966 6300
rect 7986 6280 8019 6300
rect 8039 6280 8047 6300
rect 7903 6274 8047 6280
rect 8113 6304 8151 6312
rect 8229 6308 8265 6309
rect 8113 6284 8122 6304
rect 8142 6284 8151 6304
rect 8113 6275 8151 6284
rect 8180 6300 8265 6308
rect 8180 6280 8237 6300
rect 8257 6280 8265 6300
rect 8113 6274 8150 6275
rect 8180 6274 8265 6280
rect 8331 6304 8369 6312
rect 8331 6284 8340 6304
rect 8360 6284 8369 6304
rect 8501 6302 8513 6320
rect 8531 6302 8541 6320
rect 8946 6347 8998 6536
rect 9344 6511 9383 6536
rect 10027 6549 10176 6556
rect 10027 6529 10086 6549
rect 10106 6529 10145 6549
rect 10165 6529 10176 6549
rect 10027 6521 10176 6529
rect 10243 6552 10400 6559
rect 10243 6532 10363 6552
rect 10383 6532 10400 6552
rect 10243 6522 10400 6532
rect 10243 6521 10278 6522
rect 9128 6486 9315 6510
rect 9344 6491 9739 6511
rect 9759 6491 9762 6511
rect 10243 6500 10274 6521
rect 10461 6500 10497 6610
rect 10516 6609 10553 6610
rect 10612 6609 10649 6610
rect 10572 6550 10662 6556
rect 10572 6530 10581 6550
rect 10601 6548 10662 6550
rect 10601 6530 10626 6548
rect 10572 6528 10626 6530
rect 10646 6528 10662 6548
rect 10572 6522 10662 6528
rect 10086 6499 10123 6500
rect 9344 6486 9762 6491
rect 10085 6490 10123 6499
rect 9128 6415 9165 6486
rect 9344 6485 9687 6486
rect 9344 6482 9383 6485
rect 9649 6484 9686 6485
rect 9280 6425 9311 6426
rect 9128 6395 9137 6415
rect 9157 6395 9165 6415
rect 9128 6385 9165 6395
rect 9224 6415 9311 6425
rect 9224 6395 9233 6415
rect 9253 6395 9311 6415
rect 9224 6386 9311 6395
rect 9224 6385 9261 6386
rect 8946 6329 8962 6347
rect 8980 6329 8998 6347
rect 9280 6335 9311 6386
rect 9346 6415 9383 6482
rect 10085 6470 10094 6490
rect 10114 6470 10123 6490
rect 10085 6462 10123 6470
rect 10189 6494 10274 6500
rect 10304 6499 10341 6500
rect 10189 6474 10197 6494
rect 10217 6474 10274 6494
rect 10189 6466 10274 6474
rect 10303 6490 10341 6499
rect 10303 6470 10312 6490
rect 10332 6470 10341 6490
rect 10189 6465 10225 6466
rect 10303 6462 10341 6470
rect 10407 6494 10551 6500
rect 10407 6474 10415 6494
rect 10435 6493 10523 6494
rect 10435 6475 10470 6493
rect 10488 6475 10523 6493
rect 10435 6474 10523 6475
rect 10543 6474 10551 6494
rect 10407 6466 10551 6474
rect 10407 6465 10443 6466
rect 10515 6465 10551 6466
rect 10617 6499 10654 6500
rect 10617 6498 10655 6499
rect 10617 6490 10681 6498
rect 10617 6470 10626 6490
rect 10646 6476 10681 6490
rect 10701 6476 10704 6496
rect 10646 6471 10704 6476
rect 10646 6470 10681 6471
rect 10086 6433 10123 6462
rect 10087 6431 10123 6433
rect 9498 6425 9534 6426
rect 9346 6395 9355 6415
rect 9375 6395 9383 6415
rect 9346 6385 9383 6395
rect 9442 6415 9590 6425
rect 9690 6422 9786 6424
rect 9442 6395 9451 6415
rect 9471 6395 9561 6415
rect 9581 6395 9590 6415
rect 9442 6386 9590 6395
rect 9648 6415 9786 6422
rect 9648 6395 9657 6415
rect 9677 6395 9786 6415
rect 10087 6409 10278 6431
rect 10304 6430 10341 6462
rect 10617 6458 10681 6470
rect 10721 6434 10748 6610
rect 10667 6432 10748 6434
rect 10580 6430 10748 6432
rect 10304 6404 10748 6430
rect 10414 6402 10454 6404
rect 10580 6403 10748 6404
rect 9648 6386 9786 6395
rect 10689 6401 10748 6403
rect 9442 6385 9479 6386
rect 9172 6332 9213 6333
rect 8946 6311 8998 6329
rect 9064 6325 9213 6332
rect 8501 6292 8541 6302
rect 9064 6305 9123 6325
rect 9143 6305 9182 6325
rect 9202 6305 9213 6325
rect 9064 6297 9213 6305
rect 9280 6328 9437 6335
rect 9280 6308 9400 6328
rect 9420 6308 9437 6328
rect 9280 6298 9437 6308
rect 9280 6297 9315 6298
rect 8331 6275 8369 6284
rect 9280 6276 9311 6297
rect 9498 6276 9534 6386
rect 9553 6385 9590 6386
rect 9649 6385 9686 6386
rect 9609 6326 9699 6332
rect 9609 6306 9618 6326
rect 9638 6324 9699 6326
rect 9638 6306 9663 6324
rect 9609 6304 9663 6306
rect 9683 6304 9699 6324
rect 9609 6298 9699 6304
rect 9123 6275 9160 6276
rect 8331 6274 8368 6275
rect 7792 6246 7882 6252
rect 7792 6226 7808 6246
rect 7828 6244 7882 6246
rect 7828 6226 7853 6244
rect 7792 6224 7853 6226
rect 7873 6224 7882 6244
rect 7792 6218 7882 6224
rect 7805 6164 7842 6165
rect 7901 6164 7938 6165
rect 7957 6164 7993 6274
rect 8180 6253 8211 6274
rect 9122 6266 9160 6275
rect 8176 6252 8211 6253
rect 8054 6242 8211 6252
rect 8054 6222 8071 6242
rect 8091 6222 8211 6242
rect 8054 6215 8211 6222
rect 8278 6245 8427 6253
rect 8278 6225 8289 6245
rect 8309 6225 8348 6245
rect 8368 6225 8427 6245
rect 8950 6248 8990 6258
rect 8278 6218 8427 6225
rect 8493 6221 8545 6239
rect 8278 6217 8319 6218
rect 8012 6164 8049 6165
rect 7705 6155 7843 6164
rect 7177 6144 7210 6146
rect 6806 6132 7253 6144
rect 6809 6118 7253 6132
rect 6809 6116 6977 6118
rect 6809 5938 6836 6116
rect 6876 6078 6940 6090
rect 7216 6086 7253 6118
rect 7279 6117 7470 6139
rect 7705 6135 7814 6155
rect 7834 6135 7843 6155
rect 7705 6128 7843 6135
rect 7901 6155 8049 6164
rect 7901 6135 7910 6155
rect 7930 6135 8020 6155
rect 8040 6135 8049 6155
rect 7705 6126 7801 6128
rect 7901 6125 8049 6135
rect 8108 6155 8145 6165
rect 8108 6135 8116 6155
rect 8136 6135 8145 6155
rect 7957 6124 7993 6125
rect 7434 6115 7470 6117
rect 7434 6086 7471 6115
rect 6876 6077 6911 6078
rect 6853 6072 6911 6077
rect 6853 6052 6856 6072
rect 6876 6058 6911 6072
rect 6931 6058 6940 6078
rect 6876 6050 6940 6058
rect 6902 6049 6940 6050
rect 6903 6048 6940 6049
rect 7006 6082 7042 6083
rect 7114 6082 7150 6083
rect 7006 6074 7150 6082
rect 7006 6054 7014 6074
rect 7034 6072 7122 6074
rect 7034 6054 7067 6072
rect 7006 6053 7067 6054
rect 7088 6054 7122 6072
rect 7142 6054 7150 6074
rect 7088 6053 7150 6054
rect 7006 6048 7150 6053
rect 7216 6078 7254 6086
rect 7332 6082 7368 6083
rect 7216 6058 7225 6078
rect 7245 6058 7254 6078
rect 7216 6049 7254 6058
rect 7283 6074 7368 6082
rect 7283 6054 7340 6074
rect 7360 6054 7368 6074
rect 7216 6048 7253 6049
rect 7283 6048 7368 6054
rect 7434 6078 7472 6086
rect 7434 6058 7443 6078
rect 7463 6058 7472 6078
rect 8108 6068 8145 6135
rect 8180 6164 8211 6215
rect 8493 6203 8511 6221
rect 8529 6203 8545 6221
rect 8230 6164 8267 6165
rect 8180 6155 8267 6164
rect 8180 6135 8238 6155
rect 8258 6135 8267 6155
rect 8180 6125 8267 6135
rect 8326 6155 8363 6165
rect 8326 6135 8334 6155
rect 8354 6135 8363 6155
rect 8180 6124 8211 6125
rect 7805 6065 7842 6066
rect 8108 6065 8147 6068
rect 7804 6064 8147 6065
rect 8326 6064 8363 6135
rect 7434 6049 7472 6058
rect 7729 6059 8147 6064
rect 7434 6048 7471 6049
rect 6895 6020 6985 6026
rect 6895 6000 6911 6020
rect 6931 6018 6985 6020
rect 6931 6000 6956 6018
rect 6895 5998 6956 6000
rect 6976 5998 6985 6018
rect 6895 5992 6985 5998
rect 6908 5938 6945 5939
rect 7004 5938 7041 5939
rect 7060 5938 7096 6048
rect 7283 6027 7314 6048
rect 7729 6039 7732 6059
rect 7752 6039 8147 6059
rect 8176 6040 8363 6064
rect 7279 6026 7314 6027
rect 7157 6016 7314 6026
rect 7157 5996 7174 6016
rect 7194 5996 7314 6016
rect 7157 5989 7314 5996
rect 7381 6019 7530 6027
rect 7381 5999 7392 6019
rect 7412 5999 7451 6019
rect 7471 5999 7530 6019
rect 7381 5992 7530 5999
rect 8108 6014 8147 6039
rect 8493 6014 8545 6203
rect 8950 6230 8960 6248
rect 8978 6230 8990 6248
rect 9122 6246 9131 6266
rect 9151 6246 9160 6266
rect 9122 6238 9160 6246
rect 9226 6270 9311 6276
rect 9341 6275 9378 6276
rect 9226 6250 9234 6270
rect 9254 6250 9311 6270
rect 9226 6242 9311 6250
rect 9340 6266 9378 6275
rect 9340 6246 9349 6266
rect 9369 6246 9378 6266
rect 9226 6241 9262 6242
rect 9340 6238 9378 6246
rect 9444 6270 9588 6276
rect 9444 6250 9452 6270
rect 9472 6250 9505 6270
rect 9525 6250 9560 6270
rect 9580 6250 9588 6270
rect 9444 6242 9588 6250
rect 9444 6241 9480 6242
rect 9552 6241 9588 6242
rect 9654 6275 9691 6276
rect 9654 6274 9692 6275
rect 9654 6266 9718 6274
rect 9654 6246 9663 6266
rect 9683 6252 9718 6266
rect 9738 6252 9741 6272
rect 9683 6247 9741 6252
rect 9683 6246 9718 6247
rect 8950 6174 8990 6230
rect 9123 6209 9160 6238
rect 9124 6207 9160 6209
rect 9124 6185 9315 6207
rect 9341 6206 9378 6238
rect 9654 6234 9718 6246
rect 9758 6208 9785 6386
rect 10689 6383 10718 6401
rect 9617 6206 9785 6208
rect 9341 6196 9785 6206
rect 9926 6302 10113 6326
rect 10144 6307 10537 6327
rect 10557 6307 10560 6327
rect 10144 6302 10560 6307
rect 9926 6231 9963 6302
rect 10144 6301 10485 6302
rect 10078 6241 10109 6242
rect 9926 6211 9935 6231
rect 9955 6211 9963 6231
rect 9926 6201 9963 6211
rect 10022 6231 10109 6241
rect 10022 6211 10031 6231
rect 10051 6211 10109 6231
rect 10022 6202 10109 6211
rect 10022 6201 10059 6202
rect 8947 6169 8990 6174
rect 9338 6180 9785 6196
rect 9338 6174 9366 6180
rect 9617 6179 9785 6180
rect 8947 6166 9097 6169
rect 9338 6166 9365 6174
rect 8947 6164 9365 6166
rect 8947 6146 8956 6164
rect 8974 6146 9365 6164
rect 10078 6151 10109 6202
rect 10144 6231 10181 6301
rect 10447 6300 10484 6301
rect 10296 6241 10332 6242
rect 10144 6211 10153 6231
rect 10173 6211 10181 6231
rect 10144 6201 10181 6211
rect 10240 6231 10388 6241
rect 10488 6238 10584 6240
rect 10240 6211 10249 6231
rect 10269 6211 10359 6231
rect 10379 6211 10388 6231
rect 10240 6202 10388 6211
rect 10446 6231 10584 6238
rect 10446 6211 10455 6231
rect 10475 6211 10584 6231
rect 10446 6202 10584 6211
rect 10240 6201 10277 6202
rect 9970 6148 10011 6149
rect 8947 6143 9365 6146
rect 8947 6137 8990 6143
rect 8950 6134 8990 6137
rect 9862 6141 10011 6148
rect 9347 6125 9387 6126
rect 9058 6108 9387 6125
rect 9862 6121 9921 6141
rect 9941 6121 9980 6141
rect 10000 6121 10011 6141
rect 9862 6113 10011 6121
rect 10078 6144 10235 6151
rect 10078 6124 10198 6144
rect 10218 6124 10235 6144
rect 10078 6114 10235 6124
rect 10078 6113 10113 6114
rect 8942 6065 8985 6076
rect 8942 6047 8954 6065
rect 8972 6047 8985 6065
rect 8942 6021 8985 6047
rect 9058 6021 9085 6108
rect 9347 6099 9387 6108
rect 8108 5996 8547 6014
rect 7381 5991 7422 5992
rect 7115 5938 7152 5939
rect 6808 5929 6946 5938
rect 6808 5909 6917 5929
rect 6937 5909 6946 5929
rect 6808 5902 6946 5909
rect 7004 5929 7152 5938
rect 7004 5909 7013 5929
rect 7033 5909 7123 5929
rect 7143 5909 7152 5929
rect 6808 5900 6904 5902
rect 7004 5899 7152 5909
rect 7211 5929 7248 5939
rect 7211 5909 7219 5929
rect 7239 5909 7248 5929
rect 7060 5898 7096 5899
rect 6908 5839 6945 5840
rect 7211 5839 7248 5909
rect 7283 5938 7314 5989
rect 8108 5978 8508 5996
rect 8526 5978 8547 5996
rect 8108 5972 8547 5978
rect 8114 5968 8547 5972
rect 8942 6000 9085 6021
rect 9129 6073 9163 6089
rect 9347 6079 9740 6099
rect 9760 6079 9763 6099
rect 10078 6092 10109 6113
rect 10296 6092 10332 6202
rect 10351 6201 10388 6202
rect 10447 6201 10484 6202
rect 10407 6142 10497 6148
rect 10407 6122 10416 6142
rect 10436 6140 10497 6142
rect 10436 6122 10461 6140
rect 10407 6120 10461 6122
rect 10481 6120 10497 6140
rect 10407 6114 10497 6120
rect 9921 6091 9958 6092
rect 9347 6074 9763 6079
rect 9920 6082 9958 6091
rect 9347 6073 9688 6074
rect 9129 6003 9166 6073
rect 9281 6013 9312 6014
rect 8942 5998 9079 6000
rect 8493 5966 8545 5968
rect 8942 5956 8985 5998
rect 9129 5983 9138 6003
rect 9158 5983 9166 6003
rect 9129 5973 9166 5983
rect 9225 6003 9312 6013
rect 9225 5983 9234 6003
rect 9254 5983 9312 6003
rect 9225 5974 9312 5983
rect 9225 5973 9262 5974
rect 8940 5946 8985 5956
rect 7333 5938 7370 5939
rect 7283 5929 7370 5938
rect 7283 5909 7341 5929
rect 7361 5909 7370 5929
rect 7283 5899 7370 5909
rect 7429 5929 7466 5939
rect 7429 5909 7437 5929
rect 7457 5909 7466 5929
rect 8940 5928 8949 5946
rect 8967 5928 8985 5946
rect 8940 5922 8985 5928
rect 9281 5923 9312 5974
rect 9347 6003 9384 6073
rect 9650 6072 9687 6073
rect 9920 6062 9929 6082
rect 9949 6062 9958 6082
rect 9920 6054 9958 6062
rect 10024 6086 10109 6092
rect 10139 6091 10176 6092
rect 10024 6066 10032 6086
rect 10052 6066 10109 6086
rect 10024 6058 10109 6066
rect 10138 6082 10176 6091
rect 10138 6062 10147 6082
rect 10167 6062 10176 6082
rect 10024 6057 10060 6058
rect 10138 6054 10176 6062
rect 10242 6086 10386 6092
rect 10242 6066 10250 6086
rect 10270 6067 10302 6086
rect 10323 6067 10358 6086
rect 10270 6066 10358 6067
rect 10378 6066 10386 6086
rect 10242 6058 10386 6066
rect 10242 6057 10278 6058
rect 10350 6057 10386 6058
rect 10452 6091 10489 6092
rect 10452 6090 10490 6091
rect 10452 6082 10516 6090
rect 10452 6062 10461 6082
rect 10481 6068 10516 6082
rect 10536 6068 10539 6088
rect 10481 6063 10539 6068
rect 10481 6062 10516 6063
rect 9921 6025 9958 6054
rect 9922 6023 9958 6025
rect 9499 6013 9535 6014
rect 9347 5983 9356 6003
rect 9376 5983 9384 6003
rect 9347 5973 9384 5983
rect 9443 6003 9591 6013
rect 9691 6010 9787 6012
rect 9443 5983 9452 6003
rect 9472 5983 9562 6003
rect 9582 5983 9591 6003
rect 9443 5974 9591 5983
rect 9649 6003 9787 6010
rect 9649 5983 9658 6003
rect 9678 5983 9787 6003
rect 9922 6001 10113 6023
rect 10139 6022 10176 6054
rect 10452 6050 10516 6062
rect 10556 6024 10583 6202
rect 10415 6022 10583 6024
rect 10139 5996 10583 6022
rect 9649 5974 9787 5983
rect 9443 5973 9480 5974
rect 8940 5919 8977 5922
rect 9173 5920 9214 5921
rect 7283 5898 7314 5899
rect 6907 5838 7248 5839
rect 7429 5838 7466 5909
rect 9065 5913 9214 5920
rect 8496 5901 8533 5906
rect 8487 5897 8534 5901
rect 8487 5879 8506 5897
rect 8524 5879 8534 5897
rect 9065 5893 9124 5913
rect 9144 5893 9183 5913
rect 9203 5893 9214 5913
rect 9065 5885 9214 5893
rect 9281 5916 9438 5923
rect 9281 5896 9401 5916
rect 9421 5896 9438 5916
rect 9281 5886 9438 5896
rect 9281 5885 9316 5886
rect 6832 5833 7248 5838
rect 6832 5813 6835 5833
rect 6855 5813 7248 5833
rect 7279 5814 7466 5838
rect 8091 5836 8131 5841
rect 8487 5836 8534 5879
rect 9281 5864 9312 5885
rect 9499 5864 9535 5974
rect 9554 5973 9591 5974
rect 9650 5973 9687 5974
rect 9610 5914 9700 5920
rect 9610 5894 9619 5914
rect 9639 5912 9700 5914
rect 9639 5894 9664 5912
rect 9610 5892 9664 5894
rect 9684 5892 9700 5912
rect 9610 5886 9700 5892
rect 9124 5863 9161 5864
rect 8091 5797 8534 5836
rect 8937 5855 8974 5857
rect 8937 5847 8979 5855
rect 8937 5829 8947 5847
rect 8965 5829 8979 5847
rect 8937 5820 8979 5829
rect 9123 5854 9161 5863
rect 9123 5834 9132 5854
rect 9152 5834 9161 5854
rect 9123 5826 9161 5834
rect 9227 5858 9312 5864
rect 9342 5863 9379 5864
rect 9227 5838 9235 5858
rect 9255 5838 9312 5858
rect 9227 5830 9312 5838
rect 9341 5854 9379 5863
rect 9341 5834 9350 5854
rect 9370 5834 9379 5854
rect 9227 5829 9263 5830
rect 9341 5826 9379 5834
rect 9445 5862 9589 5864
rect 9445 5858 9497 5862
rect 9445 5838 9453 5858
rect 9473 5842 9497 5858
rect 9517 5858 9589 5862
rect 9517 5842 9561 5858
rect 9473 5838 9561 5842
rect 9581 5838 9589 5858
rect 9445 5830 9589 5838
rect 9445 5829 9481 5830
rect 9553 5829 9589 5830
rect 9655 5863 9692 5864
rect 9655 5862 9693 5863
rect 9655 5854 9719 5862
rect 9655 5834 9664 5854
rect 9684 5840 9719 5854
rect 9739 5840 9742 5860
rect 9684 5835 9742 5840
rect 9684 5834 9719 5835
rect 7185 5782 7225 5790
rect 7185 5760 7193 5782
rect 7217 5760 7225 5782
rect 6891 5536 7059 5537
rect 7185 5536 7225 5760
rect 7688 5764 7856 5765
rect 8091 5764 8131 5797
rect 8487 5764 8534 5797
rect 8938 5795 8979 5820
rect 9124 5795 9161 5826
rect 9342 5795 9379 5826
rect 9655 5822 9719 5834
rect 9759 5796 9786 5974
rect 8938 5768 8987 5795
rect 9123 5769 9172 5795
rect 9341 5794 9422 5795
rect 9618 5794 9786 5796
rect 9341 5769 9786 5794
rect 9342 5768 9786 5769
rect 7688 5763 8132 5764
rect 7688 5738 8133 5763
rect 7688 5736 7856 5738
rect 8052 5737 8133 5738
rect 8302 5737 8351 5763
rect 8487 5737 8536 5764
rect 7688 5558 7715 5736
rect 7755 5698 7819 5710
rect 8095 5706 8132 5737
rect 8313 5706 8350 5737
rect 8495 5712 8536 5737
rect 8940 5735 8987 5768
rect 9343 5735 9383 5768
rect 9618 5767 9786 5768
rect 10249 5772 10289 5996
rect 10415 5995 10583 5996
rect 10249 5750 10257 5772
rect 10281 5750 10289 5772
rect 10249 5742 10289 5750
rect 7755 5697 7790 5698
rect 7732 5692 7790 5697
rect 7732 5672 7735 5692
rect 7755 5678 7790 5692
rect 7810 5678 7819 5698
rect 7755 5670 7819 5678
rect 7781 5669 7819 5670
rect 7782 5668 7819 5669
rect 7885 5702 7921 5703
rect 7993 5702 8029 5703
rect 7885 5694 8029 5702
rect 7885 5674 7893 5694
rect 7913 5690 8001 5694
rect 7913 5674 7957 5690
rect 7885 5670 7957 5674
rect 7977 5674 8001 5690
rect 8021 5674 8029 5694
rect 7977 5670 8029 5674
rect 7885 5668 8029 5670
rect 8095 5698 8133 5706
rect 8211 5702 8247 5703
rect 8095 5678 8104 5698
rect 8124 5678 8133 5698
rect 8095 5669 8133 5678
rect 8162 5694 8247 5702
rect 8162 5674 8219 5694
rect 8239 5674 8247 5694
rect 8095 5668 8132 5669
rect 8162 5668 8247 5674
rect 8313 5698 8351 5706
rect 8313 5678 8322 5698
rect 8342 5678 8351 5698
rect 8313 5669 8351 5678
rect 8495 5703 8537 5712
rect 8495 5685 8509 5703
rect 8527 5685 8537 5703
rect 8495 5677 8537 5685
rect 8500 5675 8537 5677
rect 8940 5696 9383 5735
rect 8313 5668 8350 5669
rect 7774 5640 7864 5646
rect 7774 5620 7790 5640
rect 7810 5638 7864 5640
rect 7810 5620 7835 5638
rect 7774 5618 7835 5620
rect 7855 5618 7864 5638
rect 7774 5612 7864 5618
rect 7787 5558 7824 5559
rect 7883 5558 7920 5559
rect 7939 5558 7975 5668
rect 8162 5647 8193 5668
rect 8940 5653 8987 5696
rect 9343 5691 9383 5696
rect 10008 5694 10195 5718
rect 10226 5699 10619 5719
rect 10639 5699 10642 5719
rect 10226 5694 10642 5699
rect 8158 5646 8193 5647
rect 8036 5636 8193 5646
rect 8036 5616 8053 5636
rect 8073 5616 8193 5636
rect 8036 5609 8193 5616
rect 8260 5639 8409 5647
rect 8260 5619 8271 5639
rect 8291 5619 8330 5639
rect 8350 5619 8409 5639
rect 8940 5635 8950 5653
rect 8968 5635 8987 5653
rect 8940 5631 8987 5635
rect 8941 5626 8978 5631
rect 8260 5612 8409 5619
rect 10008 5623 10045 5694
rect 10226 5693 10567 5694
rect 10160 5633 10191 5634
rect 8260 5611 8301 5612
rect 8497 5610 8534 5613
rect 7994 5558 8031 5559
rect 7687 5549 7825 5558
rect 6891 5510 7335 5536
rect 6891 5508 7059 5510
rect 6891 5330 6918 5508
rect 6958 5470 7022 5482
rect 7298 5478 7335 5510
rect 7361 5509 7552 5531
rect 7687 5529 7796 5549
rect 7816 5529 7825 5549
rect 7687 5522 7825 5529
rect 7883 5549 8031 5558
rect 7883 5529 7892 5549
rect 7912 5529 8002 5549
rect 8022 5529 8031 5549
rect 7687 5520 7783 5522
rect 7883 5519 8031 5529
rect 8090 5549 8127 5559
rect 8090 5529 8098 5549
rect 8118 5529 8127 5549
rect 7939 5518 7975 5519
rect 7516 5507 7552 5509
rect 7516 5478 7553 5507
rect 6958 5469 6993 5470
rect 6935 5464 6993 5469
rect 6935 5444 6938 5464
rect 6958 5450 6993 5464
rect 7013 5450 7022 5470
rect 6958 5442 7022 5450
rect 6984 5441 7022 5442
rect 6985 5440 7022 5441
rect 7088 5474 7124 5475
rect 7196 5474 7232 5475
rect 7088 5466 7232 5474
rect 7088 5446 7096 5466
rect 7116 5465 7204 5466
rect 7116 5446 7151 5465
rect 7172 5446 7204 5465
rect 7224 5446 7232 5466
rect 7088 5440 7232 5446
rect 7298 5470 7336 5478
rect 7414 5474 7450 5475
rect 7298 5450 7307 5470
rect 7327 5450 7336 5470
rect 7298 5441 7336 5450
rect 7365 5466 7450 5474
rect 7365 5446 7422 5466
rect 7442 5446 7450 5466
rect 7298 5440 7335 5441
rect 7365 5440 7450 5446
rect 7516 5470 7554 5478
rect 7516 5450 7525 5470
rect 7545 5450 7554 5470
rect 7787 5459 7824 5460
rect 8090 5459 8127 5529
rect 8162 5558 8193 5609
rect 8489 5604 8534 5610
rect 8489 5586 8507 5604
rect 8525 5586 8534 5604
rect 10008 5603 10017 5623
rect 10037 5603 10045 5623
rect 10008 5593 10045 5603
rect 10104 5623 10191 5633
rect 10104 5603 10113 5623
rect 10133 5603 10191 5623
rect 10104 5594 10191 5603
rect 10104 5593 10141 5594
rect 8489 5576 8534 5586
rect 8212 5558 8249 5559
rect 8162 5549 8249 5558
rect 8162 5529 8220 5549
rect 8240 5529 8249 5549
rect 8162 5519 8249 5529
rect 8308 5549 8345 5559
rect 8308 5529 8316 5549
rect 8336 5529 8345 5549
rect 8489 5534 8532 5576
rect 8929 5564 8981 5566
rect 8395 5532 8532 5534
rect 8162 5518 8193 5519
rect 8308 5459 8345 5529
rect 7786 5458 8127 5459
rect 7516 5441 7554 5450
rect 7711 5453 8127 5458
rect 7516 5440 7553 5441
rect 6977 5412 7067 5418
rect 6977 5392 6993 5412
rect 7013 5410 7067 5412
rect 7013 5392 7038 5410
rect 6977 5390 7038 5392
rect 7058 5390 7067 5410
rect 6977 5384 7067 5390
rect 6990 5330 7027 5331
rect 7086 5330 7123 5331
rect 7142 5330 7178 5440
rect 7365 5419 7396 5440
rect 7711 5433 7714 5453
rect 7734 5433 8127 5453
rect 8311 5443 8345 5459
rect 8389 5511 8532 5532
rect 8927 5560 9360 5564
rect 8927 5554 9366 5560
rect 8927 5536 8948 5554
rect 8966 5536 9366 5554
rect 10160 5543 10191 5594
rect 10226 5623 10263 5693
rect 10529 5692 10566 5693
rect 10378 5633 10414 5634
rect 10226 5603 10235 5623
rect 10255 5603 10263 5623
rect 10226 5593 10263 5603
rect 10322 5623 10470 5633
rect 10570 5630 10666 5632
rect 10322 5603 10331 5623
rect 10351 5603 10441 5623
rect 10461 5603 10470 5623
rect 10322 5594 10470 5603
rect 10528 5623 10666 5630
rect 10528 5603 10537 5623
rect 10557 5603 10666 5623
rect 10528 5594 10666 5603
rect 10322 5593 10359 5594
rect 10052 5540 10093 5541
rect 8927 5518 9366 5536
rect 8087 5424 8127 5433
rect 8389 5424 8416 5511
rect 8489 5485 8532 5511
rect 8489 5467 8502 5485
rect 8520 5467 8532 5485
rect 8489 5456 8532 5467
rect 7361 5418 7396 5419
rect 7239 5408 7396 5418
rect 7239 5388 7256 5408
rect 7276 5388 7396 5408
rect 7239 5381 7396 5388
rect 7463 5411 7612 5419
rect 7463 5391 7474 5411
rect 7494 5391 7533 5411
rect 7553 5391 7612 5411
rect 8087 5407 8416 5424
rect 8087 5406 8127 5407
rect 7463 5384 7612 5391
rect 8484 5395 8524 5398
rect 8484 5389 8527 5395
rect 8109 5386 8527 5389
rect 7463 5383 7504 5384
rect 7197 5330 7234 5331
rect 6890 5321 7028 5330
rect 6588 5146 6628 5318
rect 6890 5301 6999 5321
rect 7019 5301 7028 5321
rect 6890 5294 7028 5301
rect 7086 5321 7234 5330
rect 7086 5301 7095 5321
rect 7115 5301 7205 5321
rect 7225 5301 7234 5321
rect 6890 5292 6986 5294
rect 7086 5291 7234 5301
rect 7293 5321 7330 5331
rect 7293 5301 7301 5321
rect 7321 5301 7330 5321
rect 7142 5290 7178 5291
rect 6990 5231 7027 5232
rect 7293 5231 7330 5301
rect 7365 5330 7396 5381
rect 8109 5368 8500 5386
rect 8518 5368 8527 5386
rect 8109 5366 8527 5368
rect 8109 5358 8136 5366
rect 8377 5363 8527 5366
rect 7689 5352 7857 5353
rect 8108 5352 8136 5358
rect 7689 5336 8136 5352
rect 8484 5358 8527 5363
rect 7415 5330 7452 5331
rect 7365 5321 7452 5330
rect 7365 5301 7423 5321
rect 7443 5301 7452 5321
rect 7365 5291 7452 5301
rect 7511 5321 7548 5331
rect 7511 5301 7519 5321
rect 7539 5301 7548 5321
rect 7365 5290 7396 5291
rect 6989 5230 7330 5231
rect 7511 5230 7548 5301
rect 6914 5225 7330 5230
rect 6914 5205 6917 5225
rect 6937 5205 7330 5225
rect 7361 5206 7548 5230
rect 7689 5326 8133 5336
rect 7689 5324 7857 5326
rect 7689 5146 7716 5324
rect 7756 5286 7820 5298
rect 8096 5294 8133 5326
rect 8159 5325 8350 5347
rect 8314 5323 8350 5325
rect 8314 5294 8351 5323
rect 8484 5302 8524 5358
rect 7756 5285 7791 5286
rect 7733 5280 7791 5285
rect 7733 5260 7736 5280
rect 7756 5266 7791 5280
rect 7811 5266 7820 5286
rect 7756 5258 7820 5266
rect 7782 5257 7820 5258
rect 7783 5256 7820 5257
rect 7886 5290 7922 5291
rect 7994 5290 8030 5291
rect 7886 5282 8030 5290
rect 7886 5262 7894 5282
rect 7914 5262 7949 5282
rect 7969 5262 8002 5282
rect 8022 5262 8030 5282
rect 7886 5256 8030 5262
rect 8096 5286 8134 5294
rect 8212 5290 8248 5291
rect 8096 5266 8105 5286
rect 8125 5266 8134 5286
rect 8096 5257 8134 5266
rect 8163 5282 8248 5290
rect 8163 5262 8220 5282
rect 8240 5262 8248 5282
rect 8096 5256 8133 5257
rect 8163 5256 8248 5262
rect 8314 5286 8352 5294
rect 8314 5266 8323 5286
rect 8343 5266 8352 5286
rect 8484 5284 8496 5302
rect 8514 5284 8524 5302
rect 8929 5329 8981 5518
rect 9327 5493 9366 5518
rect 9944 5533 10093 5540
rect 9944 5513 10003 5533
rect 10023 5513 10062 5533
rect 10082 5513 10093 5533
rect 9944 5505 10093 5513
rect 10160 5536 10317 5543
rect 10160 5516 10280 5536
rect 10300 5516 10317 5536
rect 10160 5506 10317 5516
rect 10160 5505 10195 5506
rect 9111 5468 9298 5492
rect 9327 5473 9722 5493
rect 9742 5473 9745 5493
rect 10160 5484 10191 5505
rect 10378 5484 10414 5594
rect 10433 5593 10470 5594
rect 10529 5593 10566 5594
rect 10489 5534 10579 5540
rect 10489 5514 10498 5534
rect 10518 5532 10579 5534
rect 10518 5514 10543 5532
rect 10489 5512 10543 5514
rect 10563 5512 10579 5532
rect 10489 5506 10579 5512
rect 10003 5483 10040 5484
rect 9327 5468 9745 5473
rect 10002 5474 10040 5483
rect 9111 5397 9148 5468
rect 9327 5467 9670 5468
rect 9327 5464 9366 5467
rect 9632 5466 9669 5467
rect 9263 5407 9294 5408
rect 9111 5377 9120 5397
rect 9140 5377 9148 5397
rect 9111 5367 9148 5377
rect 9207 5397 9294 5407
rect 9207 5377 9216 5397
rect 9236 5377 9294 5397
rect 9207 5368 9294 5377
rect 9207 5367 9244 5368
rect 8929 5311 8945 5329
rect 8963 5311 8981 5329
rect 9263 5317 9294 5368
rect 9329 5397 9366 5464
rect 10002 5454 10011 5474
rect 10031 5454 10040 5474
rect 10002 5446 10040 5454
rect 10106 5478 10191 5484
rect 10221 5483 10258 5484
rect 10106 5458 10114 5478
rect 10134 5458 10191 5478
rect 10106 5450 10191 5458
rect 10220 5474 10258 5483
rect 10220 5454 10229 5474
rect 10249 5454 10258 5474
rect 10106 5449 10142 5450
rect 10220 5446 10258 5454
rect 10324 5478 10468 5484
rect 10324 5458 10332 5478
rect 10352 5473 10440 5478
rect 10352 5458 10388 5473
rect 10324 5456 10388 5458
rect 10407 5458 10440 5473
rect 10460 5458 10468 5478
rect 10407 5456 10468 5458
rect 10324 5450 10468 5456
rect 10324 5449 10360 5450
rect 10432 5449 10468 5450
rect 10534 5483 10571 5484
rect 10534 5482 10572 5483
rect 10534 5474 10598 5482
rect 10534 5454 10543 5474
rect 10563 5460 10598 5474
rect 10618 5460 10621 5480
rect 10563 5455 10621 5460
rect 10563 5454 10598 5455
rect 10003 5417 10040 5446
rect 10004 5415 10040 5417
rect 9481 5407 9517 5408
rect 9329 5377 9338 5397
rect 9358 5377 9366 5397
rect 9329 5367 9366 5377
rect 9425 5397 9573 5407
rect 9673 5404 9769 5406
rect 9425 5377 9434 5397
rect 9454 5377 9544 5397
rect 9564 5377 9573 5397
rect 9425 5368 9573 5377
rect 9631 5397 9769 5404
rect 9631 5377 9640 5397
rect 9660 5377 9769 5397
rect 10004 5393 10195 5415
rect 10221 5414 10258 5446
rect 10534 5442 10598 5454
rect 10638 5416 10665 5594
rect 10497 5414 10665 5416
rect 10221 5400 10665 5414
rect 10689 5437 10717 6383
rect 10689 5407 10734 5437
rect 10221 5388 10668 5400
rect 10264 5386 10297 5388
rect 9631 5368 9769 5377
rect 9425 5367 9462 5368
rect 9155 5314 9196 5315
rect 8929 5293 8981 5311
rect 9047 5307 9196 5314
rect 8484 5274 8524 5284
rect 9047 5287 9106 5307
rect 9126 5287 9165 5307
rect 9185 5287 9196 5307
rect 9047 5279 9196 5287
rect 9263 5310 9420 5317
rect 9263 5290 9383 5310
rect 9403 5290 9420 5310
rect 9263 5280 9420 5290
rect 9263 5279 9298 5280
rect 8314 5257 8352 5266
rect 9263 5258 9294 5279
rect 9481 5258 9517 5368
rect 9536 5367 9573 5368
rect 9632 5367 9669 5368
rect 9592 5308 9682 5314
rect 9592 5288 9601 5308
rect 9621 5306 9682 5308
rect 9621 5288 9646 5306
rect 9592 5286 9646 5288
rect 9666 5286 9682 5306
rect 9592 5280 9682 5286
rect 9106 5257 9143 5258
rect 8314 5256 8351 5257
rect 7775 5228 7865 5234
rect 7775 5208 7791 5228
rect 7811 5226 7865 5228
rect 7811 5208 7836 5226
rect 7775 5206 7836 5208
rect 7856 5206 7865 5226
rect 7775 5200 7865 5206
rect 7788 5146 7825 5147
rect 7884 5146 7921 5147
rect 7940 5146 7976 5256
rect 8163 5235 8194 5256
rect 9105 5248 9143 5257
rect 8159 5234 8194 5235
rect 8037 5224 8194 5234
rect 8037 5204 8054 5224
rect 8074 5204 8194 5224
rect 8037 5197 8194 5204
rect 8261 5227 8410 5235
rect 8261 5207 8272 5227
rect 8292 5207 8331 5227
rect 8351 5207 8410 5227
rect 8933 5230 8973 5240
rect 8261 5200 8410 5207
rect 8476 5203 8528 5221
rect 8261 5199 8302 5200
rect 7995 5146 8032 5147
rect 6589 5131 6628 5146
rect 7688 5137 7826 5146
rect 6589 5130 6755 5131
rect 6881 5130 6921 5132
rect 6589 5104 7031 5130
rect 6589 5102 6755 5104
rect 6253 4990 6290 4998
rect 6253 4971 6261 4990
rect 6282 4971 6290 4990
rect 6253 4965 6290 4971
rect 6589 4924 6614 5102
rect 6654 5064 6718 5076
rect 6994 5072 7031 5104
rect 7057 5103 7248 5125
rect 7688 5117 7797 5137
rect 7817 5117 7826 5137
rect 7688 5110 7826 5117
rect 7884 5137 8032 5146
rect 7884 5117 7893 5137
rect 7913 5117 8003 5137
rect 8023 5117 8032 5137
rect 7688 5108 7784 5110
rect 7884 5107 8032 5117
rect 8091 5137 8128 5147
rect 8091 5117 8099 5137
rect 8119 5117 8128 5137
rect 7940 5106 7976 5107
rect 7212 5101 7248 5103
rect 7212 5072 7249 5101
rect 6654 5063 6689 5064
rect 6631 5058 6689 5063
rect 6631 5038 6634 5058
rect 6654 5044 6689 5058
rect 6709 5044 6718 5064
rect 6654 5036 6718 5044
rect 6680 5035 6718 5036
rect 6681 5034 6718 5035
rect 6784 5068 6820 5069
rect 6892 5068 6928 5069
rect 6784 5063 6928 5068
rect 6784 5060 6846 5063
rect 6784 5040 6792 5060
rect 6812 5040 6846 5060
rect 6784 5037 6846 5040
rect 6872 5060 6928 5063
rect 6872 5040 6900 5060
rect 6920 5040 6928 5060
rect 6872 5037 6928 5040
rect 6784 5034 6928 5037
rect 6994 5064 7032 5072
rect 7110 5068 7146 5069
rect 6994 5044 7003 5064
rect 7023 5044 7032 5064
rect 6994 5035 7032 5044
rect 7061 5060 7146 5068
rect 7061 5040 7118 5060
rect 7138 5040 7146 5060
rect 6994 5034 7031 5035
rect 7061 5034 7146 5040
rect 7212 5064 7250 5072
rect 7212 5044 7221 5064
rect 7241 5044 7250 5064
rect 8091 5050 8128 5117
rect 8163 5146 8194 5197
rect 8476 5185 8494 5203
rect 8512 5185 8528 5203
rect 8213 5146 8250 5147
rect 8163 5137 8250 5146
rect 8163 5117 8221 5137
rect 8241 5117 8250 5137
rect 8163 5107 8250 5117
rect 8309 5137 8346 5147
rect 8309 5117 8317 5137
rect 8337 5117 8346 5137
rect 8163 5106 8194 5107
rect 7788 5047 7825 5048
rect 8091 5047 8130 5050
rect 7787 5046 8130 5047
rect 8309 5046 8346 5117
rect 7212 5035 7250 5044
rect 7712 5041 8130 5046
rect 7212 5034 7249 5035
rect 6673 5006 6763 5012
rect 6673 4986 6689 5006
rect 6709 5004 6763 5006
rect 6709 4986 6734 5004
rect 6673 4984 6734 4986
rect 6754 4984 6763 5004
rect 6673 4978 6763 4984
rect 6686 4924 6723 4925
rect 6782 4924 6819 4925
rect 6838 4924 6874 5034
rect 7061 5013 7092 5034
rect 7712 5021 7715 5041
rect 7735 5021 8130 5041
rect 8159 5022 8346 5046
rect 7057 5012 7092 5013
rect 6935 5002 7092 5012
rect 6935 4982 6952 5002
rect 6972 4982 7092 5002
rect 6935 4975 7092 4982
rect 7159 5005 7308 5013
rect 7159 4985 7170 5005
rect 7190 4985 7229 5005
rect 7249 4985 7308 5005
rect 7159 4978 7308 4985
rect 8091 4996 8130 5021
rect 8476 4996 8528 5185
rect 8933 5212 8943 5230
rect 8961 5212 8973 5230
rect 9105 5228 9114 5248
rect 9134 5228 9143 5248
rect 9105 5220 9143 5228
rect 9209 5252 9294 5258
rect 9324 5257 9361 5258
rect 9209 5232 9217 5252
rect 9237 5232 9294 5252
rect 9209 5224 9294 5232
rect 9323 5248 9361 5257
rect 9323 5228 9332 5248
rect 9352 5228 9361 5248
rect 9209 5223 9245 5224
rect 9323 5220 9361 5228
rect 9427 5252 9571 5258
rect 9427 5232 9435 5252
rect 9455 5232 9488 5252
rect 9508 5232 9543 5252
rect 9563 5232 9571 5252
rect 9427 5224 9571 5232
rect 9427 5223 9463 5224
rect 9535 5223 9571 5224
rect 9637 5257 9674 5258
rect 9637 5256 9675 5257
rect 9637 5248 9701 5256
rect 9637 5228 9646 5248
rect 9666 5234 9701 5248
rect 9721 5234 9724 5254
rect 9666 5229 9724 5234
rect 9666 5228 9701 5229
rect 8933 5156 8973 5212
rect 9106 5191 9143 5220
rect 9107 5189 9143 5191
rect 9107 5167 9298 5189
rect 9324 5188 9361 5220
rect 9637 5216 9701 5228
rect 9741 5190 9768 5368
rect 10626 5343 10668 5388
rect 10689 5389 10700 5407
rect 10722 5389 10734 5407
rect 10689 5383 10734 5389
rect 10690 5382 10734 5383
rect 9600 5188 9768 5190
rect 9324 5178 9768 5188
rect 9909 5284 10096 5308
rect 10127 5289 10520 5309
rect 10540 5289 10543 5309
rect 10127 5284 10543 5289
rect 9909 5213 9946 5284
rect 10127 5283 10468 5284
rect 10061 5223 10092 5224
rect 9909 5193 9918 5213
rect 9938 5193 9946 5213
rect 9909 5183 9946 5193
rect 10005 5213 10092 5223
rect 10005 5193 10014 5213
rect 10034 5193 10092 5213
rect 10005 5184 10092 5193
rect 10005 5183 10042 5184
rect 8930 5151 8973 5156
rect 9321 5162 9768 5178
rect 9321 5156 9349 5162
rect 9600 5161 9768 5162
rect 8930 5148 9080 5151
rect 9321 5148 9348 5156
rect 8930 5146 9348 5148
rect 8930 5128 8939 5146
rect 8957 5128 9348 5146
rect 10061 5133 10092 5184
rect 10127 5213 10164 5283
rect 10430 5282 10467 5283
rect 10279 5223 10315 5224
rect 10127 5193 10136 5213
rect 10156 5193 10164 5213
rect 10127 5183 10164 5193
rect 10223 5213 10371 5223
rect 10471 5220 10567 5222
rect 10223 5193 10232 5213
rect 10252 5193 10342 5213
rect 10362 5193 10371 5213
rect 10223 5184 10371 5193
rect 10429 5213 10567 5220
rect 10429 5193 10438 5213
rect 10458 5193 10567 5213
rect 10429 5184 10567 5193
rect 10223 5183 10260 5184
rect 9953 5130 9994 5131
rect 8930 5125 9348 5128
rect 8930 5119 8973 5125
rect 8933 5116 8973 5119
rect 9848 5123 9994 5130
rect 9330 5107 9370 5108
rect 9041 5090 9370 5107
rect 9848 5103 9904 5123
rect 9924 5103 9963 5123
rect 9983 5103 9994 5123
rect 9848 5095 9994 5103
rect 10061 5126 10218 5133
rect 10061 5106 10181 5126
rect 10201 5106 10218 5126
rect 10061 5096 10218 5106
rect 10061 5095 10096 5096
rect 8925 5047 8968 5058
rect 8925 5029 8937 5047
rect 8955 5029 8968 5047
rect 8925 5003 8968 5029
rect 9041 5003 9068 5090
rect 9330 5081 9370 5090
rect 8091 4978 8530 4996
rect 7159 4977 7200 4978
rect 6893 4924 6930 4925
rect 6589 4915 6724 4924
rect 6589 4895 6695 4915
rect 6715 4895 6724 4915
rect 6589 4888 6724 4895
rect 6782 4915 6930 4924
rect 6782 4895 6791 4915
rect 6811 4895 6901 4915
rect 6921 4895 6930 4915
rect 6589 4886 6682 4888
rect 6782 4885 6930 4895
rect 6989 4915 7026 4925
rect 6989 4895 6997 4915
rect 7017 4895 7026 4915
rect 6838 4884 6874 4885
rect 6686 4825 6723 4826
rect 6989 4825 7026 4895
rect 7061 4924 7092 4975
rect 8091 4960 8491 4978
rect 8509 4960 8530 4978
rect 8091 4954 8530 4960
rect 8097 4950 8530 4954
rect 8925 4982 9068 5003
rect 9112 5055 9146 5071
rect 9330 5061 9723 5081
rect 9743 5061 9746 5081
rect 10061 5074 10092 5095
rect 10279 5074 10315 5184
rect 10334 5183 10371 5184
rect 10430 5183 10467 5184
rect 10390 5124 10480 5130
rect 10390 5104 10399 5124
rect 10419 5122 10480 5124
rect 10419 5104 10444 5122
rect 10390 5102 10444 5104
rect 10464 5102 10480 5122
rect 10390 5096 10480 5102
rect 9904 5073 9941 5074
rect 9330 5056 9746 5061
rect 9903 5064 9941 5073
rect 9330 5055 9671 5056
rect 9112 4985 9149 5055
rect 9264 4995 9295 4996
rect 8925 4980 9062 4982
rect 8476 4948 8528 4950
rect 8925 4938 8968 4980
rect 9112 4965 9121 4985
rect 9141 4965 9149 4985
rect 9112 4955 9149 4965
rect 9208 4985 9295 4995
rect 9208 4965 9217 4985
rect 9237 4965 9295 4985
rect 9208 4956 9295 4965
rect 9208 4955 9245 4956
rect 8923 4928 8968 4938
rect 7111 4924 7148 4925
rect 7061 4915 7148 4924
rect 7061 4895 7119 4915
rect 7139 4895 7148 4915
rect 7061 4885 7148 4895
rect 7207 4915 7244 4925
rect 7207 4895 7215 4915
rect 7235 4895 7244 4915
rect 8923 4910 8932 4928
rect 8950 4910 8968 4928
rect 8923 4904 8968 4910
rect 9264 4905 9295 4956
rect 9330 4985 9367 5055
rect 9633 5054 9670 5055
rect 9903 5044 9912 5064
rect 9932 5044 9941 5064
rect 9903 5036 9941 5044
rect 10007 5068 10092 5074
rect 10122 5073 10159 5074
rect 10007 5048 10015 5068
rect 10035 5048 10092 5068
rect 10007 5040 10092 5048
rect 10121 5064 10159 5073
rect 10121 5044 10130 5064
rect 10150 5044 10159 5064
rect 10007 5039 10043 5040
rect 10121 5036 10159 5044
rect 10225 5068 10369 5074
rect 10225 5048 10233 5068
rect 10253 5065 10341 5068
rect 10253 5048 10288 5065
rect 10225 5047 10288 5048
rect 10307 5048 10341 5065
rect 10361 5048 10369 5068
rect 10307 5047 10369 5048
rect 10225 5040 10369 5047
rect 10225 5039 10261 5040
rect 10333 5039 10369 5040
rect 10435 5073 10472 5074
rect 10435 5072 10473 5073
rect 10495 5072 10522 5076
rect 10435 5070 10522 5072
rect 10435 5064 10499 5070
rect 10435 5044 10444 5064
rect 10464 5050 10499 5064
rect 10519 5050 10522 5070
rect 10464 5045 10522 5050
rect 10464 5044 10499 5045
rect 9904 5007 9941 5036
rect 9905 5005 9941 5007
rect 9482 4995 9518 4996
rect 9330 4965 9339 4985
rect 9359 4965 9367 4985
rect 9330 4955 9367 4965
rect 9426 4985 9574 4995
rect 9674 4992 9770 4994
rect 9426 4965 9435 4985
rect 9455 4965 9545 4985
rect 9565 4965 9574 4985
rect 9426 4956 9574 4965
rect 9632 4985 9770 4992
rect 9632 4965 9641 4985
rect 9661 4965 9770 4985
rect 9905 4983 10096 5005
rect 10122 5004 10159 5036
rect 10435 5032 10499 5044
rect 10539 5006 10566 5184
rect 10398 5004 10566 5006
rect 10122 4978 10566 5004
rect 9632 4956 9770 4965
rect 9426 4955 9463 4956
rect 8923 4901 8960 4904
rect 9156 4902 9197 4903
rect 7061 4884 7092 4885
rect 6685 4824 7026 4825
rect 7207 4824 7244 4895
rect 9048 4895 9197 4902
rect 8479 4883 8516 4888
rect 6610 4819 7026 4824
rect 6610 4799 6613 4819
rect 6633 4799 7026 4819
rect 7057 4800 7244 4824
rect 8470 4879 8517 4883
rect 8470 4861 8489 4879
rect 8507 4861 8517 4879
rect 9048 4875 9107 4895
rect 9127 4875 9166 4895
rect 9186 4875 9197 4895
rect 9048 4867 9197 4875
rect 9264 4898 9421 4905
rect 9264 4878 9384 4898
rect 9404 4878 9421 4898
rect 9264 4868 9421 4878
rect 9264 4867 9299 4868
rect 8078 4802 8116 4803
rect 8470 4802 8517 4861
rect 9264 4846 9295 4867
rect 9482 4846 9518 4956
rect 9537 4955 9574 4956
rect 9633 4955 9670 4956
rect 9593 4896 9683 4902
rect 9593 4876 9602 4896
rect 9622 4894 9683 4896
rect 9622 4876 9647 4894
rect 9593 4874 9647 4876
rect 9667 4874 9683 4894
rect 9593 4868 9683 4874
rect 9107 4845 9144 4846
rect 8920 4837 8957 4839
rect 8920 4829 8962 4837
rect 8920 4811 8930 4829
rect 8948 4811 8962 4829
rect 8920 4802 8962 4811
rect 9106 4836 9144 4845
rect 9106 4816 9115 4836
rect 9135 4816 9144 4836
rect 9106 4808 9144 4816
rect 9210 4840 9295 4846
rect 9325 4845 9362 4846
rect 9210 4820 9218 4840
rect 9238 4820 9295 4840
rect 9210 4812 9295 4820
rect 9324 4836 9362 4845
rect 9324 4816 9333 4836
rect 9353 4816 9362 4836
rect 9210 4811 9246 4812
rect 9324 4808 9362 4816
rect 9428 4844 9572 4846
rect 9428 4840 9480 4844
rect 9428 4820 9436 4840
rect 9456 4824 9480 4840
rect 9500 4840 9572 4844
rect 9500 4824 9544 4840
rect 9456 4820 9544 4824
rect 9564 4820 9572 4840
rect 9428 4812 9572 4820
rect 9428 4811 9464 4812
rect 9536 4811 9572 4812
rect 9638 4845 9675 4846
rect 9638 4844 9676 4845
rect 9638 4836 9702 4844
rect 9638 4816 9647 4836
rect 9667 4822 9702 4836
rect 9722 4822 9725 4842
rect 9667 4817 9725 4822
rect 9667 4816 9702 4817
rect 6830 4798 6895 4799
rect 4945 4720 4983 4721
rect 4544 4682 4983 4720
rect 5855 4720 5863 4742
rect 5887 4720 5895 4742
rect 5855 4712 5895 4720
rect 7166 4764 7206 4772
rect 7166 4742 7174 4764
rect 7198 4742 7206 4764
rect 8078 4764 8517 4802
rect 8078 4763 8116 4764
rect 6166 4685 6231 4686
rect 3372 4666 3407 4667
rect 3349 4661 3407 4666
rect 3349 4641 3352 4661
rect 3372 4647 3407 4661
rect 3427 4647 3436 4667
rect 3372 4639 3436 4647
rect 3398 4638 3436 4639
rect 3399 4637 3436 4638
rect 3502 4671 3538 4672
rect 3610 4671 3646 4672
rect 3502 4663 3646 4671
rect 3502 4643 3510 4663
rect 3530 4659 3618 4663
rect 3530 4643 3574 4659
rect 3502 4639 3574 4643
rect 3594 4643 3618 4659
rect 3638 4643 3646 4663
rect 3594 4639 3646 4643
rect 3502 4637 3646 4639
rect 3712 4667 3750 4675
rect 3828 4671 3864 4672
rect 3712 4647 3721 4667
rect 3741 4647 3750 4667
rect 3712 4638 3750 4647
rect 3779 4663 3864 4671
rect 3779 4643 3836 4663
rect 3856 4643 3864 4663
rect 3712 4637 3749 4638
rect 3779 4637 3864 4643
rect 3930 4667 3968 4675
rect 3930 4647 3939 4667
rect 3959 4647 3968 4667
rect 3930 4638 3968 4647
rect 4112 4672 4154 4681
rect 4112 4654 4126 4672
rect 4144 4654 4154 4672
rect 4112 4646 4154 4654
rect 4117 4644 4154 4646
rect 3930 4637 3967 4638
rect 3391 4609 3481 4615
rect 3391 4589 3407 4609
rect 3427 4607 3481 4609
rect 3427 4589 3452 4607
rect 3391 4587 3452 4589
rect 3472 4587 3481 4607
rect 3391 4581 3481 4587
rect 3404 4527 3441 4528
rect 3500 4527 3537 4528
rect 3556 4527 3592 4637
rect 3779 4616 3810 4637
rect 4544 4623 4591 4682
rect 4945 4681 4983 4682
rect 3775 4615 3810 4616
rect 3653 4605 3810 4615
rect 3653 4585 3670 4605
rect 3690 4585 3810 4605
rect 3653 4578 3810 4585
rect 3877 4608 4026 4616
rect 3877 4588 3888 4608
rect 3908 4588 3947 4608
rect 3967 4588 4026 4608
rect 4544 4605 4554 4623
rect 4572 4605 4591 4623
rect 4544 4601 4591 4605
rect 5817 4660 6004 4684
rect 6035 4665 6428 4685
rect 6448 4665 6451 4685
rect 6035 4660 6451 4665
rect 4545 4596 4582 4601
rect 3877 4581 4026 4588
rect 5817 4589 5854 4660
rect 6035 4659 6376 4660
rect 5969 4599 6000 4600
rect 3877 4580 3918 4581
rect 4114 4579 4151 4582
rect 3611 4527 3648 4528
rect 3304 4518 3442 4527
rect 2508 4479 2952 4505
rect 2508 4477 2676 4479
rect 2508 4299 2535 4477
rect 2575 4439 2639 4451
rect 2915 4447 2952 4479
rect 2978 4478 3169 4500
rect 3304 4498 3413 4518
rect 3433 4498 3442 4518
rect 3304 4491 3442 4498
rect 3500 4518 3648 4527
rect 3500 4498 3509 4518
rect 3529 4498 3619 4518
rect 3639 4498 3648 4518
rect 3304 4489 3400 4491
rect 3500 4488 3648 4498
rect 3707 4518 3744 4528
rect 3707 4498 3715 4518
rect 3735 4498 3744 4518
rect 3556 4487 3592 4488
rect 3133 4476 3169 4478
rect 3133 4447 3170 4476
rect 2575 4438 2610 4439
rect 2552 4433 2610 4438
rect 2552 4413 2555 4433
rect 2575 4419 2610 4433
rect 2630 4419 2639 4439
rect 2575 4413 2639 4419
rect 2552 4411 2639 4413
rect 2552 4407 2579 4411
rect 2601 4410 2639 4411
rect 2602 4409 2639 4410
rect 2705 4443 2741 4444
rect 2813 4443 2849 4444
rect 2705 4436 2849 4443
rect 2705 4435 2767 4436
rect 2705 4415 2713 4435
rect 2733 4418 2767 4435
rect 2786 4435 2849 4436
rect 2786 4418 2821 4435
rect 2733 4415 2821 4418
rect 2841 4415 2849 4435
rect 2705 4409 2849 4415
rect 2915 4439 2953 4447
rect 3031 4443 3067 4444
rect 2915 4419 2924 4439
rect 2944 4419 2953 4439
rect 2915 4410 2953 4419
rect 2982 4435 3067 4443
rect 2982 4415 3039 4435
rect 3059 4415 3067 4435
rect 2915 4409 2952 4410
rect 2982 4409 3067 4415
rect 3133 4439 3171 4447
rect 3133 4419 3142 4439
rect 3162 4419 3171 4439
rect 3404 4428 3441 4429
rect 3707 4428 3744 4498
rect 3779 4527 3810 4578
rect 4106 4573 4151 4579
rect 4106 4555 4124 4573
rect 4142 4555 4151 4573
rect 5817 4569 5826 4589
rect 5846 4569 5854 4589
rect 5817 4559 5854 4569
rect 5913 4589 6000 4599
rect 5913 4569 5922 4589
rect 5942 4569 6000 4589
rect 5913 4560 6000 4569
rect 5913 4559 5950 4560
rect 4106 4545 4151 4555
rect 3829 4527 3866 4528
rect 3779 4518 3866 4527
rect 3779 4498 3837 4518
rect 3857 4498 3866 4518
rect 3779 4488 3866 4498
rect 3925 4518 3962 4528
rect 3925 4498 3933 4518
rect 3953 4498 3962 4518
rect 4106 4503 4149 4545
rect 4533 4534 4585 4536
rect 4012 4501 4149 4503
rect 3779 4487 3810 4488
rect 3925 4428 3962 4498
rect 3403 4427 3744 4428
rect 3133 4410 3171 4419
rect 3328 4422 3744 4427
rect 3133 4409 3170 4410
rect 2594 4381 2684 4387
rect 2594 4361 2610 4381
rect 2630 4379 2684 4381
rect 2630 4361 2655 4379
rect 2594 4359 2655 4361
rect 2675 4359 2684 4379
rect 2594 4353 2684 4359
rect 2607 4299 2644 4300
rect 2703 4299 2740 4300
rect 2759 4299 2795 4409
rect 2982 4388 3013 4409
rect 3328 4402 3331 4422
rect 3351 4402 3744 4422
rect 3928 4412 3962 4428
rect 4006 4480 4149 4501
rect 4531 4530 4964 4534
rect 4531 4524 4970 4530
rect 4531 4506 4552 4524
rect 4570 4506 4970 4524
rect 5969 4509 6000 4560
rect 6035 4589 6072 4659
rect 6338 4658 6375 4659
rect 6187 4599 6223 4600
rect 6035 4569 6044 4589
rect 6064 4569 6072 4589
rect 6035 4559 6072 4569
rect 6131 4589 6279 4599
rect 6379 4596 6475 4598
rect 6131 4569 6140 4589
rect 6160 4569 6250 4589
rect 6270 4569 6279 4589
rect 6131 4560 6279 4569
rect 6337 4589 6475 4596
rect 6337 4569 6346 4589
rect 6366 4569 6475 4589
rect 6337 4560 6475 4569
rect 6131 4559 6168 4560
rect 5861 4506 5902 4507
rect 4531 4488 4970 4506
rect 3704 4393 3744 4402
rect 4006 4393 4033 4480
rect 4106 4454 4149 4480
rect 4106 4436 4119 4454
rect 4137 4436 4149 4454
rect 4106 4425 4149 4436
rect 2978 4387 3013 4388
rect 2856 4377 3013 4387
rect 2856 4357 2873 4377
rect 2893 4357 3013 4377
rect 2856 4350 3013 4357
rect 3080 4380 3226 4388
rect 3080 4360 3091 4380
rect 3111 4360 3150 4380
rect 3170 4360 3226 4380
rect 3704 4376 4033 4393
rect 3704 4375 3744 4376
rect 3080 4353 3226 4360
rect 4101 4364 4141 4367
rect 4101 4358 4144 4364
rect 3726 4355 4144 4358
rect 3080 4352 3121 4353
rect 2814 4299 2851 4300
rect 2507 4290 2645 4299
rect 2507 4270 2616 4290
rect 2636 4270 2645 4290
rect 2507 4263 2645 4270
rect 2703 4290 2851 4299
rect 2703 4270 2712 4290
rect 2732 4270 2822 4290
rect 2842 4270 2851 4290
rect 2507 4261 2603 4263
rect 2703 4260 2851 4270
rect 2910 4290 2947 4300
rect 2910 4270 2918 4290
rect 2938 4270 2947 4290
rect 2759 4259 2795 4260
rect 2607 4200 2644 4201
rect 2910 4200 2947 4270
rect 2982 4299 3013 4350
rect 3726 4337 4117 4355
rect 4135 4337 4144 4355
rect 3726 4335 4144 4337
rect 3726 4327 3753 4335
rect 3994 4332 4144 4335
rect 3306 4321 3474 4322
rect 3725 4321 3753 4327
rect 3306 4305 3753 4321
rect 4101 4327 4144 4332
rect 3032 4299 3069 4300
rect 2982 4290 3069 4299
rect 2982 4270 3040 4290
rect 3060 4270 3069 4290
rect 2982 4260 3069 4270
rect 3128 4290 3165 4300
rect 3128 4270 3136 4290
rect 3156 4270 3165 4290
rect 2982 4259 3013 4260
rect 2606 4199 2947 4200
rect 3128 4199 3165 4270
rect 2531 4194 2947 4199
rect 2531 4174 2534 4194
rect 2554 4174 2947 4194
rect 2978 4175 3165 4199
rect 3306 4295 3750 4305
rect 3306 4293 3474 4295
rect 2340 4100 2384 4101
rect 2340 4094 2385 4100
rect 2340 4076 2352 4094
rect 2374 4076 2385 4094
rect 2406 4095 2448 4140
rect 3306 4115 3333 4293
rect 3373 4255 3437 4267
rect 3713 4263 3750 4295
rect 3776 4294 3967 4316
rect 3931 4292 3967 4294
rect 3931 4263 3968 4292
rect 4101 4271 4141 4327
rect 3373 4254 3408 4255
rect 3350 4249 3408 4254
rect 3350 4229 3353 4249
rect 3373 4235 3408 4249
rect 3428 4235 3437 4255
rect 3373 4227 3437 4235
rect 3399 4226 3437 4227
rect 3400 4225 3437 4226
rect 3503 4259 3539 4260
rect 3611 4259 3647 4260
rect 3503 4251 3647 4259
rect 3503 4231 3511 4251
rect 3531 4231 3566 4251
rect 3586 4231 3619 4251
rect 3639 4231 3647 4251
rect 3503 4225 3647 4231
rect 3713 4255 3751 4263
rect 3829 4259 3865 4260
rect 3713 4235 3722 4255
rect 3742 4235 3751 4255
rect 3713 4226 3751 4235
rect 3780 4251 3865 4259
rect 3780 4231 3837 4251
rect 3857 4231 3865 4251
rect 3713 4225 3750 4226
rect 3780 4225 3865 4231
rect 3931 4255 3969 4263
rect 3931 4235 3940 4255
rect 3960 4235 3969 4255
rect 4101 4253 4113 4271
rect 4131 4253 4141 4271
rect 4533 4299 4585 4488
rect 4931 4463 4970 4488
rect 5753 4499 5902 4506
rect 5753 4479 5812 4499
rect 5832 4479 5871 4499
rect 5891 4479 5902 4499
rect 5753 4471 5902 4479
rect 5969 4502 6126 4509
rect 5969 4482 6089 4502
rect 6109 4482 6126 4502
rect 5969 4472 6126 4482
rect 5969 4471 6004 4472
rect 4715 4438 4902 4462
rect 4931 4443 5326 4463
rect 5346 4443 5349 4463
rect 5969 4450 6000 4471
rect 6187 4450 6223 4560
rect 6242 4559 6279 4560
rect 6338 4559 6375 4560
rect 6298 4500 6388 4506
rect 6298 4480 6307 4500
rect 6327 4498 6388 4500
rect 6327 4480 6352 4498
rect 6298 4478 6352 4480
rect 6372 4478 6388 4498
rect 6298 4472 6388 4478
rect 5812 4449 5849 4450
rect 4931 4438 5349 4443
rect 5811 4440 5849 4449
rect 4715 4367 4752 4438
rect 4931 4437 5274 4438
rect 4931 4434 4970 4437
rect 5236 4436 5273 4437
rect 4867 4377 4898 4378
rect 4715 4347 4724 4367
rect 4744 4347 4752 4367
rect 4715 4337 4752 4347
rect 4811 4367 4898 4377
rect 4811 4347 4820 4367
rect 4840 4347 4898 4367
rect 4811 4338 4898 4347
rect 4811 4337 4848 4338
rect 4533 4281 4549 4299
rect 4567 4281 4585 4299
rect 4867 4287 4898 4338
rect 4933 4367 4970 4434
rect 5811 4420 5820 4440
rect 5840 4420 5849 4440
rect 5811 4412 5849 4420
rect 5915 4444 6000 4450
rect 6030 4449 6067 4450
rect 5915 4424 5923 4444
rect 5943 4424 6000 4444
rect 5915 4416 6000 4424
rect 6029 4440 6067 4449
rect 6029 4420 6038 4440
rect 6058 4420 6067 4440
rect 5915 4415 5951 4416
rect 6029 4412 6067 4420
rect 6133 4444 6277 4450
rect 6133 4424 6141 4444
rect 6161 4438 6249 4444
rect 6161 4424 6190 4438
rect 6133 4416 6190 4424
rect 6133 4415 6169 4416
rect 6213 4424 6249 4438
rect 6269 4424 6277 4444
rect 6213 4416 6277 4424
rect 6241 4415 6277 4416
rect 6343 4449 6380 4450
rect 6343 4448 6381 4449
rect 6343 4440 6407 4448
rect 6343 4420 6352 4440
rect 6372 4426 6407 4440
rect 6427 4426 6430 4446
rect 6372 4421 6430 4426
rect 6372 4420 6407 4421
rect 5812 4383 5849 4412
rect 5813 4381 5849 4383
rect 5085 4377 5121 4378
rect 4933 4347 4942 4367
rect 4962 4347 4970 4367
rect 4933 4337 4970 4347
rect 5029 4367 5177 4377
rect 5277 4374 5373 4376
rect 5029 4347 5038 4367
rect 5058 4347 5148 4367
rect 5168 4347 5177 4367
rect 5029 4338 5177 4347
rect 5235 4367 5373 4374
rect 5235 4347 5244 4367
rect 5264 4347 5373 4367
rect 5813 4359 6004 4381
rect 6030 4380 6067 4412
rect 6343 4408 6407 4420
rect 6447 4382 6474 4560
rect 6771 4513 6808 4519
rect 6771 4494 6779 4513
rect 6800 4494 6808 4513
rect 6771 4486 6808 4494
rect 6306 4380 6474 4382
rect 6030 4354 6474 4380
rect 6140 4352 6180 4354
rect 6306 4353 6474 4354
rect 5235 4338 5373 4347
rect 6433 4348 6474 4353
rect 5029 4337 5066 4338
rect 4759 4284 4800 4285
rect 4533 4263 4585 4281
rect 4651 4277 4800 4284
rect 4101 4243 4141 4253
rect 4651 4257 4710 4277
rect 4730 4257 4769 4277
rect 4789 4257 4800 4277
rect 4651 4249 4800 4257
rect 4867 4280 5024 4287
rect 4867 4260 4987 4280
rect 5007 4260 5024 4280
rect 4867 4250 5024 4260
rect 4867 4249 4902 4250
rect 3931 4226 3969 4235
rect 4867 4228 4898 4249
rect 5085 4228 5121 4338
rect 5140 4337 5177 4338
rect 5236 4337 5273 4338
rect 5196 4278 5286 4284
rect 5196 4258 5205 4278
rect 5225 4276 5286 4278
rect 5225 4258 5250 4276
rect 5196 4256 5250 4258
rect 5270 4256 5286 4276
rect 5196 4250 5286 4256
rect 4710 4227 4747 4228
rect 3931 4225 3968 4226
rect 3392 4197 3482 4203
rect 3392 4177 3408 4197
rect 3428 4195 3482 4197
rect 3428 4177 3453 4195
rect 3392 4175 3453 4177
rect 3473 4175 3482 4195
rect 3392 4169 3482 4175
rect 3405 4115 3442 4116
rect 3501 4115 3538 4116
rect 3557 4115 3593 4225
rect 3780 4204 3811 4225
rect 4709 4218 4747 4227
rect 3776 4203 3811 4204
rect 3654 4193 3811 4203
rect 3654 4173 3671 4193
rect 3691 4173 3811 4193
rect 3654 4166 3811 4173
rect 3878 4196 4027 4204
rect 3878 4176 3889 4196
rect 3909 4176 3948 4196
rect 3968 4176 4027 4196
rect 4537 4200 4577 4210
rect 3878 4169 4027 4176
rect 4093 4172 4145 4190
rect 3878 4168 3919 4169
rect 3612 4115 3649 4116
rect 3305 4106 3443 4115
rect 2777 4095 2810 4097
rect 2406 4083 2853 4095
rect 2340 4046 2385 4076
rect 2357 3100 2385 4046
rect 2409 4069 2853 4083
rect 2409 4067 2577 4069
rect 2409 3889 2436 4067
rect 2476 4029 2540 4041
rect 2816 4037 2853 4069
rect 2879 4068 3070 4090
rect 3305 4086 3414 4106
rect 3434 4086 3443 4106
rect 3305 4079 3443 4086
rect 3501 4106 3649 4115
rect 3501 4086 3510 4106
rect 3530 4086 3620 4106
rect 3640 4086 3649 4106
rect 3305 4077 3401 4079
rect 3501 4076 3649 4086
rect 3708 4106 3745 4116
rect 3708 4086 3716 4106
rect 3736 4086 3745 4106
rect 3557 4075 3593 4076
rect 3034 4066 3070 4068
rect 3034 4037 3071 4066
rect 2476 4028 2511 4029
rect 2453 4023 2511 4028
rect 2453 4003 2456 4023
rect 2476 4009 2511 4023
rect 2531 4009 2540 4029
rect 2476 4001 2540 4009
rect 2502 4000 2540 4001
rect 2503 3999 2540 4000
rect 2606 4033 2642 4034
rect 2714 4033 2750 4034
rect 2606 4027 2750 4033
rect 2606 4025 2667 4027
rect 2606 4005 2614 4025
rect 2634 4010 2667 4025
rect 2686 4025 2750 4027
rect 2686 4010 2722 4025
rect 2634 4005 2722 4010
rect 2742 4005 2750 4025
rect 2606 3999 2750 4005
rect 2816 4029 2854 4037
rect 2932 4033 2968 4034
rect 2816 4009 2825 4029
rect 2845 4009 2854 4029
rect 2816 4000 2854 4009
rect 2883 4025 2968 4033
rect 2883 4005 2940 4025
rect 2960 4005 2968 4025
rect 2816 3999 2853 4000
rect 2883 3999 2968 4005
rect 3034 4029 3072 4037
rect 3034 4009 3043 4029
rect 3063 4009 3072 4029
rect 3708 4019 3745 4086
rect 3780 4115 3811 4166
rect 4093 4154 4111 4172
rect 4129 4154 4145 4172
rect 3830 4115 3867 4116
rect 3780 4106 3867 4115
rect 3780 4086 3838 4106
rect 3858 4086 3867 4106
rect 3780 4076 3867 4086
rect 3926 4106 3963 4116
rect 3926 4086 3934 4106
rect 3954 4086 3963 4106
rect 3780 4075 3811 4076
rect 3405 4016 3442 4017
rect 3708 4016 3747 4019
rect 3404 4015 3747 4016
rect 3926 4015 3963 4086
rect 3034 4000 3072 4009
rect 3329 4010 3747 4015
rect 3034 3999 3071 4000
rect 2495 3971 2585 3977
rect 2495 3951 2511 3971
rect 2531 3969 2585 3971
rect 2531 3951 2556 3969
rect 2495 3949 2556 3951
rect 2576 3949 2585 3969
rect 2495 3943 2585 3949
rect 2508 3889 2545 3890
rect 2604 3889 2641 3890
rect 2660 3889 2696 3999
rect 2883 3978 2914 3999
rect 3329 3990 3332 4010
rect 3352 3990 3747 4010
rect 3776 3991 3963 4015
rect 2879 3977 2914 3978
rect 2757 3967 2914 3977
rect 2757 3947 2774 3967
rect 2794 3947 2914 3967
rect 2757 3940 2914 3947
rect 2981 3970 3130 3978
rect 2981 3950 2992 3970
rect 3012 3950 3051 3970
rect 3071 3950 3130 3970
rect 2981 3943 3130 3950
rect 3708 3965 3747 3990
rect 4093 3965 4145 4154
rect 4537 4182 4547 4200
rect 4565 4182 4577 4200
rect 4709 4198 4718 4218
rect 4738 4198 4747 4218
rect 4709 4190 4747 4198
rect 4813 4222 4898 4228
rect 4928 4227 4965 4228
rect 4813 4202 4821 4222
rect 4841 4202 4898 4222
rect 4813 4194 4898 4202
rect 4927 4218 4965 4227
rect 4927 4198 4936 4218
rect 4956 4198 4965 4218
rect 4813 4193 4849 4194
rect 4927 4190 4965 4198
rect 5031 4222 5175 4228
rect 5031 4202 5039 4222
rect 5059 4202 5092 4222
rect 5112 4202 5147 4222
rect 5167 4202 5175 4222
rect 5031 4194 5175 4202
rect 5031 4193 5067 4194
rect 5139 4193 5175 4194
rect 5241 4227 5278 4228
rect 5241 4226 5279 4227
rect 5241 4218 5305 4226
rect 5241 4198 5250 4218
rect 5270 4204 5305 4218
rect 5325 4204 5328 4224
rect 5270 4199 5328 4204
rect 5270 4198 5305 4199
rect 4537 4126 4577 4182
rect 4710 4161 4747 4190
rect 4711 4159 4747 4161
rect 4711 4137 4902 4159
rect 4928 4158 4965 4190
rect 5241 4186 5305 4198
rect 5345 4160 5372 4338
rect 5204 4158 5372 4160
rect 4928 4148 5372 4158
rect 5513 4254 5700 4278
rect 5731 4259 6124 4279
rect 6144 4259 6147 4279
rect 5731 4254 6147 4259
rect 5513 4183 5550 4254
rect 5731 4253 6072 4254
rect 5665 4193 5696 4194
rect 5513 4163 5522 4183
rect 5542 4163 5550 4183
rect 5513 4153 5550 4163
rect 5609 4183 5696 4193
rect 5609 4163 5618 4183
rect 5638 4163 5696 4183
rect 5609 4154 5696 4163
rect 5609 4153 5646 4154
rect 4534 4121 4577 4126
rect 4925 4132 5372 4148
rect 4925 4126 4953 4132
rect 5204 4131 5372 4132
rect 4534 4118 4684 4121
rect 4925 4118 4952 4126
rect 4534 4116 4952 4118
rect 4534 4098 4543 4116
rect 4561 4098 4952 4116
rect 5665 4103 5696 4154
rect 5731 4183 5768 4253
rect 6034 4252 6071 4253
rect 5883 4193 5919 4194
rect 5731 4163 5740 4183
rect 5760 4163 5768 4183
rect 5731 4153 5768 4163
rect 5827 4183 5975 4193
rect 6075 4190 6171 4192
rect 5827 4163 5836 4183
rect 5856 4163 5946 4183
rect 5966 4163 5975 4183
rect 5827 4154 5975 4163
rect 6033 4183 6171 4190
rect 6033 4163 6042 4183
rect 6062 4163 6171 4183
rect 6433 4166 6473 4348
rect 6033 4154 6171 4163
rect 5827 4153 5864 4154
rect 5557 4100 5598 4101
rect 4534 4095 4952 4098
rect 4534 4089 4577 4095
rect 4537 4086 4577 4089
rect 5449 4093 5598 4100
rect 4934 4077 4974 4078
rect 4645 4060 4974 4077
rect 5449 4073 5508 4093
rect 5528 4073 5567 4093
rect 5587 4073 5598 4093
rect 5449 4065 5598 4073
rect 5665 4096 5822 4103
rect 5665 4076 5785 4096
rect 5805 4076 5822 4096
rect 5665 4066 5822 4076
rect 5665 4065 5700 4066
rect 4529 4017 4572 4028
rect 4529 3999 4541 4017
rect 4559 3999 4572 4017
rect 4529 3973 4572 3999
rect 4645 3973 4672 4060
rect 4934 4051 4974 4060
rect 3708 3947 4147 3965
rect 2981 3942 3022 3943
rect 2715 3889 2752 3890
rect 2408 3880 2546 3889
rect 2408 3860 2517 3880
rect 2537 3860 2546 3880
rect 2408 3853 2546 3860
rect 2604 3880 2752 3889
rect 2604 3860 2613 3880
rect 2633 3860 2723 3880
rect 2743 3860 2752 3880
rect 2408 3851 2504 3853
rect 2604 3850 2752 3860
rect 2811 3880 2848 3890
rect 2811 3860 2819 3880
rect 2839 3860 2848 3880
rect 2660 3849 2696 3850
rect 2508 3790 2545 3791
rect 2811 3790 2848 3860
rect 2883 3889 2914 3940
rect 3708 3929 4108 3947
rect 4126 3929 4147 3947
rect 3708 3923 4147 3929
rect 3714 3919 4147 3923
rect 4529 3952 4672 3973
rect 4716 4025 4750 4041
rect 4934 4031 5327 4051
rect 5347 4031 5350 4051
rect 5665 4044 5696 4065
rect 5883 4044 5919 4154
rect 5938 4153 5975 4154
rect 6034 4153 6071 4154
rect 5994 4094 6084 4100
rect 5994 4074 6003 4094
rect 6023 4092 6084 4094
rect 6023 4074 6048 4092
rect 5994 4072 6048 4074
rect 6068 4072 6084 4092
rect 5994 4066 6084 4072
rect 5508 4043 5545 4044
rect 4934 4026 5350 4031
rect 5507 4034 5545 4043
rect 4934 4025 5275 4026
rect 4716 3955 4753 4025
rect 4868 3965 4899 3966
rect 4529 3950 4666 3952
rect 4093 3917 4145 3919
rect 4529 3908 4572 3950
rect 4716 3935 4725 3955
rect 4745 3935 4753 3955
rect 4716 3925 4753 3935
rect 4812 3955 4899 3965
rect 4812 3935 4821 3955
rect 4841 3935 4899 3955
rect 4812 3926 4899 3935
rect 4812 3925 4849 3926
rect 4527 3898 4572 3908
rect 2933 3889 2970 3890
rect 2883 3880 2970 3889
rect 2883 3860 2941 3880
rect 2961 3860 2970 3880
rect 2883 3850 2970 3860
rect 3029 3880 3066 3890
rect 3029 3860 3037 3880
rect 3057 3860 3066 3880
rect 4527 3880 4536 3898
rect 4554 3880 4572 3898
rect 4527 3874 4572 3880
rect 4868 3875 4899 3926
rect 4934 3955 4971 4025
rect 5237 4024 5274 4025
rect 5507 4014 5516 4034
rect 5536 4014 5545 4034
rect 5507 4006 5545 4014
rect 5611 4038 5696 4044
rect 5726 4043 5763 4044
rect 5611 4018 5619 4038
rect 5639 4018 5696 4038
rect 5611 4010 5696 4018
rect 5725 4034 5763 4043
rect 5725 4014 5734 4034
rect 5754 4014 5763 4034
rect 5611 4009 5647 4010
rect 5725 4006 5763 4014
rect 5829 4038 5973 4044
rect 5829 4018 5837 4038
rect 5857 4019 5889 4038
rect 5910 4019 5945 4038
rect 5857 4018 5945 4019
rect 5965 4018 5973 4038
rect 5829 4010 5973 4018
rect 5829 4009 5865 4010
rect 5937 4009 5973 4010
rect 6039 4043 6076 4044
rect 6039 4042 6077 4043
rect 6039 4034 6103 4042
rect 6039 4014 6048 4034
rect 6068 4020 6103 4034
rect 6123 4020 6126 4040
rect 6068 4015 6126 4020
rect 6068 4014 6103 4015
rect 5508 3977 5545 4006
rect 5509 3975 5545 3977
rect 5086 3965 5122 3966
rect 4934 3935 4943 3955
rect 4963 3935 4971 3955
rect 4934 3925 4971 3935
rect 5030 3955 5178 3965
rect 5278 3962 5374 3964
rect 5030 3935 5039 3955
rect 5059 3935 5149 3955
rect 5169 3935 5178 3955
rect 5030 3926 5178 3935
rect 5236 3955 5374 3962
rect 5236 3935 5245 3955
rect 5265 3935 5374 3955
rect 5509 3953 5700 3975
rect 5726 3974 5763 4006
rect 6039 4002 6103 4014
rect 6143 3976 6170 4154
rect 6002 3974 6170 3976
rect 5726 3948 6170 3974
rect 5236 3926 5374 3935
rect 5030 3925 5067 3926
rect 4527 3871 4564 3874
rect 4760 3872 4801 3873
rect 2883 3849 2914 3850
rect 2507 3789 2848 3790
rect 3029 3789 3066 3860
rect 4652 3865 4801 3872
rect 4096 3852 4133 3857
rect 4087 3848 4134 3852
rect 4087 3830 4106 3848
rect 4124 3830 4134 3848
rect 4652 3845 4711 3865
rect 4731 3845 4770 3865
rect 4790 3845 4801 3865
rect 4652 3837 4801 3845
rect 4868 3868 5025 3875
rect 4868 3848 4988 3868
rect 5008 3848 5025 3868
rect 4868 3838 5025 3848
rect 4868 3837 4903 3838
rect 2432 3784 2848 3789
rect 2432 3764 2435 3784
rect 2455 3764 2848 3784
rect 2879 3765 3066 3789
rect 3691 3787 3731 3792
rect 4087 3787 4134 3830
rect 4868 3816 4899 3837
rect 5086 3816 5122 3926
rect 5141 3925 5178 3926
rect 5237 3925 5274 3926
rect 5197 3866 5287 3872
rect 5197 3846 5206 3866
rect 5226 3864 5287 3866
rect 5226 3846 5251 3864
rect 5197 3844 5251 3846
rect 5271 3844 5287 3864
rect 5197 3838 5287 3844
rect 4711 3815 4748 3816
rect 3691 3748 4134 3787
rect 4524 3807 4561 3809
rect 4524 3799 4566 3807
rect 4524 3781 4534 3799
rect 4552 3781 4566 3799
rect 4524 3772 4566 3781
rect 4710 3806 4748 3815
rect 4710 3786 4719 3806
rect 4739 3786 4748 3806
rect 4710 3778 4748 3786
rect 4814 3810 4899 3816
rect 4929 3815 4966 3816
rect 4814 3790 4822 3810
rect 4842 3790 4899 3810
rect 4814 3782 4899 3790
rect 4928 3806 4966 3815
rect 4928 3786 4937 3806
rect 4957 3786 4966 3806
rect 4814 3781 4850 3782
rect 4928 3778 4966 3786
rect 5032 3814 5176 3816
rect 5032 3810 5084 3814
rect 5032 3790 5040 3810
rect 5060 3794 5084 3810
rect 5104 3810 5176 3814
rect 5104 3794 5148 3810
rect 5060 3790 5148 3794
rect 5168 3790 5176 3810
rect 5032 3782 5176 3790
rect 5032 3781 5068 3782
rect 5140 3781 5176 3782
rect 5242 3815 5279 3816
rect 5242 3814 5280 3815
rect 5242 3806 5306 3814
rect 5242 3786 5251 3806
rect 5271 3792 5306 3806
rect 5326 3792 5329 3812
rect 5271 3787 5329 3792
rect 5271 3786 5306 3787
rect 2785 3733 2825 3741
rect 2785 3711 2793 3733
rect 2817 3711 2825 3733
rect 2491 3487 2659 3488
rect 2785 3487 2825 3711
rect 3288 3715 3456 3716
rect 3691 3715 3731 3748
rect 4087 3715 4134 3748
rect 4525 3747 4566 3772
rect 4711 3747 4748 3778
rect 4929 3747 4966 3778
rect 5242 3774 5306 3786
rect 5346 3748 5373 3926
rect 4525 3720 4574 3747
rect 4710 3721 4759 3747
rect 4928 3746 5009 3747
rect 5205 3746 5373 3748
rect 4928 3721 5373 3746
rect 4929 3720 5373 3721
rect 3288 3714 3732 3715
rect 3288 3689 3733 3714
rect 3288 3687 3456 3689
rect 3652 3688 3733 3689
rect 3902 3688 3951 3714
rect 4087 3688 4136 3715
rect 3288 3509 3315 3687
rect 3355 3649 3419 3661
rect 3695 3657 3732 3688
rect 3913 3657 3950 3688
rect 4095 3663 4136 3688
rect 4527 3687 4574 3720
rect 4930 3687 4970 3720
rect 5205 3719 5373 3720
rect 5836 3724 5876 3948
rect 6002 3947 6170 3948
rect 5836 3702 5844 3724
rect 5868 3702 5876 3724
rect 5836 3694 5876 3702
rect 3355 3648 3390 3649
rect 3332 3643 3390 3648
rect 3332 3623 3335 3643
rect 3355 3629 3390 3643
rect 3410 3629 3419 3649
rect 3355 3621 3419 3629
rect 3381 3620 3419 3621
rect 3382 3619 3419 3620
rect 3485 3653 3521 3654
rect 3593 3653 3629 3654
rect 3485 3645 3629 3653
rect 3485 3625 3493 3645
rect 3513 3641 3601 3645
rect 3513 3625 3557 3641
rect 3485 3621 3557 3625
rect 3577 3625 3601 3641
rect 3621 3625 3629 3645
rect 3577 3621 3629 3625
rect 3485 3619 3629 3621
rect 3695 3649 3733 3657
rect 3811 3653 3847 3654
rect 3695 3629 3704 3649
rect 3724 3629 3733 3649
rect 3695 3620 3733 3629
rect 3762 3645 3847 3653
rect 3762 3625 3819 3645
rect 3839 3625 3847 3645
rect 3695 3619 3732 3620
rect 3762 3619 3847 3625
rect 3913 3649 3951 3657
rect 3913 3629 3922 3649
rect 3942 3629 3951 3649
rect 3913 3620 3951 3629
rect 4095 3654 4137 3663
rect 4095 3636 4109 3654
rect 4127 3636 4137 3654
rect 4095 3628 4137 3636
rect 4100 3626 4137 3628
rect 4527 3648 4970 3687
rect 3913 3619 3950 3620
rect 3374 3591 3464 3597
rect 3374 3571 3390 3591
rect 3410 3589 3464 3591
rect 3410 3571 3435 3589
rect 3374 3569 3435 3571
rect 3455 3569 3464 3589
rect 3374 3563 3464 3569
rect 3387 3509 3424 3510
rect 3483 3509 3520 3510
rect 3539 3509 3575 3619
rect 3762 3598 3793 3619
rect 4527 3605 4574 3648
rect 4930 3643 4970 3648
rect 5595 3646 5782 3670
rect 5813 3651 6206 3671
rect 6226 3651 6229 3671
rect 5813 3646 6229 3651
rect 3758 3597 3793 3598
rect 3636 3587 3793 3597
rect 3636 3567 3653 3587
rect 3673 3567 3793 3587
rect 3636 3560 3793 3567
rect 3860 3590 4009 3598
rect 3860 3570 3871 3590
rect 3891 3570 3930 3590
rect 3950 3570 4009 3590
rect 4527 3587 4537 3605
rect 4555 3587 4574 3605
rect 4527 3583 4574 3587
rect 4528 3578 4565 3583
rect 3860 3563 4009 3570
rect 5595 3575 5632 3646
rect 5813 3645 6154 3646
rect 5747 3585 5778 3586
rect 3860 3562 3901 3563
rect 4097 3561 4134 3564
rect 3594 3509 3631 3510
rect 3287 3500 3425 3509
rect 2491 3461 2935 3487
rect 2491 3459 2659 3461
rect 2491 3281 2518 3459
rect 2558 3421 2622 3433
rect 2898 3429 2935 3461
rect 2961 3460 3152 3482
rect 3287 3480 3396 3500
rect 3416 3480 3425 3500
rect 3287 3473 3425 3480
rect 3483 3500 3631 3509
rect 3483 3480 3492 3500
rect 3512 3480 3602 3500
rect 3622 3480 3631 3500
rect 3287 3471 3383 3473
rect 3483 3470 3631 3480
rect 3690 3500 3727 3510
rect 3690 3480 3698 3500
rect 3718 3480 3727 3500
rect 3539 3469 3575 3470
rect 3116 3458 3152 3460
rect 3116 3429 3153 3458
rect 2558 3420 2593 3421
rect 2535 3415 2593 3420
rect 2535 3395 2538 3415
rect 2558 3401 2593 3415
rect 2613 3401 2622 3421
rect 2558 3393 2622 3401
rect 2584 3392 2622 3393
rect 2585 3391 2622 3392
rect 2688 3425 2724 3426
rect 2796 3425 2832 3426
rect 2688 3417 2832 3425
rect 2688 3397 2696 3417
rect 2716 3416 2804 3417
rect 2716 3397 2751 3416
rect 2772 3397 2804 3416
rect 2824 3397 2832 3417
rect 2688 3391 2832 3397
rect 2898 3421 2936 3429
rect 3014 3425 3050 3426
rect 2898 3401 2907 3421
rect 2927 3401 2936 3421
rect 2898 3392 2936 3401
rect 2965 3417 3050 3425
rect 2965 3397 3022 3417
rect 3042 3397 3050 3417
rect 2898 3391 2935 3392
rect 2965 3391 3050 3397
rect 3116 3421 3154 3429
rect 3116 3401 3125 3421
rect 3145 3401 3154 3421
rect 3387 3410 3424 3411
rect 3690 3410 3727 3480
rect 3762 3509 3793 3560
rect 4089 3555 4134 3561
rect 4089 3537 4107 3555
rect 4125 3537 4134 3555
rect 5595 3555 5604 3575
rect 5624 3555 5632 3575
rect 5595 3545 5632 3555
rect 5691 3575 5778 3585
rect 5691 3555 5700 3575
rect 5720 3555 5778 3575
rect 5691 3546 5778 3555
rect 5691 3545 5728 3546
rect 4089 3527 4134 3537
rect 3812 3509 3849 3510
rect 3762 3500 3849 3509
rect 3762 3480 3820 3500
rect 3840 3480 3849 3500
rect 3762 3470 3849 3480
rect 3908 3500 3945 3510
rect 3908 3480 3916 3500
rect 3936 3480 3945 3500
rect 4089 3485 4132 3527
rect 4516 3516 4568 3518
rect 3995 3483 4132 3485
rect 3762 3469 3793 3470
rect 3908 3410 3945 3480
rect 3386 3409 3727 3410
rect 3116 3392 3154 3401
rect 3311 3404 3727 3409
rect 3116 3391 3153 3392
rect 2577 3363 2667 3369
rect 2577 3343 2593 3363
rect 2613 3361 2667 3363
rect 2613 3343 2638 3361
rect 2577 3341 2638 3343
rect 2658 3341 2667 3361
rect 2577 3335 2667 3341
rect 2590 3281 2627 3282
rect 2686 3281 2723 3282
rect 2742 3281 2778 3391
rect 2965 3370 2996 3391
rect 3311 3384 3314 3404
rect 3334 3384 3727 3404
rect 3911 3394 3945 3410
rect 3989 3462 4132 3483
rect 4514 3512 4947 3516
rect 4514 3506 4953 3512
rect 4514 3488 4535 3506
rect 4553 3488 4953 3506
rect 5747 3495 5778 3546
rect 5813 3575 5850 3645
rect 6116 3644 6153 3645
rect 5965 3585 6001 3586
rect 5813 3555 5822 3575
rect 5842 3555 5850 3575
rect 5813 3545 5850 3555
rect 5909 3575 6057 3585
rect 6157 3582 6253 3584
rect 5909 3555 5918 3575
rect 5938 3555 6028 3575
rect 6048 3555 6057 3575
rect 5909 3546 6057 3555
rect 6115 3575 6253 3582
rect 6115 3555 6124 3575
rect 6144 3555 6253 3575
rect 6115 3546 6253 3555
rect 5909 3545 5946 3546
rect 5639 3492 5680 3493
rect 4514 3470 4953 3488
rect 3687 3375 3727 3384
rect 3989 3375 4016 3462
rect 4089 3436 4132 3462
rect 4089 3418 4102 3436
rect 4120 3418 4132 3436
rect 4089 3407 4132 3418
rect 2961 3369 2996 3370
rect 2839 3359 2996 3369
rect 2839 3339 2856 3359
rect 2876 3339 2996 3359
rect 2839 3332 2996 3339
rect 3063 3362 3212 3370
rect 3063 3342 3074 3362
rect 3094 3342 3133 3362
rect 3153 3342 3212 3362
rect 3687 3358 4016 3375
rect 3687 3357 3727 3358
rect 3063 3335 3212 3342
rect 4084 3346 4124 3349
rect 4084 3340 4127 3346
rect 3709 3337 4127 3340
rect 3063 3334 3104 3335
rect 2797 3281 2834 3282
rect 2490 3272 2628 3281
rect 2490 3252 2599 3272
rect 2619 3252 2628 3272
rect 2490 3245 2628 3252
rect 2686 3272 2834 3281
rect 2686 3252 2695 3272
rect 2715 3252 2805 3272
rect 2825 3252 2834 3272
rect 2490 3243 2586 3245
rect 2686 3242 2834 3252
rect 2893 3272 2930 3282
rect 2893 3252 2901 3272
rect 2921 3252 2930 3272
rect 2742 3241 2778 3242
rect 2590 3182 2627 3183
rect 2893 3182 2930 3252
rect 2965 3281 2996 3332
rect 3709 3319 4100 3337
rect 4118 3319 4127 3337
rect 3709 3317 4127 3319
rect 3709 3309 3736 3317
rect 3977 3314 4127 3317
rect 3289 3303 3457 3304
rect 3708 3303 3736 3309
rect 3289 3287 3736 3303
rect 4084 3309 4127 3314
rect 3015 3281 3052 3282
rect 2965 3272 3052 3281
rect 2965 3252 3023 3272
rect 3043 3252 3052 3272
rect 2965 3242 3052 3252
rect 3111 3272 3148 3282
rect 3111 3252 3119 3272
rect 3139 3252 3148 3272
rect 2965 3241 2996 3242
rect 2589 3181 2930 3182
rect 3111 3181 3148 3252
rect 2514 3176 2930 3181
rect 2514 3156 2517 3176
rect 2537 3156 2930 3176
rect 2961 3157 3148 3181
rect 3289 3277 3733 3287
rect 3289 3275 3457 3277
rect 2356 3082 2385 3100
rect 3289 3097 3316 3275
rect 3356 3237 3420 3249
rect 3696 3245 3733 3277
rect 3759 3276 3950 3298
rect 3914 3274 3950 3276
rect 3914 3245 3951 3274
rect 4084 3253 4124 3309
rect 3356 3236 3391 3237
rect 3333 3231 3391 3236
rect 3333 3211 3336 3231
rect 3356 3217 3391 3231
rect 3411 3217 3420 3237
rect 3356 3209 3420 3217
rect 3382 3208 3420 3209
rect 3383 3207 3420 3208
rect 3486 3241 3522 3242
rect 3594 3241 3630 3242
rect 3486 3233 3630 3241
rect 3486 3213 3494 3233
rect 3514 3213 3549 3233
rect 3569 3213 3602 3233
rect 3622 3213 3630 3233
rect 3486 3207 3630 3213
rect 3696 3237 3734 3245
rect 3812 3241 3848 3242
rect 3696 3217 3705 3237
rect 3725 3217 3734 3237
rect 3696 3208 3734 3217
rect 3763 3233 3848 3241
rect 3763 3213 3820 3233
rect 3840 3213 3848 3233
rect 3696 3207 3733 3208
rect 3763 3207 3848 3213
rect 3914 3237 3952 3245
rect 3914 3217 3923 3237
rect 3943 3217 3952 3237
rect 4084 3235 4096 3253
rect 4114 3235 4124 3253
rect 4516 3281 4568 3470
rect 4914 3445 4953 3470
rect 5531 3485 5680 3492
rect 5531 3465 5590 3485
rect 5610 3465 5649 3485
rect 5669 3465 5680 3485
rect 5531 3457 5680 3465
rect 5747 3488 5904 3495
rect 5747 3468 5867 3488
rect 5887 3468 5904 3488
rect 5747 3458 5904 3468
rect 5747 3457 5782 3458
rect 4698 3420 4885 3444
rect 4914 3425 5309 3445
rect 5329 3425 5332 3445
rect 5747 3436 5778 3457
rect 5965 3436 6001 3546
rect 6020 3545 6057 3546
rect 6116 3545 6153 3546
rect 6076 3486 6166 3492
rect 6076 3466 6085 3486
rect 6105 3484 6166 3486
rect 6105 3466 6130 3484
rect 6076 3464 6130 3466
rect 6150 3464 6166 3484
rect 6076 3458 6166 3464
rect 5590 3435 5627 3436
rect 4914 3420 5332 3425
rect 5589 3426 5627 3435
rect 4698 3349 4735 3420
rect 4914 3419 5257 3420
rect 4914 3416 4953 3419
rect 5219 3418 5256 3419
rect 4850 3359 4881 3360
rect 4698 3329 4707 3349
rect 4727 3329 4735 3349
rect 4698 3319 4735 3329
rect 4794 3349 4881 3359
rect 4794 3329 4803 3349
rect 4823 3329 4881 3349
rect 4794 3320 4881 3329
rect 4794 3319 4831 3320
rect 4516 3263 4532 3281
rect 4550 3263 4568 3281
rect 4850 3269 4881 3320
rect 4916 3349 4953 3416
rect 5589 3406 5598 3426
rect 5618 3406 5627 3426
rect 5589 3398 5627 3406
rect 5693 3430 5778 3436
rect 5808 3435 5845 3436
rect 5693 3410 5701 3430
rect 5721 3410 5778 3430
rect 5693 3402 5778 3410
rect 5807 3426 5845 3435
rect 5807 3406 5816 3426
rect 5836 3406 5845 3426
rect 5693 3401 5729 3402
rect 5807 3398 5845 3406
rect 5911 3431 6055 3436
rect 5911 3430 5973 3431
rect 5911 3410 5919 3430
rect 5939 3412 5973 3430
rect 5994 3430 6055 3431
rect 5994 3412 6027 3430
rect 5939 3410 6027 3412
rect 6047 3410 6055 3430
rect 5911 3402 6055 3410
rect 5911 3401 5947 3402
rect 6019 3401 6055 3402
rect 6121 3435 6158 3436
rect 6121 3434 6159 3435
rect 6121 3426 6185 3434
rect 6121 3406 6130 3426
rect 6150 3412 6185 3426
rect 6205 3412 6208 3432
rect 6150 3407 6208 3412
rect 6150 3406 6185 3407
rect 5590 3369 5627 3398
rect 5591 3367 5627 3369
rect 5068 3359 5104 3360
rect 4916 3329 4925 3349
rect 4945 3329 4953 3349
rect 4916 3319 4953 3329
rect 5012 3349 5160 3359
rect 5260 3356 5356 3358
rect 5012 3329 5021 3349
rect 5041 3329 5131 3349
rect 5151 3329 5160 3349
rect 5012 3320 5160 3329
rect 5218 3349 5356 3356
rect 5218 3329 5227 3349
rect 5247 3329 5356 3349
rect 5591 3345 5782 3367
rect 5808 3366 5845 3398
rect 6121 3394 6185 3406
rect 6225 3368 6252 3546
rect 6084 3366 6252 3368
rect 5808 3352 6252 3366
rect 5808 3340 6255 3352
rect 5851 3338 5884 3340
rect 5218 3320 5356 3329
rect 5012 3319 5049 3320
rect 4742 3266 4783 3267
rect 4516 3245 4568 3263
rect 4634 3259 4783 3266
rect 4084 3225 4124 3235
rect 4634 3239 4693 3259
rect 4713 3239 4752 3259
rect 4772 3239 4783 3259
rect 4634 3231 4783 3239
rect 4850 3262 5007 3269
rect 4850 3242 4970 3262
rect 4990 3242 5007 3262
rect 4850 3232 5007 3242
rect 4850 3231 4885 3232
rect 3914 3208 3952 3217
rect 4850 3210 4881 3231
rect 5068 3210 5104 3320
rect 5123 3319 5160 3320
rect 5219 3319 5256 3320
rect 5179 3260 5269 3266
rect 5179 3240 5188 3260
rect 5208 3258 5269 3260
rect 5208 3240 5233 3258
rect 5179 3238 5233 3240
rect 5253 3238 5269 3258
rect 5179 3232 5269 3238
rect 4693 3209 4730 3210
rect 3914 3207 3951 3208
rect 3375 3179 3465 3185
rect 3375 3159 3391 3179
rect 3411 3177 3465 3179
rect 3411 3159 3436 3177
rect 3375 3157 3436 3159
rect 3456 3157 3465 3177
rect 3375 3151 3465 3157
rect 3388 3097 3425 3098
rect 3484 3097 3521 3098
rect 3540 3097 3576 3207
rect 3763 3186 3794 3207
rect 4692 3200 4730 3209
rect 3759 3185 3794 3186
rect 3637 3175 3794 3185
rect 3637 3155 3654 3175
rect 3674 3155 3794 3175
rect 3637 3148 3794 3155
rect 3861 3178 4010 3186
rect 3861 3158 3872 3178
rect 3892 3158 3931 3178
rect 3951 3158 4010 3178
rect 4520 3182 4560 3192
rect 3861 3151 4010 3158
rect 4076 3154 4128 3172
rect 3861 3150 3902 3151
rect 3595 3097 3632 3098
rect 2326 3080 2385 3082
rect 3288 3088 3426 3097
rect 2326 3079 2494 3080
rect 2620 3079 2660 3081
rect 2326 3053 2770 3079
rect 2326 3051 2494 3053
rect 2326 3049 2407 3051
rect 2326 2873 2353 3049
rect 2393 3013 2457 3025
rect 2733 3021 2770 3053
rect 2796 3052 2987 3074
rect 3288 3068 3397 3088
rect 3417 3068 3426 3088
rect 3288 3061 3426 3068
rect 3484 3088 3632 3097
rect 3484 3068 3493 3088
rect 3513 3068 3603 3088
rect 3623 3068 3632 3088
rect 3288 3059 3384 3061
rect 3484 3058 3632 3068
rect 3691 3088 3728 3098
rect 3691 3068 3699 3088
rect 3719 3068 3728 3088
rect 3540 3057 3576 3058
rect 2951 3050 2987 3052
rect 2951 3021 2988 3050
rect 2393 3012 2428 3013
rect 2370 3007 2428 3012
rect 2370 2987 2373 3007
rect 2393 2993 2428 3007
rect 2448 2993 2457 3013
rect 2393 2985 2457 2993
rect 2419 2984 2457 2985
rect 2420 2983 2457 2984
rect 2523 3017 2559 3018
rect 2631 3017 2667 3018
rect 2523 3009 2667 3017
rect 2523 2989 2531 3009
rect 2551 3008 2639 3009
rect 2551 2990 2586 3008
rect 2604 2990 2639 3008
rect 2551 2989 2639 2990
rect 2659 2989 2667 3009
rect 2523 2983 2667 2989
rect 2733 3013 2771 3021
rect 2849 3017 2885 3018
rect 2733 2993 2742 3013
rect 2762 2993 2771 3013
rect 2733 2984 2771 2993
rect 2800 3009 2885 3017
rect 2800 2989 2857 3009
rect 2877 2989 2885 3009
rect 2733 2983 2770 2984
rect 2800 2983 2885 2989
rect 2951 3013 2989 3021
rect 2951 2993 2960 3013
rect 2980 2993 2989 3013
rect 3691 3001 3728 3068
rect 3763 3097 3794 3148
rect 4076 3136 4094 3154
rect 4112 3136 4128 3154
rect 3813 3097 3850 3098
rect 3763 3088 3850 3097
rect 3763 3068 3821 3088
rect 3841 3068 3850 3088
rect 3763 3058 3850 3068
rect 3909 3088 3946 3098
rect 3909 3068 3917 3088
rect 3937 3068 3946 3088
rect 3763 3057 3794 3058
rect 3388 2998 3425 2999
rect 3691 2998 3730 3001
rect 3387 2997 3730 2998
rect 3909 2997 3946 3068
rect 2951 2984 2989 2993
rect 3312 2992 3730 2997
rect 2951 2983 2988 2984
rect 2412 2955 2502 2961
rect 2412 2935 2428 2955
rect 2448 2953 2502 2955
rect 2448 2935 2473 2953
rect 2412 2933 2473 2935
rect 2493 2933 2502 2953
rect 2412 2927 2502 2933
rect 2425 2873 2462 2874
rect 2521 2873 2558 2874
rect 2577 2873 2613 2983
rect 2800 2962 2831 2983
rect 3312 2972 3315 2992
rect 3335 2972 3730 2992
rect 3759 2973 3946 2997
rect 2796 2961 2831 2962
rect 2674 2951 2831 2961
rect 2674 2931 2691 2951
rect 2711 2931 2831 2951
rect 2674 2924 2831 2931
rect 2898 2954 3047 2962
rect 2898 2934 2909 2954
rect 2929 2934 2968 2954
rect 2988 2934 3047 2954
rect 2898 2927 3047 2934
rect 3691 2947 3730 2972
rect 4076 2947 4128 3136
rect 4520 3164 4530 3182
rect 4548 3164 4560 3182
rect 4692 3180 4701 3200
rect 4721 3180 4730 3200
rect 4692 3172 4730 3180
rect 4796 3204 4881 3210
rect 4911 3209 4948 3210
rect 4796 3184 4804 3204
rect 4824 3184 4881 3204
rect 4796 3176 4881 3184
rect 4910 3200 4948 3209
rect 4910 3180 4919 3200
rect 4939 3180 4948 3200
rect 4796 3175 4832 3176
rect 4910 3172 4948 3180
rect 5014 3204 5158 3210
rect 5014 3184 5022 3204
rect 5042 3184 5075 3204
rect 5095 3184 5130 3204
rect 5150 3184 5158 3204
rect 5014 3176 5158 3184
rect 5014 3175 5050 3176
rect 5122 3175 5158 3176
rect 5224 3209 5261 3210
rect 5224 3208 5262 3209
rect 5224 3200 5288 3208
rect 5224 3180 5233 3200
rect 5253 3186 5288 3200
rect 5308 3186 5311 3206
rect 5253 3181 5311 3186
rect 5253 3180 5288 3181
rect 4520 3108 4560 3164
rect 4693 3143 4730 3172
rect 4694 3141 4730 3143
rect 4694 3119 4885 3141
rect 4911 3140 4948 3172
rect 5224 3168 5288 3180
rect 5328 3142 5355 3320
rect 6213 3295 6255 3340
rect 5187 3140 5355 3142
rect 4911 3130 5355 3140
rect 5496 3236 5683 3260
rect 5714 3241 6107 3261
rect 6127 3241 6130 3261
rect 5714 3236 6130 3241
rect 5496 3165 5533 3236
rect 5714 3235 6055 3236
rect 5648 3175 5679 3176
rect 5496 3145 5505 3165
rect 5525 3145 5533 3165
rect 5496 3135 5533 3145
rect 5592 3165 5679 3175
rect 5592 3145 5601 3165
rect 5621 3145 5679 3165
rect 5592 3136 5679 3145
rect 5592 3135 5629 3136
rect 4517 3103 4560 3108
rect 4908 3114 5355 3130
rect 4908 3108 4936 3114
rect 5187 3113 5355 3114
rect 4517 3100 4667 3103
rect 4908 3100 4935 3108
rect 4517 3098 4935 3100
rect 4517 3080 4526 3098
rect 4544 3080 4935 3098
rect 5648 3085 5679 3136
rect 5714 3165 5751 3235
rect 6017 3234 6054 3235
rect 5866 3175 5902 3176
rect 5714 3145 5723 3165
rect 5743 3145 5751 3165
rect 5714 3135 5751 3145
rect 5810 3165 5958 3175
rect 6058 3172 6154 3174
rect 5810 3145 5819 3165
rect 5839 3145 5929 3165
rect 5949 3145 5958 3165
rect 5810 3136 5958 3145
rect 6016 3165 6154 3172
rect 6016 3145 6025 3165
rect 6045 3145 6154 3165
rect 6016 3136 6154 3145
rect 5810 3135 5847 3136
rect 5540 3082 5581 3083
rect 4517 3077 4935 3080
rect 4517 3071 4560 3077
rect 4520 3068 4560 3071
rect 5435 3075 5581 3082
rect 4917 3059 4957 3060
rect 4628 3042 4957 3059
rect 5435 3055 5491 3075
rect 5511 3055 5550 3075
rect 5570 3055 5581 3075
rect 5435 3047 5581 3055
rect 5648 3078 5805 3085
rect 5648 3058 5768 3078
rect 5788 3058 5805 3078
rect 5648 3048 5805 3058
rect 5648 3047 5683 3048
rect 4512 2999 4555 3010
rect 4512 2981 4524 2999
rect 4542 2981 4555 2999
rect 4512 2955 4555 2981
rect 4628 2955 4655 3042
rect 4917 3033 4957 3042
rect 3691 2929 4130 2947
rect 2898 2926 2939 2927
rect 2632 2873 2669 2874
rect 2325 2864 2463 2873
rect 2325 2844 2434 2864
rect 2454 2844 2463 2864
rect 2325 2837 2463 2844
rect 2521 2864 2669 2873
rect 2521 2844 2530 2864
rect 2550 2844 2640 2864
rect 2660 2844 2669 2864
rect 2325 2835 2421 2837
rect 2521 2834 2669 2844
rect 2728 2864 2765 2874
rect 2728 2844 2736 2864
rect 2756 2844 2765 2864
rect 2577 2833 2613 2834
rect 2425 2774 2462 2775
rect 2728 2774 2765 2844
rect 2800 2873 2831 2924
rect 3691 2911 4091 2929
rect 4109 2911 4130 2929
rect 3691 2905 4130 2911
rect 3697 2901 4130 2905
rect 4512 2934 4655 2955
rect 4699 3007 4733 3023
rect 4917 3013 5310 3033
rect 5330 3013 5333 3033
rect 5648 3026 5679 3047
rect 5866 3026 5902 3136
rect 5921 3135 5958 3136
rect 6017 3135 6054 3136
rect 5977 3076 6067 3082
rect 5977 3056 5986 3076
rect 6006 3074 6067 3076
rect 6006 3056 6031 3074
rect 5977 3054 6031 3056
rect 6051 3054 6067 3074
rect 5977 3048 6067 3054
rect 5491 3025 5528 3026
rect 4917 3008 5333 3013
rect 5490 3016 5528 3025
rect 4917 3007 5258 3008
rect 4699 2937 4736 3007
rect 4851 2947 4882 2948
rect 4512 2932 4649 2934
rect 4076 2899 4128 2901
rect 4512 2890 4555 2932
rect 4699 2917 4708 2937
rect 4728 2917 4736 2937
rect 4699 2907 4736 2917
rect 4795 2937 4882 2947
rect 4795 2917 4804 2937
rect 4824 2917 4882 2937
rect 4795 2908 4882 2917
rect 4795 2907 4832 2908
rect 4510 2880 4555 2890
rect 2850 2873 2887 2874
rect 2800 2864 2887 2873
rect 2800 2844 2858 2864
rect 2878 2844 2887 2864
rect 2800 2834 2887 2844
rect 2946 2864 2983 2874
rect 2946 2844 2954 2864
rect 2974 2844 2983 2864
rect 4510 2862 4519 2880
rect 4537 2862 4555 2880
rect 4510 2856 4555 2862
rect 4851 2857 4882 2908
rect 4917 2937 4954 3007
rect 5220 3006 5257 3007
rect 5490 2996 5499 3016
rect 5519 2996 5528 3016
rect 5490 2988 5528 2996
rect 5594 3020 5679 3026
rect 5709 3025 5746 3026
rect 5594 3000 5602 3020
rect 5622 3000 5679 3020
rect 5594 2992 5679 3000
rect 5708 3016 5746 3025
rect 5708 2996 5717 3016
rect 5737 2996 5746 3016
rect 5594 2991 5630 2992
rect 5708 2988 5746 2996
rect 5812 3020 5956 3026
rect 5812 3000 5820 3020
rect 5840 3017 5928 3020
rect 5840 3000 5875 3017
rect 5812 2999 5875 3000
rect 5894 3000 5928 3017
rect 5948 3000 5956 3020
rect 5894 2999 5956 3000
rect 5812 2992 5956 2999
rect 5812 2991 5848 2992
rect 5920 2991 5956 2992
rect 6022 3025 6059 3026
rect 6022 3024 6060 3025
rect 6082 3024 6109 3028
rect 6022 3022 6109 3024
rect 6022 3016 6086 3022
rect 6022 2996 6031 3016
rect 6051 3002 6086 3016
rect 6106 3002 6109 3022
rect 6051 2997 6109 3002
rect 6051 2996 6086 2997
rect 5491 2959 5528 2988
rect 5492 2957 5528 2959
rect 5069 2947 5105 2948
rect 4917 2917 4926 2937
rect 4946 2917 4954 2937
rect 4917 2907 4954 2917
rect 5013 2937 5161 2947
rect 5261 2944 5357 2946
rect 5013 2917 5022 2937
rect 5042 2917 5132 2937
rect 5152 2917 5161 2937
rect 5013 2908 5161 2917
rect 5219 2937 5357 2944
rect 5219 2917 5228 2937
rect 5248 2917 5357 2937
rect 5492 2935 5683 2957
rect 5709 2956 5746 2988
rect 6022 2984 6086 2996
rect 6126 2958 6153 3136
rect 5985 2956 6153 2958
rect 5709 2930 6153 2956
rect 5219 2908 5357 2917
rect 5013 2907 5050 2908
rect 4510 2853 4547 2856
rect 4743 2854 4784 2855
rect 2800 2833 2831 2834
rect 2424 2773 2765 2774
rect 2946 2773 2983 2844
rect 4635 2847 4784 2854
rect 4079 2834 4116 2839
rect 2349 2768 2765 2773
rect 2349 2748 2352 2768
rect 2372 2748 2765 2768
rect 2796 2749 2983 2773
rect 4070 2830 4117 2834
rect 4070 2812 4089 2830
rect 4107 2812 4117 2830
rect 4635 2827 4694 2847
rect 4714 2827 4753 2847
rect 4773 2827 4784 2847
rect 4635 2819 4784 2827
rect 4851 2850 5008 2857
rect 4851 2830 4971 2850
rect 4991 2830 5008 2850
rect 4851 2820 5008 2830
rect 4851 2819 4886 2820
rect 4070 2764 4117 2812
rect 4851 2798 4882 2819
rect 5069 2798 5105 2908
rect 5124 2907 5161 2908
rect 5220 2907 5257 2908
rect 5180 2848 5270 2854
rect 5180 2828 5189 2848
rect 5209 2846 5270 2848
rect 5209 2828 5234 2846
rect 5180 2826 5234 2828
rect 5254 2826 5270 2846
rect 5180 2820 5270 2826
rect 4694 2797 4731 2798
rect 3694 2761 4117 2764
rect 2569 2747 2634 2748
rect 3672 2731 4117 2761
rect 4506 2789 4544 2791
rect 4506 2781 4549 2789
rect 4506 2763 4517 2781
rect 4535 2763 4549 2781
rect 4506 2736 4549 2763
rect 4693 2788 4731 2797
rect 4693 2768 4702 2788
rect 4722 2768 4731 2788
rect 4693 2760 4731 2768
rect 4797 2792 4882 2798
rect 4912 2797 4949 2798
rect 4797 2772 4805 2792
rect 4825 2772 4882 2792
rect 4797 2764 4882 2772
rect 4911 2788 4949 2797
rect 4911 2768 4920 2788
rect 4940 2768 4949 2788
rect 4797 2763 4833 2764
rect 4911 2760 4949 2768
rect 5015 2796 5159 2798
rect 5015 2792 5067 2796
rect 5015 2772 5023 2792
rect 5043 2776 5067 2792
rect 5087 2792 5159 2796
rect 5087 2776 5131 2792
rect 5043 2772 5131 2776
rect 5151 2772 5159 2792
rect 5015 2764 5159 2772
rect 5015 2763 5051 2764
rect 5123 2763 5159 2764
rect 5225 2797 5262 2798
rect 5225 2796 5263 2797
rect 5225 2788 5289 2796
rect 5225 2768 5234 2788
rect 5254 2774 5289 2788
rect 5309 2774 5312 2794
rect 5254 2769 5312 2774
rect 5254 2768 5289 2769
rect 2765 2715 2805 2723
rect 2765 2693 2773 2715
rect 2797 2693 2805 2715
rect 2370 2464 2407 2470
rect 2370 2445 2378 2464
rect 2399 2445 2407 2464
rect 2370 2437 2407 2445
rect 2070 2316 2077 2338
rect 2101 2316 2109 2338
rect 2070 2310 2109 2316
rect 1600 2305 1640 2307
rect 1766 2306 1934 2307
rect 1868 2305 1905 2306
rect 834 2289 972 2298
rect 628 2288 665 2289
rect 358 2235 399 2236
rect 132 2214 184 2232
rect 250 2228 399 2235
rect 250 2208 309 2228
rect 329 2208 368 2228
rect 388 2208 399 2228
rect 250 2200 399 2208
rect 466 2231 623 2238
rect 466 2211 586 2231
rect 606 2211 623 2231
rect 466 2201 623 2211
rect 466 2200 501 2201
rect 466 2179 497 2200
rect 684 2179 720 2289
rect 739 2288 776 2289
rect 835 2288 872 2289
rect 795 2229 885 2235
rect 795 2209 804 2229
rect 824 2227 885 2229
rect 824 2209 849 2227
rect 795 2207 849 2209
rect 869 2207 885 2227
rect 795 2201 885 2207
rect 309 2178 346 2179
rect 308 2169 346 2178
rect 136 2151 176 2161
rect 136 2133 146 2151
rect 164 2133 176 2151
rect 308 2149 317 2169
rect 337 2149 346 2169
rect 308 2141 346 2149
rect 412 2173 497 2179
rect 527 2178 564 2179
rect 412 2153 420 2173
rect 440 2153 497 2173
rect 412 2145 497 2153
rect 526 2169 564 2178
rect 526 2149 535 2169
rect 555 2149 564 2169
rect 412 2144 448 2145
rect 526 2141 564 2149
rect 630 2173 774 2179
rect 630 2153 638 2173
rect 658 2153 691 2173
rect 711 2153 746 2173
rect 766 2153 774 2173
rect 630 2145 774 2153
rect 630 2144 666 2145
rect 738 2144 774 2145
rect 840 2178 877 2179
rect 840 2177 878 2178
rect 840 2169 904 2177
rect 840 2149 849 2169
rect 869 2155 904 2169
rect 924 2155 927 2175
rect 869 2150 927 2155
rect 869 2149 904 2150
rect 136 2077 176 2133
rect 309 2112 346 2141
rect 310 2110 346 2112
rect 310 2088 501 2110
rect 527 2109 564 2141
rect 840 2137 904 2149
rect 944 2111 971 2289
rect 803 2109 971 2111
rect 527 2099 971 2109
rect 1112 2205 1299 2229
rect 1330 2210 1723 2230
rect 1743 2210 1746 2230
rect 1330 2205 1746 2210
rect 1112 2134 1149 2205
rect 1330 2204 1671 2205
rect 1264 2144 1295 2145
rect 1112 2114 1121 2134
rect 1141 2114 1149 2134
rect 1112 2104 1149 2114
rect 1208 2134 1295 2144
rect 1208 2114 1217 2134
rect 1237 2114 1295 2134
rect 1208 2105 1295 2114
rect 1208 2104 1245 2105
rect 133 2072 176 2077
rect 524 2083 971 2099
rect 524 2077 552 2083
rect 803 2082 971 2083
rect 133 2069 283 2072
rect 524 2069 551 2077
rect 133 2067 551 2069
rect 133 2049 142 2067
rect 160 2049 551 2067
rect 1264 2054 1295 2105
rect 1330 2134 1367 2204
rect 1633 2203 1670 2204
rect 1871 2146 1904 2305
rect 1482 2144 1518 2145
rect 1330 2114 1339 2134
rect 1359 2114 1367 2134
rect 1330 2104 1367 2114
rect 1426 2134 1574 2144
rect 1674 2141 1770 2143
rect 1426 2114 1435 2134
rect 1455 2114 1545 2134
rect 1565 2114 1574 2134
rect 1426 2105 1574 2114
rect 1632 2134 1770 2141
rect 1632 2114 1641 2134
rect 1661 2114 1770 2134
rect 1871 2142 1907 2146
rect 1871 2124 1880 2142
rect 1902 2124 1907 2142
rect 1871 2118 1907 2124
rect 1632 2105 1770 2114
rect 1426 2104 1463 2105
rect 1156 2051 1197 2052
rect 133 2046 551 2049
rect 133 2040 176 2046
rect 136 2037 176 2040
rect 1048 2044 1197 2051
rect 533 2028 573 2029
rect 244 2011 573 2028
rect 1048 2024 1107 2044
rect 1127 2024 1166 2044
rect 1186 2024 1197 2044
rect 1048 2016 1197 2024
rect 1264 2047 1421 2054
rect 1264 2027 1384 2047
rect 1404 2027 1421 2047
rect 1264 2017 1421 2027
rect 1264 2016 1299 2017
rect 128 1968 171 1979
rect 128 1950 140 1968
rect 158 1950 171 1968
rect 128 1924 171 1950
rect 244 1924 271 2011
rect 533 2002 573 2011
rect 128 1903 271 1924
rect 315 1976 349 1992
rect 533 1982 926 2002
rect 946 1982 949 2002
rect 1264 1995 1295 2016
rect 1482 1995 1518 2105
rect 1537 2104 1574 2105
rect 1633 2104 1670 2105
rect 1593 2045 1683 2051
rect 1593 2025 1602 2045
rect 1622 2043 1683 2045
rect 1622 2025 1647 2043
rect 1593 2023 1647 2025
rect 1667 2023 1683 2043
rect 1593 2017 1683 2023
rect 1107 1994 1144 1995
rect 533 1977 949 1982
rect 1106 1985 1144 1994
rect 533 1976 874 1977
rect 315 1906 352 1976
rect 467 1916 498 1917
rect 128 1901 265 1903
rect 128 1859 171 1901
rect 315 1886 324 1906
rect 344 1886 352 1906
rect 315 1876 352 1886
rect 411 1906 498 1916
rect 411 1886 420 1906
rect 440 1886 498 1906
rect 411 1877 498 1886
rect 411 1876 448 1877
rect 126 1849 171 1859
rect 126 1831 135 1849
rect 153 1831 171 1849
rect 126 1825 171 1831
rect 467 1826 498 1877
rect 533 1906 570 1976
rect 836 1975 873 1976
rect 1106 1965 1115 1985
rect 1135 1965 1144 1985
rect 1106 1957 1144 1965
rect 1210 1989 1295 1995
rect 1325 1994 1362 1995
rect 1210 1969 1218 1989
rect 1238 1969 1295 1989
rect 1210 1961 1295 1969
rect 1324 1985 1362 1994
rect 1324 1965 1333 1985
rect 1353 1965 1362 1985
rect 1210 1960 1246 1961
rect 1324 1957 1362 1965
rect 1428 1989 1572 1995
rect 1428 1969 1436 1989
rect 1456 1970 1488 1989
rect 1509 1970 1544 1989
rect 1456 1969 1544 1970
rect 1564 1969 1572 1989
rect 1428 1961 1572 1969
rect 1428 1960 1464 1961
rect 1536 1960 1572 1961
rect 1638 1994 1675 1995
rect 1638 1993 1676 1994
rect 1638 1985 1702 1993
rect 1638 1965 1647 1985
rect 1667 1971 1702 1985
rect 1722 1971 1725 1991
rect 1667 1966 1725 1971
rect 1667 1965 1702 1966
rect 1107 1928 1144 1957
rect 1108 1926 1144 1928
rect 685 1916 721 1917
rect 533 1886 542 1906
rect 562 1886 570 1906
rect 533 1876 570 1886
rect 629 1906 777 1916
rect 877 1913 973 1915
rect 629 1886 638 1906
rect 658 1886 748 1906
rect 768 1886 777 1906
rect 629 1877 777 1886
rect 835 1906 973 1913
rect 835 1886 844 1906
rect 864 1886 973 1906
rect 1108 1904 1299 1926
rect 1325 1925 1362 1957
rect 1638 1953 1702 1965
rect 1742 1927 1769 2105
rect 2374 2104 2407 2437
rect 2471 2469 2639 2470
rect 2765 2469 2805 2693
rect 3268 2697 3436 2698
rect 3672 2697 3713 2731
rect 4070 2710 4117 2731
rect 3268 2687 3713 2697
rect 3785 2695 3928 2696
rect 3268 2671 3712 2687
rect 3268 2669 3436 2671
rect 3632 2670 3712 2671
rect 3785 2670 3930 2695
rect 4072 2670 4117 2710
rect 3268 2491 3295 2669
rect 3335 2631 3399 2643
rect 3675 2639 3712 2670
rect 3893 2639 3930 2670
rect 4075 2663 4117 2670
rect 4507 2729 4549 2736
rect 4694 2729 4731 2760
rect 4912 2729 4949 2760
rect 5225 2756 5289 2768
rect 5329 2730 5356 2908
rect 4507 2689 4552 2729
rect 4694 2704 4839 2729
rect 4912 2728 4992 2729
rect 5188 2728 5356 2730
rect 4912 2712 5356 2728
rect 4696 2703 4839 2704
rect 4911 2702 5356 2712
rect 4507 2668 4554 2689
rect 4911 2668 4952 2702
rect 5188 2701 5356 2702
rect 5819 2706 5859 2930
rect 5985 2929 6153 2930
rect 6217 2962 6250 3295
rect 6217 2954 6254 2962
rect 6217 2935 6225 2954
rect 6246 2935 6254 2954
rect 6217 2929 6254 2935
rect 5819 2684 5827 2706
rect 5851 2684 5859 2706
rect 5819 2676 5859 2684
rect 3335 2630 3370 2631
rect 3312 2625 3370 2630
rect 3312 2605 3315 2625
rect 3335 2611 3370 2625
rect 3390 2611 3399 2631
rect 3335 2603 3399 2611
rect 3361 2602 3399 2603
rect 3362 2601 3399 2602
rect 3465 2635 3501 2636
rect 3573 2635 3609 2636
rect 3465 2627 3609 2635
rect 3465 2607 3473 2627
rect 3493 2623 3581 2627
rect 3493 2607 3537 2623
rect 3465 2603 3537 2607
rect 3557 2607 3581 2623
rect 3601 2607 3609 2627
rect 3557 2603 3609 2607
rect 3465 2601 3609 2603
rect 3675 2631 3713 2639
rect 3791 2635 3827 2636
rect 3675 2611 3684 2631
rect 3704 2611 3713 2631
rect 3675 2602 3713 2611
rect 3742 2627 3827 2635
rect 3742 2607 3799 2627
rect 3819 2607 3827 2627
rect 3675 2601 3712 2602
rect 3742 2601 3827 2607
rect 3893 2631 3931 2639
rect 3893 2611 3902 2631
rect 3922 2611 3931 2631
rect 3893 2602 3931 2611
rect 4075 2636 4118 2663
rect 4075 2618 4089 2636
rect 4107 2618 4118 2636
rect 4075 2610 4118 2618
rect 4080 2608 4118 2610
rect 4507 2638 4952 2668
rect 5990 2651 6055 2652
rect 4507 2635 4930 2638
rect 3893 2601 3930 2602
rect 3354 2573 3444 2579
rect 3354 2553 3370 2573
rect 3390 2571 3444 2573
rect 3390 2553 3415 2571
rect 3354 2551 3415 2553
rect 3435 2551 3444 2571
rect 3354 2545 3444 2551
rect 3367 2491 3404 2492
rect 3463 2491 3500 2492
rect 3519 2491 3555 2601
rect 3742 2580 3773 2601
rect 4507 2587 4554 2635
rect 3738 2579 3773 2580
rect 3616 2569 3773 2579
rect 3616 2549 3633 2569
rect 3653 2549 3773 2569
rect 3616 2542 3773 2549
rect 3840 2572 3989 2580
rect 3840 2552 3851 2572
rect 3871 2552 3910 2572
rect 3930 2552 3989 2572
rect 4507 2569 4517 2587
rect 4535 2569 4554 2587
rect 4507 2565 4554 2569
rect 5641 2626 5828 2650
rect 5859 2631 6252 2651
rect 6272 2631 6275 2651
rect 5859 2626 6275 2631
rect 4508 2560 4545 2565
rect 3840 2545 3989 2552
rect 5641 2555 5678 2626
rect 5859 2625 6200 2626
rect 5793 2565 5824 2566
rect 3840 2544 3881 2545
rect 4077 2543 4114 2546
rect 3574 2491 3611 2492
rect 3267 2482 3405 2491
rect 2471 2443 2915 2469
rect 2471 2441 2639 2443
rect 2471 2263 2498 2441
rect 2538 2403 2602 2415
rect 2878 2411 2915 2443
rect 2941 2442 3132 2464
rect 3267 2462 3376 2482
rect 3396 2462 3405 2482
rect 3267 2455 3405 2462
rect 3463 2482 3611 2491
rect 3463 2462 3472 2482
rect 3492 2462 3582 2482
rect 3602 2462 3611 2482
rect 3267 2453 3363 2455
rect 3463 2452 3611 2462
rect 3670 2482 3707 2492
rect 3670 2462 3678 2482
rect 3698 2462 3707 2482
rect 3519 2451 3555 2452
rect 3096 2440 3132 2442
rect 3096 2411 3133 2440
rect 2538 2402 2573 2403
rect 2515 2397 2573 2402
rect 2515 2377 2518 2397
rect 2538 2383 2573 2397
rect 2593 2383 2602 2403
rect 2538 2377 2602 2383
rect 2515 2375 2602 2377
rect 2515 2371 2542 2375
rect 2564 2374 2602 2375
rect 2565 2373 2602 2374
rect 2668 2407 2704 2408
rect 2776 2407 2812 2408
rect 2668 2400 2812 2407
rect 2668 2399 2730 2400
rect 2668 2379 2676 2399
rect 2696 2382 2730 2399
rect 2749 2399 2812 2400
rect 2749 2382 2784 2399
rect 2696 2379 2784 2382
rect 2804 2379 2812 2399
rect 2668 2373 2812 2379
rect 2878 2403 2916 2411
rect 2994 2407 3030 2408
rect 2878 2383 2887 2403
rect 2907 2383 2916 2403
rect 2878 2374 2916 2383
rect 2945 2399 3030 2407
rect 2945 2379 3002 2399
rect 3022 2379 3030 2399
rect 2878 2373 2915 2374
rect 2945 2373 3030 2379
rect 3096 2403 3134 2411
rect 3096 2383 3105 2403
rect 3125 2383 3134 2403
rect 3367 2392 3404 2393
rect 3670 2392 3707 2462
rect 3742 2491 3773 2542
rect 4069 2537 4114 2543
rect 4069 2519 4087 2537
rect 4105 2519 4114 2537
rect 5641 2535 5650 2555
rect 5670 2535 5678 2555
rect 5641 2525 5678 2535
rect 5737 2555 5824 2565
rect 5737 2535 5746 2555
rect 5766 2535 5824 2555
rect 5737 2526 5824 2535
rect 5737 2525 5774 2526
rect 4069 2509 4114 2519
rect 3792 2491 3829 2492
rect 3742 2482 3829 2491
rect 3742 2462 3800 2482
rect 3820 2462 3829 2482
rect 3742 2452 3829 2462
rect 3888 2482 3925 2492
rect 3888 2462 3896 2482
rect 3916 2462 3925 2482
rect 4069 2467 4112 2509
rect 4496 2498 4548 2500
rect 3975 2465 4112 2467
rect 3742 2451 3773 2452
rect 3888 2392 3925 2462
rect 3366 2391 3707 2392
rect 3096 2374 3134 2383
rect 3291 2386 3707 2391
rect 3096 2373 3133 2374
rect 2557 2345 2647 2351
rect 2557 2325 2573 2345
rect 2593 2343 2647 2345
rect 2593 2325 2618 2343
rect 2557 2323 2618 2325
rect 2638 2323 2647 2343
rect 2557 2317 2647 2323
rect 2570 2263 2607 2264
rect 2666 2263 2703 2264
rect 2722 2263 2758 2373
rect 2945 2352 2976 2373
rect 3291 2366 3294 2386
rect 3314 2366 3707 2386
rect 3891 2376 3925 2392
rect 3969 2444 4112 2465
rect 4494 2494 4927 2498
rect 4494 2488 4933 2494
rect 4494 2470 4515 2488
rect 4533 2470 4933 2488
rect 5793 2475 5824 2526
rect 5859 2555 5896 2625
rect 6162 2624 6199 2625
rect 6011 2565 6047 2566
rect 5859 2535 5868 2555
rect 5888 2535 5896 2555
rect 5859 2525 5896 2535
rect 5955 2555 6103 2565
rect 6203 2562 6299 2564
rect 5955 2535 5964 2555
rect 5984 2535 6074 2555
rect 6094 2535 6103 2555
rect 5955 2526 6103 2535
rect 6161 2555 6299 2562
rect 6161 2535 6170 2555
rect 6190 2535 6299 2555
rect 6161 2526 6299 2535
rect 5955 2525 5992 2526
rect 5685 2472 5726 2473
rect 4494 2452 4933 2470
rect 3667 2357 3707 2366
rect 3969 2357 3996 2444
rect 4069 2418 4112 2444
rect 4069 2400 4082 2418
rect 4100 2400 4112 2418
rect 4069 2389 4112 2400
rect 2941 2351 2976 2352
rect 2819 2341 2976 2351
rect 2819 2321 2836 2341
rect 2856 2321 2976 2341
rect 2819 2314 2976 2321
rect 3043 2344 3189 2352
rect 3043 2324 3054 2344
rect 3074 2324 3113 2344
rect 3133 2324 3189 2344
rect 3667 2340 3996 2357
rect 3667 2339 3707 2340
rect 3043 2317 3189 2324
rect 4064 2328 4104 2331
rect 4064 2322 4107 2328
rect 3689 2319 4107 2322
rect 3043 2316 3084 2317
rect 2777 2263 2814 2264
rect 2470 2254 2608 2263
rect 2470 2234 2579 2254
rect 2599 2234 2608 2254
rect 2470 2227 2608 2234
rect 2666 2254 2814 2263
rect 2666 2234 2675 2254
rect 2695 2234 2785 2254
rect 2805 2234 2814 2254
rect 2470 2225 2566 2227
rect 2666 2224 2814 2234
rect 2873 2254 2910 2264
rect 2873 2234 2881 2254
rect 2901 2234 2910 2254
rect 2722 2223 2758 2224
rect 2570 2164 2607 2165
rect 2873 2164 2910 2234
rect 2945 2263 2976 2314
rect 3689 2301 4080 2319
rect 4098 2301 4107 2319
rect 3689 2299 4107 2301
rect 3689 2291 3716 2299
rect 3957 2296 4107 2299
rect 3269 2285 3437 2286
rect 3688 2285 3716 2291
rect 3269 2269 3716 2285
rect 4064 2291 4107 2296
rect 2995 2263 3032 2264
rect 2945 2254 3032 2263
rect 2945 2234 3003 2254
rect 3023 2234 3032 2254
rect 2945 2224 3032 2234
rect 3091 2254 3128 2264
rect 3091 2234 3099 2254
rect 3119 2234 3128 2254
rect 2945 2223 2976 2224
rect 2569 2163 2910 2164
rect 3091 2163 3128 2234
rect 2494 2158 2910 2163
rect 2494 2138 2497 2158
rect 2517 2138 2910 2158
rect 2941 2139 3128 2163
rect 3269 2259 3713 2269
rect 3269 2257 3437 2259
rect 2369 2059 2411 2104
rect 3269 2079 3296 2257
rect 3336 2219 3400 2231
rect 3676 2227 3713 2259
rect 3739 2258 3930 2280
rect 3894 2256 3930 2258
rect 3894 2227 3931 2256
rect 4064 2235 4104 2291
rect 3336 2218 3371 2219
rect 3313 2213 3371 2218
rect 3313 2193 3316 2213
rect 3336 2199 3371 2213
rect 3391 2199 3400 2219
rect 3336 2191 3400 2199
rect 3362 2190 3400 2191
rect 3363 2189 3400 2190
rect 3466 2223 3502 2224
rect 3574 2223 3610 2224
rect 3466 2215 3610 2223
rect 3466 2195 3474 2215
rect 3494 2195 3529 2215
rect 3549 2195 3582 2215
rect 3602 2195 3610 2215
rect 3466 2189 3610 2195
rect 3676 2219 3714 2227
rect 3792 2223 3828 2224
rect 3676 2199 3685 2219
rect 3705 2199 3714 2219
rect 3676 2190 3714 2199
rect 3743 2215 3828 2223
rect 3743 2195 3800 2215
rect 3820 2195 3828 2215
rect 3676 2189 3713 2190
rect 3743 2189 3828 2195
rect 3894 2219 3932 2227
rect 3894 2199 3903 2219
rect 3923 2199 3932 2219
rect 4064 2217 4076 2235
rect 4094 2217 4104 2235
rect 4496 2263 4548 2452
rect 4894 2427 4933 2452
rect 5577 2465 5726 2472
rect 5577 2445 5636 2465
rect 5656 2445 5695 2465
rect 5715 2445 5726 2465
rect 5577 2437 5726 2445
rect 5793 2468 5950 2475
rect 5793 2448 5913 2468
rect 5933 2448 5950 2468
rect 5793 2438 5950 2448
rect 5793 2437 5828 2438
rect 4678 2402 4865 2426
rect 4894 2407 5289 2427
rect 5309 2407 5312 2427
rect 5793 2416 5824 2437
rect 6011 2416 6047 2526
rect 6066 2525 6103 2526
rect 6162 2525 6199 2526
rect 6122 2466 6212 2472
rect 6122 2446 6131 2466
rect 6151 2464 6212 2466
rect 6151 2446 6176 2464
rect 6122 2444 6176 2446
rect 6196 2444 6212 2464
rect 6122 2438 6212 2444
rect 5636 2415 5673 2416
rect 4894 2402 5312 2407
rect 5635 2406 5673 2415
rect 4678 2331 4715 2402
rect 4894 2401 5237 2402
rect 4894 2398 4933 2401
rect 5199 2400 5236 2401
rect 4830 2341 4861 2342
rect 4678 2311 4687 2331
rect 4707 2311 4715 2331
rect 4678 2301 4715 2311
rect 4774 2331 4861 2341
rect 4774 2311 4783 2331
rect 4803 2311 4861 2331
rect 4774 2302 4861 2311
rect 4774 2301 4811 2302
rect 4496 2245 4512 2263
rect 4530 2245 4548 2263
rect 4830 2251 4861 2302
rect 4896 2331 4933 2398
rect 5635 2386 5644 2406
rect 5664 2386 5673 2406
rect 5635 2378 5673 2386
rect 5739 2410 5824 2416
rect 5854 2415 5891 2416
rect 5739 2390 5747 2410
rect 5767 2390 5824 2410
rect 5739 2382 5824 2390
rect 5853 2406 5891 2415
rect 5853 2386 5862 2406
rect 5882 2386 5891 2406
rect 5739 2381 5775 2382
rect 5853 2378 5891 2386
rect 5957 2414 6101 2416
rect 5957 2410 6017 2414
rect 5957 2390 5965 2410
rect 5985 2392 6017 2410
rect 6040 2410 6101 2414
rect 6040 2392 6073 2410
rect 5985 2390 6073 2392
rect 6093 2390 6101 2410
rect 5957 2382 6101 2390
rect 5957 2381 5993 2382
rect 6065 2381 6101 2382
rect 6167 2415 6204 2416
rect 6167 2414 6205 2415
rect 6167 2406 6231 2414
rect 6167 2386 6176 2406
rect 6196 2392 6231 2406
rect 6251 2392 6254 2412
rect 6196 2387 6254 2392
rect 6196 2386 6231 2387
rect 5636 2349 5673 2378
rect 5637 2347 5673 2349
rect 5048 2341 5084 2342
rect 4896 2311 4905 2331
rect 4925 2311 4933 2331
rect 4896 2301 4933 2311
rect 4992 2331 5140 2341
rect 5240 2338 5336 2340
rect 4992 2311 5001 2331
rect 5021 2311 5111 2331
rect 5131 2311 5140 2331
rect 4992 2302 5140 2311
rect 5198 2331 5336 2338
rect 5198 2311 5207 2331
rect 5227 2311 5336 2331
rect 5637 2325 5828 2347
rect 5854 2346 5891 2378
rect 6167 2374 6231 2386
rect 5854 2345 6129 2346
rect 6271 2345 6298 2526
rect 5854 2320 6298 2345
rect 6434 2351 6473 4166
rect 6775 4153 6808 4486
rect 6872 4518 7040 4519
rect 7166 4518 7206 4742
rect 7669 4746 7837 4747
rect 8078 4746 8113 4763
rect 8470 4753 8517 4764
rect 7669 4720 8113 4746
rect 7669 4718 7837 4720
rect 8033 4719 8113 4720
rect 8268 4719 8335 4745
rect 8474 4719 8517 4753
rect 7669 4540 7696 4718
rect 7736 4680 7800 4692
rect 8076 4688 8113 4719
rect 8294 4688 8331 4719
rect 8476 4694 8517 4719
rect 8921 4777 8962 4802
rect 9107 4777 9144 4808
rect 9325 4777 9362 4808
rect 9638 4804 9702 4816
rect 9742 4778 9769 4956
rect 8921 4743 8964 4777
rect 9103 4751 9170 4777
rect 9325 4776 9405 4777
rect 9601 4776 9769 4778
rect 9325 4750 9769 4776
rect 8921 4732 8968 4743
rect 9325 4733 9360 4750
rect 9601 4749 9769 4750
rect 10232 4754 10272 4978
rect 10398 4977 10566 4978
rect 10630 5010 10663 5343
rect 10965 5330 11004 7145
rect 11140 7151 11584 7176
rect 11140 6970 11167 7151
rect 11309 7150 11584 7151
rect 11207 7110 11271 7122
rect 11547 7118 11584 7150
rect 11610 7149 11801 7171
rect 12102 7165 12211 7185
rect 12231 7165 12240 7185
rect 12102 7158 12240 7165
rect 12298 7185 12446 7194
rect 12298 7165 12307 7185
rect 12327 7165 12417 7185
rect 12437 7165 12446 7185
rect 12102 7156 12198 7158
rect 12298 7155 12446 7165
rect 12505 7185 12542 7195
rect 12505 7165 12513 7185
rect 12533 7165 12542 7185
rect 12354 7154 12390 7155
rect 11765 7147 11801 7149
rect 11765 7118 11802 7147
rect 11207 7109 11242 7110
rect 11184 7104 11242 7109
rect 11184 7084 11187 7104
rect 11207 7090 11242 7104
rect 11262 7090 11271 7110
rect 11207 7082 11271 7090
rect 11233 7081 11271 7082
rect 11234 7080 11271 7081
rect 11337 7114 11373 7115
rect 11445 7114 11481 7115
rect 11337 7106 11481 7114
rect 11337 7086 11345 7106
rect 11365 7104 11453 7106
rect 11365 7086 11398 7104
rect 11337 7082 11398 7086
rect 11421 7086 11453 7104
rect 11473 7086 11481 7106
rect 11421 7082 11481 7086
rect 11337 7080 11481 7082
rect 11547 7110 11585 7118
rect 11663 7114 11699 7115
rect 11547 7090 11556 7110
rect 11576 7090 11585 7110
rect 11547 7081 11585 7090
rect 11614 7106 11699 7114
rect 11614 7086 11671 7106
rect 11691 7086 11699 7106
rect 11547 7080 11584 7081
rect 11614 7080 11699 7086
rect 11765 7110 11803 7118
rect 11765 7090 11774 7110
rect 11794 7090 11803 7110
rect 12505 7098 12542 7165
rect 12577 7194 12608 7245
rect 12890 7233 12908 7251
rect 12926 7233 12942 7251
rect 12627 7194 12664 7195
rect 12577 7185 12664 7194
rect 12577 7165 12635 7185
rect 12655 7165 12664 7185
rect 12577 7155 12664 7165
rect 12723 7185 12760 7195
rect 12723 7165 12731 7185
rect 12751 7165 12760 7185
rect 12577 7154 12608 7155
rect 12202 7095 12239 7096
rect 12505 7095 12544 7098
rect 12201 7094 12544 7095
rect 12723 7094 12760 7165
rect 11765 7081 11803 7090
rect 12126 7089 12544 7094
rect 11765 7080 11802 7081
rect 11226 7052 11316 7058
rect 11226 7032 11242 7052
rect 11262 7050 11316 7052
rect 11262 7032 11287 7050
rect 11226 7030 11287 7032
rect 11307 7030 11316 7050
rect 11226 7024 11316 7030
rect 11239 6970 11276 6971
rect 11335 6970 11372 6971
rect 11391 6970 11427 7080
rect 11614 7059 11645 7080
rect 12126 7069 12129 7089
rect 12149 7069 12544 7089
rect 12573 7070 12760 7094
rect 11610 7058 11645 7059
rect 11488 7048 11645 7058
rect 11488 7028 11505 7048
rect 11525 7028 11645 7048
rect 11488 7021 11645 7028
rect 11712 7051 11861 7059
rect 11712 7031 11723 7051
rect 11743 7031 11782 7051
rect 11802 7031 11861 7051
rect 11712 7024 11861 7031
rect 12505 7044 12544 7069
rect 12890 7044 12942 7233
rect 13334 7261 13344 7279
rect 13362 7261 13374 7279
rect 13506 7277 13515 7297
rect 13535 7277 13544 7297
rect 13506 7269 13544 7277
rect 13610 7301 13695 7307
rect 13725 7306 13762 7307
rect 13610 7281 13618 7301
rect 13638 7281 13695 7301
rect 13610 7273 13695 7281
rect 13724 7297 13762 7306
rect 13724 7277 13733 7297
rect 13753 7277 13762 7297
rect 13610 7272 13646 7273
rect 13724 7269 13762 7277
rect 13828 7301 13972 7307
rect 13828 7281 13836 7301
rect 13856 7281 13889 7301
rect 13909 7281 13944 7301
rect 13964 7281 13972 7301
rect 13828 7273 13972 7281
rect 13828 7272 13864 7273
rect 13936 7272 13972 7273
rect 14038 7306 14075 7307
rect 14038 7305 14076 7306
rect 14038 7297 14102 7305
rect 14038 7277 14047 7297
rect 14067 7283 14102 7297
rect 14122 7283 14125 7303
rect 14067 7278 14125 7283
rect 14067 7277 14102 7278
rect 13334 7205 13374 7261
rect 13507 7240 13544 7269
rect 13508 7238 13544 7240
rect 13508 7216 13699 7238
rect 13725 7237 13762 7269
rect 14038 7265 14102 7277
rect 14142 7239 14169 7417
rect 15027 7392 15069 7437
rect 14001 7237 14169 7239
rect 13725 7227 14169 7237
rect 14310 7333 14497 7357
rect 14528 7338 14921 7358
rect 14941 7338 14944 7358
rect 14528 7333 14944 7338
rect 14310 7262 14347 7333
rect 14528 7332 14869 7333
rect 14462 7272 14493 7273
rect 14310 7242 14319 7262
rect 14339 7242 14347 7262
rect 14310 7232 14347 7242
rect 14406 7262 14493 7272
rect 14406 7242 14415 7262
rect 14435 7242 14493 7262
rect 14406 7233 14493 7242
rect 14406 7232 14443 7233
rect 13331 7200 13374 7205
rect 13722 7211 14169 7227
rect 13722 7205 13750 7211
rect 14001 7210 14169 7211
rect 13331 7197 13481 7200
rect 13722 7197 13749 7205
rect 13331 7195 13749 7197
rect 13331 7177 13340 7195
rect 13358 7177 13749 7195
rect 14462 7182 14493 7233
rect 14528 7262 14565 7332
rect 14831 7331 14868 7332
rect 14680 7272 14716 7273
rect 14528 7242 14537 7262
rect 14557 7242 14565 7262
rect 14528 7232 14565 7242
rect 14624 7262 14772 7272
rect 14872 7269 14968 7271
rect 14624 7242 14633 7262
rect 14653 7242 14743 7262
rect 14763 7242 14772 7262
rect 14624 7233 14772 7242
rect 14830 7262 14968 7269
rect 14830 7242 14839 7262
rect 14859 7242 14968 7262
rect 14830 7233 14968 7242
rect 14624 7232 14661 7233
rect 14354 7179 14395 7180
rect 13331 7174 13749 7177
rect 13331 7168 13374 7174
rect 13334 7165 13374 7168
rect 14249 7172 14395 7179
rect 13731 7156 13771 7157
rect 13442 7139 13771 7156
rect 14249 7152 14305 7172
rect 14325 7152 14364 7172
rect 14384 7152 14395 7172
rect 14249 7144 14395 7152
rect 14462 7175 14619 7182
rect 14462 7155 14582 7175
rect 14602 7155 14619 7175
rect 14462 7145 14619 7155
rect 14462 7144 14497 7145
rect 13326 7096 13369 7107
rect 13326 7078 13338 7096
rect 13356 7078 13369 7096
rect 13326 7052 13369 7078
rect 13442 7052 13469 7139
rect 13731 7130 13771 7139
rect 12505 7026 12944 7044
rect 11712 7023 11753 7024
rect 11446 6970 11483 6971
rect 11139 6961 11277 6970
rect 11139 6941 11248 6961
rect 11268 6941 11277 6961
rect 11139 6934 11277 6941
rect 11335 6961 11483 6970
rect 11335 6941 11344 6961
rect 11364 6941 11454 6961
rect 11474 6941 11483 6961
rect 11139 6932 11235 6934
rect 11335 6931 11483 6941
rect 11542 6961 11579 6971
rect 11542 6941 11550 6961
rect 11570 6941 11579 6961
rect 11391 6930 11427 6931
rect 11239 6871 11276 6872
rect 11542 6871 11579 6941
rect 11614 6970 11645 7021
rect 12505 7008 12905 7026
rect 12923 7008 12944 7026
rect 12505 7002 12944 7008
rect 12511 6998 12944 7002
rect 13326 7031 13469 7052
rect 13513 7104 13547 7120
rect 13731 7110 14124 7130
rect 14144 7110 14147 7130
rect 14462 7123 14493 7144
rect 14680 7123 14716 7233
rect 14735 7232 14772 7233
rect 14831 7232 14868 7233
rect 14791 7173 14881 7179
rect 14791 7153 14800 7173
rect 14820 7171 14881 7173
rect 14820 7153 14845 7171
rect 14791 7151 14845 7153
rect 14865 7151 14881 7171
rect 14791 7145 14881 7151
rect 14305 7122 14342 7123
rect 13731 7105 14147 7110
rect 14304 7113 14342 7122
rect 13731 7104 14072 7105
rect 13513 7034 13550 7104
rect 13665 7044 13696 7045
rect 13326 7029 13463 7031
rect 12890 6996 12942 6998
rect 13326 6987 13369 7029
rect 13513 7014 13522 7034
rect 13542 7014 13550 7034
rect 13513 7004 13550 7014
rect 13609 7034 13696 7044
rect 13609 7014 13618 7034
rect 13638 7014 13696 7034
rect 13609 7005 13696 7014
rect 13609 7004 13646 7005
rect 13324 6977 13369 6987
rect 11664 6970 11701 6971
rect 11614 6961 11701 6970
rect 11614 6941 11672 6961
rect 11692 6941 11701 6961
rect 11614 6931 11701 6941
rect 11760 6961 11797 6971
rect 11760 6941 11768 6961
rect 11788 6941 11797 6961
rect 13324 6959 13333 6977
rect 13351 6959 13369 6977
rect 13324 6953 13369 6959
rect 13665 6954 13696 7005
rect 13731 7034 13768 7104
rect 14034 7103 14071 7104
rect 14304 7093 14313 7113
rect 14333 7093 14342 7113
rect 14304 7085 14342 7093
rect 14408 7117 14493 7123
rect 14523 7122 14560 7123
rect 14408 7097 14416 7117
rect 14436 7097 14493 7117
rect 14408 7089 14493 7097
rect 14522 7113 14560 7122
rect 14522 7093 14531 7113
rect 14551 7093 14560 7113
rect 14408 7088 14444 7089
rect 14522 7085 14560 7093
rect 14626 7117 14770 7123
rect 14626 7097 14634 7117
rect 14654 7114 14742 7117
rect 14654 7097 14689 7114
rect 14626 7096 14689 7097
rect 14708 7097 14742 7114
rect 14762 7097 14770 7117
rect 14708 7096 14770 7097
rect 14626 7089 14770 7096
rect 14626 7088 14662 7089
rect 14734 7088 14770 7089
rect 14836 7122 14873 7123
rect 14836 7121 14874 7122
rect 14896 7121 14923 7125
rect 14836 7119 14923 7121
rect 14836 7113 14900 7119
rect 14836 7093 14845 7113
rect 14865 7099 14900 7113
rect 14920 7099 14923 7119
rect 14865 7094 14923 7099
rect 14865 7093 14900 7094
rect 14305 7056 14342 7085
rect 14306 7054 14342 7056
rect 13883 7044 13919 7045
rect 13731 7014 13740 7034
rect 13760 7014 13768 7034
rect 13731 7004 13768 7014
rect 13827 7034 13975 7044
rect 14075 7041 14171 7043
rect 13827 7014 13836 7034
rect 13856 7014 13946 7034
rect 13966 7014 13975 7034
rect 13827 7005 13975 7014
rect 14033 7034 14171 7041
rect 14033 7014 14042 7034
rect 14062 7014 14171 7034
rect 14306 7032 14497 7054
rect 14523 7053 14560 7085
rect 14836 7081 14900 7093
rect 14940 7055 14967 7233
rect 14799 7053 14967 7055
rect 14523 7027 14967 7053
rect 14033 7005 14171 7014
rect 13827 7004 13864 7005
rect 13324 6950 13361 6953
rect 13557 6951 13598 6952
rect 11614 6930 11645 6931
rect 11238 6870 11579 6871
rect 11760 6870 11797 6941
rect 13449 6944 13598 6951
rect 12893 6931 12930 6936
rect 11163 6865 11579 6870
rect 11163 6845 11166 6865
rect 11186 6845 11579 6865
rect 11610 6846 11797 6870
rect 12884 6927 12931 6931
rect 12884 6909 12903 6927
rect 12921 6909 12931 6927
rect 13449 6924 13508 6944
rect 13528 6924 13567 6944
rect 13587 6924 13598 6944
rect 13449 6916 13598 6924
rect 13665 6947 13822 6954
rect 13665 6927 13785 6947
rect 13805 6927 13822 6947
rect 13665 6917 13822 6927
rect 13665 6916 13700 6917
rect 12884 6861 12931 6909
rect 13665 6895 13696 6916
rect 13883 6895 13919 7005
rect 13938 7004 13975 7005
rect 14034 7004 14071 7005
rect 13994 6945 14084 6951
rect 13994 6925 14003 6945
rect 14023 6943 14084 6945
rect 14023 6925 14048 6943
rect 13994 6923 14048 6925
rect 14068 6923 14084 6943
rect 13994 6917 14084 6923
rect 13508 6894 13545 6895
rect 12508 6858 12931 6861
rect 11383 6844 11448 6845
rect 12486 6828 12931 6858
rect 13320 6886 13358 6888
rect 13320 6878 13363 6886
rect 13320 6860 13331 6878
rect 13349 6860 13363 6878
rect 13320 6833 13363 6860
rect 13507 6885 13545 6894
rect 13507 6865 13516 6885
rect 13536 6865 13545 6885
rect 13507 6857 13545 6865
rect 13611 6889 13696 6895
rect 13726 6894 13763 6895
rect 13611 6869 13619 6889
rect 13639 6869 13696 6889
rect 13611 6861 13696 6869
rect 13725 6885 13763 6894
rect 13725 6865 13734 6885
rect 13754 6865 13763 6885
rect 13611 6860 13647 6861
rect 13725 6857 13763 6865
rect 13829 6893 13973 6895
rect 13829 6889 13881 6893
rect 13829 6869 13837 6889
rect 13857 6873 13881 6889
rect 13901 6889 13973 6893
rect 13901 6873 13945 6889
rect 13857 6869 13945 6873
rect 13965 6869 13973 6889
rect 13829 6861 13973 6869
rect 13829 6860 13865 6861
rect 13937 6860 13973 6861
rect 14039 6894 14076 6895
rect 14039 6893 14077 6894
rect 14039 6885 14103 6893
rect 14039 6865 14048 6885
rect 14068 6871 14103 6885
rect 14123 6871 14126 6891
rect 14068 6866 14126 6871
rect 14068 6865 14103 6866
rect 11579 6812 11619 6820
rect 11579 6790 11587 6812
rect 11611 6790 11619 6812
rect 11184 6561 11221 6567
rect 11184 6542 11192 6561
rect 11213 6542 11221 6561
rect 11184 6534 11221 6542
rect 11188 6201 11221 6534
rect 11285 6566 11453 6567
rect 11579 6566 11619 6790
rect 12082 6794 12250 6795
rect 12486 6794 12527 6828
rect 12884 6807 12931 6828
rect 12082 6784 12527 6794
rect 12599 6792 12742 6793
rect 12082 6768 12526 6784
rect 12082 6766 12250 6768
rect 12446 6767 12526 6768
rect 12599 6767 12744 6792
rect 12886 6767 12931 6807
rect 12082 6588 12109 6766
rect 12149 6728 12213 6740
rect 12489 6736 12526 6767
rect 12707 6736 12744 6767
rect 12889 6760 12931 6767
rect 13321 6826 13363 6833
rect 13508 6826 13545 6857
rect 13726 6826 13763 6857
rect 14039 6853 14103 6865
rect 14143 6827 14170 7005
rect 13321 6786 13366 6826
rect 13508 6801 13653 6826
rect 13726 6825 13806 6826
rect 14002 6825 14170 6827
rect 13726 6809 14170 6825
rect 13510 6800 13653 6801
rect 13725 6799 14170 6809
rect 13321 6765 13368 6786
rect 13725 6765 13766 6799
rect 14002 6798 14170 6799
rect 14633 6803 14673 7027
rect 14799 7026 14967 7027
rect 15031 7059 15064 7392
rect 15669 7391 15696 7569
rect 15736 7531 15800 7543
rect 16076 7539 16113 7571
rect 16139 7570 16330 7592
rect 16465 7590 16574 7610
rect 16594 7590 16603 7610
rect 16465 7583 16603 7590
rect 16661 7610 16809 7619
rect 16661 7590 16670 7610
rect 16690 7590 16780 7610
rect 16800 7590 16809 7610
rect 16465 7581 16561 7583
rect 16661 7580 16809 7590
rect 16868 7610 16905 7620
rect 16868 7590 16876 7610
rect 16896 7590 16905 7610
rect 16717 7579 16753 7580
rect 16294 7568 16330 7570
rect 16294 7539 16331 7568
rect 15736 7530 15771 7531
rect 15713 7525 15771 7530
rect 15713 7505 15716 7525
rect 15736 7511 15771 7525
rect 15791 7511 15800 7531
rect 15736 7503 15800 7511
rect 15762 7502 15800 7503
rect 15763 7501 15800 7502
rect 15866 7535 15902 7536
rect 15974 7535 16010 7536
rect 15866 7527 16010 7535
rect 15866 7507 15874 7527
rect 15894 7526 15982 7527
rect 15894 7507 15929 7526
rect 15950 7507 15982 7526
rect 16002 7507 16010 7527
rect 15866 7501 16010 7507
rect 16076 7531 16114 7539
rect 16192 7535 16228 7536
rect 16076 7511 16085 7531
rect 16105 7511 16114 7531
rect 16076 7502 16114 7511
rect 16143 7527 16228 7535
rect 16143 7507 16200 7527
rect 16220 7507 16228 7527
rect 16076 7501 16113 7502
rect 16143 7501 16228 7507
rect 16294 7531 16332 7539
rect 16294 7511 16303 7531
rect 16323 7511 16332 7531
rect 16565 7520 16602 7521
rect 16868 7520 16905 7590
rect 16940 7619 16971 7670
rect 17267 7665 17312 7671
rect 17267 7647 17285 7665
rect 17303 7647 17312 7665
rect 17267 7637 17312 7647
rect 16990 7619 17027 7620
rect 16940 7610 17027 7619
rect 16940 7590 16998 7610
rect 17018 7590 17027 7610
rect 16940 7580 17027 7590
rect 17086 7610 17123 7620
rect 17086 7590 17094 7610
rect 17114 7590 17123 7610
rect 17267 7595 17310 7637
rect 17173 7593 17310 7595
rect 16940 7579 16971 7580
rect 17086 7520 17123 7590
rect 16564 7519 16905 7520
rect 16294 7502 16332 7511
rect 16489 7514 16905 7519
rect 16294 7501 16331 7502
rect 15755 7473 15845 7479
rect 15755 7453 15771 7473
rect 15791 7471 15845 7473
rect 15791 7453 15816 7471
rect 15755 7451 15816 7453
rect 15836 7451 15845 7471
rect 15755 7445 15845 7451
rect 15768 7391 15805 7392
rect 15864 7391 15901 7392
rect 15920 7391 15956 7501
rect 16143 7480 16174 7501
rect 16489 7494 16492 7514
rect 16512 7494 16905 7514
rect 17089 7504 17123 7520
rect 17167 7572 17310 7593
rect 16865 7485 16905 7494
rect 17167 7485 17194 7572
rect 17267 7546 17310 7572
rect 17267 7528 17280 7546
rect 17298 7528 17310 7546
rect 17267 7517 17310 7528
rect 16139 7479 16174 7480
rect 16017 7469 16174 7479
rect 16017 7449 16034 7469
rect 16054 7449 16174 7469
rect 16017 7442 16174 7449
rect 16241 7472 16390 7480
rect 16241 7452 16252 7472
rect 16272 7452 16311 7472
rect 16331 7452 16390 7472
rect 16865 7468 17194 7485
rect 16865 7467 16905 7468
rect 16241 7445 16390 7452
rect 17262 7456 17302 7459
rect 17262 7450 17305 7456
rect 16887 7447 17305 7450
rect 16241 7444 16282 7445
rect 15975 7391 16012 7392
rect 15668 7382 15806 7391
rect 15531 7372 15567 7378
rect 15531 7354 15536 7372
rect 15558 7354 15567 7372
rect 15531 7350 15567 7354
rect 15668 7362 15777 7382
rect 15797 7362 15806 7382
rect 15668 7355 15806 7362
rect 15864 7382 16012 7391
rect 15864 7362 15873 7382
rect 15893 7362 15983 7382
rect 16003 7362 16012 7382
rect 15668 7353 15764 7355
rect 15864 7352 16012 7362
rect 16071 7382 16108 7392
rect 16071 7362 16079 7382
rect 16099 7362 16108 7382
rect 15920 7351 15956 7352
rect 15534 7191 15567 7350
rect 15768 7292 15805 7293
rect 16071 7292 16108 7362
rect 16143 7391 16174 7442
rect 16887 7429 17278 7447
rect 17296 7429 17305 7447
rect 16887 7427 17305 7429
rect 16887 7419 16914 7427
rect 17155 7424 17305 7427
rect 16467 7413 16635 7414
rect 16886 7413 16914 7419
rect 16467 7397 16914 7413
rect 17262 7419 17305 7424
rect 16193 7391 16230 7392
rect 16143 7382 16230 7391
rect 16143 7362 16201 7382
rect 16221 7362 16230 7382
rect 16143 7352 16230 7362
rect 16289 7382 16326 7392
rect 16289 7362 16297 7382
rect 16317 7362 16326 7382
rect 16143 7351 16174 7352
rect 15767 7291 16108 7292
rect 16289 7291 16326 7362
rect 15692 7286 16108 7291
rect 15692 7266 15695 7286
rect 15715 7266 16108 7286
rect 16139 7267 16326 7291
rect 16467 7387 16911 7397
rect 16467 7385 16635 7387
rect 16467 7207 16494 7385
rect 16534 7347 16598 7359
rect 16874 7355 16911 7387
rect 16937 7386 17128 7408
rect 17092 7384 17128 7386
rect 17092 7355 17129 7384
rect 17262 7363 17302 7419
rect 16534 7346 16569 7347
rect 16511 7341 16569 7346
rect 16511 7321 16514 7341
rect 16534 7327 16569 7341
rect 16589 7327 16598 7347
rect 16534 7319 16598 7327
rect 16560 7318 16598 7319
rect 16561 7317 16598 7318
rect 16664 7351 16700 7352
rect 16772 7351 16808 7352
rect 16664 7343 16808 7351
rect 16664 7323 16672 7343
rect 16692 7323 16727 7343
rect 16747 7323 16780 7343
rect 16800 7323 16808 7343
rect 16664 7317 16808 7323
rect 16874 7347 16912 7355
rect 16990 7351 17026 7352
rect 16874 7327 16883 7347
rect 16903 7327 16912 7347
rect 16874 7318 16912 7327
rect 16941 7343 17026 7351
rect 16941 7323 16998 7343
rect 17018 7323 17026 7343
rect 16874 7317 16911 7318
rect 16941 7317 17026 7323
rect 17092 7347 17130 7355
rect 17092 7327 17101 7347
rect 17121 7327 17130 7347
rect 17262 7345 17274 7363
rect 17292 7345 17302 7363
rect 17262 7335 17302 7345
rect 17092 7318 17130 7327
rect 17092 7317 17129 7318
rect 16553 7289 16643 7295
rect 16553 7269 16569 7289
rect 16589 7287 16643 7289
rect 16589 7269 16614 7287
rect 16553 7267 16614 7269
rect 16634 7267 16643 7287
rect 16553 7261 16643 7267
rect 16566 7207 16603 7208
rect 16662 7207 16699 7208
rect 16718 7207 16754 7317
rect 16941 7296 16972 7317
rect 16937 7295 16972 7296
rect 16815 7285 16972 7295
rect 16815 7265 16832 7285
rect 16852 7265 16972 7285
rect 16815 7258 16972 7265
rect 17039 7288 17188 7296
rect 17039 7268 17050 7288
rect 17070 7268 17109 7288
rect 17129 7268 17188 7288
rect 17039 7261 17188 7268
rect 17254 7264 17306 7282
rect 17039 7260 17080 7261
rect 16773 7207 16810 7208
rect 16466 7198 16604 7207
rect 15533 7190 15570 7191
rect 15504 7189 15672 7190
rect 15798 7189 15838 7191
rect 15329 7180 15368 7186
rect 15329 7158 15337 7180
rect 15361 7158 15368 7180
rect 15031 7051 15068 7059
rect 15031 7032 15039 7051
rect 15060 7032 15068 7051
rect 15031 7026 15068 7032
rect 14633 6781 14641 6803
rect 14665 6781 14673 6803
rect 14633 6773 14673 6781
rect 12149 6727 12184 6728
rect 12126 6722 12184 6727
rect 12126 6702 12129 6722
rect 12149 6708 12184 6722
rect 12204 6708 12213 6728
rect 12149 6700 12213 6708
rect 12175 6699 12213 6700
rect 12176 6698 12213 6699
rect 12279 6732 12315 6733
rect 12387 6732 12423 6733
rect 12279 6724 12423 6732
rect 12279 6704 12287 6724
rect 12307 6720 12395 6724
rect 12307 6704 12351 6720
rect 12279 6700 12351 6704
rect 12371 6704 12395 6720
rect 12415 6704 12423 6724
rect 12371 6700 12423 6704
rect 12279 6698 12423 6700
rect 12489 6728 12527 6736
rect 12605 6732 12641 6733
rect 12489 6708 12498 6728
rect 12518 6708 12527 6728
rect 12489 6699 12527 6708
rect 12556 6724 12641 6732
rect 12556 6704 12613 6724
rect 12633 6704 12641 6724
rect 12489 6698 12526 6699
rect 12556 6698 12641 6704
rect 12707 6728 12745 6736
rect 12707 6708 12716 6728
rect 12736 6708 12745 6728
rect 12707 6699 12745 6708
rect 12889 6733 12932 6760
rect 12889 6715 12903 6733
rect 12921 6715 12932 6733
rect 12889 6707 12932 6715
rect 12894 6705 12932 6707
rect 13321 6735 13766 6765
rect 14804 6748 14869 6749
rect 13321 6732 13744 6735
rect 12707 6698 12744 6699
rect 12168 6670 12258 6676
rect 12168 6650 12184 6670
rect 12204 6668 12258 6670
rect 12204 6650 12229 6668
rect 12168 6648 12229 6650
rect 12249 6648 12258 6668
rect 12168 6642 12258 6648
rect 12181 6588 12218 6589
rect 12277 6588 12314 6589
rect 12333 6588 12369 6698
rect 12556 6677 12587 6698
rect 13321 6684 13368 6732
rect 12552 6676 12587 6677
rect 12430 6666 12587 6676
rect 12430 6646 12447 6666
rect 12467 6646 12587 6666
rect 12430 6639 12587 6646
rect 12654 6669 12803 6677
rect 12654 6649 12665 6669
rect 12685 6649 12724 6669
rect 12744 6649 12803 6669
rect 13321 6666 13331 6684
rect 13349 6666 13368 6684
rect 13321 6662 13368 6666
rect 14455 6723 14642 6747
rect 14673 6728 15066 6748
rect 15086 6728 15089 6748
rect 14673 6723 15089 6728
rect 13322 6657 13359 6662
rect 12654 6642 12803 6649
rect 14455 6652 14492 6723
rect 14673 6722 15014 6723
rect 14607 6662 14638 6663
rect 12654 6641 12695 6642
rect 12891 6640 12928 6643
rect 12388 6588 12425 6589
rect 12081 6579 12219 6588
rect 11285 6540 11729 6566
rect 11285 6538 11453 6540
rect 11285 6360 11312 6538
rect 11352 6500 11416 6512
rect 11692 6508 11729 6540
rect 11755 6539 11946 6561
rect 12081 6559 12190 6579
rect 12210 6559 12219 6579
rect 12081 6552 12219 6559
rect 12277 6579 12425 6588
rect 12277 6559 12286 6579
rect 12306 6559 12396 6579
rect 12416 6559 12425 6579
rect 12081 6550 12177 6552
rect 12277 6549 12425 6559
rect 12484 6579 12521 6589
rect 12484 6559 12492 6579
rect 12512 6559 12521 6579
rect 12333 6548 12369 6549
rect 11910 6537 11946 6539
rect 11910 6508 11947 6537
rect 11352 6499 11387 6500
rect 11329 6494 11387 6499
rect 11329 6474 11332 6494
rect 11352 6480 11387 6494
rect 11407 6480 11416 6500
rect 11352 6474 11416 6480
rect 11329 6472 11416 6474
rect 11329 6468 11356 6472
rect 11378 6471 11416 6472
rect 11379 6470 11416 6471
rect 11482 6504 11518 6505
rect 11590 6504 11626 6505
rect 11482 6497 11626 6504
rect 11482 6496 11544 6497
rect 11482 6476 11490 6496
rect 11510 6479 11544 6496
rect 11563 6496 11626 6497
rect 11563 6479 11598 6496
rect 11510 6476 11598 6479
rect 11618 6476 11626 6496
rect 11482 6470 11626 6476
rect 11692 6500 11730 6508
rect 11808 6504 11844 6505
rect 11692 6480 11701 6500
rect 11721 6480 11730 6500
rect 11692 6471 11730 6480
rect 11759 6496 11844 6504
rect 11759 6476 11816 6496
rect 11836 6476 11844 6496
rect 11692 6470 11729 6471
rect 11759 6470 11844 6476
rect 11910 6500 11948 6508
rect 11910 6480 11919 6500
rect 11939 6480 11948 6500
rect 12181 6489 12218 6490
rect 12484 6489 12521 6559
rect 12556 6588 12587 6639
rect 12883 6634 12928 6640
rect 12883 6616 12901 6634
rect 12919 6616 12928 6634
rect 14455 6632 14464 6652
rect 14484 6632 14492 6652
rect 14455 6622 14492 6632
rect 14551 6652 14638 6662
rect 14551 6632 14560 6652
rect 14580 6632 14638 6652
rect 14551 6623 14638 6632
rect 14551 6622 14588 6623
rect 12883 6606 12928 6616
rect 12606 6588 12643 6589
rect 12556 6579 12643 6588
rect 12556 6559 12614 6579
rect 12634 6559 12643 6579
rect 12556 6549 12643 6559
rect 12702 6579 12739 6589
rect 12702 6559 12710 6579
rect 12730 6559 12739 6579
rect 12883 6564 12926 6606
rect 13310 6595 13362 6597
rect 12789 6562 12926 6564
rect 12556 6548 12587 6549
rect 12702 6489 12739 6559
rect 12180 6488 12521 6489
rect 11910 6471 11948 6480
rect 12105 6483 12521 6488
rect 11910 6470 11947 6471
rect 11371 6442 11461 6448
rect 11371 6422 11387 6442
rect 11407 6440 11461 6442
rect 11407 6422 11432 6440
rect 11371 6420 11432 6422
rect 11452 6420 11461 6440
rect 11371 6414 11461 6420
rect 11384 6360 11421 6361
rect 11480 6360 11517 6361
rect 11536 6360 11572 6470
rect 11759 6449 11790 6470
rect 12105 6463 12108 6483
rect 12128 6463 12521 6483
rect 12705 6473 12739 6489
rect 12783 6541 12926 6562
rect 13308 6591 13741 6595
rect 13308 6585 13747 6591
rect 13308 6567 13329 6585
rect 13347 6567 13747 6585
rect 14607 6572 14638 6623
rect 14673 6652 14710 6722
rect 14976 6721 15013 6722
rect 14825 6662 14861 6663
rect 14673 6632 14682 6652
rect 14702 6632 14710 6652
rect 14673 6622 14710 6632
rect 14769 6652 14917 6662
rect 15017 6659 15113 6661
rect 14769 6632 14778 6652
rect 14798 6632 14888 6652
rect 14908 6632 14917 6652
rect 14769 6623 14917 6632
rect 14975 6652 15113 6659
rect 14975 6632 14984 6652
rect 15004 6632 15113 6652
rect 14975 6623 15113 6632
rect 14769 6622 14806 6623
rect 14499 6569 14540 6570
rect 13308 6549 13747 6567
rect 12481 6454 12521 6463
rect 12783 6454 12810 6541
rect 12883 6515 12926 6541
rect 12883 6497 12896 6515
rect 12914 6497 12926 6515
rect 12883 6486 12926 6497
rect 11755 6448 11790 6449
rect 11633 6438 11790 6448
rect 11633 6418 11650 6438
rect 11670 6418 11790 6438
rect 11633 6411 11790 6418
rect 11857 6441 12003 6449
rect 11857 6421 11868 6441
rect 11888 6421 11927 6441
rect 11947 6421 12003 6441
rect 12481 6437 12810 6454
rect 12481 6436 12521 6437
rect 11857 6414 12003 6421
rect 12878 6425 12918 6428
rect 12878 6419 12921 6425
rect 12503 6416 12921 6419
rect 11857 6413 11898 6414
rect 11591 6360 11628 6361
rect 11284 6351 11422 6360
rect 11284 6331 11393 6351
rect 11413 6331 11422 6351
rect 11284 6324 11422 6331
rect 11480 6351 11628 6360
rect 11480 6331 11489 6351
rect 11509 6331 11599 6351
rect 11619 6331 11628 6351
rect 11284 6322 11380 6324
rect 11480 6321 11628 6331
rect 11687 6351 11724 6361
rect 11687 6331 11695 6351
rect 11715 6331 11724 6351
rect 11536 6320 11572 6321
rect 11384 6261 11421 6262
rect 11687 6261 11724 6331
rect 11759 6360 11790 6411
rect 12503 6398 12894 6416
rect 12912 6398 12921 6416
rect 12503 6396 12921 6398
rect 12503 6388 12530 6396
rect 12771 6393 12921 6396
rect 12083 6382 12251 6383
rect 12502 6382 12530 6388
rect 12083 6366 12530 6382
rect 12878 6388 12921 6393
rect 11809 6360 11846 6361
rect 11759 6351 11846 6360
rect 11759 6331 11817 6351
rect 11837 6331 11846 6351
rect 11759 6321 11846 6331
rect 11905 6351 11942 6361
rect 11905 6331 11913 6351
rect 11933 6331 11942 6351
rect 11759 6320 11790 6321
rect 11383 6260 11724 6261
rect 11905 6260 11942 6331
rect 11308 6255 11724 6260
rect 11308 6235 11311 6255
rect 11331 6235 11724 6255
rect 11755 6236 11942 6260
rect 12083 6356 12527 6366
rect 12083 6354 12251 6356
rect 11183 6156 11225 6201
rect 12083 6176 12110 6354
rect 12150 6316 12214 6328
rect 12490 6324 12527 6356
rect 12553 6355 12744 6377
rect 12708 6353 12744 6355
rect 12708 6324 12745 6353
rect 12878 6332 12918 6388
rect 12150 6315 12185 6316
rect 12127 6310 12185 6315
rect 12127 6290 12130 6310
rect 12150 6296 12185 6310
rect 12205 6296 12214 6316
rect 12150 6288 12214 6296
rect 12176 6287 12214 6288
rect 12177 6286 12214 6287
rect 12280 6320 12316 6321
rect 12388 6320 12424 6321
rect 12280 6312 12424 6320
rect 12280 6292 12288 6312
rect 12308 6292 12343 6312
rect 12363 6292 12396 6312
rect 12416 6292 12424 6312
rect 12280 6286 12424 6292
rect 12490 6316 12528 6324
rect 12606 6320 12642 6321
rect 12490 6296 12499 6316
rect 12519 6296 12528 6316
rect 12490 6287 12528 6296
rect 12557 6312 12642 6320
rect 12557 6292 12614 6312
rect 12634 6292 12642 6312
rect 12490 6286 12527 6287
rect 12557 6286 12642 6292
rect 12708 6316 12746 6324
rect 12708 6296 12717 6316
rect 12737 6296 12746 6316
rect 12878 6314 12890 6332
rect 12908 6314 12918 6332
rect 13310 6360 13362 6549
rect 13708 6524 13747 6549
rect 14391 6562 14540 6569
rect 14391 6542 14450 6562
rect 14470 6542 14509 6562
rect 14529 6542 14540 6562
rect 14391 6534 14540 6542
rect 14607 6565 14764 6572
rect 14607 6545 14727 6565
rect 14747 6545 14764 6565
rect 14607 6535 14764 6545
rect 14607 6534 14642 6535
rect 13492 6499 13679 6523
rect 13708 6504 14103 6524
rect 14123 6504 14126 6524
rect 14607 6513 14638 6534
rect 14825 6513 14861 6623
rect 14880 6622 14917 6623
rect 14976 6622 15013 6623
rect 14936 6563 15026 6569
rect 14936 6543 14945 6563
rect 14965 6561 15026 6563
rect 14965 6543 14990 6561
rect 14936 6541 14990 6543
rect 15010 6541 15026 6561
rect 14936 6535 15026 6541
rect 14450 6512 14487 6513
rect 13708 6499 14126 6504
rect 14449 6503 14487 6512
rect 13492 6428 13529 6499
rect 13708 6498 14051 6499
rect 13708 6495 13747 6498
rect 14013 6497 14050 6498
rect 13644 6438 13675 6439
rect 13492 6408 13501 6428
rect 13521 6408 13529 6428
rect 13492 6398 13529 6408
rect 13588 6428 13675 6438
rect 13588 6408 13597 6428
rect 13617 6408 13675 6428
rect 13588 6399 13675 6408
rect 13588 6398 13625 6399
rect 13310 6342 13326 6360
rect 13344 6342 13362 6360
rect 13644 6348 13675 6399
rect 13710 6428 13747 6495
rect 14449 6483 14458 6503
rect 14478 6483 14487 6503
rect 14449 6475 14487 6483
rect 14553 6507 14638 6513
rect 14668 6512 14705 6513
rect 14553 6487 14561 6507
rect 14581 6487 14638 6507
rect 14553 6479 14638 6487
rect 14667 6503 14705 6512
rect 14667 6483 14676 6503
rect 14696 6483 14705 6503
rect 14553 6478 14589 6479
rect 14667 6475 14705 6483
rect 14771 6507 14915 6513
rect 14771 6487 14779 6507
rect 14799 6506 14887 6507
rect 14799 6488 14834 6506
rect 14852 6488 14887 6506
rect 14799 6487 14887 6488
rect 14907 6487 14915 6507
rect 14771 6479 14915 6487
rect 14771 6478 14807 6479
rect 14879 6478 14915 6479
rect 14981 6512 15018 6513
rect 14981 6511 15019 6512
rect 14981 6503 15045 6511
rect 14981 6483 14990 6503
rect 15010 6489 15045 6503
rect 15065 6489 15068 6509
rect 15010 6484 15068 6489
rect 15010 6483 15045 6484
rect 14450 6446 14487 6475
rect 14451 6444 14487 6446
rect 13862 6438 13898 6439
rect 13710 6408 13719 6428
rect 13739 6408 13747 6428
rect 13710 6398 13747 6408
rect 13806 6428 13954 6438
rect 14054 6435 14150 6437
rect 13806 6408 13815 6428
rect 13835 6408 13925 6428
rect 13945 6408 13954 6428
rect 13806 6399 13954 6408
rect 14012 6428 14150 6435
rect 14012 6408 14021 6428
rect 14041 6408 14150 6428
rect 14451 6422 14642 6444
rect 14668 6443 14705 6475
rect 14981 6471 15045 6483
rect 15085 6447 15112 6623
rect 15031 6445 15112 6447
rect 14944 6443 15112 6445
rect 14668 6417 15112 6443
rect 14778 6415 14818 6417
rect 14944 6416 15112 6417
rect 14012 6399 14150 6408
rect 15053 6414 15112 6416
rect 13806 6398 13843 6399
rect 13536 6345 13577 6346
rect 13310 6324 13362 6342
rect 13428 6338 13577 6345
rect 12878 6304 12918 6314
rect 13428 6318 13487 6338
rect 13507 6318 13546 6338
rect 13566 6318 13577 6338
rect 13428 6310 13577 6318
rect 13644 6341 13801 6348
rect 13644 6321 13764 6341
rect 13784 6321 13801 6341
rect 13644 6311 13801 6321
rect 13644 6310 13679 6311
rect 12708 6287 12746 6296
rect 13644 6289 13675 6310
rect 13862 6289 13898 6399
rect 13917 6398 13954 6399
rect 14013 6398 14050 6399
rect 13973 6339 14063 6345
rect 13973 6319 13982 6339
rect 14002 6337 14063 6339
rect 14002 6319 14027 6337
rect 13973 6317 14027 6319
rect 14047 6317 14063 6337
rect 13973 6311 14063 6317
rect 13487 6288 13524 6289
rect 12708 6286 12745 6287
rect 12169 6258 12259 6264
rect 12169 6238 12185 6258
rect 12205 6256 12259 6258
rect 12205 6238 12230 6256
rect 12169 6236 12230 6238
rect 12250 6236 12259 6256
rect 12169 6230 12259 6236
rect 12182 6176 12219 6177
rect 12278 6176 12315 6177
rect 12334 6176 12370 6286
rect 12557 6265 12588 6286
rect 13486 6279 13524 6288
rect 12553 6264 12588 6265
rect 12431 6254 12588 6264
rect 12431 6234 12448 6254
rect 12468 6234 12588 6254
rect 12431 6227 12588 6234
rect 12655 6257 12804 6265
rect 12655 6237 12666 6257
rect 12686 6237 12725 6257
rect 12745 6237 12804 6257
rect 13314 6261 13354 6271
rect 12655 6230 12804 6237
rect 12870 6233 12922 6251
rect 12655 6229 12696 6230
rect 12389 6176 12426 6177
rect 12082 6167 12220 6176
rect 11554 6156 11587 6158
rect 11183 6144 11630 6156
rect 11186 6130 11630 6144
rect 11186 6128 11354 6130
rect 11186 5950 11213 6128
rect 11253 6090 11317 6102
rect 11593 6098 11630 6130
rect 11656 6129 11847 6151
rect 12082 6147 12191 6167
rect 12211 6147 12220 6167
rect 12082 6140 12220 6147
rect 12278 6167 12426 6176
rect 12278 6147 12287 6167
rect 12307 6147 12397 6167
rect 12417 6147 12426 6167
rect 12082 6138 12178 6140
rect 12278 6137 12426 6147
rect 12485 6167 12522 6177
rect 12485 6147 12493 6167
rect 12513 6147 12522 6167
rect 12334 6136 12370 6137
rect 11811 6127 11847 6129
rect 11811 6098 11848 6127
rect 11253 6089 11288 6090
rect 11230 6084 11288 6089
rect 11230 6064 11233 6084
rect 11253 6070 11288 6084
rect 11308 6070 11317 6090
rect 11253 6062 11317 6070
rect 11279 6061 11317 6062
rect 11280 6060 11317 6061
rect 11383 6094 11419 6095
rect 11491 6094 11527 6095
rect 11383 6086 11527 6094
rect 11383 6066 11391 6086
rect 11411 6084 11499 6086
rect 11411 6066 11444 6084
rect 11383 6065 11444 6066
rect 11465 6066 11499 6084
rect 11519 6066 11527 6086
rect 11465 6065 11527 6066
rect 11383 6060 11527 6065
rect 11593 6090 11631 6098
rect 11709 6094 11745 6095
rect 11593 6070 11602 6090
rect 11622 6070 11631 6090
rect 11593 6061 11631 6070
rect 11660 6086 11745 6094
rect 11660 6066 11717 6086
rect 11737 6066 11745 6086
rect 11593 6060 11630 6061
rect 11660 6060 11745 6066
rect 11811 6090 11849 6098
rect 11811 6070 11820 6090
rect 11840 6070 11849 6090
rect 12485 6080 12522 6147
rect 12557 6176 12588 6227
rect 12870 6215 12888 6233
rect 12906 6215 12922 6233
rect 12607 6176 12644 6177
rect 12557 6167 12644 6176
rect 12557 6147 12615 6167
rect 12635 6147 12644 6167
rect 12557 6137 12644 6147
rect 12703 6167 12740 6177
rect 12703 6147 12711 6167
rect 12731 6147 12740 6167
rect 12557 6136 12588 6137
rect 12182 6077 12219 6078
rect 12485 6077 12524 6080
rect 12181 6076 12524 6077
rect 12703 6076 12740 6147
rect 11811 6061 11849 6070
rect 12106 6071 12524 6076
rect 11811 6060 11848 6061
rect 11272 6032 11362 6038
rect 11272 6012 11288 6032
rect 11308 6030 11362 6032
rect 11308 6012 11333 6030
rect 11272 6010 11333 6012
rect 11353 6010 11362 6030
rect 11272 6004 11362 6010
rect 11285 5950 11322 5951
rect 11381 5950 11418 5951
rect 11437 5950 11473 6060
rect 11660 6039 11691 6060
rect 12106 6051 12109 6071
rect 12129 6051 12524 6071
rect 12553 6052 12740 6076
rect 11656 6038 11691 6039
rect 11534 6028 11691 6038
rect 11534 6008 11551 6028
rect 11571 6008 11691 6028
rect 11534 6001 11691 6008
rect 11758 6031 11907 6039
rect 11758 6011 11769 6031
rect 11789 6011 11828 6031
rect 11848 6011 11907 6031
rect 11758 6004 11907 6011
rect 12485 6026 12524 6051
rect 12870 6026 12922 6215
rect 13314 6243 13324 6261
rect 13342 6243 13354 6261
rect 13486 6259 13495 6279
rect 13515 6259 13524 6279
rect 13486 6251 13524 6259
rect 13590 6283 13675 6289
rect 13705 6288 13742 6289
rect 13590 6263 13598 6283
rect 13618 6263 13675 6283
rect 13590 6255 13675 6263
rect 13704 6279 13742 6288
rect 13704 6259 13713 6279
rect 13733 6259 13742 6279
rect 13590 6254 13626 6255
rect 13704 6251 13742 6259
rect 13808 6283 13952 6289
rect 13808 6263 13816 6283
rect 13836 6263 13869 6283
rect 13889 6263 13924 6283
rect 13944 6263 13952 6283
rect 13808 6255 13952 6263
rect 13808 6254 13844 6255
rect 13916 6254 13952 6255
rect 14018 6288 14055 6289
rect 14018 6287 14056 6288
rect 14018 6279 14082 6287
rect 14018 6259 14027 6279
rect 14047 6265 14082 6279
rect 14102 6265 14105 6285
rect 14047 6260 14105 6265
rect 14047 6259 14082 6260
rect 13314 6187 13354 6243
rect 13487 6222 13524 6251
rect 13488 6220 13524 6222
rect 13488 6198 13679 6220
rect 13705 6219 13742 6251
rect 14018 6247 14082 6259
rect 14122 6221 14149 6399
rect 15053 6396 15082 6414
rect 13981 6219 14149 6221
rect 13705 6209 14149 6219
rect 14290 6315 14477 6339
rect 14508 6320 14901 6340
rect 14921 6320 14924 6340
rect 14508 6315 14924 6320
rect 14290 6244 14327 6315
rect 14508 6314 14849 6315
rect 14442 6254 14473 6255
rect 14290 6224 14299 6244
rect 14319 6224 14327 6244
rect 14290 6214 14327 6224
rect 14386 6244 14473 6254
rect 14386 6224 14395 6244
rect 14415 6224 14473 6244
rect 14386 6215 14473 6224
rect 14386 6214 14423 6215
rect 13311 6182 13354 6187
rect 13702 6193 14149 6209
rect 13702 6187 13730 6193
rect 13981 6192 14149 6193
rect 13311 6179 13461 6182
rect 13702 6179 13729 6187
rect 13311 6177 13729 6179
rect 13311 6159 13320 6177
rect 13338 6159 13729 6177
rect 14442 6164 14473 6215
rect 14508 6244 14545 6314
rect 14811 6313 14848 6314
rect 14660 6254 14696 6255
rect 14508 6224 14517 6244
rect 14537 6224 14545 6244
rect 14508 6214 14545 6224
rect 14604 6244 14752 6254
rect 14852 6251 14948 6253
rect 14604 6224 14613 6244
rect 14633 6224 14723 6244
rect 14743 6224 14752 6244
rect 14604 6215 14752 6224
rect 14810 6244 14948 6251
rect 14810 6224 14819 6244
rect 14839 6224 14948 6244
rect 14810 6215 14948 6224
rect 14604 6214 14641 6215
rect 14334 6161 14375 6162
rect 13311 6156 13729 6159
rect 13311 6150 13354 6156
rect 13314 6147 13354 6150
rect 14226 6154 14375 6161
rect 13711 6138 13751 6139
rect 13422 6121 13751 6138
rect 14226 6134 14285 6154
rect 14305 6134 14344 6154
rect 14364 6134 14375 6154
rect 14226 6126 14375 6134
rect 14442 6157 14599 6164
rect 14442 6137 14562 6157
rect 14582 6137 14599 6157
rect 14442 6127 14599 6137
rect 14442 6126 14477 6127
rect 13306 6078 13349 6089
rect 13306 6060 13318 6078
rect 13336 6060 13349 6078
rect 13306 6034 13349 6060
rect 13422 6034 13449 6121
rect 13711 6112 13751 6121
rect 12485 6008 12924 6026
rect 11758 6003 11799 6004
rect 11492 5950 11529 5951
rect 11185 5941 11323 5950
rect 11185 5921 11294 5941
rect 11314 5921 11323 5941
rect 11185 5914 11323 5921
rect 11381 5941 11529 5950
rect 11381 5921 11390 5941
rect 11410 5921 11500 5941
rect 11520 5921 11529 5941
rect 11185 5912 11281 5914
rect 11381 5911 11529 5921
rect 11588 5941 11625 5951
rect 11588 5921 11596 5941
rect 11616 5921 11625 5941
rect 11437 5910 11473 5911
rect 11285 5851 11322 5852
rect 11588 5851 11625 5921
rect 11660 5950 11691 6001
rect 12485 5990 12885 6008
rect 12903 5990 12924 6008
rect 12485 5984 12924 5990
rect 12491 5980 12924 5984
rect 13306 6013 13449 6034
rect 13493 6086 13527 6102
rect 13711 6092 14104 6112
rect 14124 6092 14127 6112
rect 14442 6105 14473 6126
rect 14660 6105 14696 6215
rect 14715 6214 14752 6215
rect 14811 6214 14848 6215
rect 14771 6155 14861 6161
rect 14771 6135 14780 6155
rect 14800 6153 14861 6155
rect 14800 6135 14825 6153
rect 14771 6133 14825 6135
rect 14845 6133 14861 6153
rect 14771 6127 14861 6133
rect 14285 6104 14322 6105
rect 13711 6087 14127 6092
rect 14284 6095 14322 6104
rect 13711 6086 14052 6087
rect 13493 6016 13530 6086
rect 13645 6026 13676 6027
rect 13306 6011 13443 6013
rect 12870 5978 12922 5980
rect 13306 5969 13349 6011
rect 13493 5996 13502 6016
rect 13522 5996 13530 6016
rect 13493 5986 13530 5996
rect 13589 6016 13676 6026
rect 13589 5996 13598 6016
rect 13618 5996 13676 6016
rect 13589 5987 13676 5996
rect 13589 5986 13626 5987
rect 13304 5959 13349 5969
rect 11710 5950 11747 5951
rect 11660 5941 11747 5950
rect 11660 5921 11718 5941
rect 11738 5921 11747 5941
rect 11660 5911 11747 5921
rect 11806 5941 11843 5951
rect 11806 5921 11814 5941
rect 11834 5921 11843 5941
rect 13304 5941 13313 5959
rect 13331 5941 13349 5959
rect 13304 5935 13349 5941
rect 13645 5936 13676 5987
rect 13711 6016 13748 6086
rect 14014 6085 14051 6086
rect 14284 6075 14293 6095
rect 14313 6075 14322 6095
rect 14284 6067 14322 6075
rect 14388 6099 14473 6105
rect 14503 6104 14540 6105
rect 14388 6079 14396 6099
rect 14416 6079 14473 6099
rect 14388 6071 14473 6079
rect 14502 6095 14540 6104
rect 14502 6075 14511 6095
rect 14531 6075 14540 6095
rect 14388 6070 14424 6071
rect 14502 6067 14540 6075
rect 14606 6099 14750 6105
rect 14606 6079 14614 6099
rect 14634 6080 14666 6099
rect 14687 6080 14722 6099
rect 14634 6079 14722 6080
rect 14742 6079 14750 6099
rect 14606 6071 14750 6079
rect 14606 6070 14642 6071
rect 14714 6070 14750 6071
rect 14816 6104 14853 6105
rect 14816 6103 14854 6104
rect 14816 6095 14880 6103
rect 14816 6075 14825 6095
rect 14845 6081 14880 6095
rect 14900 6081 14903 6101
rect 14845 6076 14903 6081
rect 14845 6075 14880 6076
rect 14285 6038 14322 6067
rect 14286 6036 14322 6038
rect 13863 6026 13899 6027
rect 13711 5996 13720 6016
rect 13740 5996 13748 6016
rect 13711 5986 13748 5996
rect 13807 6016 13955 6026
rect 14055 6023 14151 6025
rect 13807 5996 13816 6016
rect 13836 5996 13926 6016
rect 13946 5996 13955 6016
rect 13807 5987 13955 5996
rect 14013 6016 14151 6023
rect 14013 5996 14022 6016
rect 14042 5996 14151 6016
rect 14286 6014 14477 6036
rect 14503 6035 14540 6067
rect 14816 6063 14880 6075
rect 14920 6037 14947 6215
rect 14779 6035 14947 6037
rect 14503 6009 14947 6035
rect 14013 5987 14151 5996
rect 13807 5986 13844 5987
rect 13304 5932 13341 5935
rect 13537 5933 13578 5934
rect 11660 5910 11691 5911
rect 11284 5850 11625 5851
rect 11806 5850 11843 5921
rect 13429 5926 13578 5933
rect 12873 5913 12910 5918
rect 12864 5909 12911 5913
rect 12864 5891 12883 5909
rect 12901 5891 12911 5909
rect 13429 5906 13488 5926
rect 13508 5906 13547 5926
rect 13567 5906 13578 5926
rect 13429 5898 13578 5906
rect 13645 5929 13802 5936
rect 13645 5909 13765 5929
rect 13785 5909 13802 5929
rect 13645 5899 13802 5909
rect 13645 5898 13680 5899
rect 11209 5845 11625 5850
rect 11209 5825 11212 5845
rect 11232 5825 11625 5845
rect 11656 5826 11843 5850
rect 12468 5848 12508 5853
rect 12864 5848 12911 5891
rect 13645 5877 13676 5898
rect 13863 5877 13899 5987
rect 13918 5986 13955 5987
rect 14014 5986 14051 5987
rect 13974 5927 14064 5933
rect 13974 5907 13983 5927
rect 14003 5925 14064 5927
rect 14003 5907 14028 5925
rect 13974 5905 14028 5907
rect 14048 5905 14064 5925
rect 13974 5899 14064 5905
rect 13488 5876 13525 5877
rect 12468 5809 12911 5848
rect 13301 5868 13338 5870
rect 13301 5860 13343 5868
rect 13301 5842 13311 5860
rect 13329 5842 13343 5860
rect 13301 5833 13343 5842
rect 13487 5867 13525 5876
rect 13487 5847 13496 5867
rect 13516 5847 13525 5867
rect 13487 5839 13525 5847
rect 13591 5871 13676 5877
rect 13706 5876 13743 5877
rect 13591 5851 13599 5871
rect 13619 5851 13676 5871
rect 13591 5843 13676 5851
rect 13705 5867 13743 5876
rect 13705 5847 13714 5867
rect 13734 5847 13743 5867
rect 13591 5842 13627 5843
rect 13705 5839 13743 5847
rect 13809 5875 13953 5877
rect 13809 5871 13861 5875
rect 13809 5851 13817 5871
rect 13837 5855 13861 5871
rect 13881 5871 13953 5875
rect 13881 5855 13925 5871
rect 13837 5851 13925 5855
rect 13945 5851 13953 5871
rect 13809 5843 13953 5851
rect 13809 5842 13845 5843
rect 13917 5842 13953 5843
rect 14019 5876 14056 5877
rect 14019 5875 14057 5876
rect 14019 5867 14083 5875
rect 14019 5847 14028 5867
rect 14048 5853 14083 5867
rect 14103 5853 14106 5873
rect 14048 5848 14106 5853
rect 14048 5847 14083 5848
rect 11562 5794 11602 5802
rect 11562 5772 11570 5794
rect 11594 5772 11602 5794
rect 11268 5548 11436 5549
rect 11562 5548 11602 5772
rect 12065 5776 12233 5777
rect 12468 5776 12508 5809
rect 12864 5776 12911 5809
rect 13302 5808 13343 5833
rect 13488 5808 13525 5839
rect 13706 5808 13743 5839
rect 14019 5835 14083 5847
rect 14123 5809 14150 5987
rect 13302 5781 13351 5808
rect 13487 5782 13536 5808
rect 13705 5807 13786 5808
rect 13982 5807 14150 5809
rect 13705 5782 14150 5807
rect 13706 5781 14150 5782
rect 12065 5775 12509 5776
rect 12065 5750 12510 5775
rect 12065 5748 12233 5750
rect 12429 5749 12510 5750
rect 12679 5749 12728 5775
rect 12864 5749 12913 5776
rect 12065 5570 12092 5748
rect 12132 5710 12196 5722
rect 12472 5718 12509 5749
rect 12690 5718 12727 5749
rect 12872 5724 12913 5749
rect 13304 5748 13351 5781
rect 13707 5748 13747 5781
rect 13982 5780 14150 5781
rect 14613 5785 14653 6009
rect 14779 6008 14947 6009
rect 14613 5763 14621 5785
rect 14645 5763 14653 5785
rect 14613 5755 14653 5763
rect 12132 5709 12167 5710
rect 12109 5704 12167 5709
rect 12109 5684 12112 5704
rect 12132 5690 12167 5704
rect 12187 5690 12196 5710
rect 12132 5682 12196 5690
rect 12158 5681 12196 5682
rect 12159 5680 12196 5681
rect 12262 5714 12298 5715
rect 12370 5714 12406 5715
rect 12262 5706 12406 5714
rect 12262 5686 12270 5706
rect 12290 5702 12378 5706
rect 12290 5686 12334 5702
rect 12262 5682 12334 5686
rect 12354 5686 12378 5702
rect 12398 5686 12406 5706
rect 12354 5682 12406 5686
rect 12262 5680 12406 5682
rect 12472 5710 12510 5718
rect 12588 5714 12624 5715
rect 12472 5690 12481 5710
rect 12501 5690 12510 5710
rect 12472 5681 12510 5690
rect 12539 5706 12624 5714
rect 12539 5686 12596 5706
rect 12616 5686 12624 5706
rect 12472 5680 12509 5681
rect 12539 5680 12624 5686
rect 12690 5710 12728 5718
rect 12690 5690 12699 5710
rect 12719 5690 12728 5710
rect 12690 5681 12728 5690
rect 12872 5715 12914 5724
rect 12872 5697 12886 5715
rect 12904 5697 12914 5715
rect 12872 5689 12914 5697
rect 12877 5687 12914 5689
rect 13304 5709 13747 5748
rect 12690 5680 12727 5681
rect 12151 5652 12241 5658
rect 12151 5632 12167 5652
rect 12187 5650 12241 5652
rect 12187 5632 12212 5650
rect 12151 5630 12212 5632
rect 12232 5630 12241 5650
rect 12151 5624 12241 5630
rect 12164 5570 12201 5571
rect 12260 5570 12297 5571
rect 12316 5570 12352 5680
rect 12539 5659 12570 5680
rect 13304 5666 13351 5709
rect 13707 5704 13747 5709
rect 14372 5707 14559 5731
rect 14590 5712 14983 5732
rect 15003 5712 15006 5732
rect 14590 5707 15006 5712
rect 12535 5658 12570 5659
rect 12413 5648 12570 5658
rect 12413 5628 12430 5648
rect 12450 5628 12570 5648
rect 12413 5621 12570 5628
rect 12637 5651 12786 5659
rect 12637 5631 12648 5651
rect 12668 5631 12707 5651
rect 12727 5631 12786 5651
rect 13304 5648 13314 5666
rect 13332 5648 13351 5666
rect 13304 5644 13351 5648
rect 13305 5639 13342 5644
rect 12637 5624 12786 5631
rect 14372 5636 14409 5707
rect 14590 5706 14931 5707
rect 14524 5646 14555 5647
rect 12637 5623 12678 5624
rect 12874 5622 12911 5625
rect 12371 5570 12408 5571
rect 12064 5561 12202 5570
rect 11268 5522 11712 5548
rect 11268 5520 11436 5522
rect 11268 5342 11295 5520
rect 11335 5482 11399 5494
rect 11675 5490 11712 5522
rect 11738 5521 11929 5543
rect 12064 5541 12173 5561
rect 12193 5541 12202 5561
rect 12064 5534 12202 5541
rect 12260 5561 12408 5570
rect 12260 5541 12269 5561
rect 12289 5541 12379 5561
rect 12399 5541 12408 5561
rect 12064 5532 12160 5534
rect 12260 5531 12408 5541
rect 12467 5561 12504 5571
rect 12467 5541 12475 5561
rect 12495 5541 12504 5561
rect 12316 5530 12352 5531
rect 11893 5519 11929 5521
rect 11893 5490 11930 5519
rect 11335 5481 11370 5482
rect 11312 5476 11370 5481
rect 11312 5456 11315 5476
rect 11335 5462 11370 5476
rect 11390 5462 11399 5482
rect 11335 5454 11399 5462
rect 11361 5453 11399 5454
rect 11362 5452 11399 5453
rect 11465 5486 11501 5487
rect 11573 5486 11609 5487
rect 11465 5478 11609 5486
rect 11465 5458 11473 5478
rect 11493 5477 11581 5478
rect 11493 5458 11528 5477
rect 11549 5458 11581 5477
rect 11601 5458 11609 5478
rect 11465 5452 11609 5458
rect 11675 5482 11713 5490
rect 11791 5486 11827 5487
rect 11675 5462 11684 5482
rect 11704 5462 11713 5482
rect 11675 5453 11713 5462
rect 11742 5478 11827 5486
rect 11742 5458 11799 5478
rect 11819 5458 11827 5478
rect 11675 5452 11712 5453
rect 11742 5452 11827 5458
rect 11893 5482 11931 5490
rect 11893 5462 11902 5482
rect 11922 5462 11931 5482
rect 12164 5471 12201 5472
rect 12467 5471 12504 5541
rect 12539 5570 12570 5621
rect 12866 5616 12911 5622
rect 12866 5598 12884 5616
rect 12902 5598 12911 5616
rect 14372 5616 14381 5636
rect 14401 5616 14409 5636
rect 14372 5606 14409 5616
rect 14468 5636 14555 5646
rect 14468 5616 14477 5636
rect 14497 5616 14555 5636
rect 14468 5607 14555 5616
rect 14468 5606 14505 5607
rect 12866 5588 12911 5598
rect 12589 5570 12626 5571
rect 12539 5561 12626 5570
rect 12539 5541 12597 5561
rect 12617 5541 12626 5561
rect 12539 5531 12626 5541
rect 12685 5561 12722 5571
rect 12685 5541 12693 5561
rect 12713 5541 12722 5561
rect 12866 5546 12909 5588
rect 13293 5577 13345 5579
rect 12772 5544 12909 5546
rect 12539 5530 12570 5531
rect 12685 5471 12722 5541
rect 12163 5470 12504 5471
rect 11893 5453 11931 5462
rect 12088 5465 12504 5470
rect 11893 5452 11930 5453
rect 11354 5424 11444 5430
rect 11354 5404 11370 5424
rect 11390 5422 11444 5424
rect 11390 5404 11415 5422
rect 11354 5402 11415 5404
rect 11435 5402 11444 5422
rect 11354 5396 11444 5402
rect 11367 5342 11404 5343
rect 11463 5342 11500 5343
rect 11519 5342 11555 5452
rect 11742 5431 11773 5452
rect 12088 5445 12091 5465
rect 12111 5445 12504 5465
rect 12688 5455 12722 5471
rect 12766 5523 12909 5544
rect 13291 5573 13724 5577
rect 13291 5567 13730 5573
rect 13291 5549 13312 5567
rect 13330 5549 13730 5567
rect 14524 5556 14555 5607
rect 14590 5636 14627 5706
rect 14893 5705 14930 5706
rect 14742 5646 14778 5647
rect 14590 5616 14599 5636
rect 14619 5616 14627 5636
rect 14590 5606 14627 5616
rect 14686 5636 14834 5646
rect 14934 5643 15030 5645
rect 14686 5616 14695 5636
rect 14715 5616 14805 5636
rect 14825 5616 14834 5636
rect 14686 5607 14834 5616
rect 14892 5636 15030 5643
rect 14892 5616 14901 5636
rect 14921 5616 15030 5636
rect 14892 5607 15030 5616
rect 14686 5606 14723 5607
rect 14416 5553 14457 5554
rect 13291 5531 13730 5549
rect 12464 5436 12504 5445
rect 12766 5436 12793 5523
rect 12866 5497 12909 5523
rect 12866 5479 12879 5497
rect 12897 5479 12909 5497
rect 12866 5468 12909 5479
rect 11738 5430 11773 5431
rect 11616 5420 11773 5430
rect 11616 5400 11633 5420
rect 11653 5400 11773 5420
rect 11616 5393 11773 5400
rect 11840 5423 11989 5431
rect 11840 5403 11851 5423
rect 11871 5403 11910 5423
rect 11930 5403 11989 5423
rect 12464 5419 12793 5436
rect 12464 5418 12504 5419
rect 11840 5396 11989 5403
rect 12861 5407 12901 5410
rect 12861 5401 12904 5407
rect 12486 5398 12904 5401
rect 11840 5395 11881 5396
rect 11574 5342 11611 5343
rect 11267 5333 11405 5342
rect 10965 5158 11005 5330
rect 11267 5313 11376 5333
rect 11396 5313 11405 5333
rect 11267 5306 11405 5313
rect 11463 5333 11611 5342
rect 11463 5313 11472 5333
rect 11492 5313 11582 5333
rect 11602 5313 11611 5333
rect 11267 5304 11363 5306
rect 11463 5303 11611 5313
rect 11670 5333 11707 5343
rect 11670 5313 11678 5333
rect 11698 5313 11707 5333
rect 11519 5302 11555 5303
rect 11367 5243 11404 5244
rect 11670 5243 11707 5313
rect 11742 5342 11773 5393
rect 12486 5380 12877 5398
rect 12895 5380 12904 5398
rect 12486 5378 12904 5380
rect 12486 5370 12513 5378
rect 12754 5375 12904 5378
rect 12066 5364 12234 5365
rect 12485 5364 12513 5370
rect 12066 5348 12513 5364
rect 12861 5370 12904 5375
rect 11792 5342 11829 5343
rect 11742 5333 11829 5342
rect 11742 5313 11800 5333
rect 11820 5313 11829 5333
rect 11742 5303 11829 5313
rect 11888 5333 11925 5343
rect 11888 5313 11896 5333
rect 11916 5313 11925 5333
rect 11742 5302 11773 5303
rect 11366 5242 11707 5243
rect 11888 5242 11925 5313
rect 11291 5237 11707 5242
rect 11291 5217 11294 5237
rect 11314 5217 11707 5237
rect 11738 5218 11925 5242
rect 12066 5338 12510 5348
rect 12066 5336 12234 5338
rect 12066 5158 12093 5336
rect 12133 5298 12197 5310
rect 12473 5306 12510 5338
rect 12536 5337 12727 5359
rect 12691 5335 12727 5337
rect 12691 5306 12728 5335
rect 12861 5314 12901 5370
rect 12133 5297 12168 5298
rect 12110 5292 12168 5297
rect 12110 5272 12113 5292
rect 12133 5278 12168 5292
rect 12188 5278 12197 5298
rect 12133 5270 12197 5278
rect 12159 5269 12197 5270
rect 12160 5268 12197 5269
rect 12263 5302 12299 5303
rect 12371 5302 12407 5303
rect 12263 5294 12407 5302
rect 12263 5274 12271 5294
rect 12291 5274 12326 5294
rect 12346 5274 12379 5294
rect 12399 5274 12407 5294
rect 12263 5268 12407 5274
rect 12473 5298 12511 5306
rect 12589 5302 12625 5303
rect 12473 5278 12482 5298
rect 12502 5278 12511 5298
rect 12473 5269 12511 5278
rect 12540 5294 12625 5302
rect 12540 5274 12597 5294
rect 12617 5274 12625 5294
rect 12473 5268 12510 5269
rect 12540 5268 12625 5274
rect 12691 5298 12729 5306
rect 12691 5278 12700 5298
rect 12720 5278 12729 5298
rect 12861 5296 12873 5314
rect 12891 5296 12901 5314
rect 13293 5342 13345 5531
rect 13691 5506 13730 5531
rect 14308 5546 14457 5553
rect 14308 5526 14367 5546
rect 14387 5526 14426 5546
rect 14446 5526 14457 5546
rect 14308 5518 14457 5526
rect 14524 5549 14681 5556
rect 14524 5529 14644 5549
rect 14664 5529 14681 5549
rect 14524 5519 14681 5529
rect 14524 5518 14559 5519
rect 13475 5481 13662 5505
rect 13691 5486 14086 5506
rect 14106 5486 14109 5506
rect 14524 5497 14555 5518
rect 14742 5497 14778 5607
rect 14797 5606 14834 5607
rect 14893 5606 14930 5607
rect 14853 5547 14943 5553
rect 14853 5527 14862 5547
rect 14882 5545 14943 5547
rect 14882 5527 14907 5545
rect 14853 5525 14907 5527
rect 14927 5525 14943 5545
rect 14853 5519 14943 5525
rect 14367 5496 14404 5497
rect 13691 5481 14109 5486
rect 14366 5487 14404 5496
rect 13475 5410 13512 5481
rect 13691 5480 14034 5481
rect 13691 5477 13730 5480
rect 13996 5479 14033 5480
rect 13627 5420 13658 5421
rect 13475 5390 13484 5410
rect 13504 5390 13512 5410
rect 13475 5380 13512 5390
rect 13571 5410 13658 5420
rect 13571 5390 13580 5410
rect 13600 5390 13658 5410
rect 13571 5381 13658 5390
rect 13571 5380 13608 5381
rect 13293 5324 13309 5342
rect 13327 5324 13345 5342
rect 13627 5330 13658 5381
rect 13693 5410 13730 5477
rect 14366 5467 14375 5487
rect 14395 5467 14404 5487
rect 14366 5459 14404 5467
rect 14470 5491 14555 5497
rect 14585 5496 14622 5497
rect 14470 5471 14478 5491
rect 14498 5471 14555 5491
rect 14470 5463 14555 5471
rect 14584 5487 14622 5496
rect 14584 5467 14593 5487
rect 14613 5467 14622 5487
rect 14470 5462 14506 5463
rect 14584 5459 14622 5467
rect 14688 5491 14832 5497
rect 14688 5471 14696 5491
rect 14716 5486 14804 5491
rect 14716 5471 14752 5486
rect 14688 5469 14752 5471
rect 14771 5471 14804 5486
rect 14824 5471 14832 5491
rect 14771 5469 14832 5471
rect 14688 5463 14832 5469
rect 14688 5462 14724 5463
rect 14796 5462 14832 5463
rect 14898 5496 14935 5497
rect 14898 5495 14936 5496
rect 14898 5487 14962 5495
rect 14898 5467 14907 5487
rect 14927 5473 14962 5487
rect 14982 5473 14985 5493
rect 14927 5468 14985 5473
rect 14927 5467 14962 5468
rect 14367 5430 14404 5459
rect 14368 5428 14404 5430
rect 13845 5420 13881 5421
rect 13693 5390 13702 5410
rect 13722 5390 13730 5410
rect 13693 5380 13730 5390
rect 13789 5410 13937 5420
rect 14037 5417 14133 5419
rect 13789 5390 13798 5410
rect 13818 5390 13908 5410
rect 13928 5390 13937 5410
rect 13789 5381 13937 5390
rect 13995 5410 14133 5417
rect 13995 5390 14004 5410
rect 14024 5390 14133 5410
rect 14368 5406 14559 5428
rect 14585 5427 14622 5459
rect 14898 5455 14962 5467
rect 15002 5429 15029 5607
rect 14861 5427 15029 5429
rect 14585 5413 15029 5427
rect 15053 5450 15081 6396
rect 15053 5420 15098 5450
rect 14585 5401 15032 5413
rect 14628 5399 14661 5401
rect 13995 5381 14133 5390
rect 13789 5380 13826 5381
rect 13519 5327 13560 5328
rect 13293 5306 13345 5324
rect 13411 5320 13560 5327
rect 12861 5286 12901 5296
rect 13411 5300 13470 5320
rect 13490 5300 13529 5320
rect 13549 5300 13560 5320
rect 13411 5292 13560 5300
rect 13627 5323 13784 5330
rect 13627 5303 13747 5323
rect 13767 5303 13784 5323
rect 13627 5293 13784 5303
rect 13627 5292 13662 5293
rect 12691 5269 12729 5278
rect 13627 5271 13658 5292
rect 13845 5271 13881 5381
rect 13900 5380 13937 5381
rect 13996 5380 14033 5381
rect 13956 5321 14046 5327
rect 13956 5301 13965 5321
rect 13985 5319 14046 5321
rect 13985 5301 14010 5319
rect 13956 5299 14010 5301
rect 14030 5299 14046 5319
rect 13956 5293 14046 5299
rect 13470 5270 13507 5271
rect 12691 5268 12728 5269
rect 12152 5240 12242 5246
rect 12152 5220 12168 5240
rect 12188 5238 12242 5240
rect 12188 5220 12213 5238
rect 12152 5218 12213 5220
rect 12233 5218 12242 5238
rect 12152 5212 12242 5218
rect 12165 5158 12202 5159
rect 12261 5158 12298 5159
rect 12317 5158 12353 5268
rect 12540 5247 12571 5268
rect 13469 5261 13507 5270
rect 12536 5246 12571 5247
rect 12414 5236 12571 5246
rect 12414 5216 12431 5236
rect 12451 5216 12571 5236
rect 12414 5209 12571 5216
rect 12638 5239 12787 5247
rect 12638 5219 12649 5239
rect 12669 5219 12708 5239
rect 12728 5219 12787 5239
rect 13297 5243 13337 5253
rect 12638 5212 12787 5219
rect 12853 5215 12905 5233
rect 12638 5211 12679 5212
rect 12372 5158 12409 5159
rect 10966 5143 11005 5158
rect 12065 5149 12203 5158
rect 10966 5142 11132 5143
rect 11258 5142 11298 5144
rect 10966 5116 11408 5142
rect 10966 5114 11132 5116
rect 10630 5002 10667 5010
rect 10630 4983 10638 5002
rect 10659 4983 10667 5002
rect 10630 4977 10667 4983
rect 10966 4936 10991 5114
rect 11031 5076 11095 5088
rect 11371 5084 11408 5116
rect 11434 5115 11625 5137
rect 12065 5129 12174 5149
rect 12194 5129 12203 5149
rect 12065 5122 12203 5129
rect 12261 5149 12409 5158
rect 12261 5129 12270 5149
rect 12290 5129 12380 5149
rect 12400 5129 12409 5149
rect 12065 5120 12161 5122
rect 12261 5119 12409 5129
rect 12468 5149 12505 5159
rect 12468 5129 12476 5149
rect 12496 5129 12505 5149
rect 12317 5118 12353 5119
rect 11589 5113 11625 5115
rect 11589 5084 11626 5113
rect 11031 5075 11066 5076
rect 11008 5070 11066 5075
rect 11008 5050 11011 5070
rect 11031 5056 11066 5070
rect 11086 5056 11095 5076
rect 11031 5048 11095 5056
rect 11057 5047 11095 5048
rect 11058 5046 11095 5047
rect 11161 5080 11197 5081
rect 11269 5080 11305 5081
rect 11161 5075 11305 5080
rect 11161 5072 11223 5075
rect 11161 5052 11169 5072
rect 11189 5052 11223 5072
rect 11161 5049 11223 5052
rect 11249 5072 11305 5075
rect 11249 5052 11277 5072
rect 11297 5052 11305 5072
rect 11249 5049 11305 5052
rect 11161 5046 11305 5049
rect 11371 5076 11409 5084
rect 11487 5080 11523 5081
rect 11371 5056 11380 5076
rect 11400 5056 11409 5076
rect 11371 5047 11409 5056
rect 11438 5072 11523 5080
rect 11438 5052 11495 5072
rect 11515 5052 11523 5072
rect 11371 5046 11408 5047
rect 11438 5046 11523 5052
rect 11589 5076 11627 5084
rect 11589 5056 11598 5076
rect 11618 5056 11627 5076
rect 12468 5062 12505 5129
rect 12540 5158 12571 5209
rect 12853 5197 12871 5215
rect 12889 5197 12905 5215
rect 12590 5158 12627 5159
rect 12540 5149 12627 5158
rect 12540 5129 12598 5149
rect 12618 5129 12627 5149
rect 12540 5119 12627 5129
rect 12686 5149 12723 5159
rect 12686 5129 12694 5149
rect 12714 5129 12723 5149
rect 12540 5118 12571 5119
rect 12165 5059 12202 5060
rect 12468 5059 12507 5062
rect 12164 5058 12507 5059
rect 12686 5058 12723 5129
rect 11589 5047 11627 5056
rect 12089 5053 12507 5058
rect 11589 5046 11626 5047
rect 11050 5018 11140 5024
rect 11050 4998 11066 5018
rect 11086 5016 11140 5018
rect 11086 4998 11111 5016
rect 11050 4996 11111 4998
rect 11131 4996 11140 5016
rect 11050 4990 11140 4996
rect 11063 4936 11100 4937
rect 11159 4936 11196 4937
rect 11215 4936 11251 5046
rect 11438 5025 11469 5046
rect 12089 5033 12092 5053
rect 12112 5033 12507 5053
rect 12536 5034 12723 5058
rect 11434 5024 11469 5025
rect 11312 5014 11469 5024
rect 11312 4994 11329 5014
rect 11349 4994 11469 5014
rect 11312 4987 11469 4994
rect 11536 5017 11685 5025
rect 11536 4997 11547 5017
rect 11567 4997 11606 5017
rect 11626 4997 11685 5017
rect 11536 4990 11685 4997
rect 12468 5008 12507 5033
rect 12853 5008 12905 5197
rect 13297 5225 13307 5243
rect 13325 5225 13337 5243
rect 13469 5241 13478 5261
rect 13498 5241 13507 5261
rect 13469 5233 13507 5241
rect 13573 5265 13658 5271
rect 13688 5270 13725 5271
rect 13573 5245 13581 5265
rect 13601 5245 13658 5265
rect 13573 5237 13658 5245
rect 13687 5261 13725 5270
rect 13687 5241 13696 5261
rect 13716 5241 13725 5261
rect 13573 5236 13609 5237
rect 13687 5233 13725 5241
rect 13791 5265 13935 5271
rect 13791 5245 13799 5265
rect 13819 5245 13852 5265
rect 13872 5245 13907 5265
rect 13927 5245 13935 5265
rect 13791 5237 13935 5245
rect 13791 5236 13827 5237
rect 13899 5236 13935 5237
rect 14001 5270 14038 5271
rect 14001 5269 14039 5270
rect 14001 5261 14065 5269
rect 14001 5241 14010 5261
rect 14030 5247 14065 5261
rect 14085 5247 14088 5267
rect 14030 5242 14088 5247
rect 14030 5241 14065 5242
rect 13297 5169 13337 5225
rect 13470 5204 13507 5233
rect 13471 5202 13507 5204
rect 13471 5180 13662 5202
rect 13688 5201 13725 5233
rect 14001 5229 14065 5241
rect 14105 5203 14132 5381
rect 14990 5356 15032 5401
rect 15053 5402 15064 5420
rect 15086 5402 15098 5420
rect 15053 5396 15098 5402
rect 15054 5395 15098 5396
rect 13964 5201 14132 5203
rect 13688 5191 14132 5201
rect 14273 5297 14460 5321
rect 14491 5302 14884 5322
rect 14904 5302 14907 5322
rect 14491 5297 14907 5302
rect 14273 5226 14310 5297
rect 14491 5296 14832 5297
rect 14425 5236 14456 5237
rect 14273 5206 14282 5226
rect 14302 5206 14310 5226
rect 14273 5196 14310 5206
rect 14369 5226 14456 5236
rect 14369 5206 14378 5226
rect 14398 5206 14456 5226
rect 14369 5197 14456 5206
rect 14369 5196 14406 5197
rect 13294 5164 13337 5169
rect 13685 5175 14132 5191
rect 13685 5169 13713 5175
rect 13964 5174 14132 5175
rect 13294 5161 13444 5164
rect 13685 5161 13712 5169
rect 13294 5159 13712 5161
rect 13294 5141 13303 5159
rect 13321 5141 13712 5159
rect 14425 5146 14456 5197
rect 14491 5226 14528 5296
rect 14794 5295 14831 5296
rect 14643 5236 14679 5237
rect 14491 5206 14500 5226
rect 14520 5206 14528 5226
rect 14491 5196 14528 5206
rect 14587 5226 14735 5236
rect 14835 5233 14931 5235
rect 14587 5206 14596 5226
rect 14616 5206 14706 5226
rect 14726 5206 14735 5226
rect 14587 5197 14735 5206
rect 14793 5226 14931 5233
rect 14793 5206 14802 5226
rect 14822 5206 14931 5226
rect 14793 5197 14931 5206
rect 14587 5196 14624 5197
rect 14317 5143 14358 5144
rect 13294 5138 13712 5141
rect 13294 5132 13337 5138
rect 13297 5129 13337 5132
rect 14212 5136 14358 5143
rect 13694 5120 13734 5121
rect 13405 5103 13734 5120
rect 14212 5116 14268 5136
rect 14288 5116 14327 5136
rect 14347 5116 14358 5136
rect 14212 5108 14358 5116
rect 14425 5139 14582 5146
rect 14425 5119 14545 5139
rect 14565 5119 14582 5139
rect 14425 5109 14582 5119
rect 14425 5108 14460 5109
rect 13289 5060 13332 5071
rect 13289 5042 13301 5060
rect 13319 5042 13332 5060
rect 13289 5016 13332 5042
rect 13405 5016 13432 5103
rect 13694 5094 13734 5103
rect 12468 4990 12907 5008
rect 11536 4989 11577 4990
rect 11270 4936 11307 4937
rect 10966 4927 11101 4936
rect 10966 4907 11072 4927
rect 11092 4907 11101 4927
rect 10966 4900 11101 4907
rect 11159 4927 11307 4936
rect 11159 4907 11168 4927
rect 11188 4907 11278 4927
rect 11298 4907 11307 4927
rect 10966 4898 11059 4900
rect 11159 4897 11307 4907
rect 11366 4927 11403 4937
rect 11366 4907 11374 4927
rect 11394 4907 11403 4927
rect 11215 4896 11251 4897
rect 11063 4837 11100 4838
rect 11366 4837 11403 4907
rect 11438 4936 11469 4987
rect 12468 4972 12868 4990
rect 12886 4972 12907 4990
rect 12468 4966 12907 4972
rect 12474 4962 12907 4966
rect 13289 4995 13432 5016
rect 13476 5068 13510 5084
rect 13694 5074 14087 5094
rect 14107 5074 14110 5094
rect 14425 5087 14456 5108
rect 14643 5087 14679 5197
rect 14698 5196 14735 5197
rect 14794 5196 14831 5197
rect 14754 5137 14844 5143
rect 14754 5117 14763 5137
rect 14783 5135 14844 5137
rect 14783 5117 14808 5135
rect 14754 5115 14808 5117
rect 14828 5115 14844 5135
rect 14754 5109 14844 5115
rect 14268 5086 14305 5087
rect 13694 5069 14110 5074
rect 14267 5077 14305 5086
rect 13694 5068 14035 5069
rect 13476 4998 13513 5068
rect 13628 5008 13659 5009
rect 13289 4993 13426 4995
rect 12853 4960 12905 4962
rect 13289 4951 13332 4993
rect 13476 4978 13485 4998
rect 13505 4978 13513 4998
rect 13476 4968 13513 4978
rect 13572 4998 13659 5008
rect 13572 4978 13581 4998
rect 13601 4978 13659 4998
rect 13572 4969 13659 4978
rect 13572 4968 13609 4969
rect 13287 4941 13332 4951
rect 11488 4936 11525 4937
rect 11438 4927 11525 4936
rect 11438 4907 11496 4927
rect 11516 4907 11525 4927
rect 11438 4897 11525 4907
rect 11584 4927 11621 4937
rect 11584 4907 11592 4927
rect 11612 4907 11621 4927
rect 13287 4923 13296 4941
rect 13314 4923 13332 4941
rect 13287 4917 13332 4923
rect 13628 4918 13659 4969
rect 13694 4998 13731 5068
rect 13997 5067 14034 5068
rect 14267 5057 14276 5077
rect 14296 5057 14305 5077
rect 14267 5049 14305 5057
rect 14371 5081 14456 5087
rect 14486 5086 14523 5087
rect 14371 5061 14379 5081
rect 14399 5061 14456 5081
rect 14371 5053 14456 5061
rect 14485 5077 14523 5086
rect 14485 5057 14494 5077
rect 14514 5057 14523 5077
rect 14371 5052 14407 5053
rect 14485 5049 14523 5057
rect 14589 5081 14733 5087
rect 14589 5061 14597 5081
rect 14617 5078 14705 5081
rect 14617 5061 14652 5078
rect 14589 5060 14652 5061
rect 14671 5061 14705 5078
rect 14725 5061 14733 5081
rect 14671 5060 14733 5061
rect 14589 5053 14733 5060
rect 14589 5052 14625 5053
rect 14697 5052 14733 5053
rect 14799 5086 14836 5087
rect 14799 5085 14837 5086
rect 14859 5085 14886 5089
rect 14799 5083 14886 5085
rect 14799 5077 14863 5083
rect 14799 5057 14808 5077
rect 14828 5063 14863 5077
rect 14883 5063 14886 5083
rect 14828 5058 14886 5063
rect 14828 5057 14863 5058
rect 14268 5020 14305 5049
rect 14269 5018 14305 5020
rect 13846 5008 13882 5009
rect 13694 4978 13703 4998
rect 13723 4978 13731 4998
rect 13694 4968 13731 4978
rect 13790 4998 13938 5008
rect 14038 5005 14134 5007
rect 13790 4978 13799 4998
rect 13819 4978 13909 4998
rect 13929 4978 13938 4998
rect 13790 4969 13938 4978
rect 13996 4998 14134 5005
rect 13996 4978 14005 4998
rect 14025 4978 14134 4998
rect 14269 4996 14460 5018
rect 14486 5017 14523 5049
rect 14799 5045 14863 5057
rect 14903 5019 14930 5197
rect 14762 5017 14930 5019
rect 14486 4991 14930 5017
rect 13996 4969 14134 4978
rect 13790 4968 13827 4969
rect 13287 4914 13324 4917
rect 13520 4915 13561 4916
rect 11438 4896 11469 4897
rect 11062 4836 11403 4837
rect 11584 4836 11621 4907
rect 13412 4908 13561 4915
rect 12856 4895 12893 4900
rect 10987 4831 11403 4836
rect 10987 4811 10990 4831
rect 11010 4811 11403 4831
rect 11434 4812 11621 4836
rect 12847 4891 12894 4895
rect 12847 4873 12866 4891
rect 12884 4873 12894 4891
rect 13412 4888 13471 4908
rect 13491 4888 13530 4908
rect 13550 4888 13561 4908
rect 13412 4880 13561 4888
rect 13628 4911 13785 4918
rect 13628 4891 13748 4911
rect 13768 4891 13785 4911
rect 13628 4881 13785 4891
rect 13628 4880 13663 4881
rect 12455 4814 12493 4815
rect 12847 4814 12894 4873
rect 13628 4859 13659 4880
rect 13846 4859 13882 4969
rect 13901 4968 13938 4969
rect 13997 4968 14034 4969
rect 13957 4909 14047 4915
rect 13957 4889 13966 4909
rect 13986 4907 14047 4909
rect 13986 4889 14011 4907
rect 13957 4887 14011 4889
rect 14031 4887 14047 4907
rect 13957 4881 14047 4887
rect 13471 4858 13508 4859
rect 13284 4850 13321 4852
rect 13284 4842 13326 4850
rect 13284 4824 13294 4842
rect 13312 4824 13326 4842
rect 13284 4815 13326 4824
rect 13470 4849 13508 4858
rect 13470 4829 13479 4849
rect 13499 4829 13508 4849
rect 13470 4821 13508 4829
rect 13574 4853 13659 4859
rect 13689 4858 13726 4859
rect 13574 4833 13582 4853
rect 13602 4833 13659 4853
rect 13574 4825 13659 4833
rect 13688 4849 13726 4858
rect 13688 4829 13697 4849
rect 13717 4829 13726 4849
rect 13574 4824 13610 4825
rect 13688 4821 13726 4829
rect 13792 4857 13936 4859
rect 13792 4853 13844 4857
rect 13792 4833 13800 4853
rect 13820 4837 13844 4853
rect 13864 4853 13936 4857
rect 13864 4837 13908 4853
rect 13820 4833 13908 4837
rect 13928 4833 13936 4853
rect 13792 4825 13936 4833
rect 13792 4824 13828 4825
rect 13900 4824 13936 4825
rect 14002 4858 14039 4859
rect 14002 4857 14040 4858
rect 14002 4849 14066 4857
rect 14002 4829 14011 4849
rect 14031 4835 14066 4849
rect 14086 4835 14089 4855
rect 14031 4830 14089 4835
rect 14031 4829 14066 4830
rect 11207 4810 11272 4811
rect 9322 4732 9360 4733
rect 8921 4694 9360 4732
rect 10232 4732 10240 4754
rect 10264 4732 10272 4754
rect 10232 4724 10272 4732
rect 11543 4776 11583 4784
rect 11543 4754 11551 4776
rect 11575 4754 11583 4776
rect 12455 4776 12894 4814
rect 12455 4775 12493 4776
rect 10543 4697 10608 4698
rect 7736 4679 7771 4680
rect 7713 4674 7771 4679
rect 7713 4654 7716 4674
rect 7736 4660 7771 4674
rect 7791 4660 7800 4680
rect 7736 4652 7800 4660
rect 7762 4651 7800 4652
rect 7763 4650 7800 4651
rect 7866 4684 7902 4685
rect 7974 4684 8010 4685
rect 7866 4676 8010 4684
rect 7866 4656 7874 4676
rect 7894 4672 7982 4676
rect 7894 4656 7938 4672
rect 7866 4652 7938 4656
rect 7958 4656 7982 4672
rect 8002 4656 8010 4676
rect 7958 4652 8010 4656
rect 7866 4650 8010 4652
rect 8076 4680 8114 4688
rect 8192 4684 8228 4685
rect 8076 4660 8085 4680
rect 8105 4660 8114 4680
rect 8076 4651 8114 4660
rect 8143 4676 8228 4684
rect 8143 4656 8200 4676
rect 8220 4656 8228 4676
rect 8076 4650 8113 4651
rect 8143 4650 8228 4656
rect 8294 4680 8332 4688
rect 8294 4660 8303 4680
rect 8323 4660 8332 4680
rect 8294 4651 8332 4660
rect 8476 4685 8518 4694
rect 8476 4667 8490 4685
rect 8508 4667 8518 4685
rect 8476 4659 8518 4667
rect 8481 4657 8518 4659
rect 8294 4650 8331 4651
rect 7755 4622 7845 4628
rect 7755 4602 7771 4622
rect 7791 4620 7845 4622
rect 7791 4602 7816 4620
rect 7755 4600 7816 4602
rect 7836 4600 7845 4620
rect 7755 4594 7845 4600
rect 7768 4540 7805 4541
rect 7864 4540 7901 4541
rect 7920 4540 7956 4650
rect 8143 4629 8174 4650
rect 8921 4635 8968 4694
rect 9322 4693 9360 4694
rect 8139 4628 8174 4629
rect 8017 4618 8174 4628
rect 8017 4598 8034 4618
rect 8054 4598 8174 4618
rect 8017 4591 8174 4598
rect 8241 4621 8390 4629
rect 8241 4601 8252 4621
rect 8272 4601 8311 4621
rect 8331 4601 8390 4621
rect 8921 4617 8931 4635
rect 8949 4617 8968 4635
rect 8921 4613 8968 4617
rect 10194 4672 10381 4696
rect 10412 4677 10805 4697
rect 10825 4677 10828 4697
rect 10412 4672 10828 4677
rect 8922 4608 8959 4613
rect 8241 4594 8390 4601
rect 10194 4601 10231 4672
rect 10412 4671 10753 4672
rect 10346 4611 10377 4612
rect 8241 4593 8282 4594
rect 8478 4592 8515 4595
rect 7975 4540 8012 4541
rect 7668 4531 7806 4540
rect 6872 4492 7316 4518
rect 6872 4490 7040 4492
rect 6872 4312 6899 4490
rect 6939 4452 7003 4464
rect 7279 4460 7316 4492
rect 7342 4491 7533 4513
rect 7668 4511 7777 4531
rect 7797 4511 7806 4531
rect 7668 4504 7806 4511
rect 7864 4531 8012 4540
rect 7864 4511 7873 4531
rect 7893 4511 7983 4531
rect 8003 4511 8012 4531
rect 7668 4502 7764 4504
rect 7864 4501 8012 4511
rect 8071 4531 8108 4541
rect 8071 4511 8079 4531
rect 8099 4511 8108 4531
rect 7920 4500 7956 4501
rect 7497 4489 7533 4491
rect 7497 4460 7534 4489
rect 6939 4451 6974 4452
rect 6916 4446 6974 4451
rect 6916 4426 6919 4446
rect 6939 4432 6974 4446
rect 6994 4432 7003 4452
rect 6939 4426 7003 4432
rect 6916 4424 7003 4426
rect 6916 4420 6943 4424
rect 6965 4423 7003 4424
rect 6966 4422 7003 4423
rect 7069 4456 7105 4457
rect 7177 4456 7213 4457
rect 7069 4449 7213 4456
rect 7069 4448 7131 4449
rect 7069 4428 7077 4448
rect 7097 4431 7131 4448
rect 7150 4448 7213 4449
rect 7150 4431 7185 4448
rect 7097 4428 7185 4431
rect 7205 4428 7213 4448
rect 7069 4422 7213 4428
rect 7279 4452 7317 4460
rect 7395 4456 7431 4457
rect 7279 4432 7288 4452
rect 7308 4432 7317 4452
rect 7279 4423 7317 4432
rect 7346 4448 7431 4456
rect 7346 4428 7403 4448
rect 7423 4428 7431 4448
rect 7279 4422 7316 4423
rect 7346 4422 7431 4428
rect 7497 4452 7535 4460
rect 7497 4432 7506 4452
rect 7526 4432 7535 4452
rect 7768 4441 7805 4442
rect 8071 4441 8108 4511
rect 8143 4540 8174 4591
rect 8470 4586 8515 4592
rect 8470 4568 8488 4586
rect 8506 4568 8515 4586
rect 10194 4581 10203 4601
rect 10223 4581 10231 4601
rect 10194 4571 10231 4581
rect 10290 4601 10377 4611
rect 10290 4581 10299 4601
rect 10319 4581 10377 4601
rect 10290 4572 10377 4581
rect 10290 4571 10327 4572
rect 8470 4558 8515 4568
rect 8193 4540 8230 4541
rect 8143 4531 8230 4540
rect 8143 4511 8201 4531
rect 8221 4511 8230 4531
rect 8143 4501 8230 4511
rect 8289 4531 8326 4541
rect 8289 4511 8297 4531
rect 8317 4511 8326 4531
rect 8470 4516 8513 4558
rect 8910 4546 8962 4548
rect 8376 4514 8513 4516
rect 8143 4500 8174 4501
rect 8289 4441 8326 4511
rect 7767 4440 8108 4441
rect 7497 4423 7535 4432
rect 7692 4435 8108 4440
rect 7497 4422 7534 4423
rect 6958 4394 7048 4400
rect 6958 4374 6974 4394
rect 6994 4392 7048 4394
rect 6994 4374 7019 4392
rect 6958 4372 7019 4374
rect 7039 4372 7048 4392
rect 6958 4366 7048 4372
rect 6971 4312 7008 4313
rect 7067 4312 7104 4313
rect 7123 4312 7159 4422
rect 7346 4401 7377 4422
rect 7692 4415 7695 4435
rect 7715 4415 8108 4435
rect 8292 4425 8326 4441
rect 8370 4493 8513 4514
rect 8908 4542 9341 4546
rect 8908 4536 9347 4542
rect 8908 4518 8929 4536
rect 8947 4518 9347 4536
rect 10346 4521 10377 4572
rect 10412 4601 10449 4671
rect 10715 4670 10752 4671
rect 10564 4611 10600 4612
rect 10412 4581 10421 4601
rect 10441 4581 10449 4601
rect 10412 4571 10449 4581
rect 10508 4601 10656 4611
rect 10756 4608 10852 4610
rect 10508 4581 10517 4601
rect 10537 4581 10627 4601
rect 10647 4581 10656 4601
rect 10508 4572 10656 4581
rect 10714 4601 10852 4608
rect 10714 4581 10723 4601
rect 10743 4581 10852 4601
rect 10714 4572 10852 4581
rect 10508 4571 10545 4572
rect 10238 4518 10279 4519
rect 8908 4500 9347 4518
rect 8068 4406 8108 4415
rect 8370 4406 8397 4493
rect 8470 4467 8513 4493
rect 8470 4449 8483 4467
rect 8501 4449 8513 4467
rect 8470 4438 8513 4449
rect 7342 4400 7377 4401
rect 7220 4390 7377 4400
rect 7220 4370 7237 4390
rect 7257 4370 7377 4390
rect 7220 4363 7377 4370
rect 7444 4393 7590 4401
rect 7444 4373 7455 4393
rect 7475 4373 7514 4393
rect 7534 4373 7590 4393
rect 8068 4389 8397 4406
rect 8068 4388 8108 4389
rect 7444 4366 7590 4373
rect 8465 4377 8505 4380
rect 8465 4371 8508 4377
rect 8090 4368 8508 4371
rect 7444 4365 7485 4366
rect 7178 4312 7215 4313
rect 6871 4303 7009 4312
rect 6871 4283 6980 4303
rect 7000 4283 7009 4303
rect 6871 4276 7009 4283
rect 7067 4303 7215 4312
rect 7067 4283 7076 4303
rect 7096 4283 7186 4303
rect 7206 4283 7215 4303
rect 6871 4274 6967 4276
rect 7067 4273 7215 4283
rect 7274 4303 7311 4313
rect 7274 4283 7282 4303
rect 7302 4283 7311 4303
rect 7123 4272 7159 4273
rect 6971 4213 7008 4214
rect 7274 4213 7311 4283
rect 7346 4312 7377 4363
rect 8090 4350 8481 4368
rect 8499 4350 8508 4368
rect 8090 4348 8508 4350
rect 8090 4340 8117 4348
rect 8358 4345 8508 4348
rect 7670 4334 7838 4335
rect 8089 4334 8117 4340
rect 7670 4318 8117 4334
rect 8465 4340 8508 4345
rect 7396 4312 7433 4313
rect 7346 4303 7433 4312
rect 7346 4283 7404 4303
rect 7424 4283 7433 4303
rect 7346 4273 7433 4283
rect 7492 4303 7529 4313
rect 7492 4283 7500 4303
rect 7520 4283 7529 4303
rect 7346 4272 7377 4273
rect 6970 4212 7311 4213
rect 7492 4212 7529 4283
rect 6895 4207 7311 4212
rect 6895 4187 6898 4207
rect 6918 4187 7311 4207
rect 7342 4188 7529 4212
rect 7670 4308 8114 4318
rect 7670 4306 7838 4308
rect 6704 4113 6748 4114
rect 6704 4107 6749 4113
rect 6704 4089 6716 4107
rect 6738 4089 6749 4107
rect 6770 4108 6812 4153
rect 7670 4128 7697 4306
rect 7737 4268 7801 4280
rect 8077 4276 8114 4308
rect 8140 4307 8331 4329
rect 8295 4305 8331 4307
rect 8295 4276 8332 4305
rect 8465 4284 8505 4340
rect 7737 4267 7772 4268
rect 7714 4262 7772 4267
rect 7714 4242 7717 4262
rect 7737 4248 7772 4262
rect 7792 4248 7801 4268
rect 7737 4240 7801 4248
rect 7763 4239 7801 4240
rect 7764 4238 7801 4239
rect 7867 4272 7903 4273
rect 7975 4272 8011 4273
rect 7867 4264 8011 4272
rect 7867 4244 7875 4264
rect 7895 4244 7930 4264
rect 7950 4244 7983 4264
rect 8003 4244 8011 4264
rect 7867 4238 8011 4244
rect 8077 4268 8115 4276
rect 8193 4272 8229 4273
rect 8077 4248 8086 4268
rect 8106 4248 8115 4268
rect 8077 4239 8115 4248
rect 8144 4264 8229 4272
rect 8144 4244 8201 4264
rect 8221 4244 8229 4264
rect 8077 4238 8114 4239
rect 8144 4238 8229 4244
rect 8295 4268 8333 4276
rect 8295 4248 8304 4268
rect 8324 4248 8333 4268
rect 8465 4266 8477 4284
rect 8495 4266 8505 4284
rect 8910 4311 8962 4500
rect 9308 4475 9347 4500
rect 10130 4511 10279 4518
rect 10130 4491 10189 4511
rect 10209 4491 10248 4511
rect 10268 4491 10279 4511
rect 10130 4483 10279 4491
rect 10346 4514 10503 4521
rect 10346 4494 10466 4514
rect 10486 4494 10503 4514
rect 10346 4484 10503 4494
rect 10346 4483 10381 4484
rect 9092 4450 9279 4474
rect 9308 4455 9703 4475
rect 9723 4455 9726 4475
rect 10346 4462 10377 4483
rect 10564 4462 10600 4572
rect 10619 4571 10656 4572
rect 10715 4571 10752 4572
rect 10675 4512 10765 4518
rect 10675 4492 10684 4512
rect 10704 4510 10765 4512
rect 10704 4492 10729 4510
rect 10675 4490 10729 4492
rect 10749 4490 10765 4510
rect 10675 4484 10765 4490
rect 10189 4461 10226 4462
rect 9308 4450 9726 4455
rect 10188 4452 10226 4461
rect 9092 4379 9129 4450
rect 9308 4449 9651 4450
rect 9308 4446 9347 4449
rect 9613 4448 9650 4449
rect 9244 4389 9275 4390
rect 9092 4359 9101 4379
rect 9121 4359 9129 4379
rect 9092 4349 9129 4359
rect 9188 4379 9275 4389
rect 9188 4359 9197 4379
rect 9217 4359 9275 4379
rect 9188 4350 9275 4359
rect 9188 4349 9225 4350
rect 8910 4293 8926 4311
rect 8944 4293 8962 4311
rect 9244 4299 9275 4350
rect 9310 4379 9347 4446
rect 10188 4432 10197 4452
rect 10217 4432 10226 4452
rect 10188 4424 10226 4432
rect 10292 4456 10377 4462
rect 10407 4461 10444 4462
rect 10292 4436 10300 4456
rect 10320 4436 10377 4456
rect 10292 4428 10377 4436
rect 10406 4452 10444 4461
rect 10406 4432 10415 4452
rect 10435 4432 10444 4452
rect 10292 4427 10328 4428
rect 10406 4424 10444 4432
rect 10510 4456 10654 4462
rect 10510 4436 10518 4456
rect 10538 4450 10626 4456
rect 10538 4436 10567 4450
rect 10510 4428 10567 4436
rect 10510 4427 10546 4428
rect 10590 4436 10626 4450
rect 10646 4436 10654 4456
rect 10590 4428 10654 4436
rect 10618 4427 10654 4428
rect 10720 4461 10757 4462
rect 10720 4460 10758 4461
rect 10720 4452 10784 4460
rect 10720 4432 10729 4452
rect 10749 4438 10784 4452
rect 10804 4438 10807 4458
rect 10749 4433 10807 4438
rect 10749 4432 10784 4433
rect 10189 4395 10226 4424
rect 10190 4393 10226 4395
rect 9462 4389 9498 4390
rect 9310 4359 9319 4379
rect 9339 4359 9347 4379
rect 9310 4349 9347 4359
rect 9406 4379 9554 4389
rect 9654 4386 9750 4388
rect 9406 4359 9415 4379
rect 9435 4359 9525 4379
rect 9545 4359 9554 4379
rect 9406 4350 9554 4359
rect 9612 4379 9750 4386
rect 9612 4359 9621 4379
rect 9641 4359 9750 4379
rect 10190 4371 10381 4393
rect 10407 4392 10444 4424
rect 10720 4420 10784 4432
rect 10824 4394 10851 4572
rect 11148 4525 11185 4531
rect 11148 4506 11156 4525
rect 11177 4506 11185 4525
rect 11148 4498 11185 4506
rect 10683 4392 10851 4394
rect 10407 4366 10851 4392
rect 10517 4364 10557 4366
rect 10683 4365 10851 4366
rect 9612 4350 9750 4359
rect 10810 4360 10851 4365
rect 9406 4349 9443 4350
rect 9136 4296 9177 4297
rect 8910 4275 8962 4293
rect 9028 4289 9177 4296
rect 8465 4256 8505 4266
rect 9028 4269 9087 4289
rect 9107 4269 9146 4289
rect 9166 4269 9177 4289
rect 9028 4261 9177 4269
rect 9244 4292 9401 4299
rect 9244 4272 9364 4292
rect 9384 4272 9401 4292
rect 9244 4262 9401 4272
rect 9244 4261 9279 4262
rect 8295 4239 8333 4248
rect 9244 4240 9275 4261
rect 9462 4240 9498 4350
rect 9517 4349 9554 4350
rect 9613 4349 9650 4350
rect 9573 4290 9663 4296
rect 9573 4270 9582 4290
rect 9602 4288 9663 4290
rect 9602 4270 9627 4288
rect 9573 4268 9627 4270
rect 9647 4268 9663 4288
rect 9573 4262 9663 4268
rect 9087 4239 9124 4240
rect 8295 4238 8332 4239
rect 7756 4210 7846 4216
rect 7756 4190 7772 4210
rect 7792 4208 7846 4210
rect 7792 4190 7817 4208
rect 7756 4188 7817 4190
rect 7837 4188 7846 4208
rect 7756 4182 7846 4188
rect 7769 4128 7806 4129
rect 7865 4128 7902 4129
rect 7921 4128 7957 4238
rect 8144 4217 8175 4238
rect 9086 4230 9124 4239
rect 8140 4216 8175 4217
rect 8018 4206 8175 4216
rect 8018 4186 8035 4206
rect 8055 4186 8175 4206
rect 8018 4179 8175 4186
rect 8242 4209 8391 4217
rect 8242 4189 8253 4209
rect 8273 4189 8312 4209
rect 8332 4189 8391 4209
rect 8914 4212 8954 4222
rect 8242 4182 8391 4189
rect 8457 4185 8509 4203
rect 8242 4181 8283 4182
rect 7976 4128 8013 4129
rect 7669 4119 7807 4128
rect 7141 4108 7174 4110
rect 6770 4096 7217 4108
rect 6704 4059 6749 4089
rect 6721 3113 6749 4059
rect 6773 4082 7217 4096
rect 6773 4080 6941 4082
rect 6773 3902 6800 4080
rect 6840 4042 6904 4054
rect 7180 4050 7217 4082
rect 7243 4081 7434 4103
rect 7669 4099 7778 4119
rect 7798 4099 7807 4119
rect 7669 4092 7807 4099
rect 7865 4119 8013 4128
rect 7865 4099 7874 4119
rect 7894 4099 7984 4119
rect 8004 4099 8013 4119
rect 7669 4090 7765 4092
rect 7865 4089 8013 4099
rect 8072 4119 8109 4129
rect 8072 4099 8080 4119
rect 8100 4099 8109 4119
rect 7921 4088 7957 4089
rect 7398 4079 7434 4081
rect 7398 4050 7435 4079
rect 6840 4041 6875 4042
rect 6817 4036 6875 4041
rect 6817 4016 6820 4036
rect 6840 4022 6875 4036
rect 6895 4022 6904 4042
rect 6840 4014 6904 4022
rect 6866 4013 6904 4014
rect 6867 4012 6904 4013
rect 6970 4046 7006 4047
rect 7078 4046 7114 4047
rect 6970 4040 7114 4046
rect 6970 4038 7031 4040
rect 6970 4018 6978 4038
rect 6998 4023 7031 4038
rect 7050 4038 7114 4040
rect 7050 4023 7086 4038
rect 6998 4018 7086 4023
rect 7106 4018 7114 4038
rect 6970 4012 7114 4018
rect 7180 4042 7218 4050
rect 7296 4046 7332 4047
rect 7180 4022 7189 4042
rect 7209 4022 7218 4042
rect 7180 4013 7218 4022
rect 7247 4038 7332 4046
rect 7247 4018 7304 4038
rect 7324 4018 7332 4038
rect 7180 4012 7217 4013
rect 7247 4012 7332 4018
rect 7398 4042 7436 4050
rect 7398 4022 7407 4042
rect 7427 4022 7436 4042
rect 8072 4032 8109 4099
rect 8144 4128 8175 4179
rect 8457 4167 8475 4185
rect 8493 4167 8509 4185
rect 8194 4128 8231 4129
rect 8144 4119 8231 4128
rect 8144 4099 8202 4119
rect 8222 4099 8231 4119
rect 8144 4089 8231 4099
rect 8290 4119 8327 4129
rect 8290 4099 8298 4119
rect 8318 4099 8327 4119
rect 8144 4088 8175 4089
rect 7769 4029 7806 4030
rect 8072 4029 8111 4032
rect 7768 4028 8111 4029
rect 8290 4028 8327 4099
rect 7398 4013 7436 4022
rect 7693 4023 8111 4028
rect 7398 4012 7435 4013
rect 6859 3984 6949 3990
rect 6859 3964 6875 3984
rect 6895 3982 6949 3984
rect 6895 3964 6920 3982
rect 6859 3962 6920 3964
rect 6940 3962 6949 3982
rect 6859 3956 6949 3962
rect 6872 3902 6909 3903
rect 6968 3902 7005 3903
rect 7024 3902 7060 4012
rect 7247 3991 7278 4012
rect 7693 4003 7696 4023
rect 7716 4003 8111 4023
rect 8140 4004 8327 4028
rect 7243 3990 7278 3991
rect 7121 3980 7278 3990
rect 7121 3960 7138 3980
rect 7158 3960 7278 3980
rect 7121 3953 7278 3960
rect 7345 3983 7494 3991
rect 7345 3963 7356 3983
rect 7376 3963 7415 3983
rect 7435 3963 7494 3983
rect 7345 3956 7494 3963
rect 8072 3978 8111 4003
rect 8457 3978 8509 4167
rect 8914 4194 8924 4212
rect 8942 4194 8954 4212
rect 9086 4210 9095 4230
rect 9115 4210 9124 4230
rect 9086 4202 9124 4210
rect 9190 4234 9275 4240
rect 9305 4239 9342 4240
rect 9190 4214 9198 4234
rect 9218 4214 9275 4234
rect 9190 4206 9275 4214
rect 9304 4230 9342 4239
rect 9304 4210 9313 4230
rect 9333 4210 9342 4230
rect 9190 4205 9226 4206
rect 9304 4202 9342 4210
rect 9408 4234 9552 4240
rect 9408 4214 9416 4234
rect 9436 4214 9469 4234
rect 9489 4214 9524 4234
rect 9544 4214 9552 4234
rect 9408 4206 9552 4214
rect 9408 4205 9444 4206
rect 9516 4205 9552 4206
rect 9618 4239 9655 4240
rect 9618 4238 9656 4239
rect 9618 4230 9682 4238
rect 9618 4210 9627 4230
rect 9647 4216 9682 4230
rect 9702 4216 9705 4236
rect 9647 4211 9705 4216
rect 9647 4210 9682 4211
rect 8914 4138 8954 4194
rect 9087 4173 9124 4202
rect 9088 4171 9124 4173
rect 9088 4149 9279 4171
rect 9305 4170 9342 4202
rect 9618 4198 9682 4210
rect 9722 4172 9749 4350
rect 9581 4170 9749 4172
rect 9305 4160 9749 4170
rect 9890 4266 10077 4290
rect 10108 4271 10501 4291
rect 10521 4271 10524 4291
rect 10108 4266 10524 4271
rect 9890 4195 9927 4266
rect 10108 4265 10449 4266
rect 10042 4205 10073 4206
rect 9890 4175 9899 4195
rect 9919 4175 9927 4195
rect 9890 4165 9927 4175
rect 9986 4195 10073 4205
rect 9986 4175 9995 4195
rect 10015 4175 10073 4195
rect 9986 4166 10073 4175
rect 9986 4165 10023 4166
rect 8911 4133 8954 4138
rect 9302 4144 9749 4160
rect 9302 4138 9330 4144
rect 9581 4143 9749 4144
rect 8911 4130 9061 4133
rect 9302 4130 9329 4138
rect 8911 4128 9329 4130
rect 8911 4110 8920 4128
rect 8938 4110 9329 4128
rect 10042 4115 10073 4166
rect 10108 4195 10145 4265
rect 10411 4264 10448 4265
rect 10260 4205 10296 4206
rect 10108 4175 10117 4195
rect 10137 4175 10145 4195
rect 10108 4165 10145 4175
rect 10204 4195 10352 4205
rect 10452 4202 10548 4204
rect 10204 4175 10213 4195
rect 10233 4175 10323 4195
rect 10343 4175 10352 4195
rect 10204 4166 10352 4175
rect 10410 4195 10548 4202
rect 10410 4175 10419 4195
rect 10439 4175 10548 4195
rect 10810 4178 10850 4360
rect 10410 4166 10548 4175
rect 10204 4165 10241 4166
rect 9934 4112 9975 4113
rect 8911 4107 9329 4110
rect 8911 4101 8954 4107
rect 8914 4098 8954 4101
rect 9826 4105 9975 4112
rect 9311 4089 9351 4090
rect 9022 4072 9351 4089
rect 9826 4085 9885 4105
rect 9905 4085 9944 4105
rect 9964 4085 9975 4105
rect 9826 4077 9975 4085
rect 10042 4108 10199 4115
rect 10042 4088 10162 4108
rect 10182 4088 10199 4108
rect 10042 4078 10199 4088
rect 10042 4077 10077 4078
rect 8906 4029 8949 4040
rect 8906 4011 8918 4029
rect 8936 4011 8949 4029
rect 8906 3985 8949 4011
rect 9022 3985 9049 4072
rect 9311 4063 9351 4072
rect 8072 3960 8511 3978
rect 7345 3955 7386 3956
rect 7079 3902 7116 3903
rect 6772 3893 6910 3902
rect 6772 3873 6881 3893
rect 6901 3873 6910 3893
rect 6772 3866 6910 3873
rect 6968 3893 7116 3902
rect 6968 3873 6977 3893
rect 6997 3873 7087 3893
rect 7107 3873 7116 3893
rect 6772 3864 6868 3866
rect 6968 3863 7116 3873
rect 7175 3893 7212 3903
rect 7175 3873 7183 3893
rect 7203 3873 7212 3893
rect 7024 3862 7060 3863
rect 6872 3803 6909 3804
rect 7175 3803 7212 3873
rect 7247 3902 7278 3953
rect 8072 3942 8472 3960
rect 8490 3942 8511 3960
rect 8072 3936 8511 3942
rect 8078 3932 8511 3936
rect 8906 3964 9049 3985
rect 9093 4037 9127 4053
rect 9311 4043 9704 4063
rect 9724 4043 9727 4063
rect 10042 4056 10073 4077
rect 10260 4056 10296 4166
rect 10315 4165 10352 4166
rect 10411 4165 10448 4166
rect 10371 4106 10461 4112
rect 10371 4086 10380 4106
rect 10400 4104 10461 4106
rect 10400 4086 10425 4104
rect 10371 4084 10425 4086
rect 10445 4084 10461 4104
rect 10371 4078 10461 4084
rect 9885 4055 9922 4056
rect 9311 4038 9727 4043
rect 9884 4046 9922 4055
rect 9311 4037 9652 4038
rect 9093 3967 9130 4037
rect 9245 3977 9276 3978
rect 8906 3962 9043 3964
rect 8457 3930 8509 3932
rect 8906 3920 8949 3962
rect 9093 3947 9102 3967
rect 9122 3947 9130 3967
rect 9093 3937 9130 3947
rect 9189 3967 9276 3977
rect 9189 3947 9198 3967
rect 9218 3947 9276 3967
rect 9189 3938 9276 3947
rect 9189 3937 9226 3938
rect 8904 3910 8949 3920
rect 7297 3902 7334 3903
rect 7247 3893 7334 3902
rect 7247 3873 7305 3893
rect 7325 3873 7334 3893
rect 7247 3863 7334 3873
rect 7393 3893 7430 3903
rect 7393 3873 7401 3893
rect 7421 3873 7430 3893
rect 8904 3892 8913 3910
rect 8931 3892 8949 3910
rect 8904 3886 8949 3892
rect 9245 3887 9276 3938
rect 9311 3967 9348 4037
rect 9614 4036 9651 4037
rect 9884 4026 9893 4046
rect 9913 4026 9922 4046
rect 9884 4018 9922 4026
rect 9988 4050 10073 4056
rect 10103 4055 10140 4056
rect 9988 4030 9996 4050
rect 10016 4030 10073 4050
rect 9988 4022 10073 4030
rect 10102 4046 10140 4055
rect 10102 4026 10111 4046
rect 10131 4026 10140 4046
rect 9988 4021 10024 4022
rect 10102 4018 10140 4026
rect 10206 4050 10350 4056
rect 10206 4030 10214 4050
rect 10234 4031 10266 4050
rect 10287 4031 10322 4050
rect 10234 4030 10322 4031
rect 10342 4030 10350 4050
rect 10206 4022 10350 4030
rect 10206 4021 10242 4022
rect 10314 4021 10350 4022
rect 10416 4055 10453 4056
rect 10416 4054 10454 4055
rect 10416 4046 10480 4054
rect 10416 4026 10425 4046
rect 10445 4032 10480 4046
rect 10500 4032 10503 4052
rect 10445 4027 10503 4032
rect 10445 4026 10480 4027
rect 9885 3989 9922 4018
rect 9886 3987 9922 3989
rect 9463 3977 9499 3978
rect 9311 3947 9320 3967
rect 9340 3947 9348 3967
rect 9311 3937 9348 3947
rect 9407 3967 9555 3977
rect 9655 3974 9751 3976
rect 9407 3947 9416 3967
rect 9436 3947 9526 3967
rect 9546 3947 9555 3967
rect 9407 3938 9555 3947
rect 9613 3967 9751 3974
rect 9613 3947 9622 3967
rect 9642 3947 9751 3967
rect 9886 3965 10077 3987
rect 10103 3986 10140 4018
rect 10416 4014 10480 4026
rect 10520 3988 10547 4166
rect 10379 3986 10547 3988
rect 10103 3960 10547 3986
rect 9613 3938 9751 3947
rect 9407 3937 9444 3938
rect 8904 3883 8941 3886
rect 9137 3884 9178 3885
rect 7247 3862 7278 3863
rect 6871 3802 7212 3803
rect 7393 3802 7430 3873
rect 9029 3877 9178 3884
rect 8460 3865 8497 3870
rect 8451 3861 8498 3865
rect 8451 3843 8470 3861
rect 8488 3843 8498 3861
rect 9029 3857 9088 3877
rect 9108 3857 9147 3877
rect 9167 3857 9178 3877
rect 9029 3849 9178 3857
rect 9245 3880 9402 3887
rect 9245 3860 9365 3880
rect 9385 3860 9402 3880
rect 9245 3850 9402 3860
rect 9245 3849 9280 3850
rect 6796 3797 7212 3802
rect 6796 3777 6799 3797
rect 6819 3777 7212 3797
rect 7243 3778 7430 3802
rect 8055 3800 8095 3805
rect 8451 3800 8498 3843
rect 9245 3828 9276 3849
rect 9463 3828 9499 3938
rect 9518 3937 9555 3938
rect 9614 3937 9651 3938
rect 9574 3878 9664 3884
rect 9574 3858 9583 3878
rect 9603 3876 9664 3878
rect 9603 3858 9628 3876
rect 9574 3856 9628 3858
rect 9648 3856 9664 3876
rect 9574 3850 9664 3856
rect 9088 3827 9125 3828
rect 8055 3761 8498 3800
rect 8901 3819 8938 3821
rect 8901 3811 8943 3819
rect 8901 3793 8911 3811
rect 8929 3793 8943 3811
rect 8901 3784 8943 3793
rect 9087 3818 9125 3827
rect 9087 3798 9096 3818
rect 9116 3798 9125 3818
rect 9087 3790 9125 3798
rect 9191 3822 9276 3828
rect 9306 3827 9343 3828
rect 9191 3802 9199 3822
rect 9219 3802 9276 3822
rect 9191 3794 9276 3802
rect 9305 3818 9343 3827
rect 9305 3798 9314 3818
rect 9334 3798 9343 3818
rect 9191 3793 9227 3794
rect 9305 3790 9343 3798
rect 9409 3826 9553 3828
rect 9409 3822 9461 3826
rect 9409 3802 9417 3822
rect 9437 3806 9461 3822
rect 9481 3822 9553 3826
rect 9481 3806 9525 3822
rect 9437 3802 9525 3806
rect 9545 3802 9553 3822
rect 9409 3794 9553 3802
rect 9409 3793 9445 3794
rect 9517 3793 9553 3794
rect 9619 3827 9656 3828
rect 9619 3826 9657 3827
rect 9619 3818 9683 3826
rect 9619 3798 9628 3818
rect 9648 3804 9683 3818
rect 9703 3804 9706 3824
rect 9648 3799 9706 3804
rect 9648 3798 9683 3799
rect 7149 3746 7189 3754
rect 7149 3724 7157 3746
rect 7181 3724 7189 3746
rect 6855 3500 7023 3501
rect 7149 3500 7189 3724
rect 7652 3728 7820 3729
rect 8055 3728 8095 3761
rect 8451 3728 8498 3761
rect 8902 3759 8943 3784
rect 9088 3759 9125 3790
rect 9306 3759 9343 3790
rect 9619 3786 9683 3798
rect 9723 3760 9750 3938
rect 8902 3732 8951 3759
rect 9087 3733 9136 3759
rect 9305 3758 9386 3759
rect 9582 3758 9750 3760
rect 9305 3733 9750 3758
rect 9306 3732 9750 3733
rect 7652 3727 8096 3728
rect 7652 3702 8097 3727
rect 7652 3700 7820 3702
rect 8016 3701 8097 3702
rect 8266 3701 8315 3727
rect 8451 3701 8500 3728
rect 7652 3522 7679 3700
rect 7719 3662 7783 3674
rect 8059 3670 8096 3701
rect 8277 3670 8314 3701
rect 8459 3676 8500 3701
rect 8904 3699 8951 3732
rect 9307 3699 9347 3732
rect 9582 3731 9750 3732
rect 10213 3736 10253 3960
rect 10379 3959 10547 3960
rect 10213 3714 10221 3736
rect 10245 3714 10253 3736
rect 10213 3706 10253 3714
rect 7719 3661 7754 3662
rect 7696 3656 7754 3661
rect 7696 3636 7699 3656
rect 7719 3642 7754 3656
rect 7774 3642 7783 3662
rect 7719 3634 7783 3642
rect 7745 3633 7783 3634
rect 7746 3632 7783 3633
rect 7849 3666 7885 3667
rect 7957 3666 7993 3667
rect 7849 3658 7993 3666
rect 7849 3638 7857 3658
rect 7877 3654 7965 3658
rect 7877 3638 7921 3654
rect 7849 3634 7921 3638
rect 7941 3638 7965 3654
rect 7985 3638 7993 3658
rect 7941 3634 7993 3638
rect 7849 3632 7993 3634
rect 8059 3662 8097 3670
rect 8175 3666 8211 3667
rect 8059 3642 8068 3662
rect 8088 3642 8097 3662
rect 8059 3633 8097 3642
rect 8126 3658 8211 3666
rect 8126 3638 8183 3658
rect 8203 3638 8211 3658
rect 8059 3632 8096 3633
rect 8126 3632 8211 3638
rect 8277 3662 8315 3670
rect 8277 3642 8286 3662
rect 8306 3642 8315 3662
rect 8277 3633 8315 3642
rect 8459 3667 8501 3676
rect 8459 3649 8473 3667
rect 8491 3649 8501 3667
rect 8459 3641 8501 3649
rect 8464 3639 8501 3641
rect 8904 3660 9347 3699
rect 8277 3632 8314 3633
rect 7738 3604 7828 3610
rect 7738 3584 7754 3604
rect 7774 3602 7828 3604
rect 7774 3584 7799 3602
rect 7738 3582 7799 3584
rect 7819 3582 7828 3602
rect 7738 3576 7828 3582
rect 7751 3522 7788 3523
rect 7847 3522 7884 3523
rect 7903 3522 7939 3632
rect 8126 3611 8157 3632
rect 8904 3617 8951 3660
rect 9307 3655 9347 3660
rect 9972 3658 10159 3682
rect 10190 3663 10583 3683
rect 10603 3663 10606 3683
rect 10190 3658 10606 3663
rect 8122 3610 8157 3611
rect 8000 3600 8157 3610
rect 8000 3580 8017 3600
rect 8037 3580 8157 3600
rect 8000 3573 8157 3580
rect 8224 3603 8373 3611
rect 8224 3583 8235 3603
rect 8255 3583 8294 3603
rect 8314 3583 8373 3603
rect 8904 3599 8914 3617
rect 8932 3599 8951 3617
rect 8904 3595 8951 3599
rect 8905 3590 8942 3595
rect 8224 3576 8373 3583
rect 9972 3587 10009 3658
rect 10190 3657 10531 3658
rect 10124 3597 10155 3598
rect 8224 3575 8265 3576
rect 8461 3574 8498 3577
rect 7958 3522 7995 3523
rect 7651 3513 7789 3522
rect 6855 3474 7299 3500
rect 6855 3472 7023 3474
rect 6855 3294 6882 3472
rect 6922 3434 6986 3446
rect 7262 3442 7299 3474
rect 7325 3473 7516 3495
rect 7651 3493 7760 3513
rect 7780 3493 7789 3513
rect 7651 3486 7789 3493
rect 7847 3513 7995 3522
rect 7847 3493 7856 3513
rect 7876 3493 7966 3513
rect 7986 3493 7995 3513
rect 7651 3484 7747 3486
rect 7847 3483 7995 3493
rect 8054 3513 8091 3523
rect 8054 3493 8062 3513
rect 8082 3493 8091 3513
rect 7903 3482 7939 3483
rect 7480 3471 7516 3473
rect 7480 3442 7517 3471
rect 6922 3433 6957 3434
rect 6899 3428 6957 3433
rect 6899 3408 6902 3428
rect 6922 3414 6957 3428
rect 6977 3414 6986 3434
rect 6922 3406 6986 3414
rect 6948 3405 6986 3406
rect 6949 3404 6986 3405
rect 7052 3438 7088 3439
rect 7160 3438 7196 3439
rect 7052 3430 7196 3438
rect 7052 3410 7060 3430
rect 7080 3429 7168 3430
rect 7080 3410 7115 3429
rect 7136 3410 7168 3429
rect 7188 3410 7196 3430
rect 7052 3404 7196 3410
rect 7262 3434 7300 3442
rect 7378 3438 7414 3439
rect 7262 3414 7271 3434
rect 7291 3414 7300 3434
rect 7262 3405 7300 3414
rect 7329 3430 7414 3438
rect 7329 3410 7386 3430
rect 7406 3410 7414 3430
rect 7262 3404 7299 3405
rect 7329 3404 7414 3410
rect 7480 3434 7518 3442
rect 7480 3414 7489 3434
rect 7509 3414 7518 3434
rect 7751 3423 7788 3424
rect 8054 3423 8091 3493
rect 8126 3522 8157 3573
rect 8453 3568 8498 3574
rect 8453 3550 8471 3568
rect 8489 3550 8498 3568
rect 9972 3567 9981 3587
rect 10001 3567 10009 3587
rect 9972 3557 10009 3567
rect 10068 3587 10155 3597
rect 10068 3567 10077 3587
rect 10097 3567 10155 3587
rect 10068 3558 10155 3567
rect 10068 3557 10105 3558
rect 8453 3540 8498 3550
rect 8176 3522 8213 3523
rect 8126 3513 8213 3522
rect 8126 3493 8184 3513
rect 8204 3493 8213 3513
rect 8126 3483 8213 3493
rect 8272 3513 8309 3523
rect 8272 3493 8280 3513
rect 8300 3493 8309 3513
rect 8453 3498 8496 3540
rect 8893 3528 8945 3530
rect 8359 3496 8496 3498
rect 8126 3482 8157 3483
rect 8272 3423 8309 3493
rect 7750 3422 8091 3423
rect 7480 3405 7518 3414
rect 7675 3417 8091 3422
rect 7480 3404 7517 3405
rect 6941 3376 7031 3382
rect 6941 3356 6957 3376
rect 6977 3374 7031 3376
rect 6977 3356 7002 3374
rect 6941 3354 7002 3356
rect 7022 3354 7031 3374
rect 6941 3348 7031 3354
rect 6954 3294 6991 3295
rect 7050 3294 7087 3295
rect 7106 3294 7142 3404
rect 7329 3383 7360 3404
rect 7675 3397 7678 3417
rect 7698 3397 8091 3417
rect 8275 3407 8309 3423
rect 8353 3475 8496 3496
rect 8891 3524 9324 3528
rect 8891 3518 9330 3524
rect 8891 3500 8912 3518
rect 8930 3500 9330 3518
rect 10124 3507 10155 3558
rect 10190 3587 10227 3657
rect 10493 3656 10530 3657
rect 10342 3597 10378 3598
rect 10190 3567 10199 3587
rect 10219 3567 10227 3587
rect 10190 3557 10227 3567
rect 10286 3587 10434 3597
rect 10534 3594 10630 3596
rect 10286 3567 10295 3587
rect 10315 3567 10405 3587
rect 10425 3567 10434 3587
rect 10286 3558 10434 3567
rect 10492 3587 10630 3594
rect 10492 3567 10501 3587
rect 10521 3567 10630 3587
rect 10492 3558 10630 3567
rect 10286 3557 10323 3558
rect 10016 3504 10057 3505
rect 8891 3482 9330 3500
rect 8051 3388 8091 3397
rect 8353 3388 8380 3475
rect 8453 3449 8496 3475
rect 8453 3431 8466 3449
rect 8484 3431 8496 3449
rect 8453 3420 8496 3431
rect 7325 3382 7360 3383
rect 7203 3372 7360 3382
rect 7203 3352 7220 3372
rect 7240 3352 7360 3372
rect 7203 3345 7360 3352
rect 7427 3375 7576 3383
rect 7427 3355 7438 3375
rect 7458 3355 7497 3375
rect 7517 3355 7576 3375
rect 8051 3371 8380 3388
rect 8051 3370 8091 3371
rect 7427 3348 7576 3355
rect 8448 3359 8488 3362
rect 8448 3353 8491 3359
rect 8073 3350 8491 3353
rect 7427 3347 7468 3348
rect 7161 3294 7198 3295
rect 6854 3285 6992 3294
rect 6854 3265 6963 3285
rect 6983 3265 6992 3285
rect 6854 3258 6992 3265
rect 7050 3285 7198 3294
rect 7050 3265 7059 3285
rect 7079 3265 7169 3285
rect 7189 3265 7198 3285
rect 6854 3256 6950 3258
rect 7050 3255 7198 3265
rect 7257 3285 7294 3295
rect 7257 3265 7265 3285
rect 7285 3265 7294 3285
rect 7106 3254 7142 3255
rect 6954 3195 6991 3196
rect 7257 3195 7294 3265
rect 7329 3294 7360 3345
rect 8073 3332 8464 3350
rect 8482 3332 8491 3350
rect 8073 3330 8491 3332
rect 8073 3322 8100 3330
rect 8341 3327 8491 3330
rect 7653 3316 7821 3317
rect 8072 3316 8100 3322
rect 7653 3300 8100 3316
rect 8448 3322 8491 3327
rect 7379 3294 7416 3295
rect 7329 3285 7416 3294
rect 7329 3265 7387 3285
rect 7407 3265 7416 3285
rect 7329 3255 7416 3265
rect 7475 3285 7512 3295
rect 7475 3265 7483 3285
rect 7503 3265 7512 3285
rect 7329 3254 7360 3255
rect 6953 3194 7294 3195
rect 7475 3194 7512 3265
rect 6878 3189 7294 3194
rect 6878 3169 6881 3189
rect 6901 3169 7294 3189
rect 7325 3170 7512 3194
rect 7653 3290 8097 3300
rect 7653 3288 7821 3290
rect 6720 3095 6749 3113
rect 7653 3110 7680 3288
rect 7720 3250 7784 3262
rect 8060 3258 8097 3290
rect 8123 3289 8314 3311
rect 8278 3287 8314 3289
rect 8278 3258 8315 3287
rect 8448 3266 8488 3322
rect 7720 3249 7755 3250
rect 7697 3244 7755 3249
rect 7697 3224 7700 3244
rect 7720 3230 7755 3244
rect 7775 3230 7784 3250
rect 7720 3222 7784 3230
rect 7746 3221 7784 3222
rect 7747 3220 7784 3221
rect 7850 3254 7886 3255
rect 7958 3254 7994 3255
rect 7850 3246 7994 3254
rect 7850 3226 7858 3246
rect 7878 3226 7913 3246
rect 7933 3226 7966 3246
rect 7986 3226 7994 3246
rect 7850 3220 7994 3226
rect 8060 3250 8098 3258
rect 8176 3254 8212 3255
rect 8060 3230 8069 3250
rect 8089 3230 8098 3250
rect 8060 3221 8098 3230
rect 8127 3246 8212 3254
rect 8127 3226 8184 3246
rect 8204 3226 8212 3246
rect 8060 3220 8097 3221
rect 8127 3220 8212 3226
rect 8278 3250 8316 3258
rect 8278 3230 8287 3250
rect 8307 3230 8316 3250
rect 8448 3248 8460 3266
rect 8478 3248 8488 3266
rect 8893 3293 8945 3482
rect 9291 3457 9330 3482
rect 9908 3497 10057 3504
rect 9908 3477 9967 3497
rect 9987 3477 10026 3497
rect 10046 3477 10057 3497
rect 9908 3469 10057 3477
rect 10124 3500 10281 3507
rect 10124 3480 10244 3500
rect 10264 3480 10281 3500
rect 10124 3470 10281 3480
rect 10124 3469 10159 3470
rect 9075 3432 9262 3456
rect 9291 3437 9686 3457
rect 9706 3437 9709 3457
rect 10124 3448 10155 3469
rect 10342 3448 10378 3558
rect 10397 3557 10434 3558
rect 10493 3557 10530 3558
rect 10453 3498 10543 3504
rect 10453 3478 10462 3498
rect 10482 3496 10543 3498
rect 10482 3478 10507 3496
rect 10453 3476 10507 3478
rect 10527 3476 10543 3496
rect 10453 3470 10543 3476
rect 9967 3447 10004 3448
rect 9291 3432 9709 3437
rect 9966 3438 10004 3447
rect 9075 3361 9112 3432
rect 9291 3431 9634 3432
rect 9291 3428 9330 3431
rect 9596 3430 9633 3431
rect 9227 3371 9258 3372
rect 9075 3341 9084 3361
rect 9104 3341 9112 3361
rect 9075 3331 9112 3341
rect 9171 3361 9258 3371
rect 9171 3341 9180 3361
rect 9200 3341 9258 3361
rect 9171 3332 9258 3341
rect 9171 3331 9208 3332
rect 8893 3275 8909 3293
rect 8927 3275 8945 3293
rect 9227 3281 9258 3332
rect 9293 3361 9330 3428
rect 9966 3418 9975 3438
rect 9995 3418 10004 3438
rect 9966 3410 10004 3418
rect 10070 3442 10155 3448
rect 10185 3447 10222 3448
rect 10070 3422 10078 3442
rect 10098 3422 10155 3442
rect 10070 3414 10155 3422
rect 10184 3438 10222 3447
rect 10184 3418 10193 3438
rect 10213 3418 10222 3438
rect 10070 3413 10106 3414
rect 10184 3410 10222 3418
rect 10288 3443 10432 3448
rect 10288 3442 10350 3443
rect 10288 3422 10296 3442
rect 10316 3424 10350 3442
rect 10371 3442 10432 3443
rect 10371 3424 10404 3442
rect 10316 3422 10404 3424
rect 10424 3422 10432 3442
rect 10288 3414 10432 3422
rect 10288 3413 10324 3414
rect 10396 3413 10432 3414
rect 10498 3447 10535 3448
rect 10498 3446 10536 3447
rect 10498 3438 10562 3446
rect 10498 3418 10507 3438
rect 10527 3424 10562 3438
rect 10582 3424 10585 3444
rect 10527 3419 10585 3424
rect 10527 3418 10562 3419
rect 9967 3381 10004 3410
rect 9968 3379 10004 3381
rect 9445 3371 9481 3372
rect 9293 3341 9302 3361
rect 9322 3341 9330 3361
rect 9293 3331 9330 3341
rect 9389 3361 9537 3371
rect 9637 3368 9733 3370
rect 9389 3341 9398 3361
rect 9418 3341 9508 3361
rect 9528 3341 9537 3361
rect 9389 3332 9537 3341
rect 9595 3361 9733 3368
rect 9595 3341 9604 3361
rect 9624 3341 9733 3361
rect 9968 3357 10159 3379
rect 10185 3378 10222 3410
rect 10498 3406 10562 3418
rect 10602 3380 10629 3558
rect 10461 3378 10629 3380
rect 10185 3364 10629 3378
rect 10185 3352 10632 3364
rect 10228 3350 10261 3352
rect 9595 3332 9733 3341
rect 9389 3331 9426 3332
rect 9119 3278 9160 3279
rect 8893 3257 8945 3275
rect 9011 3271 9160 3278
rect 8448 3238 8488 3248
rect 9011 3251 9070 3271
rect 9090 3251 9129 3271
rect 9149 3251 9160 3271
rect 9011 3243 9160 3251
rect 9227 3274 9384 3281
rect 9227 3254 9347 3274
rect 9367 3254 9384 3274
rect 9227 3244 9384 3254
rect 9227 3243 9262 3244
rect 8278 3221 8316 3230
rect 9227 3222 9258 3243
rect 9445 3222 9481 3332
rect 9500 3331 9537 3332
rect 9596 3331 9633 3332
rect 9556 3272 9646 3278
rect 9556 3252 9565 3272
rect 9585 3270 9646 3272
rect 9585 3252 9610 3270
rect 9556 3250 9610 3252
rect 9630 3250 9646 3270
rect 9556 3244 9646 3250
rect 9070 3221 9107 3222
rect 8278 3220 8315 3221
rect 7739 3192 7829 3198
rect 7739 3172 7755 3192
rect 7775 3190 7829 3192
rect 7775 3172 7800 3190
rect 7739 3170 7800 3172
rect 7820 3170 7829 3190
rect 7739 3164 7829 3170
rect 7752 3110 7789 3111
rect 7848 3110 7885 3111
rect 7904 3110 7940 3220
rect 8127 3199 8158 3220
rect 9069 3212 9107 3221
rect 8123 3198 8158 3199
rect 8001 3188 8158 3198
rect 8001 3168 8018 3188
rect 8038 3168 8158 3188
rect 8001 3161 8158 3168
rect 8225 3191 8374 3199
rect 8225 3171 8236 3191
rect 8256 3171 8295 3191
rect 8315 3171 8374 3191
rect 8897 3194 8937 3204
rect 8225 3164 8374 3171
rect 8440 3167 8492 3185
rect 8225 3163 8266 3164
rect 7959 3110 7996 3111
rect 6690 3093 6749 3095
rect 7652 3101 7790 3110
rect 6690 3092 6858 3093
rect 6984 3092 7024 3094
rect 6690 3066 7134 3092
rect 6690 3064 6858 3066
rect 6690 3062 6771 3064
rect 6690 2886 6717 3062
rect 6757 3026 6821 3038
rect 7097 3034 7134 3066
rect 7160 3065 7351 3087
rect 7652 3081 7761 3101
rect 7781 3081 7790 3101
rect 7652 3074 7790 3081
rect 7848 3101 7996 3110
rect 7848 3081 7857 3101
rect 7877 3081 7967 3101
rect 7987 3081 7996 3101
rect 7652 3072 7748 3074
rect 7848 3071 7996 3081
rect 8055 3101 8092 3111
rect 8055 3081 8063 3101
rect 8083 3081 8092 3101
rect 7904 3070 7940 3071
rect 7315 3063 7351 3065
rect 7315 3034 7352 3063
rect 6757 3025 6792 3026
rect 6734 3020 6792 3025
rect 6734 3000 6737 3020
rect 6757 3006 6792 3020
rect 6812 3006 6821 3026
rect 6757 2998 6821 3006
rect 6783 2997 6821 2998
rect 6784 2996 6821 2997
rect 6887 3030 6923 3031
rect 6995 3030 7031 3031
rect 6887 3022 7031 3030
rect 6887 3002 6895 3022
rect 6915 3021 7003 3022
rect 6915 3003 6950 3021
rect 6968 3003 7003 3021
rect 6915 3002 7003 3003
rect 7023 3002 7031 3022
rect 6887 2996 7031 3002
rect 7097 3026 7135 3034
rect 7213 3030 7249 3031
rect 7097 3006 7106 3026
rect 7126 3006 7135 3026
rect 7097 2997 7135 3006
rect 7164 3022 7249 3030
rect 7164 3002 7221 3022
rect 7241 3002 7249 3022
rect 7097 2996 7134 2997
rect 7164 2996 7249 3002
rect 7315 3026 7353 3034
rect 7315 3006 7324 3026
rect 7344 3006 7353 3026
rect 8055 3014 8092 3081
rect 8127 3110 8158 3161
rect 8440 3149 8458 3167
rect 8476 3149 8492 3167
rect 8177 3110 8214 3111
rect 8127 3101 8214 3110
rect 8127 3081 8185 3101
rect 8205 3081 8214 3101
rect 8127 3071 8214 3081
rect 8273 3101 8310 3111
rect 8273 3081 8281 3101
rect 8301 3081 8310 3101
rect 8127 3070 8158 3071
rect 7752 3011 7789 3012
rect 8055 3011 8094 3014
rect 7751 3010 8094 3011
rect 8273 3010 8310 3081
rect 7315 2997 7353 3006
rect 7676 3005 8094 3010
rect 7315 2996 7352 2997
rect 6776 2968 6866 2974
rect 6776 2948 6792 2968
rect 6812 2966 6866 2968
rect 6812 2948 6837 2966
rect 6776 2946 6837 2948
rect 6857 2946 6866 2966
rect 6776 2940 6866 2946
rect 6789 2886 6826 2887
rect 6885 2886 6922 2887
rect 6941 2886 6977 2996
rect 7164 2975 7195 2996
rect 7676 2985 7679 3005
rect 7699 2985 8094 3005
rect 8123 2986 8310 3010
rect 7160 2974 7195 2975
rect 7038 2964 7195 2974
rect 7038 2944 7055 2964
rect 7075 2944 7195 2964
rect 7038 2937 7195 2944
rect 7262 2967 7411 2975
rect 7262 2947 7273 2967
rect 7293 2947 7332 2967
rect 7352 2947 7411 2967
rect 7262 2940 7411 2947
rect 8055 2960 8094 2985
rect 8440 2960 8492 3149
rect 8897 3176 8907 3194
rect 8925 3176 8937 3194
rect 9069 3192 9078 3212
rect 9098 3192 9107 3212
rect 9069 3184 9107 3192
rect 9173 3216 9258 3222
rect 9288 3221 9325 3222
rect 9173 3196 9181 3216
rect 9201 3196 9258 3216
rect 9173 3188 9258 3196
rect 9287 3212 9325 3221
rect 9287 3192 9296 3212
rect 9316 3192 9325 3212
rect 9173 3187 9209 3188
rect 9287 3184 9325 3192
rect 9391 3216 9535 3222
rect 9391 3196 9399 3216
rect 9419 3196 9452 3216
rect 9472 3196 9507 3216
rect 9527 3196 9535 3216
rect 9391 3188 9535 3196
rect 9391 3187 9427 3188
rect 9499 3187 9535 3188
rect 9601 3221 9638 3222
rect 9601 3220 9639 3221
rect 9601 3212 9665 3220
rect 9601 3192 9610 3212
rect 9630 3198 9665 3212
rect 9685 3198 9688 3218
rect 9630 3193 9688 3198
rect 9630 3192 9665 3193
rect 8897 3120 8937 3176
rect 9070 3155 9107 3184
rect 9071 3153 9107 3155
rect 9071 3131 9262 3153
rect 9288 3152 9325 3184
rect 9601 3180 9665 3192
rect 9705 3154 9732 3332
rect 10590 3307 10632 3352
rect 9564 3152 9732 3154
rect 9288 3142 9732 3152
rect 9873 3248 10060 3272
rect 10091 3253 10484 3273
rect 10504 3253 10507 3273
rect 10091 3248 10507 3253
rect 9873 3177 9910 3248
rect 10091 3247 10432 3248
rect 10025 3187 10056 3188
rect 9873 3157 9882 3177
rect 9902 3157 9910 3177
rect 9873 3147 9910 3157
rect 9969 3177 10056 3187
rect 9969 3157 9978 3177
rect 9998 3157 10056 3177
rect 9969 3148 10056 3157
rect 9969 3147 10006 3148
rect 8894 3115 8937 3120
rect 9285 3126 9732 3142
rect 9285 3120 9313 3126
rect 9564 3125 9732 3126
rect 8894 3112 9044 3115
rect 9285 3112 9312 3120
rect 8894 3110 9312 3112
rect 8894 3092 8903 3110
rect 8921 3092 9312 3110
rect 10025 3097 10056 3148
rect 10091 3177 10128 3247
rect 10394 3246 10431 3247
rect 10243 3187 10279 3188
rect 10091 3157 10100 3177
rect 10120 3157 10128 3177
rect 10091 3147 10128 3157
rect 10187 3177 10335 3187
rect 10435 3184 10531 3186
rect 10187 3157 10196 3177
rect 10216 3157 10306 3177
rect 10326 3157 10335 3177
rect 10187 3148 10335 3157
rect 10393 3177 10531 3184
rect 10393 3157 10402 3177
rect 10422 3157 10531 3177
rect 10393 3148 10531 3157
rect 10187 3147 10224 3148
rect 9917 3094 9958 3095
rect 8894 3089 9312 3092
rect 8894 3083 8937 3089
rect 8897 3080 8937 3083
rect 9812 3087 9958 3094
rect 9294 3071 9334 3072
rect 9005 3054 9334 3071
rect 9812 3067 9868 3087
rect 9888 3067 9927 3087
rect 9947 3067 9958 3087
rect 9812 3059 9958 3067
rect 10025 3090 10182 3097
rect 10025 3070 10145 3090
rect 10165 3070 10182 3090
rect 10025 3060 10182 3070
rect 10025 3059 10060 3060
rect 8889 3011 8932 3022
rect 8889 2993 8901 3011
rect 8919 2993 8932 3011
rect 8889 2967 8932 2993
rect 9005 2967 9032 3054
rect 9294 3045 9334 3054
rect 8055 2942 8494 2960
rect 7262 2939 7303 2940
rect 6996 2886 7033 2887
rect 6689 2877 6827 2886
rect 6689 2857 6798 2877
rect 6818 2857 6827 2877
rect 6689 2850 6827 2857
rect 6885 2877 7033 2886
rect 6885 2857 6894 2877
rect 6914 2857 7004 2877
rect 7024 2857 7033 2877
rect 6689 2848 6785 2850
rect 6885 2847 7033 2857
rect 7092 2877 7129 2887
rect 7092 2857 7100 2877
rect 7120 2857 7129 2877
rect 6941 2846 6977 2847
rect 6789 2787 6826 2788
rect 7092 2787 7129 2857
rect 7164 2886 7195 2937
rect 8055 2924 8455 2942
rect 8473 2924 8494 2942
rect 8055 2918 8494 2924
rect 8061 2914 8494 2918
rect 8889 2946 9032 2967
rect 9076 3019 9110 3035
rect 9294 3025 9687 3045
rect 9707 3025 9710 3045
rect 10025 3038 10056 3059
rect 10243 3038 10279 3148
rect 10298 3147 10335 3148
rect 10394 3147 10431 3148
rect 10354 3088 10444 3094
rect 10354 3068 10363 3088
rect 10383 3086 10444 3088
rect 10383 3068 10408 3086
rect 10354 3066 10408 3068
rect 10428 3066 10444 3086
rect 10354 3060 10444 3066
rect 9868 3037 9905 3038
rect 9294 3020 9710 3025
rect 9867 3028 9905 3037
rect 9294 3019 9635 3020
rect 9076 2949 9113 3019
rect 9228 2959 9259 2960
rect 8889 2944 9026 2946
rect 8440 2912 8492 2914
rect 8889 2902 8932 2944
rect 9076 2929 9085 2949
rect 9105 2929 9113 2949
rect 9076 2919 9113 2929
rect 9172 2949 9259 2959
rect 9172 2929 9181 2949
rect 9201 2929 9259 2949
rect 9172 2920 9259 2929
rect 9172 2919 9209 2920
rect 8887 2892 8932 2902
rect 7214 2886 7251 2887
rect 7164 2877 7251 2886
rect 7164 2857 7222 2877
rect 7242 2857 7251 2877
rect 7164 2847 7251 2857
rect 7310 2877 7347 2887
rect 7310 2857 7318 2877
rect 7338 2857 7347 2877
rect 8887 2874 8896 2892
rect 8914 2874 8932 2892
rect 8887 2868 8932 2874
rect 9228 2869 9259 2920
rect 9294 2949 9331 3019
rect 9597 3018 9634 3019
rect 9867 3008 9876 3028
rect 9896 3008 9905 3028
rect 9867 3000 9905 3008
rect 9971 3032 10056 3038
rect 10086 3037 10123 3038
rect 9971 3012 9979 3032
rect 9999 3012 10056 3032
rect 9971 3004 10056 3012
rect 10085 3028 10123 3037
rect 10085 3008 10094 3028
rect 10114 3008 10123 3028
rect 9971 3003 10007 3004
rect 10085 3000 10123 3008
rect 10189 3032 10333 3038
rect 10189 3012 10197 3032
rect 10217 3029 10305 3032
rect 10217 3012 10252 3029
rect 10189 3011 10252 3012
rect 10271 3012 10305 3029
rect 10325 3012 10333 3032
rect 10271 3011 10333 3012
rect 10189 3004 10333 3011
rect 10189 3003 10225 3004
rect 10297 3003 10333 3004
rect 10399 3037 10436 3038
rect 10399 3036 10437 3037
rect 10459 3036 10486 3040
rect 10399 3034 10486 3036
rect 10399 3028 10463 3034
rect 10399 3008 10408 3028
rect 10428 3014 10463 3028
rect 10483 3014 10486 3034
rect 10428 3009 10486 3014
rect 10428 3008 10463 3009
rect 9868 2971 9905 3000
rect 9869 2969 9905 2971
rect 9446 2959 9482 2960
rect 9294 2929 9303 2949
rect 9323 2929 9331 2949
rect 9294 2919 9331 2929
rect 9390 2949 9538 2959
rect 9638 2956 9734 2958
rect 9390 2929 9399 2949
rect 9419 2929 9509 2949
rect 9529 2929 9538 2949
rect 9390 2920 9538 2929
rect 9596 2949 9734 2956
rect 9596 2929 9605 2949
rect 9625 2929 9734 2949
rect 9869 2947 10060 2969
rect 10086 2968 10123 3000
rect 10399 2996 10463 3008
rect 10503 2970 10530 3148
rect 10362 2968 10530 2970
rect 10086 2942 10530 2968
rect 9596 2920 9734 2929
rect 9390 2919 9427 2920
rect 8887 2865 8924 2868
rect 9120 2866 9161 2867
rect 7164 2846 7195 2847
rect 6788 2786 7129 2787
rect 7310 2786 7347 2857
rect 9012 2859 9161 2866
rect 8443 2847 8480 2852
rect 6713 2781 7129 2786
rect 6713 2761 6716 2781
rect 6736 2761 7129 2781
rect 7160 2762 7347 2786
rect 8434 2843 8481 2847
rect 8434 2825 8453 2843
rect 8471 2825 8481 2843
rect 9012 2839 9071 2859
rect 9091 2839 9130 2859
rect 9150 2839 9161 2859
rect 9012 2831 9161 2839
rect 9228 2862 9385 2869
rect 9228 2842 9348 2862
rect 9368 2842 9385 2862
rect 9228 2832 9385 2842
rect 9228 2831 9263 2832
rect 8434 2777 8481 2825
rect 9228 2810 9259 2831
rect 9446 2810 9482 2920
rect 9501 2919 9538 2920
rect 9597 2919 9634 2920
rect 9557 2860 9647 2866
rect 9557 2840 9566 2860
rect 9586 2858 9647 2860
rect 9586 2840 9611 2858
rect 9557 2838 9611 2840
rect 9631 2838 9647 2858
rect 9557 2832 9647 2838
rect 9071 2809 9108 2810
rect 8058 2774 8481 2777
rect 6933 2760 6998 2761
rect 8036 2744 8481 2774
rect 8883 2801 8921 2803
rect 8883 2793 8926 2801
rect 8883 2775 8894 2793
rect 8912 2775 8926 2793
rect 8883 2748 8926 2775
rect 9070 2800 9108 2809
rect 9070 2780 9079 2800
rect 9099 2780 9108 2800
rect 9070 2772 9108 2780
rect 9174 2804 9259 2810
rect 9289 2809 9326 2810
rect 9174 2784 9182 2804
rect 9202 2784 9259 2804
rect 9174 2776 9259 2784
rect 9288 2800 9326 2809
rect 9288 2780 9297 2800
rect 9317 2780 9326 2800
rect 9174 2775 9210 2776
rect 9288 2772 9326 2780
rect 9392 2808 9536 2810
rect 9392 2804 9444 2808
rect 9392 2784 9400 2804
rect 9420 2788 9444 2804
rect 9464 2804 9536 2808
rect 9464 2788 9508 2804
rect 9420 2784 9508 2788
rect 9528 2784 9536 2804
rect 9392 2776 9536 2784
rect 9392 2775 9428 2776
rect 9500 2775 9536 2776
rect 9602 2809 9639 2810
rect 9602 2808 9640 2809
rect 9602 2800 9666 2808
rect 9602 2780 9611 2800
rect 9631 2786 9666 2800
rect 9686 2786 9689 2806
rect 9631 2781 9689 2786
rect 9631 2780 9666 2781
rect 7129 2728 7169 2736
rect 7129 2706 7137 2728
rect 7161 2706 7169 2728
rect 6734 2477 6771 2483
rect 6734 2458 6742 2477
rect 6763 2458 6771 2477
rect 6734 2450 6771 2458
rect 6434 2329 6441 2351
rect 6465 2329 6473 2351
rect 6434 2323 6473 2329
rect 5964 2318 6004 2320
rect 6130 2319 6298 2320
rect 6232 2318 6269 2319
rect 5198 2302 5336 2311
rect 4992 2301 5029 2302
rect 4722 2248 4763 2249
rect 4496 2227 4548 2245
rect 4614 2241 4763 2248
rect 4064 2207 4104 2217
rect 4614 2221 4673 2241
rect 4693 2221 4732 2241
rect 4752 2221 4763 2241
rect 4614 2213 4763 2221
rect 4830 2244 4987 2251
rect 4830 2224 4950 2244
rect 4970 2224 4987 2244
rect 4830 2214 4987 2224
rect 4830 2213 4865 2214
rect 3894 2190 3932 2199
rect 4830 2192 4861 2213
rect 5048 2192 5084 2302
rect 5103 2301 5140 2302
rect 5199 2301 5236 2302
rect 5159 2242 5249 2248
rect 5159 2222 5168 2242
rect 5188 2240 5249 2242
rect 5188 2222 5213 2240
rect 5159 2220 5213 2222
rect 5233 2220 5249 2240
rect 5159 2214 5249 2220
rect 4673 2191 4710 2192
rect 3894 2189 3931 2190
rect 3355 2161 3445 2167
rect 3355 2141 3371 2161
rect 3391 2159 3445 2161
rect 3391 2141 3416 2159
rect 3355 2139 3416 2141
rect 3436 2139 3445 2159
rect 3355 2133 3445 2139
rect 3368 2079 3405 2080
rect 3464 2079 3501 2080
rect 3520 2079 3556 2189
rect 3743 2168 3774 2189
rect 4672 2182 4710 2191
rect 3739 2167 3774 2168
rect 3617 2157 3774 2167
rect 3617 2137 3634 2157
rect 3654 2137 3774 2157
rect 3617 2130 3774 2137
rect 3841 2160 3990 2168
rect 3841 2140 3852 2160
rect 3872 2140 3911 2160
rect 3931 2140 3990 2160
rect 4500 2164 4540 2174
rect 3841 2133 3990 2140
rect 4056 2136 4108 2154
rect 3841 2132 3882 2133
rect 3575 2079 3612 2080
rect 3268 2070 3406 2079
rect 2740 2059 2773 2061
rect 2369 2047 2816 2059
rect 1601 1925 1769 1927
rect 1325 1899 1769 1925
rect 835 1877 973 1886
rect 629 1876 666 1877
rect 126 1822 163 1825
rect 359 1823 400 1824
rect 251 1816 400 1823
rect 251 1796 310 1816
rect 330 1796 369 1816
rect 389 1796 400 1816
rect 251 1788 400 1796
rect 467 1819 624 1826
rect 467 1799 587 1819
rect 607 1799 624 1819
rect 467 1789 624 1799
rect 467 1788 502 1789
rect 467 1767 498 1788
rect 685 1767 721 1877
rect 740 1876 777 1877
rect 836 1876 873 1877
rect 796 1817 886 1823
rect 796 1797 805 1817
rect 825 1815 886 1817
rect 825 1797 850 1815
rect 796 1795 850 1797
rect 870 1795 886 1815
rect 796 1789 886 1795
rect 310 1766 347 1767
rect 123 1758 160 1760
rect 123 1750 165 1758
rect 123 1732 133 1750
rect 151 1732 165 1750
rect 123 1723 165 1732
rect 309 1757 347 1766
rect 309 1737 318 1757
rect 338 1737 347 1757
rect 309 1729 347 1737
rect 413 1761 498 1767
rect 528 1766 565 1767
rect 413 1741 421 1761
rect 441 1741 498 1761
rect 413 1733 498 1741
rect 527 1757 565 1766
rect 527 1737 536 1757
rect 556 1737 565 1757
rect 413 1732 449 1733
rect 527 1729 565 1737
rect 631 1765 775 1767
rect 631 1761 683 1765
rect 631 1741 639 1761
rect 659 1745 683 1761
rect 703 1761 775 1765
rect 703 1745 747 1761
rect 659 1741 747 1745
rect 767 1741 775 1761
rect 631 1733 775 1741
rect 631 1732 667 1733
rect 739 1732 775 1733
rect 841 1766 878 1767
rect 841 1765 879 1766
rect 841 1757 905 1765
rect 841 1737 850 1757
rect 870 1743 905 1757
rect 925 1743 928 1763
rect 870 1738 928 1743
rect 870 1737 905 1738
rect 124 1698 165 1723
rect 310 1698 347 1729
rect 528 1698 565 1729
rect 841 1725 905 1737
rect 945 1699 972 1877
rect 124 1671 173 1698
rect 309 1672 358 1698
rect 527 1697 608 1698
rect 804 1697 972 1699
rect 527 1672 972 1697
rect 528 1671 972 1672
rect 126 1638 173 1671
rect 529 1638 569 1671
rect 804 1670 972 1671
rect 1435 1675 1475 1899
rect 1601 1898 1769 1899
rect 2372 2033 2816 2047
rect 2372 2031 2540 2033
rect 2372 1853 2399 2031
rect 2439 1993 2503 2005
rect 2779 2001 2816 2033
rect 2842 2032 3033 2054
rect 3268 2050 3377 2070
rect 3397 2050 3406 2070
rect 3268 2043 3406 2050
rect 3464 2070 3612 2079
rect 3464 2050 3473 2070
rect 3493 2050 3583 2070
rect 3603 2050 3612 2070
rect 3268 2041 3364 2043
rect 3464 2040 3612 2050
rect 3671 2070 3708 2080
rect 3671 2050 3679 2070
rect 3699 2050 3708 2070
rect 3520 2039 3556 2040
rect 2997 2030 3033 2032
rect 2997 2001 3034 2030
rect 2439 1992 2474 1993
rect 2416 1987 2474 1992
rect 2416 1967 2419 1987
rect 2439 1973 2474 1987
rect 2494 1973 2503 1993
rect 2439 1965 2503 1973
rect 2465 1964 2503 1965
rect 2466 1963 2503 1964
rect 2569 1997 2605 1998
rect 2677 1997 2713 1998
rect 2569 1989 2713 1997
rect 2569 1969 2577 1989
rect 2597 1987 2685 1989
rect 2597 1969 2630 1987
rect 2569 1968 2630 1969
rect 2651 1969 2685 1987
rect 2705 1969 2713 1989
rect 2651 1968 2713 1969
rect 2569 1963 2713 1968
rect 2779 1993 2817 2001
rect 2895 1997 2931 1998
rect 2779 1973 2788 1993
rect 2808 1973 2817 1993
rect 2779 1964 2817 1973
rect 2846 1989 2931 1997
rect 2846 1969 2903 1989
rect 2923 1969 2931 1989
rect 2779 1963 2816 1964
rect 2846 1963 2931 1969
rect 2997 1993 3035 2001
rect 2997 1973 3006 1993
rect 3026 1973 3035 1993
rect 3671 1983 3708 2050
rect 3743 2079 3774 2130
rect 4056 2118 4074 2136
rect 4092 2118 4108 2136
rect 3793 2079 3830 2080
rect 3743 2070 3830 2079
rect 3743 2050 3801 2070
rect 3821 2050 3830 2070
rect 3743 2040 3830 2050
rect 3889 2070 3926 2080
rect 3889 2050 3897 2070
rect 3917 2050 3926 2070
rect 3743 2039 3774 2040
rect 3368 1980 3405 1981
rect 3671 1980 3710 1983
rect 3367 1979 3710 1980
rect 3889 1979 3926 2050
rect 2997 1964 3035 1973
rect 3292 1974 3710 1979
rect 2997 1963 3034 1964
rect 2458 1935 2548 1941
rect 2458 1915 2474 1935
rect 2494 1933 2548 1935
rect 2494 1915 2519 1933
rect 2458 1913 2519 1915
rect 2539 1913 2548 1933
rect 2458 1907 2548 1913
rect 2471 1853 2508 1854
rect 2567 1853 2604 1854
rect 2623 1853 2659 1963
rect 2846 1942 2877 1963
rect 3292 1954 3295 1974
rect 3315 1954 3710 1974
rect 3739 1955 3926 1979
rect 2842 1941 2877 1942
rect 2720 1931 2877 1941
rect 2720 1911 2737 1931
rect 2757 1911 2877 1931
rect 2720 1904 2877 1911
rect 2944 1934 3093 1942
rect 2944 1914 2955 1934
rect 2975 1914 3014 1934
rect 3034 1914 3093 1934
rect 2944 1907 3093 1914
rect 3671 1929 3710 1954
rect 4056 1929 4108 2118
rect 4500 2146 4510 2164
rect 4528 2146 4540 2164
rect 4672 2162 4681 2182
rect 4701 2162 4710 2182
rect 4672 2154 4710 2162
rect 4776 2186 4861 2192
rect 4891 2191 4928 2192
rect 4776 2166 4784 2186
rect 4804 2166 4861 2186
rect 4776 2158 4861 2166
rect 4890 2182 4928 2191
rect 4890 2162 4899 2182
rect 4919 2162 4928 2182
rect 4776 2157 4812 2158
rect 4890 2154 4928 2162
rect 4994 2186 5138 2192
rect 4994 2166 5002 2186
rect 5022 2166 5055 2186
rect 5075 2166 5110 2186
rect 5130 2166 5138 2186
rect 4994 2158 5138 2166
rect 4994 2157 5030 2158
rect 5102 2157 5138 2158
rect 5204 2191 5241 2192
rect 5204 2190 5242 2191
rect 5204 2182 5268 2190
rect 5204 2162 5213 2182
rect 5233 2168 5268 2182
rect 5288 2168 5291 2188
rect 5233 2163 5291 2168
rect 5233 2162 5268 2163
rect 4500 2090 4540 2146
rect 4673 2125 4710 2154
rect 4674 2123 4710 2125
rect 4674 2101 4865 2123
rect 4891 2122 4928 2154
rect 5204 2150 5268 2162
rect 5308 2124 5335 2302
rect 5167 2122 5335 2124
rect 4891 2112 5335 2122
rect 5476 2218 5663 2242
rect 5694 2223 6087 2243
rect 6107 2223 6110 2243
rect 5694 2218 6110 2223
rect 5476 2147 5513 2218
rect 5694 2217 6035 2218
rect 5628 2157 5659 2158
rect 5476 2127 5485 2147
rect 5505 2127 5513 2147
rect 5476 2117 5513 2127
rect 5572 2147 5659 2157
rect 5572 2127 5581 2147
rect 5601 2127 5659 2147
rect 5572 2118 5659 2127
rect 5572 2117 5609 2118
rect 4497 2085 4540 2090
rect 4888 2096 5335 2112
rect 4888 2090 4916 2096
rect 5167 2095 5335 2096
rect 4497 2082 4647 2085
rect 4888 2082 4915 2090
rect 4497 2080 4915 2082
rect 4497 2062 4506 2080
rect 4524 2062 4915 2080
rect 5628 2067 5659 2118
rect 5694 2147 5731 2217
rect 5997 2216 6034 2217
rect 6235 2159 6268 2318
rect 5846 2157 5882 2158
rect 5694 2127 5703 2147
rect 5723 2127 5731 2147
rect 5694 2117 5731 2127
rect 5790 2147 5938 2157
rect 6038 2154 6134 2156
rect 5790 2127 5799 2147
rect 5819 2127 5909 2147
rect 5929 2127 5938 2147
rect 5790 2118 5938 2127
rect 5996 2147 6134 2154
rect 5996 2127 6005 2147
rect 6025 2127 6134 2147
rect 6235 2155 6271 2159
rect 6235 2137 6244 2155
rect 6266 2137 6271 2155
rect 6235 2131 6271 2137
rect 5996 2118 6134 2127
rect 5790 2117 5827 2118
rect 5520 2064 5561 2065
rect 4497 2059 4915 2062
rect 4497 2053 4540 2059
rect 4500 2050 4540 2053
rect 5412 2057 5561 2064
rect 4897 2041 4937 2042
rect 4608 2024 4937 2041
rect 5412 2037 5471 2057
rect 5491 2037 5530 2057
rect 5550 2037 5561 2057
rect 5412 2029 5561 2037
rect 5628 2060 5785 2067
rect 5628 2040 5748 2060
rect 5768 2040 5785 2060
rect 5628 2030 5785 2040
rect 5628 2029 5663 2030
rect 4492 1981 4535 1992
rect 4492 1963 4504 1981
rect 4522 1963 4535 1981
rect 4492 1937 4535 1963
rect 4608 1937 4635 2024
rect 4897 2015 4937 2024
rect 3671 1911 4110 1929
rect 2944 1906 2985 1907
rect 2678 1853 2715 1854
rect 2371 1844 2509 1853
rect 2371 1824 2480 1844
rect 2500 1824 2509 1844
rect 2371 1817 2509 1824
rect 2567 1844 2715 1853
rect 2567 1824 2576 1844
rect 2596 1824 2686 1844
rect 2706 1824 2715 1844
rect 2371 1815 2467 1817
rect 2567 1814 2715 1824
rect 2774 1844 2811 1854
rect 2774 1824 2782 1844
rect 2802 1824 2811 1844
rect 2623 1813 2659 1814
rect 2471 1754 2508 1755
rect 2774 1754 2811 1824
rect 2846 1853 2877 1904
rect 3671 1893 4071 1911
rect 4089 1893 4110 1911
rect 3671 1887 4110 1893
rect 3677 1883 4110 1887
rect 4492 1916 4635 1937
rect 4679 1989 4713 2005
rect 4897 1995 5290 2015
rect 5310 1995 5313 2015
rect 5628 2008 5659 2029
rect 5846 2008 5882 2118
rect 5901 2117 5938 2118
rect 5997 2117 6034 2118
rect 5957 2058 6047 2064
rect 5957 2038 5966 2058
rect 5986 2056 6047 2058
rect 5986 2038 6011 2056
rect 5957 2036 6011 2038
rect 6031 2036 6047 2056
rect 5957 2030 6047 2036
rect 5471 2007 5508 2008
rect 4897 1990 5313 1995
rect 5470 1998 5508 2007
rect 4897 1989 5238 1990
rect 4679 1919 4716 1989
rect 4831 1929 4862 1930
rect 4492 1914 4629 1916
rect 4056 1881 4108 1883
rect 4492 1872 4535 1914
rect 4679 1899 4688 1919
rect 4708 1899 4716 1919
rect 4679 1889 4716 1899
rect 4775 1919 4862 1929
rect 4775 1899 4784 1919
rect 4804 1899 4862 1919
rect 4775 1890 4862 1899
rect 4775 1889 4812 1890
rect 4490 1862 4535 1872
rect 2896 1853 2933 1854
rect 2846 1844 2933 1853
rect 2846 1824 2904 1844
rect 2924 1824 2933 1844
rect 2846 1814 2933 1824
rect 2992 1844 3029 1854
rect 2992 1824 3000 1844
rect 3020 1824 3029 1844
rect 4490 1844 4499 1862
rect 4517 1844 4535 1862
rect 4490 1838 4535 1844
rect 4831 1839 4862 1890
rect 4897 1919 4934 1989
rect 5200 1988 5237 1989
rect 5470 1978 5479 1998
rect 5499 1978 5508 1998
rect 5470 1970 5508 1978
rect 5574 2002 5659 2008
rect 5689 2007 5726 2008
rect 5574 1982 5582 2002
rect 5602 1982 5659 2002
rect 5574 1974 5659 1982
rect 5688 1998 5726 2007
rect 5688 1978 5697 1998
rect 5717 1978 5726 1998
rect 5574 1973 5610 1974
rect 5688 1970 5726 1978
rect 5792 2002 5936 2008
rect 5792 1982 5800 2002
rect 5820 1983 5852 2002
rect 5873 1983 5908 2002
rect 5820 1982 5908 1983
rect 5928 1982 5936 2002
rect 5792 1974 5936 1982
rect 5792 1973 5828 1974
rect 5900 1973 5936 1974
rect 6002 2007 6039 2008
rect 6002 2006 6040 2007
rect 6002 1998 6066 2006
rect 6002 1978 6011 1998
rect 6031 1984 6066 1998
rect 6086 1984 6089 2004
rect 6031 1979 6089 1984
rect 6031 1978 6066 1979
rect 5471 1941 5508 1970
rect 5472 1939 5508 1941
rect 5049 1929 5085 1930
rect 4897 1899 4906 1919
rect 4926 1899 4934 1919
rect 4897 1889 4934 1899
rect 4993 1919 5141 1929
rect 5241 1926 5337 1928
rect 4993 1899 5002 1919
rect 5022 1899 5112 1919
rect 5132 1899 5141 1919
rect 4993 1890 5141 1899
rect 5199 1919 5337 1926
rect 5199 1899 5208 1919
rect 5228 1899 5337 1919
rect 5472 1917 5663 1939
rect 5689 1938 5726 1970
rect 6002 1966 6066 1978
rect 6106 1940 6133 2118
rect 6738 2117 6771 2450
rect 6835 2482 7003 2483
rect 7129 2482 7169 2706
rect 7632 2710 7800 2711
rect 8036 2710 8077 2744
rect 8434 2723 8481 2744
rect 7632 2700 8077 2710
rect 8149 2708 8292 2709
rect 7632 2684 8076 2700
rect 7632 2682 7800 2684
rect 7996 2683 8076 2684
rect 8149 2683 8294 2708
rect 8436 2683 8481 2723
rect 7632 2504 7659 2682
rect 7699 2644 7763 2656
rect 8039 2652 8076 2683
rect 8257 2652 8294 2683
rect 8439 2676 8481 2683
rect 8884 2741 8926 2748
rect 9071 2741 9108 2772
rect 9289 2741 9326 2772
rect 9602 2768 9666 2780
rect 9706 2742 9733 2920
rect 8884 2701 8929 2741
rect 9071 2716 9216 2741
rect 9289 2740 9369 2741
rect 9565 2740 9733 2742
rect 9289 2724 9733 2740
rect 9073 2715 9216 2716
rect 9288 2714 9733 2724
rect 8884 2680 8931 2701
rect 9288 2680 9329 2714
rect 9565 2713 9733 2714
rect 10196 2718 10236 2942
rect 10362 2941 10530 2942
rect 10594 2974 10627 3307
rect 10594 2966 10631 2974
rect 10594 2947 10602 2966
rect 10623 2947 10631 2966
rect 10594 2941 10631 2947
rect 10196 2696 10204 2718
rect 10228 2696 10236 2718
rect 10196 2688 10236 2696
rect 7699 2643 7734 2644
rect 7676 2638 7734 2643
rect 7676 2618 7679 2638
rect 7699 2624 7734 2638
rect 7754 2624 7763 2644
rect 7699 2616 7763 2624
rect 7725 2615 7763 2616
rect 7726 2614 7763 2615
rect 7829 2648 7865 2649
rect 7937 2648 7973 2649
rect 7829 2640 7973 2648
rect 7829 2620 7837 2640
rect 7857 2636 7945 2640
rect 7857 2620 7901 2636
rect 7829 2616 7901 2620
rect 7921 2620 7945 2636
rect 7965 2620 7973 2640
rect 7921 2616 7973 2620
rect 7829 2614 7973 2616
rect 8039 2644 8077 2652
rect 8155 2648 8191 2649
rect 8039 2624 8048 2644
rect 8068 2624 8077 2644
rect 8039 2615 8077 2624
rect 8106 2640 8191 2648
rect 8106 2620 8163 2640
rect 8183 2620 8191 2640
rect 8039 2614 8076 2615
rect 8106 2614 8191 2620
rect 8257 2644 8295 2652
rect 8257 2624 8266 2644
rect 8286 2624 8295 2644
rect 8257 2615 8295 2624
rect 8439 2649 8482 2676
rect 8439 2631 8453 2649
rect 8471 2631 8482 2649
rect 8439 2623 8482 2631
rect 8444 2621 8482 2623
rect 8884 2650 9329 2680
rect 10367 2663 10432 2664
rect 8884 2647 9307 2650
rect 8257 2614 8294 2615
rect 7718 2586 7808 2592
rect 7718 2566 7734 2586
rect 7754 2584 7808 2586
rect 7754 2566 7779 2584
rect 7718 2564 7779 2566
rect 7799 2564 7808 2584
rect 7718 2558 7808 2564
rect 7731 2504 7768 2505
rect 7827 2504 7864 2505
rect 7883 2504 7919 2614
rect 8106 2593 8137 2614
rect 8884 2599 8931 2647
rect 8102 2592 8137 2593
rect 7980 2582 8137 2592
rect 7980 2562 7997 2582
rect 8017 2562 8137 2582
rect 7980 2555 8137 2562
rect 8204 2585 8353 2593
rect 8204 2565 8215 2585
rect 8235 2565 8274 2585
rect 8294 2565 8353 2585
rect 8884 2581 8894 2599
rect 8912 2581 8931 2599
rect 8884 2577 8931 2581
rect 10018 2638 10205 2662
rect 10236 2643 10629 2663
rect 10649 2643 10652 2663
rect 10236 2638 10652 2643
rect 8885 2572 8922 2577
rect 8204 2558 8353 2565
rect 10018 2567 10055 2638
rect 10236 2637 10577 2638
rect 10170 2577 10201 2578
rect 8204 2557 8245 2558
rect 8441 2556 8478 2559
rect 7938 2504 7975 2505
rect 7631 2495 7769 2504
rect 6835 2456 7279 2482
rect 6835 2454 7003 2456
rect 6835 2276 6862 2454
rect 6902 2416 6966 2428
rect 7242 2424 7279 2456
rect 7305 2455 7496 2477
rect 7631 2475 7740 2495
rect 7760 2475 7769 2495
rect 7631 2468 7769 2475
rect 7827 2495 7975 2504
rect 7827 2475 7836 2495
rect 7856 2475 7946 2495
rect 7966 2475 7975 2495
rect 7631 2466 7727 2468
rect 7827 2465 7975 2475
rect 8034 2495 8071 2505
rect 8034 2475 8042 2495
rect 8062 2475 8071 2495
rect 7883 2464 7919 2465
rect 7460 2453 7496 2455
rect 7460 2424 7497 2453
rect 6902 2415 6937 2416
rect 6879 2410 6937 2415
rect 6879 2390 6882 2410
rect 6902 2396 6937 2410
rect 6957 2396 6966 2416
rect 6902 2390 6966 2396
rect 6879 2388 6966 2390
rect 6879 2384 6906 2388
rect 6928 2387 6966 2388
rect 6929 2386 6966 2387
rect 7032 2420 7068 2421
rect 7140 2420 7176 2421
rect 7032 2413 7176 2420
rect 7032 2412 7094 2413
rect 7032 2392 7040 2412
rect 7060 2395 7094 2412
rect 7113 2412 7176 2413
rect 7113 2395 7148 2412
rect 7060 2392 7148 2395
rect 7168 2392 7176 2412
rect 7032 2386 7176 2392
rect 7242 2416 7280 2424
rect 7358 2420 7394 2421
rect 7242 2396 7251 2416
rect 7271 2396 7280 2416
rect 7242 2387 7280 2396
rect 7309 2412 7394 2420
rect 7309 2392 7366 2412
rect 7386 2392 7394 2412
rect 7242 2386 7279 2387
rect 7309 2386 7394 2392
rect 7460 2416 7498 2424
rect 7460 2396 7469 2416
rect 7489 2396 7498 2416
rect 7731 2405 7768 2406
rect 8034 2405 8071 2475
rect 8106 2504 8137 2555
rect 8433 2550 8478 2556
rect 8433 2532 8451 2550
rect 8469 2532 8478 2550
rect 10018 2547 10027 2567
rect 10047 2547 10055 2567
rect 10018 2537 10055 2547
rect 10114 2567 10201 2577
rect 10114 2547 10123 2567
rect 10143 2547 10201 2567
rect 10114 2538 10201 2547
rect 10114 2537 10151 2538
rect 8433 2522 8478 2532
rect 8156 2504 8193 2505
rect 8106 2495 8193 2504
rect 8106 2475 8164 2495
rect 8184 2475 8193 2495
rect 8106 2465 8193 2475
rect 8252 2495 8289 2505
rect 8252 2475 8260 2495
rect 8280 2475 8289 2495
rect 8433 2480 8476 2522
rect 8873 2510 8925 2512
rect 8339 2478 8476 2480
rect 8106 2464 8137 2465
rect 8252 2405 8289 2475
rect 7730 2404 8071 2405
rect 7460 2387 7498 2396
rect 7655 2399 8071 2404
rect 7460 2386 7497 2387
rect 6921 2358 7011 2364
rect 6921 2338 6937 2358
rect 6957 2356 7011 2358
rect 6957 2338 6982 2356
rect 6921 2336 6982 2338
rect 7002 2336 7011 2356
rect 6921 2330 7011 2336
rect 6934 2276 6971 2277
rect 7030 2276 7067 2277
rect 7086 2276 7122 2386
rect 7309 2365 7340 2386
rect 7655 2379 7658 2399
rect 7678 2379 8071 2399
rect 8255 2389 8289 2405
rect 8333 2457 8476 2478
rect 8871 2506 9304 2510
rect 8871 2500 9310 2506
rect 8871 2482 8892 2500
rect 8910 2482 9310 2500
rect 10170 2487 10201 2538
rect 10236 2567 10273 2637
rect 10539 2636 10576 2637
rect 10388 2577 10424 2578
rect 10236 2547 10245 2567
rect 10265 2547 10273 2567
rect 10236 2537 10273 2547
rect 10332 2567 10480 2577
rect 10580 2574 10676 2576
rect 10332 2547 10341 2567
rect 10361 2547 10451 2567
rect 10471 2547 10480 2567
rect 10332 2538 10480 2547
rect 10538 2567 10676 2574
rect 10538 2547 10547 2567
rect 10567 2547 10676 2567
rect 10538 2538 10676 2547
rect 10332 2537 10369 2538
rect 10062 2484 10103 2485
rect 8871 2464 9310 2482
rect 8031 2370 8071 2379
rect 8333 2370 8360 2457
rect 8433 2431 8476 2457
rect 8433 2413 8446 2431
rect 8464 2413 8476 2431
rect 8433 2402 8476 2413
rect 7305 2364 7340 2365
rect 7183 2354 7340 2364
rect 7183 2334 7200 2354
rect 7220 2334 7340 2354
rect 7183 2327 7340 2334
rect 7407 2357 7553 2365
rect 7407 2337 7418 2357
rect 7438 2337 7477 2357
rect 7497 2337 7553 2357
rect 8031 2353 8360 2370
rect 8031 2352 8071 2353
rect 7407 2330 7553 2337
rect 8428 2341 8468 2344
rect 8428 2335 8471 2341
rect 8053 2332 8471 2335
rect 7407 2329 7448 2330
rect 7141 2276 7178 2277
rect 6834 2267 6972 2276
rect 6834 2247 6943 2267
rect 6963 2247 6972 2267
rect 6834 2240 6972 2247
rect 7030 2267 7178 2276
rect 7030 2247 7039 2267
rect 7059 2247 7149 2267
rect 7169 2247 7178 2267
rect 6834 2238 6930 2240
rect 7030 2237 7178 2247
rect 7237 2267 7274 2277
rect 7237 2247 7245 2267
rect 7265 2247 7274 2267
rect 7086 2236 7122 2237
rect 6934 2177 6971 2178
rect 7237 2177 7274 2247
rect 7309 2276 7340 2327
rect 8053 2314 8444 2332
rect 8462 2314 8471 2332
rect 8053 2312 8471 2314
rect 8053 2304 8080 2312
rect 8321 2309 8471 2312
rect 7633 2298 7801 2299
rect 8052 2298 8080 2304
rect 7633 2282 8080 2298
rect 8428 2304 8471 2309
rect 7359 2276 7396 2277
rect 7309 2267 7396 2276
rect 7309 2247 7367 2267
rect 7387 2247 7396 2267
rect 7309 2237 7396 2247
rect 7455 2267 7492 2277
rect 7455 2247 7463 2267
rect 7483 2247 7492 2267
rect 7309 2236 7340 2237
rect 6933 2176 7274 2177
rect 7455 2176 7492 2247
rect 6858 2171 7274 2176
rect 6858 2151 6861 2171
rect 6881 2151 7274 2171
rect 7305 2152 7492 2176
rect 7633 2272 8077 2282
rect 7633 2270 7801 2272
rect 6733 2072 6775 2117
rect 7633 2092 7660 2270
rect 7700 2232 7764 2244
rect 8040 2240 8077 2272
rect 8103 2271 8294 2293
rect 8258 2269 8294 2271
rect 8258 2240 8295 2269
rect 8428 2248 8468 2304
rect 7700 2231 7735 2232
rect 7677 2226 7735 2231
rect 7677 2206 7680 2226
rect 7700 2212 7735 2226
rect 7755 2212 7764 2232
rect 7700 2204 7764 2212
rect 7726 2203 7764 2204
rect 7727 2202 7764 2203
rect 7830 2236 7866 2237
rect 7938 2236 7974 2237
rect 7830 2228 7974 2236
rect 7830 2208 7838 2228
rect 7858 2208 7893 2228
rect 7913 2208 7946 2228
rect 7966 2208 7974 2228
rect 7830 2202 7974 2208
rect 8040 2232 8078 2240
rect 8156 2236 8192 2237
rect 8040 2212 8049 2232
rect 8069 2212 8078 2232
rect 8040 2203 8078 2212
rect 8107 2228 8192 2236
rect 8107 2208 8164 2228
rect 8184 2208 8192 2228
rect 8040 2202 8077 2203
rect 8107 2202 8192 2208
rect 8258 2232 8296 2240
rect 8258 2212 8267 2232
rect 8287 2212 8296 2232
rect 8428 2230 8440 2248
rect 8458 2230 8468 2248
rect 8873 2275 8925 2464
rect 9271 2439 9310 2464
rect 9954 2477 10103 2484
rect 9954 2457 10013 2477
rect 10033 2457 10072 2477
rect 10092 2457 10103 2477
rect 9954 2449 10103 2457
rect 10170 2480 10327 2487
rect 10170 2460 10290 2480
rect 10310 2460 10327 2480
rect 10170 2450 10327 2460
rect 10170 2449 10205 2450
rect 9055 2414 9242 2438
rect 9271 2419 9666 2439
rect 9686 2419 9689 2439
rect 10170 2428 10201 2449
rect 10388 2428 10424 2538
rect 10443 2537 10480 2538
rect 10539 2537 10576 2538
rect 10499 2478 10589 2484
rect 10499 2458 10508 2478
rect 10528 2476 10589 2478
rect 10528 2458 10553 2476
rect 10499 2456 10553 2458
rect 10573 2456 10589 2476
rect 10499 2450 10589 2456
rect 10013 2427 10050 2428
rect 9271 2414 9689 2419
rect 10012 2418 10050 2427
rect 9055 2343 9092 2414
rect 9271 2413 9614 2414
rect 9271 2410 9310 2413
rect 9576 2412 9613 2413
rect 9207 2353 9238 2354
rect 9055 2323 9064 2343
rect 9084 2323 9092 2343
rect 9055 2313 9092 2323
rect 9151 2343 9238 2353
rect 9151 2323 9160 2343
rect 9180 2323 9238 2343
rect 9151 2314 9238 2323
rect 9151 2313 9188 2314
rect 8873 2257 8889 2275
rect 8907 2257 8925 2275
rect 9207 2263 9238 2314
rect 9273 2343 9310 2410
rect 10012 2398 10021 2418
rect 10041 2398 10050 2418
rect 10012 2390 10050 2398
rect 10116 2422 10201 2428
rect 10231 2427 10268 2428
rect 10116 2402 10124 2422
rect 10144 2402 10201 2422
rect 10116 2394 10201 2402
rect 10230 2418 10268 2427
rect 10230 2398 10239 2418
rect 10259 2398 10268 2418
rect 10116 2393 10152 2394
rect 10230 2390 10268 2398
rect 10334 2426 10478 2428
rect 10334 2422 10394 2426
rect 10334 2402 10342 2422
rect 10362 2404 10394 2422
rect 10417 2422 10478 2426
rect 10417 2404 10450 2422
rect 10362 2402 10450 2404
rect 10470 2402 10478 2422
rect 10334 2394 10478 2402
rect 10334 2393 10370 2394
rect 10442 2393 10478 2394
rect 10544 2427 10581 2428
rect 10544 2426 10582 2427
rect 10544 2418 10608 2426
rect 10544 2398 10553 2418
rect 10573 2404 10608 2418
rect 10628 2404 10631 2424
rect 10573 2399 10631 2404
rect 10573 2398 10608 2399
rect 10013 2361 10050 2390
rect 10014 2359 10050 2361
rect 9425 2353 9461 2354
rect 9273 2323 9282 2343
rect 9302 2323 9310 2343
rect 9273 2313 9310 2323
rect 9369 2343 9517 2353
rect 9617 2350 9713 2352
rect 9369 2323 9378 2343
rect 9398 2323 9488 2343
rect 9508 2323 9517 2343
rect 9369 2314 9517 2323
rect 9575 2343 9713 2350
rect 9575 2323 9584 2343
rect 9604 2323 9713 2343
rect 10014 2337 10205 2359
rect 10231 2358 10268 2390
rect 10544 2386 10608 2398
rect 10231 2357 10506 2358
rect 10648 2357 10675 2538
rect 10231 2332 10675 2357
rect 10811 2363 10850 4178
rect 11152 4165 11185 4498
rect 11249 4530 11417 4531
rect 11543 4530 11583 4754
rect 12046 4758 12214 4759
rect 12455 4758 12490 4775
rect 12847 4765 12894 4776
rect 12046 4732 12490 4758
rect 12046 4730 12214 4732
rect 12410 4731 12490 4732
rect 12645 4731 12712 4757
rect 12851 4731 12894 4765
rect 12046 4552 12073 4730
rect 12113 4692 12177 4704
rect 12453 4700 12490 4731
rect 12671 4700 12708 4731
rect 12853 4706 12894 4731
rect 13285 4790 13326 4815
rect 13471 4790 13508 4821
rect 13689 4790 13726 4821
rect 14002 4817 14066 4829
rect 14106 4791 14133 4969
rect 13285 4756 13328 4790
rect 13467 4764 13534 4790
rect 13689 4789 13769 4790
rect 13965 4789 14133 4791
rect 13689 4763 14133 4789
rect 13285 4745 13332 4756
rect 13689 4746 13724 4763
rect 13965 4762 14133 4763
rect 14596 4767 14636 4991
rect 14762 4990 14930 4991
rect 14994 5023 15027 5356
rect 15329 5343 15368 7158
rect 15504 7164 15948 7189
rect 15504 6983 15531 7164
rect 15673 7163 15948 7164
rect 15571 7123 15635 7135
rect 15911 7131 15948 7163
rect 15974 7162 16165 7184
rect 16466 7178 16575 7198
rect 16595 7178 16604 7198
rect 16466 7171 16604 7178
rect 16662 7198 16810 7207
rect 16662 7178 16671 7198
rect 16691 7178 16781 7198
rect 16801 7178 16810 7198
rect 16466 7169 16562 7171
rect 16662 7168 16810 7178
rect 16869 7198 16906 7208
rect 16869 7178 16877 7198
rect 16897 7178 16906 7198
rect 16718 7167 16754 7168
rect 16129 7160 16165 7162
rect 16129 7131 16166 7160
rect 15571 7122 15606 7123
rect 15548 7117 15606 7122
rect 15548 7097 15551 7117
rect 15571 7103 15606 7117
rect 15626 7103 15635 7123
rect 15571 7095 15635 7103
rect 15597 7094 15635 7095
rect 15598 7093 15635 7094
rect 15701 7127 15737 7128
rect 15809 7127 15845 7128
rect 15701 7119 15845 7127
rect 15701 7099 15709 7119
rect 15729 7117 15817 7119
rect 15729 7099 15762 7117
rect 15701 7095 15762 7099
rect 15785 7099 15817 7117
rect 15837 7099 15845 7119
rect 15785 7095 15845 7099
rect 15701 7093 15845 7095
rect 15911 7123 15949 7131
rect 16027 7127 16063 7128
rect 15911 7103 15920 7123
rect 15940 7103 15949 7123
rect 15911 7094 15949 7103
rect 15978 7119 16063 7127
rect 15978 7099 16035 7119
rect 16055 7099 16063 7119
rect 15911 7093 15948 7094
rect 15978 7093 16063 7099
rect 16129 7123 16167 7131
rect 16129 7103 16138 7123
rect 16158 7103 16167 7123
rect 16869 7111 16906 7178
rect 16941 7207 16972 7258
rect 17254 7246 17272 7264
rect 17290 7246 17306 7264
rect 16991 7207 17028 7208
rect 16941 7198 17028 7207
rect 16941 7178 16999 7198
rect 17019 7178 17028 7198
rect 16941 7168 17028 7178
rect 17087 7198 17124 7208
rect 17087 7178 17095 7198
rect 17115 7178 17124 7198
rect 16941 7167 16972 7168
rect 16566 7108 16603 7109
rect 16869 7108 16908 7111
rect 16565 7107 16908 7108
rect 17087 7107 17124 7178
rect 16129 7094 16167 7103
rect 16490 7102 16908 7107
rect 16129 7093 16166 7094
rect 15590 7065 15680 7071
rect 15590 7045 15606 7065
rect 15626 7063 15680 7065
rect 15626 7045 15651 7063
rect 15590 7043 15651 7045
rect 15671 7043 15680 7063
rect 15590 7037 15680 7043
rect 15603 6983 15640 6984
rect 15699 6983 15736 6984
rect 15755 6983 15791 7093
rect 15978 7072 16009 7093
rect 16490 7082 16493 7102
rect 16513 7082 16908 7102
rect 16937 7083 17124 7107
rect 15974 7071 16009 7072
rect 15852 7061 16009 7071
rect 15852 7041 15869 7061
rect 15889 7041 16009 7061
rect 15852 7034 16009 7041
rect 16076 7064 16225 7072
rect 16076 7044 16087 7064
rect 16107 7044 16146 7064
rect 16166 7044 16225 7064
rect 16076 7037 16225 7044
rect 16869 7057 16908 7082
rect 17254 7057 17306 7246
rect 16869 7039 17308 7057
rect 16076 7036 16117 7037
rect 15810 6983 15847 6984
rect 15503 6974 15641 6983
rect 15503 6954 15612 6974
rect 15632 6954 15641 6974
rect 15503 6947 15641 6954
rect 15699 6974 15847 6983
rect 15699 6954 15708 6974
rect 15728 6954 15818 6974
rect 15838 6954 15847 6974
rect 15503 6945 15599 6947
rect 15699 6944 15847 6954
rect 15906 6974 15943 6984
rect 15906 6954 15914 6974
rect 15934 6954 15943 6974
rect 15755 6943 15791 6944
rect 15603 6884 15640 6885
rect 15906 6884 15943 6954
rect 15978 6983 16009 7034
rect 16869 7021 17269 7039
rect 17287 7021 17308 7039
rect 16869 7015 17308 7021
rect 16875 7011 17308 7015
rect 17254 7009 17306 7011
rect 16028 6983 16065 6984
rect 15978 6974 16065 6983
rect 15978 6954 16036 6974
rect 16056 6954 16065 6974
rect 15978 6944 16065 6954
rect 16124 6974 16161 6984
rect 16124 6954 16132 6974
rect 16152 6954 16161 6974
rect 15978 6943 16009 6944
rect 15602 6883 15943 6884
rect 16124 6883 16161 6954
rect 17257 6944 17294 6949
rect 15527 6878 15943 6883
rect 15527 6858 15530 6878
rect 15550 6858 15943 6878
rect 15974 6859 16161 6883
rect 17248 6940 17295 6944
rect 17248 6922 17267 6940
rect 17285 6922 17295 6940
rect 17248 6874 17295 6922
rect 16872 6871 17295 6874
rect 15747 6857 15812 6858
rect 16850 6841 17295 6871
rect 15943 6825 15983 6833
rect 15943 6803 15951 6825
rect 15975 6803 15983 6825
rect 15548 6574 15585 6580
rect 15548 6555 15556 6574
rect 15577 6555 15585 6574
rect 15548 6547 15585 6555
rect 15552 6214 15585 6547
rect 15649 6579 15817 6580
rect 15943 6579 15983 6803
rect 16446 6807 16614 6808
rect 16850 6807 16891 6841
rect 17248 6820 17295 6841
rect 16446 6797 16891 6807
rect 16963 6805 17106 6806
rect 16446 6781 16890 6797
rect 16446 6779 16614 6781
rect 16810 6780 16890 6781
rect 16963 6780 17108 6805
rect 17250 6780 17295 6820
rect 16446 6601 16473 6779
rect 16513 6741 16577 6753
rect 16853 6749 16890 6780
rect 17071 6749 17108 6780
rect 17253 6773 17295 6780
rect 16513 6740 16548 6741
rect 16490 6735 16548 6740
rect 16490 6715 16493 6735
rect 16513 6721 16548 6735
rect 16568 6721 16577 6741
rect 16513 6713 16577 6721
rect 16539 6712 16577 6713
rect 16540 6711 16577 6712
rect 16643 6745 16679 6746
rect 16751 6745 16787 6746
rect 16643 6737 16787 6745
rect 16643 6717 16651 6737
rect 16671 6733 16759 6737
rect 16671 6717 16715 6733
rect 16643 6713 16715 6717
rect 16735 6717 16759 6733
rect 16779 6717 16787 6737
rect 16735 6713 16787 6717
rect 16643 6711 16787 6713
rect 16853 6741 16891 6749
rect 16969 6745 17005 6746
rect 16853 6721 16862 6741
rect 16882 6721 16891 6741
rect 16853 6712 16891 6721
rect 16920 6737 17005 6745
rect 16920 6717 16977 6737
rect 16997 6717 17005 6737
rect 16853 6711 16890 6712
rect 16920 6711 17005 6717
rect 17071 6741 17109 6749
rect 17071 6721 17080 6741
rect 17100 6721 17109 6741
rect 17071 6712 17109 6721
rect 17253 6746 17296 6773
rect 17253 6728 17267 6746
rect 17285 6728 17296 6746
rect 17253 6720 17296 6728
rect 17258 6718 17296 6720
rect 17071 6711 17108 6712
rect 16532 6683 16622 6689
rect 16532 6663 16548 6683
rect 16568 6681 16622 6683
rect 16568 6663 16593 6681
rect 16532 6661 16593 6663
rect 16613 6661 16622 6681
rect 16532 6655 16622 6661
rect 16545 6601 16582 6602
rect 16641 6601 16678 6602
rect 16697 6601 16733 6711
rect 16920 6690 16951 6711
rect 16916 6689 16951 6690
rect 16794 6679 16951 6689
rect 16794 6659 16811 6679
rect 16831 6659 16951 6679
rect 16794 6652 16951 6659
rect 17018 6682 17167 6690
rect 17018 6662 17029 6682
rect 17049 6662 17088 6682
rect 17108 6662 17167 6682
rect 17018 6655 17167 6662
rect 17018 6654 17059 6655
rect 17255 6653 17292 6656
rect 16752 6601 16789 6602
rect 16445 6592 16583 6601
rect 15649 6553 16093 6579
rect 15649 6551 15817 6553
rect 15649 6373 15676 6551
rect 15716 6513 15780 6525
rect 16056 6521 16093 6553
rect 16119 6552 16310 6574
rect 16445 6572 16554 6592
rect 16574 6572 16583 6592
rect 16445 6565 16583 6572
rect 16641 6592 16789 6601
rect 16641 6572 16650 6592
rect 16670 6572 16760 6592
rect 16780 6572 16789 6592
rect 16445 6563 16541 6565
rect 16641 6562 16789 6572
rect 16848 6592 16885 6602
rect 16848 6572 16856 6592
rect 16876 6572 16885 6592
rect 16697 6561 16733 6562
rect 16274 6550 16310 6552
rect 16274 6521 16311 6550
rect 15716 6512 15751 6513
rect 15693 6507 15751 6512
rect 15693 6487 15696 6507
rect 15716 6493 15751 6507
rect 15771 6493 15780 6513
rect 15716 6487 15780 6493
rect 15693 6485 15780 6487
rect 15693 6481 15720 6485
rect 15742 6484 15780 6485
rect 15743 6483 15780 6484
rect 15846 6517 15882 6518
rect 15954 6517 15990 6518
rect 15846 6510 15990 6517
rect 15846 6509 15908 6510
rect 15846 6489 15854 6509
rect 15874 6492 15908 6509
rect 15927 6509 15990 6510
rect 15927 6492 15962 6509
rect 15874 6489 15962 6492
rect 15982 6489 15990 6509
rect 15846 6483 15990 6489
rect 16056 6513 16094 6521
rect 16172 6517 16208 6518
rect 16056 6493 16065 6513
rect 16085 6493 16094 6513
rect 16056 6484 16094 6493
rect 16123 6509 16208 6517
rect 16123 6489 16180 6509
rect 16200 6489 16208 6509
rect 16056 6483 16093 6484
rect 16123 6483 16208 6489
rect 16274 6513 16312 6521
rect 16274 6493 16283 6513
rect 16303 6493 16312 6513
rect 16545 6502 16582 6503
rect 16848 6502 16885 6572
rect 16920 6601 16951 6652
rect 17247 6647 17292 6653
rect 17247 6629 17265 6647
rect 17283 6629 17292 6647
rect 17247 6619 17292 6629
rect 16970 6601 17007 6602
rect 16920 6592 17007 6601
rect 16920 6572 16978 6592
rect 16998 6572 17007 6592
rect 16920 6562 17007 6572
rect 17066 6592 17103 6602
rect 17066 6572 17074 6592
rect 17094 6572 17103 6592
rect 17247 6577 17290 6619
rect 17153 6575 17290 6577
rect 16920 6561 16951 6562
rect 17066 6502 17103 6572
rect 16544 6501 16885 6502
rect 16274 6484 16312 6493
rect 16469 6496 16885 6501
rect 16274 6483 16311 6484
rect 15735 6455 15825 6461
rect 15735 6435 15751 6455
rect 15771 6453 15825 6455
rect 15771 6435 15796 6453
rect 15735 6433 15796 6435
rect 15816 6433 15825 6453
rect 15735 6427 15825 6433
rect 15748 6373 15785 6374
rect 15844 6373 15881 6374
rect 15900 6373 15936 6483
rect 16123 6462 16154 6483
rect 16469 6476 16472 6496
rect 16492 6476 16885 6496
rect 17069 6486 17103 6502
rect 17147 6554 17290 6575
rect 16845 6467 16885 6476
rect 17147 6467 17174 6554
rect 17247 6528 17290 6554
rect 17247 6510 17260 6528
rect 17278 6510 17290 6528
rect 17247 6499 17290 6510
rect 16119 6461 16154 6462
rect 15997 6451 16154 6461
rect 15997 6431 16014 6451
rect 16034 6431 16154 6451
rect 15997 6424 16154 6431
rect 16221 6454 16367 6462
rect 16221 6434 16232 6454
rect 16252 6434 16291 6454
rect 16311 6434 16367 6454
rect 16845 6450 17174 6467
rect 16845 6449 16885 6450
rect 16221 6427 16367 6434
rect 17242 6438 17282 6441
rect 17242 6432 17285 6438
rect 16867 6429 17285 6432
rect 16221 6426 16262 6427
rect 15955 6373 15992 6374
rect 15648 6364 15786 6373
rect 15648 6344 15757 6364
rect 15777 6344 15786 6364
rect 15648 6337 15786 6344
rect 15844 6364 15992 6373
rect 15844 6344 15853 6364
rect 15873 6344 15963 6364
rect 15983 6344 15992 6364
rect 15648 6335 15744 6337
rect 15844 6334 15992 6344
rect 16051 6364 16088 6374
rect 16051 6344 16059 6364
rect 16079 6344 16088 6364
rect 15900 6333 15936 6334
rect 15748 6274 15785 6275
rect 16051 6274 16088 6344
rect 16123 6373 16154 6424
rect 16867 6411 17258 6429
rect 17276 6411 17285 6429
rect 16867 6409 17285 6411
rect 16867 6401 16894 6409
rect 17135 6406 17285 6409
rect 16447 6395 16615 6396
rect 16866 6395 16894 6401
rect 16447 6379 16894 6395
rect 17242 6401 17285 6406
rect 16173 6373 16210 6374
rect 16123 6364 16210 6373
rect 16123 6344 16181 6364
rect 16201 6344 16210 6364
rect 16123 6334 16210 6344
rect 16269 6364 16306 6374
rect 16269 6344 16277 6364
rect 16297 6344 16306 6364
rect 16123 6333 16154 6334
rect 15747 6273 16088 6274
rect 16269 6273 16306 6344
rect 15672 6268 16088 6273
rect 15672 6248 15675 6268
rect 15695 6248 16088 6268
rect 16119 6249 16306 6273
rect 16447 6369 16891 6379
rect 16447 6367 16615 6369
rect 15547 6169 15589 6214
rect 16447 6189 16474 6367
rect 16514 6329 16578 6341
rect 16854 6337 16891 6369
rect 16917 6368 17108 6390
rect 17072 6366 17108 6368
rect 17072 6337 17109 6366
rect 17242 6345 17282 6401
rect 16514 6328 16549 6329
rect 16491 6323 16549 6328
rect 16491 6303 16494 6323
rect 16514 6309 16549 6323
rect 16569 6309 16578 6329
rect 16514 6301 16578 6309
rect 16540 6300 16578 6301
rect 16541 6299 16578 6300
rect 16644 6333 16680 6334
rect 16752 6333 16788 6334
rect 16644 6325 16788 6333
rect 16644 6305 16652 6325
rect 16672 6305 16707 6325
rect 16727 6305 16760 6325
rect 16780 6305 16788 6325
rect 16644 6299 16788 6305
rect 16854 6329 16892 6337
rect 16970 6333 17006 6334
rect 16854 6309 16863 6329
rect 16883 6309 16892 6329
rect 16854 6300 16892 6309
rect 16921 6325 17006 6333
rect 16921 6305 16978 6325
rect 16998 6305 17006 6325
rect 16854 6299 16891 6300
rect 16921 6299 17006 6305
rect 17072 6329 17110 6337
rect 17072 6309 17081 6329
rect 17101 6309 17110 6329
rect 17242 6327 17254 6345
rect 17272 6327 17282 6345
rect 17242 6317 17282 6327
rect 17072 6300 17110 6309
rect 17072 6299 17109 6300
rect 16533 6271 16623 6277
rect 16533 6251 16549 6271
rect 16569 6269 16623 6271
rect 16569 6251 16594 6269
rect 16533 6249 16594 6251
rect 16614 6249 16623 6269
rect 16533 6243 16623 6249
rect 16546 6189 16583 6190
rect 16642 6189 16679 6190
rect 16698 6189 16734 6299
rect 16921 6278 16952 6299
rect 16917 6277 16952 6278
rect 16795 6267 16952 6277
rect 16795 6247 16812 6267
rect 16832 6247 16952 6267
rect 16795 6240 16952 6247
rect 17019 6270 17168 6278
rect 17019 6250 17030 6270
rect 17050 6250 17089 6270
rect 17109 6250 17168 6270
rect 17019 6243 17168 6250
rect 17234 6246 17286 6264
rect 17019 6242 17060 6243
rect 16753 6189 16790 6190
rect 16446 6180 16584 6189
rect 15918 6169 15951 6171
rect 15547 6157 15994 6169
rect 15550 6143 15994 6157
rect 15550 6141 15718 6143
rect 15550 5963 15577 6141
rect 15617 6103 15681 6115
rect 15957 6111 15994 6143
rect 16020 6142 16211 6164
rect 16446 6160 16555 6180
rect 16575 6160 16584 6180
rect 16446 6153 16584 6160
rect 16642 6180 16790 6189
rect 16642 6160 16651 6180
rect 16671 6160 16761 6180
rect 16781 6160 16790 6180
rect 16446 6151 16542 6153
rect 16642 6150 16790 6160
rect 16849 6180 16886 6190
rect 16849 6160 16857 6180
rect 16877 6160 16886 6180
rect 16698 6149 16734 6150
rect 16175 6140 16211 6142
rect 16175 6111 16212 6140
rect 15617 6102 15652 6103
rect 15594 6097 15652 6102
rect 15594 6077 15597 6097
rect 15617 6083 15652 6097
rect 15672 6083 15681 6103
rect 15617 6075 15681 6083
rect 15643 6074 15681 6075
rect 15644 6073 15681 6074
rect 15747 6107 15783 6108
rect 15855 6107 15891 6108
rect 15747 6099 15891 6107
rect 15747 6079 15755 6099
rect 15775 6097 15863 6099
rect 15775 6079 15808 6097
rect 15747 6078 15808 6079
rect 15829 6079 15863 6097
rect 15883 6079 15891 6099
rect 15829 6078 15891 6079
rect 15747 6073 15891 6078
rect 15957 6103 15995 6111
rect 16073 6107 16109 6108
rect 15957 6083 15966 6103
rect 15986 6083 15995 6103
rect 15957 6074 15995 6083
rect 16024 6099 16109 6107
rect 16024 6079 16081 6099
rect 16101 6079 16109 6099
rect 15957 6073 15994 6074
rect 16024 6073 16109 6079
rect 16175 6103 16213 6111
rect 16175 6083 16184 6103
rect 16204 6083 16213 6103
rect 16849 6093 16886 6160
rect 16921 6189 16952 6240
rect 17234 6228 17252 6246
rect 17270 6228 17286 6246
rect 16971 6189 17008 6190
rect 16921 6180 17008 6189
rect 16921 6160 16979 6180
rect 16999 6160 17008 6180
rect 16921 6150 17008 6160
rect 17067 6180 17104 6190
rect 17067 6160 17075 6180
rect 17095 6160 17104 6180
rect 16921 6149 16952 6150
rect 16546 6090 16583 6091
rect 16849 6090 16888 6093
rect 16545 6089 16888 6090
rect 17067 6089 17104 6160
rect 16175 6074 16213 6083
rect 16470 6084 16888 6089
rect 16175 6073 16212 6074
rect 15636 6045 15726 6051
rect 15636 6025 15652 6045
rect 15672 6043 15726 6045
rect 15672 6025 15697 6043
rect 15636 6023 15697 6025
rect 15717 6023 15726 6043
rect 15636 6017 15726 6023
rect 15649 5963 15686 5964
rect 15745 5963 15782 5964
rect 15801 5963 15837 6073
rect 16024 6052 16055 6073
rect 16470 6064 16473 6084
rect 16493 6064 16888 6084
rect 16917 6065 17104 6089
rect 16020 6051 16055 6052
rect 15898 6041 16055 6051
rect 15898 6021 15915 6041
rect 15935 6021 16055 6041
rect 15898 6014 16055 6021
rect 16122 6044 16271 6052
rect 16122 6024 16133 6044
rect 16153 6024 16192 6044
rect 16212 6024 16271 6044
rect 16122 6017 16271 6024
rect 16849 6039 16888 6064
rect 17234 6039 17286 6228
rect 16849 6021 17288 6039
rect 16122 6016 16163 6017
rect 15856 5963 15893 5964
rect 15549 5954 15687 5963
rect 15549 5934 15658 5954
rect 15678 5934 15687 5954
rect 15549 5927 15687 5934
rect 15745 5954 15893 5963
rect 15745 5934 15754 5954
rect 15774 5934 15864 5954
rect 15884 5934 15893 5954
rect 15549 5925 15645 5927
rect 15745 5924 15893 5934
rect 15952 5954 15989 5964
rect 15952 5934 15960 5954
rect 15980 5934 15989 5954
rect 15801 5923 15837 5924
rect 15649 5864 15686 5865
rect 15952 5864 15989 5934
rect 16024 5963 16055 6014
rect 16849 6003 17249 6021
rect 17267 6003 17288 6021
rect 16849 5997 17288 6003
rect 16855 5993 17288 5997
rect 17234 5991 17286 5993
rect 16074 5963 16111 5964
rect 16024 5954 16111 5963
rect 16024 5934 16082 5954
rect 16102 5934 16111 5954
rect 16024 5924 16111 5934
rect 16170 5954 16207 5964
rect 16170 5934 16178 5954
rect 16198 5934 16207 5954
rect 16024 5923 16055 5924
rect 15648 5863 15989 5864
rect 16170 5863 16207 5934
rect 17237 5926 17274 5931
rect 17228 5922 17275 5926
rect 17228 5904 17247 5922
rect 17265 5904 17275 5922
rect 15573 5858 15989 5863
rect 15573 5838 15576 5858
rect 15596 5838 15989 5858
rect 16020 5839 16207 5863
rect 16832 5861 16872 5866
rect 17228 5861 17275 5904
rect 16832 5822 17275 5861
rect 15926 5807 15966 5815
rect 15926 5785 15934 5807
rect 15958 5785 15966 5807
rect 15632 5561 15800 5562
rect 15926 5561 15966 5785
rect 16429 5789 16597 5790
rect 16832 5789 16872 5822
rect 17228 5789 17275 5822
rect 16429 5788 16873 5789
rect 16429 5763 16874 5788
rect 16429 5761 16597 5763
rect 16793 5762 16874 5763
rect 17043 5762 17092 5788
rect 17228 5762 17277 5789
rect 16429 5583 16456 5761
rect 16496 5723 16560 5735
rect 16836 5731 16873 5762
rect 17054 5731 17091 5762
rect 17236 5737 17277 5762
rect 16496 5722 16531 5723
rect 16473 5717 16531 5722
rect 16473 5697 16476 5717
rect 16496 5703 16531 5717
rect 16551 5703 16560 5723
rect 16496 5695 16560 5703
rect 16522 5694 16560 5695
rect 16523 5693 16560 5694
rect 16626 5727 16662 5728
rect 16734 5727 16770 5728
rect 16626 5719 16770 5727
rect 16626 5699 16634 5719
rect 16654 5715 16742 5719
rect 16654 5699 16698 5715
rect 16626 5695 16698 5699
rect 16718 5699 16742 5715
rect 16762 5699 16770 5719
rect 16718 5695 16770 5699
rect 16626 5693 16770 5695
rect 16836 5723 16874 5731
rect 16952 5727 16988 5728
rect 16836 5703 16845 5723
rect 16865 5703 16874 5723
rect 16836 5694 16874 5703
rect 16903 5719 16988 5727
rect 16903 5699 16960 5719
rect 16980 5699 16988 5719
rect 16836 5693 16873 5694
rect 16903 5693 16988 5699
rect 17054 5723 17092 5731
rect 17054 5703 17063 5723
rect 17083 5703 17092 5723
rect 17054 5694 17092 5703
rect 17236 5728 17278 5737
rect 17236 5710 17250 5728
rect 17268 5710 17278 5728
rect 17236 5702 17278 5710
rect 17241 5700 17278 5702
rect 17054 5693 17091 5694
rect 16515 5665 16605 5671
rect 16515 5645 16531 5665
rect 16551 5663 16605 5665
rect 16551 5645 16576 5663
rect 16515 5643 16576 5645
rect 16596 5643 16605 5663
rect 16515 5637 16605 5643
rect 16528 5583 16565 5584
rect 16624 5583 16661 5584
rect 16680 5583 16716 5693
rect 16903 5672 16934 5693
rect 16899 5671 16934 5672
rect 16777 5661 16934 5671
rect 16777 5641 16794 5661
rect 16814 5641 16934 5661
rect 16777 5634 16934 5641
rect 17001 5664 17150 5672
rect 17001 5644 17012 5664
rect 17032 5644 17071 5664
rect 17091 5644 17150 5664
rect 17001 5637 17150 5644
rect 17001 5636 17042 5637
rect 17238 5635 17275 5638
rect 16735 5583 16772 5584
rect 16428 5574 16566 5583
rect 15632 5535 16076 5561
rect 15632 5533 15800 5535
rect 15632 5355 15659 5533
rect 15699 5495 15763 5507
rect 16039 5503 16076 5535
rect 16102 5534 16293 5556
rect 16428 5554 16537 5574
rect 16557 5554 16566 5574
rect 16428 5547 16566 5554
rect 16624 5574 16772 5583
rect 16624 5554 16633 5574
rect 16653 5554 16743 5574
rect 16763 5554 16772 5574
rect 16428 5545 16524 5547
rect 16624 5544 16772 5554
rect 16831 5574 16868 5584
rect 16831 5554 16839 5574
rect 16859 5554 16868 5574
rect 16680 5543 16716 5544
rect 16257 5532 16293 5534
rect 16257 5503 16294 5532
rect 15699 5494 15734 5495
rect 15676 5489 15734 5494
rect 15676 5469 15679 5489
rect 15699 5475 15734 5489
rect 15754 5475 15763 5495
rect 15699 5467 15763 5475
rect 15725 5466 15763 5467
rect 15726 5465 15763 5466
rect 15829 5499 15865 5500
rect 15937 5499 15973 5500
rect 15829 5491 15973 5499
rect 15829 5471 15837 5491
rect 15857 5490 15945 5491
rect 15857 5471 15892 5490
rect 15913 5471 15945 5490
rect 15965 5471 15973 5491
rect 15829 5465 15973 5471
rect 16039 5495 16077 5503
rect 16155 5499 16191 5500
rect 16039 5475 16048 5495
rect 16068 5475 16077 5495
rect 16039 5466 16077 5475
rect 16106 5491 16191 5499
rect 16106 5471 16163 5491
rect 16183 5471 16191 5491
rect 16039 5465 16076 5466
rect 16106 5465 16191 5471
rect 16257 5495 16295 5503
rect 16257 5475 16266 5495
rect 16286 5475 16295 5495
rect 16528 5484 16565 5485
rect 16831 5484 16868 5554
rect 16903 5583 16934 5634
rect 17230 5629 17275 5635
rect 17230 5611 17248 5629
rect 17266 5611 17275 5629
rect 17230 5601 17275 5611
rect 16953 5583 16990 5584
rect 16903 5574 16990 5583
rect 16903 5554 16961 5574
rect 16981 5554 16990 5574
rect 16903 5544 16990 5554
rect 17049 5574 17086 5584
rect 17049 5554 17057 5574
rect 17077 5554 17086 5574
rect 17230 5559 17273 5601
rect 17136 5557 17273 5559
rect 16903 5543 16934 5544
rect 17049 5484 17086 5554
rect 16527 5483 16868 5484
rect 16257 5466 16295 5475
rect 16452 5478 16868 5483
rect 16257 5465 16294 5466
rect 15718 5437 15808 5443
rect 15718 5417 15734 5437
rect 15754 5435 15808 5437
rect 15754 5417 15779 5435
rect 15718 5415 15779 5417
rect 15799 5415 15808 5435
rect 15718 5409 15808 5415
rect 15731 5355 15768 5356
rect 15827 5355 15864 5356
rect 15883 5355 15919 5465
rect 16106 5444 16137 5465
rect 16452 5458 16455 5478
rect 16475 5458 16868 5478
rect 17052 5468 17086 5484
rect 17130 5536 17273 5557
rect 16828 5449 16868 5458
rect 17130 5449 17157 5536
rect 17230 5510 17273 5536
rect 17230 5492 17243 5510
rect 17261 5492 17273 5510
rect 17230 5481 17273 5492
rect 16102 5443 16137 5444
rect 15980 5433 16137 5443
rect 15980 5413 15997 5433
rect 16017 5413 16137 5433
rect 15980 5406 16137 5413
rect 16204 5436 16353 5444
rect 16204 5416 16215 5436
rect 16235 5416 16274 5436
rect 16294 5416 16353 5436
rect 16828 5432 17157 5449
rect 16828 5431 16868 5432
rect 16204 5409 16353 5416
rect 17225 5420 17265 5423
rect 17225 5414 17268 5420
rect 16850 5411 17268 5414
rect 16204 5408 16245 5409
rect 15938 5355 15975 5356
rect 15631 5346 15769 5355
rect 15329 5171 15369 5343
rect 15631 5326 15740 5346
rect 15760 5326 15769 5346
rect 15631 5319 15769 5326
rect 15827 5346 15975 5355
rect 15827 5326 15836 5346
rect 15856 5326 15946 5346
rect 15966 5326 15975 5346
rect 15631 5317 15727 5319
rect 15827 5316 15975 5326
rect 16034 5346 16071 5356
rect 16034 5326 16042 5346
rect 16062 5326 16071 5346
rect 15883 5315 15919 5316
rect 15731 5256 15768 5257
rect 16034 5256 16071 5326
rect 16106 5355 16137 5406
rect 16850 5393 17241 5411
rect 17259 5393 17268 5411
rect 16850 5391 17268 5393
rect 16850 5383 16877 5391
rect 17118 5388 17268 5391
rect 16430 5377 16598 5378
rect 16849 5377 16877 5383
rect 16430 5361 16877 5377
rect 17225 5383 17268 5388
rect 16156 5355 16193 5356
rect 16106 5346 16193 5355
rect 16106 5326 16164 5346
rect 16184 5326 16193 5346
rect 16106 5316 16193 5326
rect 16252 5346 16289 5356
rect 16252 5326 16260 5346
rect 16280 5326 16289 5346
rect 16106 5315 16137 5316
rect 15730 5255 16071 5256
rect 16252 5255 16289 5326
rect 15655 5250 16071 5255
rect 15655 5230 15658 5250
rect 15678 5230 16071 5250
rect 16102 5231 16289 5255
rect 16430 5351 16874 5361
rect 16430 5349 16598 5351
rect 16430 5171 16457 5349
rect 16497 5311 16561 5323
rect 16837 5319 16874 5351
rect 16900 5350 17091 5372
rect 17055 5348 17091 5350
rect 17055 5319 17092 5348
rect 17225 5327 17265 5383
rect 16497 5310 16532 5311
rect 16474 5305 16532 5310
rect 16474 5285 16477 5305
rect 16497 5291 16532 5305
rect 16552 5291 16561 5311
rect 16497 5283 16561 5291
rect 16523 5282 16561 5283
rect 16524 5281 16561 5282
rect 16627 5315 16663 5316
rect 16735 5315 16771 5316
rect 16627 5307 16771 5315
rect 16627 5287 16635 5307
rect 16655 5287 16690 5307
rect 16710 5287 16743 5307
rect 16763 5287 16771 5307
rect 16627 5281 16771 5287
rect 16837 5311 16875 5319
rect 16953 5315 16989 5316
rect 16837 5291 16846 5311
rect 16866 5291 16875 5311
rect 16837 5282 16875 5291
rect 16904 5307 16989 5315
rect 16904 5287 16961 5307
rect 16981 5287 16989 5307
rect 16837 5281 16874 5282
rect 16904 5281 16989 5287
rect 17055 5311 17093 5319
rect 17055 5291 17064 5311
rect 17084 5291 17093 5311
rect 17225 5309 17237 5327
rect 17255 5309 17265 5327
rect 17225 5299 17265 5309
rect 17055 5282 17093 5291
rect 17055 5281 17092 5282
rect 16516 5253 16606 5259
rect 16516 5233 16532 5253
rect 16552 5251 16606 5253
rect 16552 5233 16577 5251
rect 16516 5231 16577 5233
rect 16597 5231 16606 5251
rect 16516 5225 16606 5231
rect 16529 5171 16566 5172
rect 16625 5171 16662 5172
rect 16681 5171 16717 5281
rect 16904 5260 16935 5281
rect 16900 5259 16935 5260
rect 16778 5249 16935 5259
rect 16778 5229 16795 5249
rect 16815 5229 16935 5249
rect 16778 5222 16935 5229
rect 17002 5252 17151 5260
rect 17002 5232 17013 5252
rect 17033 5232 17072 5252
rect 17092 5232 17151 5252
rect 17002 5225 17151 5232
rect 17217 5228 17269 5246
rect 17002 5224 17043 5225
rect 16736 5171 16773 5172
rect 15330 5156 15369 5171
rect 16429 5162 16567 5171
rect 15330 5155 15496 5156
rect 15622 5155 15662 5157
rect 15330 5129 15772 5155
rect 15330 5127 15496 5129
rect 14994 5015 15031 5023
rect 14994 4996 15002 5015
rect 15023 4996 15031 5015
rect 14994 4990 15031 4996
rect 15330 4949 15355 5127
rect 15395 5089 15459 5101
rect 15735 5097 15772 5129
rect 15798 5128 15989 5150
rect 16429 5142 16538 5162
rect 16558 5142 16567 5162
rect 16429 5135 16567 5142
rect 16625 5162 16773 5171
rect 16625 5142 16634 5162
rect 16654 5142 16744 5162
rect 16764 5142 16773 5162
rect 16429 5133 16525 5135
rect 16625 5132 16773 5142
rect 16832 5162 16869 5172
rect 16832 5142 16840 5162
rect 16860 5142 16869 5162
rect 16681 5131 16717 5132
rect 15953 5126 15989 5128
rect 15953 5097 15990 5126
rect 15395 5088 15430 5089
rect 15372 5083 15430 5088
rect 15372 5063 15375 5083
rect 15395 5069 15430 5083
rect 15450 5069 15459 5089
rect 15395 5061 15459 5069
rect 15421 5060 15459 5061
rect 15422 5059 15459 5060
rect 15525 5093 15561 5094
rect 15633 5093 15669 5094
rect 15525 5088 15669 5093
rect 15525 5085 15587 5088
rect 15525 5065 15533 5085
rect 15553 5065 15587 5085
rect 15525 5062 15587 5065
rect 15613 5085 15669 5088
rect 15613 5065 15641 5085
rect 15661 5065 15669 5085
rect 15613 5062 15669 5065
rect 15525 5059 15669 5062
rect 15735 5089 15773 5097
rect 15851 5093 15887 5094
rect 15735 5069 15744 5089
rect 15764 5069 15773 5089
rect 15735 5060 15773 5069
rect 15802 5085 15887 5093
rect 15802 5065 15859 5085
rect 15879 5065 15887 5085
rect 15735 5059 15772 5060
rect 15802 5059 15887 5065
rect 15953 5089 15991 5097
rect 15953 5069 15962 5089
rect 15982 5069 15991 5089
rect 16832 5075 16869 5142
rect 16904 5171 16935 5222
rect 17217 5210 17235 5228
rect 17253 5210 17269 5228
rect 16954 5171 16991 5172
rect 16904 5162 16991 5171
rect 16904 5142 16962 5162
rect 16982 5142 16991 5162
rect 16904 5132 16991 5142
rect 17050 5162 17087 5172
rect 17050 5142 17058 5162
rect 17078 5142 17087 5162
rect 16904 5131 16935 5132
rect 16529 5072 16566 5073
rect 16832 5072 16871 5075
rect 16528 5071 16871 5072
rect 17050 5071 17087 5142
rect 15953 5060 15991 5069
rect 16453 5066 16871 5071
rect 15953 5059 15990 5060
rect 15414 5031 15504 5037
rect 15414 5011 15430 5031
rect 15450 5029 15504 5031
rect 15450 5011 15475 5029
rect 15414 5009 15475 5011
rect 15495 5009 15504 5029
rect 15414 5003 15504 5009
rect 15427 4949 15464 4950
rect 15523 4949 15560 4950
rect 15579 4949 15615 5059
rect 15802 5038 15833 5059
rect 16453 5046 16456 5066
rect 16476 5046 16871 5066
rect 16900 5047 17087 5071
rect 15798 5037 15833 5038
rect 15676 5027 15833 5037
rect 15676 5007 15693 5027
rect 15713 5007 15833 5027
rect 15676 5000 15833 5007
rect 15900 5030 16049 5038
rect 15900 5010 15911 5030
rect 15931 5010 15970 5030
rect 15990 5010 16049 5030
rect 15900 5003 16049 5010
rect 16832 5021 16871 5046
rect 17217 5021 17269 5210
rect 16832 5003 17271 5021
rect 15900 5002 15941 5003
rect 15634 4949 15671 4950
rect 15330 4940 15465 4949
rect 15330 4920 15436 4940
rect 15456 4920 15465 4940
rect 15330 4913 15465 4920
rect 15523 4940 15671 4949
rect 15523 4920 15532 4940
rect 15552 4920 15642 4940
rect 15662 4920 15671 4940
rect 15330 4911 15423 4913
rect 15523 4910 15671 4920
rect 15730 4940 15767 4950
rect 15730 4920 15738 4940
rect 15758 4920 15767 4940
rect 15579 4909 15615 4910
rect 15427 4850 15464 4851
rect 15730 4850 15767 4920
rect 15802 4949 15833 5000
rect 16832 4985 17232 5003
rect 17250 4985 17271 5003
rect 16832 4979 17271 4985
rect 16838 4975 17271 4979
rect 17217 4973 17269 4975
rect 15852 4949 15889 4950
rect 15802 4940 15889 4949
rect 15802 4920 15860 4940
rect 15880 4920 15889 4940
rect 15802 4910 15889 4920
rect 15948 4940 15985 4950
rect 15948 4920 15956 4940
rect 15976 4920 15985 4940
rect 15802 4909 15833 4910
rect 15426 4849 15767 4850
rect 15948 4849 15985 4920
rect 17220 4908 17257 4913
rect 15351 4844 15767 4849
rect 15351 4824 15354 4844
rect 15374 4824 15767 4844
rect 15798 4825 15985 4849
rect 17211 4904 17258 4908
rect 17211 4886 17230 4904
rect 17248 4886 17258 4904
rect 16819 4827 16857 4828
rect 17211 4827 17258 4886
rect 15571 4823 15636 4824
rect 13686 4745 13724 4746
rect 13285 4707 13724 4745
rect 14596 4745 14604 4767
rect 14628 4745 14636 4767
rect 14596 4737 14636 4745
rect 15907 4789 15947 4797
rect 15907 4767 15915 4789
rect 15939 4767 15947 4789
rect 16819 4789 17258 4827
rect 16819 4788 16857 4789
rect 14907 4710 14972 4711
rect 12113 4691 12148 4692
rect 12090 4686 12148 4691
rect 12090 4666 12093 4686
rect 12113 4672 12148 4686
rect 12168 4672 12177 4692
rect 12113 4664 12177 4672
rect 12139 4663 12177 4664
rect 12140 4662 12177 4663
rect 12243 4696 12279 4697
rect 12351 4696 12387 4697
rect 12243 4688 12387 4696
rect 12243 4668 12251 4688
rect 12271 4684 12359 4688
rect 12271 4668 12315 4684
rect 12243 4664 12315 4668
rect 12335 4668 12359 4684
rect 12379 4668 12387 4688
rect 12335 4664 12387 4668
rect 12243 4662 12387 4664
rect 12453 4692 12491 4700
rect 12569 4696 12605 4697
rect 12453 4672 12462 4692
rect 12482 4672 12491 4692
rect 12453 4663 12491 4672
rect 12520 4688 12605 4696
rect 12520 4668 12577 4688
rect 12597 4668 12605 4688
rect 12453 4662 12490 4663
rect 12520 4662 12605 4668
rect 12671 4692 12709 4700
rect 12671 4672 12680 4692
rect 12700 4672 12709 4692
rect 12671 4663 12709 4672
rect 12853 4697 12895 4706
rect 12853 4679 12867 4697
rect 12885 4679 12895 4697
rect 12853 4671 12895 4679
rect 12858 4669 12895 4671
rect 12671 4662 12708 4663
rect 12132 4634 12222 4640
rect 12132 4614 12148 4634
rect 12168 4632 12222 4634
rect 12168 4614 12193 4632
rect 12132 4612 12193 4614
rect 12213 4612 12222 4632
rect 12132 4606 12222 4612
rect 12145 4552 12182 4553
rect 12241 4552 12278 4553
rect 12297 4552 12333 4662
rect 12520 4641 12551 4662
rect 13285 4648 13332 4707
rect 13686 4706 13724 4707
rect 12516 4640 12551 4641
rect 12394 4630 12551 4640
rect 12394 4610 12411 4630
rect 12431 4610 12551 4630
rect 12394 4603 12551 4610
rect 12618 4633 12767 4641
rect 12618 4613 12629 4633
rect 12649 4613 12688 4633
rect 12708 4613 12767 4633
rect 13285 4630 13295 4648
rect 13313 4630 13332 4648
rect 13285 4626 13332 4630
rect 14558 4685 14745 4709
rect 14776 4690 15169 4710
rect 15189 4690 15192 4710
rect 14776 4685 15192 4690
rect 13286 4621 13323 4626
rect 12618 4606 12767 4613
rect 14558 4614 14595 4685
rect 14776 4684 15117 4685
rect 14710 4624 14741 4625
rect 12618 4605 12659 4606
rect 12855 4604 12892 4607
rect 12352 4552 12389 4553
rect 12045 4543 12183 4552
rect 11249 4504 11693 4530
rect 11249 4502 11417 4504
rect 11249 4324 11276 4502
rect 11316 4464 11380 4476
rect 11656 4472 11693 4504
rect 11719 4503 11910 4525
rect 12045 4523 12154 4543
rect 12174 4523 12183 4543
rect 12045 4516 12183 4523
rect 12241 4543 12389 4552
rect 12241 4523 12250 4543
rect 12270 4523 12360 4543
rect 12380 4523 12389 4543
rect 12045 4514 12141 4516
rect 12241 4513 12389 4523
rect 12448 4543 12485 4553
rect 12448 4523 12456 4543
rect 12476 4523 12485 4543
rect 12297 4512 12333 4513
rect 11874 4501 11910 4503
rect 11874 4472 11911 4501
rect 11316 4463 11351 4464
rect 11293 4458 11351 4463
rect 11293 4438 11296 4458
rect 11316 4444 11351 4458
rect 11371 4444 11380 4464
rect 11316 4438 11380 4444
rect 11293 4436 11380 4438
rect 11293 4432 11320 4436
rect 11342 4435 11380 4436
rect 11343 4434 11380 4435
rect 11446 4468 11482 4469
rect 11554 4468 11590 4469
rect 11446 4461 11590 4468
rect 11446 4460 11508 4461
rect 11446 4440 11454 4460
rect 11474 4443 11508 4460
rect 11527 4460 11590 4461
rect 11527 4443 11562 4460
rect 11474 4440 11562 4443
rect 11582 4440 11590 4460
rect 11446 4434 11590 4440
rect 11656 4464 11694 4472
rect 11772 4468 11808 4469
rect 11656 4444 11665 4464
rect 11685 4444 11694 4464
rect 11656 4435 11694 4444
rect 11723 4460 11808 4468
rect 11723 4440 11780 4460
rect 11800 4440 11808 4460
rect 11656 4434 11693 4435
rect 11723 4434 11808 4440
rect 11874 4464 11912 4472
rect 11874 4444 11883 4464
rect 11903 4444 11912 4464
rect 12145 4453 12182 4454
rect 12448 4453 12485 4523
rect 12520 4552 12551 4603
rect 12847 4598 12892 4604
rect 12847 4580 12865 4598
rect 12883 4580 12892 4598
rect 14558 4594 14567 4614
rect 14587 4594 14595 4614
rect 14558 4584 14595 4594
rect 14654 4614 14741 4624
rect 14654 4594 14663 4614
rect 14683 4594 14741 4614
rect 14654 4585 14741 4594
rect 14654 4584 14691 4585
rect 12847 4570 12892 4580
rect 12570 4552 12607 4553
rect 12520 4543 12607 4552
rect 12520 4523 12578 4543
rect 12598 4523 12607 4543
rect 12520 4513 12607 4523
rect 12666 4543 12703 4553
rect 12666 4523 12674 4543
rect 12694 4523 12703 4543
rect 12847 4528 12890 4570
rect 13274 4559 13326 4561
rect 12753 4526 12890 4528
rect 12520 4512 12551 4513
rect 12666 4453 12703 4523
rect 12144 4452 12485 4453
rect 11874 4435 11912 4444
rect 12069 4447 12485 4452
rect 11874 4434 11911 4435
rect 11335 4406 11425 4412
rect 11335 4386 11351 4406
rect 11371 4404 11425 4406
rect 11371 4386 11396 4404
rect 11335 4384 11396 4386
rect 11416 4384 11425 4404
rect 11335 4378 11425 4384
rect 11348 4324 11385 4325
rect 11444 4324 11481 4325
rect 11500 4324 11536 4434
rect 11723 4413 11754 4434
rect 12069 4427 12072 4447
rect 12092 4427 12485 4447
rect 12669 4437 12703 4453
rect 12747 4505 12890 4526
rect 13272 4555 13705 4559
rect 13272 4549 13711 4555
rect 13272 4531 13293 4549
rect 13311 4531 13711 4549
rect 14710 4534 14741 4585
rect 14776 4614 14813 4684
rect 15079 4683 15116 4684
rect 14928 4624 14964 4625
rect 14776 4594 14785 4614
rect 14805 4594 14813 4614
rect 14776 4584 14813 4594
rect 14872 4614 15020 4624
rect 15120 4621 15216 4623
rect 14872 4594 14881 4614
rect 14901 4594 14991 4614
rect 15011 4594 15020 4614
rect 14872 4585 15020 4594
rect 15078 4614 15216 4621
rect 15078 4594 15087 4614
rect 15107 4594 15216 4614
rect 15078 4585 15216 4594
rect 14872 4584 14909 4585
rect 14602 4531 14643 4532
rect 13272 4513 13711 4531
rect 12445 4418 12485 4427
rect 12747 4418 12774 4505
rect 12847 4479 12890 4505
rect 12847 4461 12860 4479
rect 12878 4461 12890 4479
rect 12847 4450 12890 4461
rect 11719 4412 11754 4413
rect 11597 4402 11754 4412
rect 11597 4382 11614 4402
rect 11634 4382 11754 4402
rect 11597 4375 11754 4382
rect 11821 4405 11967 4413
rect 11821 4385 11832 4405
rect 11852 4385 11891 4405
rect 11911 4385 11967 4405
rect 12445 4401 12774 4418
rect 12445 4400 12485 4401
rect 11821 4378 11967 4385
rect 12842 4389 12882 4392
rect 12842 4383 12885 4389
rect 12467 4380 12885 4383
rect 11821 4377 11862 4378
rect 11555 4324 11592 4325
rect 11248 4315 11386 4324
rect 11248 4295 11357 4315
rect 11377 4295 11386 4315
rect 11248 4288 11386 4295
rect 11444 4315 11592 4324
rect 11444 4295 11453 4315
rect 11473 4295 11563 4315
rect 11583 4295 11592 4315
rect 11248 4286 11344 4288
rect 11444 4285 11592 4295
rect 11651 4315 11688 4325
rect 11651 4295 11659 4315
rect 11679 4295 11688 4315
rect 11500 4284 11536 4285
rect 11348 4225 11385 4226
rect 11651 4225 11688 4295
rect 11723 4324 11754 4375
rect 12467 4362 12858 4380
rect 12876 4362 12885 4380
rect 12467 4360 12885 4362
rect 12467 4352 12494 4360
rect 12735 4357 12885 4360
rect 12047 4346 12215 4347
rect 12466 4346 12494 4352
rect 12047 4330 12494 4346
rect 12842 4352 12885 4357
rect 11773 4324 11810 4325
rect 11723 4315 11810 4324
rect 11723 4295 11781 4315
rect 11801 4295 11810 4315
rect 11723 4285 11810 4295
rect 11869 4315 11906 4325
rect 11869 4295 11877 4315
rect 11897 4295 11906 4315
rect 11723 4284 11754 4285
rect 11347 4224 11688 4225
rect 11869 4224 11906 4295
rect 11272 4219 11688 4224
rect 11272 4199 11275 4219
rect 11295 4199 11688 4219
rect 11719 4200 11906 4224
rect 12047 4320 12491 4330
rect 12047 4318 12215 4320
rect 11081 4125 11125 4126
rect 11081 4119 11126 4125
rect 11081 4101 11093 4119
rect 11115 4101 11126 4119
rect 11147 4120 11189 4165
rect 12047 4140 12074 4318
rect 12114 4280 12178 4292
rect 12454 4288 12491 4320
rect 12517 4319 12708 4341
rect 12672 4317 12708 4319
rect 12672 4288 12709 4317
rect 12842 4296 12882 4352
rect 12114 4279 12149 4280
rect 12091 4274 12149 4279
rect 12091 4254 12094 4274
rect 12114 4260 12149 4274
rect 12169 4260 12178 4280
rect 12114 4252 12178 4260
rect 12140 4251 12178 4252
rect 12141 4250 12178 4251
rect 12244 4284 12280 4285
rect 12352 4284 12388 4285
rect 12244 4276 12388 4284
rect 12244 4256 12252 4276
rect 12272 4256 12307 4276
rect 12327 4256 12360 4276
rect 12380 4256 12388 4276
rect 12244 4250 12388 4256
rect 12454 4280 12492 4288
rect 12570 4284 12606 4285
rect 12454 4260 12463 4280
rect 12483 4260 12492 4280
rect 12454 4251 12492 4260
rect 12521 4276 12606 4284
rect 12521 4256 12578 4276
rect 12598 4256 12606 4276
rect 12454 4250 12491 4251
rect 12521 4250 12606 4256
rect 12672 4280 12710 4288
rect 12672 4260 12681 4280
rect 12701 4260 12710 4280
rect 12842 4278 12854 4296
rect 12872 4278 12882 4296
rect 13274 4324 13326 4513
rect 13672 4488 13711 4513
rect 14494 4524 14643 4531
rect 14494 4504 14553 4524
rect 14573 4504 14612 4524
rect 14632 4504 14643 4524
rect 14494 4496 14643 4504
rect 14710 4527 14867 4534
rect 14710 4507 14830 4527
rect 14850 4507 14867 4527
rect 14710 4497 14867 4507
rect 14710 4496 14745 4497
rect 13456 4463 13643 4487
rect 13672 4468 14067 4488
rect 14087 4468 14090 4488
rect 14710 4475 14741 4496
rect 14928 4475 14964 4585
rect 14983 4584 15020 4585
rect 15079 4584 15116 4585
rect 15039 4525 15129 4531
rect 15039 4505 15048 4525
rect 15068 4523 15129 4525
rect 15068 4505 15093 4523
rect 15039 4503 15093 4505
rect 15113 4503 15129 4523
rect 15039 4497 15129 4503
rect 14553 4474 14590 4475
rect 13672 4463 14090 4468
rect 14552 4465 14590 4474
rect 13456 4392 13493 4463
rect 13672 4462 14015 4463
rect 13672 4459 13711 4462
rect 13977 4461 14014 4462
rect 13608 4402 13639 4403
rect 13456 4372 13465 4392
rect 13485 4372 13493 4392
rect 13456 4362 13493 4372
rect 13552 4392 13639 4402
rect 13552 4372 13561 4392
rect 13581 4372 13639 4392
rect 13552 4363 13639 4372
rect 13552 4362 13589 4363
rect 13274 4306 13290 4324
rect 13308 4306 13326 4324
rect 13608 4312 13639 4363
rect 13674 4392 13711 4459
rect 14552 4445 14561 4465
rect 14581 4445 14590 4465
rect 14552 4437 14590 4445
rect 14656 4469 14741 4475
rect 14771 4474 14808 4475
rect 14656 4449 14664 4469
rect 14684 4449 14741 4469
rect 14656 4441 14741 4449
rect 14770 4465 14808 4474
rect 14770 4445 14779 4465
rect 14799 4445 14808 4465
rect 14656 4440 14692 4441
rect 14770 4437 14808 4445
rect 14874 4469 15018 4475
rect 14874 4449 14882 4469
rect 14902 4463 14990 4469
rect 14902 4449 14931 4463
rect 14874 4441 14931 4449
rect 14874 4440 14910 4441
rect 14954 4449 14990 4463
rect 15010 4449 15018 4469
rect 14954 4441 15018 4449
rect 14982 4440 15018 4441
rect 15084 4474 15121 4475
rect 15084 4473 15122 4474
rect 15084 4465 15148 4473
rect 15084 4445 15093 4465
rect 15113 4451 15148 4465
rect 15168 4451 15171 4471
rect 15113 4446 15171 4451
rect 15113 4445 15148 4446
rect 14553 4408 14590 4437
rect 14554 4406 14590 4408
rect 13826 4402 13862 4403
rect 13674 4372 13683 4392
rect 13703 4372 13711 4392
rect 13674 4362 13711 4372
rect 13770 4392 13918 4402
rect 14018 4399 14114 4401
rect 13770 4372 13779 4392
rect 13799 4372 13889 4392
rect 13909 4372 13918 4392
rect 13770 4363 13918 4372
rect 13976 4392 14114 4399
rect 13976 4372 13985 4392
rect 14005 4372 14114 4392
rect 14554 4384 14745 4406
rect 14771 4405 14808 4437
rect 15084 4433 15148 4445
rect 15188 4407 15215 4585
rect 15512 4538 15549 4544
rect 15512 4519 15520 4538
rect 15541 4519 15549 4538
rect 15512 4511 15549 4519
rect 15047 4405 15215 4407
rect 14771 4379 15215 4405
rect 14881 4377 14921 4379
rect 15047 4378 15215 4379
rect 13976 4363 14114 4372
rect 15174 4373 15215 4378
rect 13770 4362 13807 4363
rect 13500 4309 13541 4310
rect 13274 4288 13326 4306
rect 13392 4302 13541 4309
rect 12842 4268 12882 4278
rect 13392 4282 13451 4302
rect 13471 4282 13510 4302
rect 13530 4282 13541 4302
rect 13392 4274 13541 4282
rect 13608 4305 13765 4312
rect 13608 4285 13728 4305
rect 13748 4285 13765 4305
rect 13608 4275 13765 4285
rect 13608 4274 13643 4275
rect 12672 4251 12710 4260
rect 13608 4253 13639 4274
rect 13826 4253 13862 4363
rect 13881 4362 13918 4363
rect 13977 4362 14014 4363
rect 13937 4303 14027 4309
rect 13937 4283 13946 4303
rect 13966 4301 14027 4303
rect 13966 4283 13991 4301
rect 13937 4281 13991 4283
rect 14011 4281 14027 4301
rect 13937 4275 14027 4281
rect 13451 4252 13488 4253
rect 12672 4250 12709 4251
rect 12133 4222 12223 4228
rect 12133 4202 12149 4222
rect 12169 4220 12223 4222
rect 12169 4202 12194 4220
rect 12133 4200 12194 4202
rect 12214 4200 12223 4220
rect 12133 4194 12223 4200
rect 12146 4140 12183 4141
rect 12242 4140 12279 4141
rect 12298 4140 12334 4250
rect 12521 4229 12552 4250
rect 13450 4243 13488 4252
rect 12517 4228 12552 4229
rect 12395 4218 12552 4228
rect 12395 4198 12412 4218
rect 12432 4198 12552 4218
rect 12395 4191 12552 4198
rect 12619 4221 12768 4229
rect 12619 4201 12630 4221
rect 12650 4201 12689 4221
rect 12709 4201 12768 4221
rect 13278 4225 13318 4235
rect 12619 4194 12768 4201
rect 12834 4197 12886 4215
rect 12619 4193 12660 4194
rect 12353 4140 12390 4141
rect 12046 4131 12184 4140
rect 11518 4120 11551 4122
rect 11147 4108 11594 4120
rect 11081 4071 11126 4101
rect 11098 3125 11126 4071
rect 11150 4094 11594 4108
rect 11150 4092 11318 4094
rect 11150 3914 11177 4092
rect 11217 4054 11281 4066
rect 11557 4062 11594 4094
rect 11620 4093 11811 4115
rect 12046 4111 12155 4131
rect 12175 4111 12184 4131
rect 12046 4104 12184 4111
rect 12242 4131 12390 4140
rect 12242 4111 12251 4131
rect 12271 4111 12361 4131
rect 12381 4111 12390 4131
rect 12046 4102 12142 4104
rect 12242 4101 12390 4111
rect 12449 4131 12486 4141
rect 12449 4111 12457 4131
rect 12477 4111 12486 4131
rect 12298 4100 12334 4101
rect 11775 4091 11811 4093
rect 11775 4062 11812 4091
rect 11217 4053 11252 4054
rect 11194 4048 11252 4053
rect 11194 4028 11197 4048
rect 11217 4034 11252 4048
rect 11272 4034 11281 4054
rect 11217 4026 11281 4034
rect 11243 4025 11281 4026
rect 11244 4024 11281 4025
rect 11347 4058 11383 4059
rect 11455 4058 11491 4059
rect 11347 4052 11491 4058
rect 11347 4050 11408 4052
rect 11347 4030 11355 4050
rect 11375 4035 11408 4050
rect 11427 4050 11491 4052
rect 11427 4035 11463 4050
rect 11375 4030 11463 4035
rect 11483 4030 11491 4050
rect 11347 4024 11491 4030
rect 11557 4054 11595 4062
rect 11673 4058 11709 4059
rect 11557 4034 11566 4054
rect 11586 4034 11595 4054
rect 11557 4025 11595 4034
rect 11624 4050 11709 4058
rect 11624 4030 11681 4050
rect 11701 4030 11709 4050
rect 11557 4024 11594 4025
rect 11624 4024 11709 4030
rect 11775 4054 11813 4062
rect 11775 4034 11784 4054
rect 11804 4034 11813 4054
rect 12449 4044 12486 4111
rect 12521 4140 12552 4191
rect 12834 4179 12852 4197
rect 12870 4179 12886 4197
rect 12571 4140 12608 4141
rect 12521 4131 12608 4140
rect 12521 4111 12579 4131
rect 12599 4111 12608 4131
rect 12521 4101 12608 4111
rect 12667 4131 12704 4141
rect 12667 4111 12675 4131
rect 12695 4111 12704 4131
rect 12521 4100 12552 4101
rect 12146 4041 12183 4042
rect 12449 4041 12488 4044
rect 12145 4040 12488 4041
rect 12667 4040 12704 4111
rect 11775 4025 11813 4034
rect 12070 4035 12488 4040
rect 11775 4024 11812 4025
rect 11236 3996 11326 4002
rect 11236 3976 11252 3996
rect 11272 3994 11326 3996
rect 11272 3976 11297 3994
rect 11236 3974 11297 3976
rect 11317 3974 11326 3994
rect 11236 3968 11326 3974
rect 11249 3914 11286 3915
rect 11345 3914 11382 3915
rect 11401 3914 11437 4024
rect 11624 4003 11655 4024
rect 12070 4015 12073 4035
rect 12093 4015 12488 4035
rect 12517 4016 12704 4040
rect 11620 4002 11655 4003
rect 11498 3992 11655 4002
rect 11498 3972 11515 3992
rect 11535 3972 11655 3992
rect 11498 3965 11655 3972
rect 11722 3995 11871 4003
rect 11722 3975 11733 3995
rect 11753 3975 11792 3995
rect 11812 3975 11871 3995
rect 11722 3968 11871 3975
rect 12449 3990 12488 4015
rect 12834 3990 12886 4179
rect 13278 4207 13288 4225
rect 13306 4207 13318 4225
rect 13450 4223 13459 4243
rect 13479 4223 13488 4243
rect 13450 4215 13488 4223
rect 13554 4247 13639 4253
rect 13669 4252 13706 4253
rect 13554 4227 13562 4247
rect 13582 4227 13639 4247
rect 13554 4219 13639 4227
rect 13668 4243 13706 4252
rect 13668 4223 13677 4243
rect 13697 4223 13706 4243
rect 13554 4218 13590 4219
rect 13668 4215 13706 4223
rect 13772 4247 13916 4253
rect 13772 4227 13780 4247
rect 13800 4227 13833 4247
rect 13853 4227 13888 4247
rect 13908 4227 13916 4247
rect 13772 4219 13916 4227
rect 13772 4218 13808 4219
rect 13880 4218 13916 4219
rect 13982 4252 14019 4253
rect 13982 4251 14020 4252
rect 13982 4243 14046 4251
rect 13982 4223 13991 4243
rect 14011 4229 14046 4243
rect 14066 4229 14069 4249
rect 14011 4224 14069 4229
rect 14011 4223 14046 4224
rect 13278 4151 13318 4207
rect 13451 4186 13488 4215
rect 13452 4184 13488 4186
rect 13452 4162 13643 4184
rect 13669 4183 13706 4215
rect 13982 4211 14046 4223
rect 14086 4185 14113 4363
rect 13945 4183 14113 4185
rect 13669 4173 14113 4183
rect 14254 4279 14441 4303
rect 14472 4284 14865 4304
rect 14885 4284 14888 4304
rect 14472 4279 14888 4284
rect 14254 4208 14291 4279
rect 14472 4278 14813 4279
rect 14406 4218 14437 4219
rect 14254 4188 14263 4208
rect 14283 4188 14291 4208
rect 14254 4178 14291 4188
rect 14350 4208 14437 4218
rect 14350 4188 14359 4208
rect 14379 4188 14437 4208
rect 14350 4179 14437 4188
rect 14350 4178 14387 4179
rect 13275 4146 13318 4151
rect 13666 4157 14113 4173
rect 13666 4151 13694 4157
rect 13945 4156 14113 4157
rect 13275 4143 13425 4146
rect 13666 4143 13693 4151
rect 13275 4141 13693 4143
rect 13275 4123 13284 4141
rect 13302 4123 13693 4141
rect 14406 4128 14437 4179
rect 14472 4208 14509 4278
rect 14775 4277 14812 4278
rect 14624 4218 14660 4219
rect 14472 4188 14481 4208
rect 14501 4188 14509 4208
rect 14472 4178 14509 4188
rect 14568 4208 14716 4218
rect 14816 4215 14912 4217
rect 14568 4188 14577 4208
rect 14597 4188 14687 4208
rect 14707 4188 14716 4208
rect 14568 4179 14716 4188
rect 14774 4208 14912 4215
rect 14774 4188 14783 4208
rect 14803 4188 14912 4208
rect 15174 4191 15214 4373
rect 14774 4179 14912 4188
rect 14568 4178 14605 4179
rect 14298 4125 14339 4126
rect 13275 4120 13693 4123
rect 13275 4114 13318 4120
rect 13278 4111 13318 4114
rect 14190 4118 14339 4125
rect 13675 4102 13715 4103
rect 13386 4085 13715 4102
rect 14190 4098 14249 4118
rect 14269 4098 14308 4118
rect 14328 4098 14339 4118
rect 14190 4090 14339 4098
rect 14406 4121 14563 4128
rect 14406 4101 14526 4121
rect 14546 4101 14563 4121
rect 14406 4091 14563 4101
rect 14406 4090 14441 4091
rect 13270 4042 13313 4053
rect 13270 4024 13282 4042
rect 13300 4024 13313 4042
rect 13270 3998 13313 4024
rect 13386 3998 13413 4085
rect 13675 4076 13715 4085
rect 12449 3972 12888 3990
rect 11722 3967 11763 3968
rect 11456 3914 11493 3915
rect 11149 3905 11287 3914
rect 11149 3885 11258 3905
rect 11278 3885 11287 3905
rect 11149 3878 11287 3885
rect 11345 3905 11493 3914
rect 11345 3885 11354 3905
rect 11374 3885 11464 3905
rect 11484 3885 11493 3905
rect 11149 3876 11245 3878
rect 11345 3875 11493 3885
rect 11552 3905 11589 3915
rect 11552 3885 11560 3905
rect 11580 3885 11589 3905
rect 11401 3874 11437 3875
rect 11249 3815 11286 3816
rect 11552 3815 11589 3885
rect 11624 3914 11655 3965
rect 12449 3954 12849 3972
rect 12867 3954 12888 3972
rect 12449 3948 12888 3954
rect 12455 3944 12888 3948
rect 13270 3977 13413 3998
rect 13457 4050 13491 4066
rect 13675 4056 14068 4076
rect 14088 4056 14091 4076
rect 14406 4069 14437 4090
rect 14624 4069 14660 4179
rect 14679 4178 14716 4179
rect 14775 4178 14812 4179
rect 14735 4119 14825 4125
rect 14735 4099 14744 4119
rect 14764 4117 14825 4119
rect 14764 4099 14789 4117
rect 14735 4097 14789 4099
rect 14809 4097 14825 4117
rect 14735 4091 14825 4097
rect 14249 4068 14286 4069
rect 13675 4051 14091 4056
rect 14248 4059 14286 4068
rect 13675 4050 14016 4051
rect 13457 3980 13494 4050
rect 13609 3990 13640 3991
rect 13270 3975 13407 3977
rect 12834 3942 12886 3944
rect 13270 3933 13313 3975
rect 13457 3960 13466 3980
rect 13486 3960 13494 3980
rect 13457 3950 13494 3960
rect 13553 3980 13640 3990
rect 13553 3960 13562 3980
rect 13582 3960 13640 3980
rect 13553 3951 13640 3960
rect 13553 3950 13590 3951
rect 13268 3923 13313 3933
rect 11674 3914 11711 3915
rect 11624 3905 11711 3914
rect 11624 3885 11682 3905
rect 11702 3885 11711 3905
rect 11624 3875 11711 3885
rect 11770 3905 11807 3915
rect 11770 3885 11778 3905
rect 11798 3885 11807 3905
rect 13268 3905 13277 3923
rect 13295 3905 13313 3923
rect 13268 3899 13313 3905
rect 13609 3900 13640 3951
rect 13675 3980 13712 4050
rect 13978 4049 14015 4050
rect 14248 4039 14257 4059
rect 14277 4039 14286 4059
rect 14248 4031 14286 4039
rect 14352 4063 14437 4069
rect 14467 4068 14504 4069
rect 14352 4043 14360 4063
rect 14380 4043 14437 4063
rect 14352 4035 14437 4043
rect 14466 4059 14504 4068
rect 14466 4039 14475 4059
rect 14495 4039 14504 4059
rect 14352 4034 14388 4035
rect 14466 4031 14504 4039
rect 14570 4063 14714 4069
rect 14570 4043 14578 4063
rect 14598 4044 14630 4063
rect 14651 4044 14686 4063
rect 14598 4043 14686 4044
rect 14706 4043 14714 4063
rect 14570 4035 14714 4043
rect 14570 4034 14606 4035
rect 14678 4034 14714 4035
rect 14780 4068 14817 4069
rect 14780 4067 14818 4068
rect 14780 4059 14844 4067
rect 14780 4039 14789 4059
rect 14809 4045 14844 4059
rect 14864 4045 14867 4065
rect 14809 4040 14867 4045
rect 14809 4039 14844 4040
rect 14249 4002 14286 4031
rect 14250 4000 14286 4002
rect 13827 3990 13863 3991
rect 13675 3960 13684 3980
rect 13704 3960 13712 3980
rect 13675 3950 13712 3960
rect 13771 3980 13919 3990
rect 14019 3987 14115 3989
rect 13771 3960 13780 3980
rect 13800 3960 13890 3980
rect 13910 3960 13919 3980
rect 13771 3951 13919 3960
rect 13977 3980 14115 3987
rect 13977 3960 13986 3980
rect 14006 3960 14115 3980
rect 14250 3978 14441 4000
rect 14467 3999 14504 4031
rect 14780 4027 14844 4039
rect 14884 4001 14911 4179
rect 14743 3999 14911 4001
rect 14467 3973 14911 3999
rect 13977 3951 14115 3960
rect 13771 3950 13808 3951
rect 13268 3896 13305 3899
rect 13501 3897 13542 3898
rect 11624 3874 11655 3875
rect 11248 3814 11589 3815
rect 11770 3814 11807 3885
rect 13393 3890 13542 3897
rect 12837 3877 12874 3882
rect 12828 3873 12875 3877
rect 12828 3855 12847 3873
rect 12865 3855 12875 3873
rect 13393 3870 13452 3890
rect 13472 3870 13511 3890
rect 13531 3870 13542 3890
rect 13393 3862 13542 3870
rect 13609 3893 13766 3900
rect 13609 3873 13729 3893
rect 13749 3873 13766 3893
rect 13609 3863 13766 3873
rect 13609 3862 13644 3863
rect 11173 3809 11589 3814
rect 11173 3789 11176 3809
rect 11196 3789 11589 3809
rect 11620 3790 11807 3814
rect 12432 3812 12472 3817
rect 12828 3812 12875 3855
rect 13609 3841 13640 3862
rect 13827 3841 13863 3951
rect 13882 3950 13919 3951
rect 13978 3950 14015 3951
rect 13938 3891 14028 3897
rect 13938 3871 13947 3891
rect 13967 3889 14028 3891
rect 13967 3871 13992 3889
rect 13938 3869 13992 3871
rect 14012 3869 14028 3889
rect 13938 3863 14028 3869
rect 13452 3840 13489 3841
rect 12432 3773 12875 3812
rect 13265 3832 13302 3834
rect 13265 3824 13307 3832
rect 13265 3806 13275 3824
rect 13293 3806 13307 3824
rect 13265 3797 13307 3806
rect 13451 3831 13489 3840
rect 13451 3811 13460 3831
rect 13480 3811 13489 3831
rect 13451 3803 13489 3811
rect 13555 3835 13640 3841
rect 13670 3840 13707 3841
rect 13555 3815 13563 3835
rect 13583 3815 13640 3835
rect 13555 3807 13640 3815
rect 13669 3831 13707 3840
rect 13669 3811 13678 3831
rect 13698 3811 13707 3831
rect 13555 3806 13591 3807
rect 13669 3803 13707 3811
rect 13773 3839 13917 3841
rect 13773 3835 13825 3839
rect 13773 3815 13781 3835
rect 13801 3819 13825 3835
rect 13845 3835 13917 3839
rect 13845 3819 13889 3835
rect 13801 3815 13889 3819
rect 13909 3815 13917 3835
rect 13773 3807 13917 3815
rect 13773 3806 13809 3807
rect 13881 3806 13917 3807
rect 13983 3840 14020 3841
rect 13983 3839 14021 3840
rect 13983 3831 14047 3839
rect 13983 3811 13992 3831
rect 14012 3817 14047 3831
rect 14067 3817 14070 3837
rect 14012 3812 14070 3817
rect 14012 3811 14047 3812
rect 11526 3758 11566 3766
rect 11526 3736 11534 3758
rect 11558 3736 11566 3758
rect 11232 3512 11400 3513
rect 11526 3512 11566 3736
rect 12029 3740 12197 3741
rect 12432 3740 12472 3773
rect 12828 3740 12875 3773
rect 13266 3772 13307 3797
rect 13452 3772 13489 3803
rect 13670 3772 13707 3803
rect 13983 3799 14047 3811
rect 14087 3773 14114 3951
rect 13266 3745 13315 3772
rect 13451 3746 13500 3772
rect 13669 3771 13750 3772
rect 13946 3771 14114 3773
rect 13669 3746 14114 3771
rect 13670 3745 14114 3746
rect 12029 3739 12473 3740
rect 12029 3714 12474 3739
rect 12029 3712 12197 3714
rect 12393 3713 12474 3714
rect 12643 3713 12692 3739
rect 12828 3713 12877 3740
rect 12029 3534 12056 3712
rect 12096 3674 12160 3686
rect 12436 3682 12473 3713
rect 12654 3682 12691 3713
rect 12836 3688 12877 3713
rect 13268 3712 13315 3745
rect 13671 3712 13711 3745
rect 13946 3744 14114 3745
rect 14577 3749 14617 3973
rect 14743 3972 14911 3973
rect 14577 3727 14585 3749
rect 14609 3727 14617 3749
rect 14577 3719 14617 3727
rect 12096 3673 12131 3674
rect 12073 3668 12131 3673
rect 12073 3648 12076 3668
rect 12096 3654 12131 3668
rect 12151 3654 12160 3674
rect 12096 3646 12160 3654
rect 12122 3645 12160 3646
rect 12123 3644 12160 3645
rect 12226 3678 12262 3679
rect 12334 3678 12370 3679
rect 12226 3670 12370 3678
rect 12226 3650 12234 3670
rect 12254 3666 12342 3670
rect 12254 3650 12298 3666
rect 12226 3646 12298 3650
rect 12318 3650 12342 3666
rect 12362 3650 12370 3670
rect 12318 3646 12370 3650
rect 12226 3644 12370 3646
rect 12436 3674 12474 3682
rect 12552 3678 12588 3679
rect 12436 3654 12445 3674
rect 12465 3654 12474 3674
rect 12436 3645 12474 3654
rect 12503 3670 12588 3678
rect 12503 3650 12560 3670
rect 12580 3650 12588 3670
rect 12436 3644 12473 3645
rect 12503 3644 12588 3650
rect 12654 3674 12692 3682
rect 12654 3654 12663 3674
rect 12683 3654 12692 3674
rect 12654 3645 12692 3654
rect 12836 3679 12878 3688
rect 12836 3661 12850 3679
rect 12868 3661 12878 3679
rect 12836 3653 12878 3661
rect 12841 3651 12878 3653
rect 13268 3673 13711 3712
rect 12654 3644 12691 3645
rect 12115 3616 12205 3622
rect 12115 3596 12131 3616
rect 12151 3614 12205 3616
rect 12151 3596 12176 3614
rect 12115 3594 12176 3596
rect 12196 3594 12205 3614
rect 12115 3588 12205 3594
rect 12128 3534 12165 3535
rect 12224 3534 12261 3535
rect 12280 3534 12316 3644
rect 12503 3623 12534 3644
rect 13268 3630 13315 3673
rect 13671 3668 13711 3673
rect 14336 3671 14523 3695
rect 14554 3676 14947 3696
rect 14967 3676 14970 3696
rect 14554 3671 14970 3676
rect 12499 3622 12534 3623
rect 12377 3612 12534 3622
rect 12377 3592 12394 3612
rect 12414 3592 12534 3612
rect 12377 3585 12534 3592
rect 12601 3615 12750 3623
rect 12601 3595 12612 3615
rect 12632 3595 12671 3615
rect 12691 3595 12750 3615
rect 13268 3612 13278 3630
rect 13296 3612 13315 3630
rect 13268 3608 13315 3612
rect 13269 3603 13306 3608
rect 12601 3588 12750 3595
rect 14336 3600 14373 3671
rect 14554 3670 14895 3671
rect 14488 3610 14519 3611
rect 12601 3587 12642 3588
rect 12838 3586 12875 3589
rect 12335 3534 12372 3535
rect 12028 3525 12166 3534
rect 11232 3486 11676 3512
rect 11232 3484 11400 3486
rect 11232 3306 11259 3484
rect 11299 3446 11363 3458
rect 11639 3454 11676 3486
rect 11702 3485 11893 3507
rect 12028 3505 12137 3525
rect 12157 3505 12166 3525
rect 12028 3498 12166 3505
rect 12224 3525 12372 3534
rect 12224 3505 12233 3525
rect 12253 3505 12343 3525
rect 12363 3505 12372 3525
rect 12028 3496 12124 3498
rect 12224 3495 12372 3505
rect 12431 3525 12468 3535
rect 12431 3505 12439 3525
rect 12459 3505 12468 3525
rect 12280 3494 12316 3495
rect 11857 3483 11893 3485
rect 11857 3454 11894 3483
rect 11299 3445 11334 3446
rect 11276 3440 11334 3445
rect 11276 3420 11279 3440
rect 11299 3426 11334 3440
rect 11354 3426 11363 3446
rect 11299 3418 11363 3426
rect 11325 3417 11363 3418
rect 11326 3416 11363 3417
rect 11429 3450 11465 3451
rect 11537 3450 11573 3451
rect 11429 3442 11573 3450
rect 11429 3422 11437 3442
rect 11457 3441 11545 3442
rect 11457 3422 11492 3441
rect 11513 3422 11545 3441
rect 11565 3422 11573 3442
rect 11429 3416 11573 3422
rect 11639 3446 11677 3454
rect 11755 3450 11791 3451
rect 11639 3426 11648 3446
rect 11668 3426 11677 3446
rect 11639 3417 11677 3426
rect 11706 3442 11791 3450
rect 11706 3422 11763 3442
rect 11783 3422 11791 3442
rect 11639 3416 11676 3417
rect 11706 3416 11791 3422
rect 11857 3446 11895 3454
rect 11857 3426 11866 3446
rect 11886 3426 11895 3446
rect 12128 3435 12165 3436
rect 12431 3435 12468 3505
rect 12503 3534 12534 3585
rect 12830 3580 12875 3586
rect 12830 3562 12848 3580
rect 12866 3562 12875 3580
rect 14336 3580 14345 3600
rect 14365 3580 14373 3600
rect 14336 3570 14373 3580
rect 14432 3600 14519 3610
rect 14432 3580 14441 3600
rect 14461 3580 14519 3600
rect 14432 3571 14519 3580
rect 14432 3570 14469 3571
rect 12830 3552 12875 3562
rect 12553 3534 12590 3535
rect 12503 3525 12590 3534
rect 12503 3505 12561 3525
rect 12581 3505 12590 3525
rect 12503 3495 12590 3505
rect 12649 3525 12686 3535
rect 12649 3505 12657 3525
rect 12677 3505 12686 3525
rect 12830 3510 12873 3552
rect 13257 3541 13309 3543
rect 12736 3508 12873 3510
rect 12503 3494 12534 3495
rect 12649 3435 12686 3505
rect 12127 3434 12468 3435
rect 11857 3417 11895 3426
rect 12052 3429 12468 3434
rect 11857 3416 11894 3417
rect 11318 3388 11408 3394
rect 11318 3368 11334 3388
rect 11354 3386 11408 3388
rect 11354 3368 11379 3386
rect 11318 3366 11379 3368
rect 11399 3366 11408 3386
rect 11318 3360 11408 3366
rect 11331 3306 11368 3307
rect 11427 3306 11464 3307
rect 11483 3306 11519 3416
rect 11706 3395 11737 3416
rect 12052 3409 12055 3429
rect 12075 3409 12468 3429
rect 12652 3419 12686 3435
rect 12730 3487 12873 3508
rect 13255 3537 13688 3541
rect 13255 3531 13694 3537
rect 13255 3513 13276 3531
rect 13294 3513 13694 3531
rect 14488 3520 14519 3571
rect 14554 3600 14591 3670
rect 14857 3669 14894 3670
rect 14706 3610 14742 3611
rect 14554 3580 14563 3600
rect 14583 3580 14591 3600
rect 14554 3570 14591 3580
rect 14650 3600 14798 3610
rect 14898 3607 14994 3609
rect 14650 3580 14659 3600
rect 14679 3580 14769 3600
rect 14789 3580 14798 3600
rect 14650 3571 14798 3580
rect 14856 3600 14994 3607
rect 14856 3580 14865 3600
rect 14885 3580 14994 3600
rect 14856 3571 14994 3580
rect 14650 3570 14687 3571
rect 14380 3517 14421 3518
rect 13255 3495 13694 3513
rect 12428 3400 12468 3409
rect 12730 3400 12757 3487
rect 12830 3461 12873 3487
rect 12830 3443 12843 3461
rect 12861 3443 12873 3461
rect 12830 3432 12873 3443
rect 11702 3394 11737 3395
rect 11580 3384 11737 3394
rect 11580 3364 11597 3384
rect 11617 3364 11737 3384
rect 11580 3357 11737 3364
rect 11804 3387 11953 3395
rect 11804 3367 11815 3387
rect 11835 3367 11874 3387
rect 11894 3367 11953 3387
rect 12428 3383 12757 3400
rect 12428 3382 12468 3383
rect 11804 3360 11953 3367
rect 12825 3371 12865 3374
rect 12825 3365 12868 3371
rect 12450 3362 12868 3365
rect 11804 3359 11845 3360
rect 11538 3306 11575 3307
rect 11231 3297 11369 3306
rect 11231 3277 11340 3297
rect 11360 3277 11369 3297
rect 11231 3270 11369 3277
rect 11427 3297 11575 3306
rect 11427 3277 11436 3297
rect 11456 3277 11546 3297
rect 11566 3277 11575 3297
rect 11231 3268 11327 3270
rect 11427 3267 11575 3277
rect 11634 3297 11671 3307
rect 11634 3277 11642 3297
rect 11662 3277 11671 3297
rect 11483 3266 11519 3267
rect 11331 3207 11368 3208
rect 11634 3207 11671 3277
rect 11706 3306 11737 3357
rect 12450 3344 12841 3362
rect 12859 3344 12868 3362
rect 12450 3342 12868 3344
rect 12450 3334 12477 3342
rect 12718 3339 12868 3342
rect 12030 3328 12198 3329
rect 12449 3328 12477 3334
rect 12030 3312 12477 3328
rect 12825 3334 12868 3339
rect 11756 3306 11793 3307
rect 11706 3297 11793 3306
rect 11706 3277 11764 3297
rect 11784 3277 11793 3297
rect 11706 3267 11793 3277
rect 11852 3297 11889 3307
rect 11852 3277 11860 3297
rect 11880 3277 11889 3297
rect 11706 3266 11737 3267
rect 11330 3206 11671 3207
rect 11852 3206 11889 3277
rect 11255 3201 11671 3206
rect 11255 3181 11258 3201
rect 11278 3181 11671 3201
rect 11702 3182 11889 3206
rect 12030 3302 12474 3312
rect 12030 3300 12198 3302
rect 11097 3107 11126 3125
rect 12030 3122 12057 3300
rect 12097 3262 12161 3274
rect 12437 3270 12474 3302
rect 12500 3301 12691 3323
rect 12655 3299 12691 3301
rect 12655 3270 12692 3299
rect 12825 3278 12865 3334
rect 12097 3261 12132 3262
rect 12074 3256 12132 3261
rect 12074 3236 12077 3256
rect 12097 3242 12132 3256
rect 12152 3242 12161 3262
rect 12097 3234 12161 3242
rect 12123 3233 12161 3234
rect 12124 3232 12161 3233
rect 12227 3266 12263 3267
rect 12335 3266 12371 3267
rect 12227 3258 12371 3266
rect 12227 3238 12235 3258
rect 12255 3238 12290 3258
rect 12310 3238 12343 3258
rect 12363 3238 12371 3258
rect 12227 3232 12371 3238
rect 12437 3262 12475 3270
rect 12553 3266 12589 3267
rect 12437 3242 12446 3262
rect 12466 3242 12475 3262
rect 12437 3233 12475 3242
rect 12504 3258 12589 3266
rect 12504 3238 12561 3258
rect 12581 3238 12589 3258
rect 12437 3232 12474 3233
rect 12504 3232 12589 3238
rect 12655 3262 12693 3270
rect 12655 3242 12664 3262
rect 12684 3242 12693 3262
rect 12825 3260 12837 3278
rect 12855 3260 12865 3278
rect 13257 3306 13309 3495
rect 13655 3470 13694 3495
rect 14272 3510 14421 3517
rect 14272 3490 14331 3510
rect 14351 3490 14390 3510
rect 14410 3490 14421 3510
rect 14272 3482 14421 3490
rect 14488 3513 14645 3520
rect 14488 3493 14608 3513
rect 14628 3493 14645 3513
rect 14488 3483 14645 3493
rect 14488 3482 14523 3483
rect 13439 3445 13626 3469
rect 13655 3450 14050 3470
rect 14070 3450 14073 3470
rect 14488 3461 14519 3482
rect 14706 3461 14742 3571
rect 14761 3570 14798 3571
rect 14857 3570 14894 3571
rect 14817 3511 14907 3517
rect 14817 3491 14826 3511
rect 14846 3509 14907 3511
rect 14846 3491 14871 3509
rect 14817 3489 14871 3491
rect 14891 3489 14907 3509
rect 14817 3483 14907 3489
rect 14331 3460 14368 3461
rect 13655 3445 14073 3450
rect 14330 3451 14368 3460
rect 13439 3374 13476 3445
rect 13655 3444 13998 3445
rect 13655 3441 13694 3444
rect 13960 3443 13997 3444
rect 13591 3384 13622 3385
rect 13439 3354 13448 3374
rect 13468 3354 13476 3374
rect 13439 3344 13476 3354
rect 13535 3374 13622 3384
rect 13535 3354 13544 3374
rect 13564 3354 13622 3374
rect 13535 3345 13622 3354
rect 13535 3344 13572 3345
rect 13257 3288 13273 3306
rect 13291 3288 13309 3306
rect 13591 3294 13622 3345
rect 13657 3374 13694 3441
rect 14330 3431 14339 3451
rect 14359 3431 14368 3451
rect 14330 3423 14368 3431
rect 14434 3455 14519 3461
rect 14549 3460 14586 3461
rect 14434 3435 14442 3455
rect 14462 3435 14519 3455
rect 14434 3427 14519 3435
rect 14548 3451 14586 3460
rect 14548 3431 14557 3451
rect 14577 3431 14586 3451
rect 14434 3426 14470 3427
rect 14548 3423 14586 3431
rect 14652 3456 14796 3461
rect 14652 3455 14714 3456
rect 14652 3435 14660 3455
rect 14680 3437 14714 3455
rect 14735 3455 14796 3456
rect 14735 3437 14768 3455
rect 14680 3435 14768 3437
rect 14788 3435 14796 3455
rect 14652 3427 14796 3435
rect 14652 3426 14688 3427
rect 14760 3426 14796 3427
rect 14862 3460 14899 3461
rect 14862 3459 14900 3460
rect 14862 3451 14926 3459
rect 14862 3431 14871 3451
rect 14891 3437 14926 3451
rect 14946 3437 14949 3457
rect 14891 3432 14949 3437
rect 14891 3431 14926 3432
rect 14331 3394 14368 3423
rect 14332 3392 14368 3394
rect 13809 3384 13845 3385
rect 13657 3354 13666 3374
rect 13686 3354 13694 3374
rect 13657 3344 13694 3354
rect 13753 3374 13901 3384
rect 14001 3381 14097 3383
rect 13753 3354 13762 3374
rect 13782 3354 13872 3374
rect 13892 3354 13901 3374
rect 13753 3345 13901 3354
rect 13959 3374 14097 3381
rect 13959 3354 13968 3374
rect 13988 3354 14097 3374
rect 14332 3370 14523 3392
rect 14549 3391 14586 3423
rect 14862 3419 14926 3431
rect 14966 3393 14993 3571
rect 14825 3391 14993 3393
rect 14549 3377 14993 3391
rect 14549 3365 14996 3377
rect 14592 3363 14625 3365
rect 13959 3345 14097 3354
rect 13753 3344 13790 3345
rect 13483 3291 13524 3292
rect 13257 3270 13309 3288
rect 13375 3284 13524 3291
rect 12825 3250 12865 3260
rect 13375 3264 13434 3284
rect 13454 3264 13493 3284
rect 13513 3264 13524 3284
rect 13375 3256 13524 3264
rect 13591 3287 13748 3294
rect 13591 3267 13711 3287
rect 13731 3267 13748 3287
rect 13591 3257 13748 3267
rect 13591 3256 13626 3257
rect 12655 3233 12693 3242
rect 13591 3235 13622 3256
rect 13809 3235 13845 3345
rect 13864 3344 13901 3345
rect 13960 3344 13997 3345
rect 13920 3285 14010 3291
rect 13920 3265 13929 3285
rect 13949 3283 14010 3285
rect 13949 3265 13974 3283
rect 13920 3263 13974 3265
rect 13994 3263 14010 3283
rect 13920 3257 14010 3263
rect 13434 3234 13471 3235
rect 12655 3232 12692 3233
rect 12116 3204 12206 3210
rect 12116 3184 12132 3204
rect 12152 3202 12206 3204
rect 12152 3184 12177 3202
rect 12116 3182 12177 3184
rect 12197 3182 12206 3202
rect 12116 3176 12206 3182
rect 12129 3122 12166 3123
rect 12225 3122 12262 3123
rect 12281 3122 12317 3232
rect 12504 3211 12535 3232
rect 13433 3225 13471 3234
rect 12500 3210 12535 3211
rect 12378 3200 12535 3210
rect 12378 3180 12395 3200
rect 12415 3180 12535 3200
rect 12378 3173 12535 3180
rect 12602 3203 12751 3211
rect 12602 3183 12613 3203
rect 12633 3183 12672 3203
rect 12692 3183 12751 3203
rect 13261 3207 13301 3217
rect 12602 3176 12751 3183
rect 12817 3179 12869 3197
rect 12602 3175 12643 3176
rect 12336 3122 12373 3123
rect 11067 3105 11126 3107
rect 12029 3113 12167 3122
rect 11067 3104 11235 3105
rect 11361 3104 11401 3106
rect 11067 3078 11511 3104
rect 11067 3076 11235 3078
rect 11067 3074 11148 3076
rect 11067 2898 11094 3074
rect 11134 3038 11198 3050
rect 11474 3046 11511 3078
rect 11537 3077 11728 3099
rect 12029 3093 12138 3113
rect 12158 3093 12167 3113
rect 12029 3086 12167 3093
rect 12225 3113 12373 3122
rect 12225 3093 12234 3113
rect 12254 3093 12344 3113
rect 12364 3093 12373 3113
rect 12029 3084 12125 3086
rect 12225 3083 12373 3093
rect 12432 3113 12469 3123
rect 12432 3093 12440 3113
rect 12460 3093 12469 3113
rect 12281 3082 12317 3083
rect 11692 3075 11728 3077
rect 11692 3046 11729 3075
rect 11134 3037 11169 3038
rect 11111 3032 11169 3037
rect 11111 3012 11114 3032
rect 11134 3018 11169 3032
rect 11189 3018 11198 3038
rect 11134 3010 11198 3018
rect 11160 3009 11198 3010
rect 11161 3008 11198 3009
rect 11264 3042 11300 3043
rect 11372 3042 11408 3043
rect 11264 3034 11408 3042
rect 11264 3014 11272 3034
rect 11292 3033 11380 3034
rect 11292 3015 11327 3033
rect 11345 3015 11380 3033
rect 11292 3014 11380 3015
rect 11400 3014 11408 3034
rect 11264 3008 11408 3014
rect 11474 3038 11512 3046
rect 11590 3042 11626 3043
rect 11474 3018 11483 3038
rect 11503 3018 11512 3038
rect 11474 3009 11512 3018
rect 11541 3034 11626 3042
rect 11541 3014 11598 3034
rect 11618 3014 11626 3034
rect 11474 3008 11511 3009
rect 11541 3008 11626 3014
rect 11692 3038 11730 3046
rect 11692 3018 11701 3038
rect 11721 3018 11730 3038
rect 12432 3026 12469 3093
rect 12504 3122 12535 3173
rect 12817 3161 12835 3179
rect 12853 3161 12869 3179
rect 12554 3122 12591 3123
rect 12504 3113 12591 3122
rect 12504 3093 12562 3113
rect 12582 3093 12591 3113
rect 12504 3083 12591 3093
rect 12650 3113 12687 3123
rect 12650 3093 12658 3113
rect 12678 3093 12687 3113
rect 12504 3082 12535 3083
rect 12129 3023 12166 3024
rect 12432 3023 12471 3026
rect 12128 3022 12471 3023
rect 12650 3022 12687 3093
rect 11692 3009 11730 3018
rect 12053 3017 12471 3022
rect 11692 3008 11729 3009
rect 11153 2980 11243 2986
rect 11153 2960 11169 2980
rect 11189 2978 11243 2980
rect 11189 2960 11214 2978
rect 11153 2958 11214 2960
rect 11234 2958 11243 2978
rect 11153 2952 11243 2958
rect 11166 2898 11203 2899
rect 11262 2898 11299 2899
rect 11318 2898 11354 3008
rect 11541 2987 11572 3008
rect 12053 2997 12056 3017
rect 12076 2997 12471 3017
rect 12500 2998 12687 3022
rect 11537 2986 11572 2987
rect 11415 2976 11572 2986
rect 11415 2956 11432 2976
rect 11452 2956 11572 2976
rect 11415 2949 11572 2956
rect 11639 2979 11788 2987
rect 11639 2959 11650 2979
rect 11670 2959 11709 2979
rect 11729 2959 11788 2979
rect 11639 2952 11788 2959
rect 12432 2972 12471 2997
rect 12817 2972 12869 3161
rect 13261 3189 13271 3207
rect 13289 3189 13301 3207
rect 13433 3205 13442 3225
rect 13462 3205 13471 3225
rect 13433 3197 13471 3205
rect 13537 3229 13622 3235
rect 13652 3234 13689 3235
rect 13537 3209 13545 3229
rect 13565 3209 13622 3229
rect 13537 3201 13622 3209
rect 13651 3225 13689 3234
rect 13651 3205 13660 3225
rect 13680 3205 13689 3225
rect 13537 3200 13573 3201
rect 13651 3197 13689 3205
rect 13755 3229 13899 3235
rect 13755 3209 13763 3229
rect 13783 3209 13816 3229
rect 13836 3209 13871 3229
rect 13891 3209 13899 3229
rect 13755 3201 13899 3209
rect 13755 3200 13791 3201
rect 13863 3200 13899 3201
rect 13965 3234 14002 3235
rect 13965 3233 14003 3234
rect 13965 3225 14029 3233
rect 13965 3205 13974 3225
rect 13994 3211 14029 3225
rect 14049 3211 14052 3231
rect 13994 3206 14052 3211
rect 13994 3205 14029 3206
rect 13261 3133 13301 3189
rect 13434 3168 13471 3197
rect 13435 3166 13471 3168
rect 13435 3144 13626 3166
rect 13652 3165 13689 3197
rect 13965 3193 14029 3205
rect 14069 3167 14096 3345
rect 14954 3320 14996 3365
rect 13928 3165 14096 3167
rect 13652 3155 14096 3165
rect 14237 3261 14424 3285
rect 14455 3266 14848 3286
rect 14868 3266 14871 3286
rect 14455 3261 14871 3266
rect 14237 3190 14274 3261
rect 14455 3260 14796 3261
rect 14389 3200 14420 3201
rect 14237 3170 14246 3190
rect 14266 3170 14274 3190
rect 14237 3160 14274 3170
rect 14333 3190 14420 3200
rect 14333 3170 14342 3190
rect 14362 3170 14420 3190
rect 14333 3161 14420 3170
rect 14333 3160 14370 3161
rect 13258 3128 13301 3133
rect 13649 3139 14096 3155
rect 13649 3133 13677 3139
rect 13928 3138 14096 3139
rect 13258 3125 13408 3128
rect 13649 3125 13676 3133
rect 13258 3123 13676 3125
rect 13258 3105 13267 3123
rect 13285 3105 13676 3123
rect 14389 3110 14420 3161
rect 14455 3190 14492 3260
rect 14758 3259 14795 3260
rect 14607 3200 14643 3201
rect 14455 3170 14464 3190
rect 14484 3170 14492 3190
rect 14455 3160 14492 3170
rect 14551 3190 14699 3200
rect 14799 3197 14895 3199
rect 14551 3170 14560 3190
rect 14580 3170 14670 3190
rect 14690 3170 14699 3190
rect 14551 3161 14699 3170
rect 14757 3190 14895 3197
rect 14757 3170 14766 3190
rect 14786 3170 14895 3190
rect 14757 3161 14895 3170
rect 14551 3160 14588 3161
rect 14281 3107 14322 3108
rect 13258 3102 13676 3105
rect 13258 3096 13301 3102
rect 13261 3093 13301 3096
rect 14176 3100 14322 3107
rect 13658 3084 13698 3085
rect 13369 3067 13698 3084
rect 14176 3080 14232 3100
rect 14252 3080 14291 3100
rect 14311 3080 14322 3100
rect 14176 3072 14322 3080
rect 14389 3103 14546 3110
rect 14389 3083 14509 3103
rect 14529 3083 14546 3103
rect 14389 3073 14546 3083
rect 14389 3072 14424 3073
rect 13253 3024 13296 3035
rect 13253 3006 13265 3024
rect 13283 3006 13296 3024
rect 13253 2980 13296 3006
rect 13369 2980 13396 3067
rect 13658 3058 13698 3067
rect 12432 2954 12871 2972
rect 11639 2951 11680 2952
rect 11373 2898 11410 2899
rect 11066 2889 11204 2898
rect 11066 2869 11175 2889
rect 11195 2869 11204 2889
rect 11066 2862 11204 2869
rect 11262 2889 11410 2898
rect 11262 2869 11271 2889
rect 11291 2869 11381 2889
rect 11401 2869 11410 2889
rect 11066 2860 11162 2862
rect 11262 2859 11410 2869
rect 11469 2889 11506 2899
rect 11469 2869 11477 2889
rect 11497 2869 11506 2889
rect 11318 2858 11354 2859
rect 11166 2799 11203 2800
rect 11469 2799 11506 2869
rect 11541 2898 11572 2949
rect 12432 2936 12832 2954
rect 12850 2936 12871 2954
rect 12432 2930 12871 2936
rect 12438 2926 12871 2930
rect 13253 2959 13396 2980
rect 13440 3032 13474 3048
rect 13658 3038 14051 3058
rect 14071 3038 14074 3058
rect 14389 3051 14420 3072
rect 14607 3051 14643 3161
rect 14662 3160 14699 3161
rect 14758 3160 14795 3161
rect 14718 3101 14808 3107
rect 14718 3081 14727 3101
rect 14747 3099 14808 3101
rect 14747 3081 14772 3099
rect 14718 3079 14772 3081
rect 14792 3079 14808 3099
rect 14718 3073 14808 3079
rect 14232 3050 14269 3051
rect 13658 3033 14074 3038
rect 14231 3041 14269 3050
rect 13658 3032 13999 3033
rect 13440 2962 13477 3032
rect 13592 2972 13623 2973
rect 13253 2957 13390 2959
rect 12817 2924 12869 2926
rect 13253 2915 13296 2957
rect 13440 2942 13449 2962
rect 13469 2942 13477 2962
rect 13440 2932 13477 2942
rect 13536 2962 13623 2972
rect 13536 2942 13545 2962
rect 13565 2942 13623 2962
rect 13536 2933 13623 2942
rect 13536 2932 13573 2933
rect 13251 2905 13296 2915
rect 11591 2898 11628 2899
rect 11541 2889 11628 2898
rect 11541 2869 11599 2889
rect 11619 2869 11628 2889
rect 11541 2859 11628 2869
rect 11687 2889 11724 2899
rect 11687 2869 11695 2889
rect 11715 2869 11724 2889
rect 13251 2887 13260 2905
rect 13278 2887 13296 2905
rect 13251 2881 13296 2887
rect 13592 2882 13623 2933
rect 13658 2962 13695 3032
rect 13961 3031 13998 3032
rect 14231 3021 14240 3041
rect 14260 3021 14269 3041
rect 14231 3013 14269 3021
rect 14335 3045 14420 3051
rect 14450 3050 14487 3051
rect 14335 3025 14343 3045
rect 14363 3025 14420 3045
rect 14335 3017 14420 3025
rect 14449 3041 14487 3050
rect 14449 3021 14458 3041
rect 14478 3021 14487 3041
rect 14335 3016 14371 3017
rect 14449 3013 14487 3021
rect 14553 3045 14697 3051
rect 14553 3025 14561 3045
rect 14581 3042 14669 3045
rect 14581 3025 14616 3042
rect 14553 3024 14616 3025
rect 14635 3025 14669 3042
rect 14689 3025 14697 3045
rect 14635 3024 14697 3025
rect 14553 3017 14697 3024
rect 14553 3016 14589 3017
rect 14661 3016 14697 3017
rect 14763 3050 14800 3051
rect 14763 3049 14801 3050
rect 14823 3049 14850 3053
rect 14763 3047 14850 3049
rect 14763 3041 14827 3047
rect 14763 3021 14772 3041
rect 14792 3027 14827 3041
rect 14847 3027 14850 3047
rect 14792 3022 14850 3027
rect 14792 3021 14827 3022
rect 14232 2984 14269 3013
rect 14233 2982 14269 2984
rect 13810 2972 13846 2973
rect 13658 2942 13667 2962
rect 13687 2942 13695 2962
rect 13658 2932 13695 2942
rect 13754 2962 13902 2972
rect 14002 2969 14098 2971
rect 13754 2942 13763 2962
rect 13783 2942 13873 2962
rect 13893 2942 13902 2962
rect 13754 2933 13902 2942
rect 13960 2962 14098 2969
rect 13960 2942 13969 2962
rect 13989 2942 14098 2962
rect 14233 2960 14424 2982
rect 14450 2981 14487 3013
rect 14763 3009 14827 3021
rect 14867 2983 14894 3161
rect 14726 2981 14894 2983
rect 14450 2955 14894 2981
rect 13960 2933 14098 2942
rect 13754 2932 13791 2933
rect 13251 2878 13288 2881
rect 13484 2879 13525 2880
rect 11541 2858 11572 2859
rect 11165 2798 11506 2799
rect 11687 2798 11724 2869
rect 13376 2872 13525 2879
rect 12820 2859 12857 2864
rect 11090 2793 11506 2798
rect 11090 2773 11093 2793
rect 11113 2773 11506 2793
rect 11537 2774 11724 2798
rect 12811 2855 12858 2859
rect 12811 2837 12830 2855
rect 12848 2837 12858 2855
rect 13376 2852 13435 2872
rect 13455 2852 13494 2872
rect 13514 2852 13525 2872
rect 13376 2844 13525 2852
rect 13592 2875 13749 2882
rect 13592 2855 13712 2875
rect 13732 2855 13749 2875
rect 13592 2845 13749 2855
rect 13592 2844 13627 2845
rect 12811 2789 12858 2837
rect 13592 2823 13623 2844
rect 13810 2823 13846 2933
rect 13865 2932 13902 2933
rect 13961 2932 13998 2933
rect 13921 2873 14011 2879
rect 13921 2853 13930 2873
rect 13950 2871 14011 2873
rect 13950 2853 13975 2871
rect 13921 2851 13975 2853
rect 13995 2851 14011 2871
rect 13921 2845 14011 2851
rect 13435 2822 13472 2823
rect 12435 2786 12858 2789
rect 11310 2772 11375 2773
rect 12413 2756 12858 2786
rect 13247 2814 13285 2816
rect 13247 2806 13290 2814
rect 13247 2788 13258 2806
rect 13276 2788 13290 2806
rect 13247 2761 13290 2788
rect 13434 2813 13472 2822
rect 13434 2793 13443 2813
rect 13463 2793 13472 2813
rect 13434 2785 13472 2793
rect 13538 2817 13623 2823
rect 13653 2822 13690 2823
rect 13538 2797 13546 2817
rect 13566 2797 13623 2817
rect 13538 2789 13623 2797
rect 13652 2813 13690 2822
rect 13652 2793 13661 2813
rect 13681 2793 13690 2813
rect 13538 2788 13574 2789
rect 13652 2785 13690 2793
rect 13756 2821 13900 2823
rect 13756 2817 13808 2821
rect 13756 2797 13764 2817
rect 13784 2801 13808 2817
rect 13828 2817 13900 2821
rect 13828 2801 13872 2817
rect 13784 2797 13872 2801
rect 13892 2797 13900 2817
rect 13756 2789 13900 2797
rect 13756 2788 13792 2789
rect 13864 2788 13900 2789
rect 13966 2822 14003 2823
rect 13966 2821 14004 2822
rect 13966 2813 14030 2821
rect 13966 2793 13975 2813
rect 13995 2799 14030 2813
rect 14050 2799 14053 2819
rect 13995 2794 14053 2799
rect 13995 2793 14030 2794
rect 11506 2740 11546 2748
rect 11506 2718 11514 2740
rect 11538 2718 11546 2740
rect 11111 2489 11148 2495
rect 11111 2470 11119 2489
rect 11140 2470 11148 2489
rect 11111 2462 11148 2470
rect 10811 2341 10818 2363
rect 10842 2341 10850 2363
rect 10811 2335 10850 2341
rect 10341 2330 10381 2332
rect 10507 2331 10675 2332
rect 10609 2330 10646 2331
rect 9575 2314 9713 2323
rect 9369 2313 9406 2314
rect 9099 2260 9140 2261
rect 8873 2239 8925 2257
rect 8991 2253 9140 2260
rect 8428 2220 8468 2230
rect 8991 2233 9050 2253
rect 9070 2233 9109 2253
rect 9129 2233 9140 2253
rect 8991 2225 9140 2233
rect 9207 2256 9364 2263
rect 9207 2236 9327 2256
rect 9347 2236 9364 2256
rect 9207 2226 9364 2236
rect 9207 2225 9242 2226
rect 8258 2203 8296 2212
rect 9207 2204 9238 2225
rect 9425 2204 9461 2314
rect 9480 2313 9517 2314
rect 9576 2313 9613 2314
rect 9536 2254 9626 2260
rect 9536 2234 9545 2254
rect 9565 2252 9626 2254
rect 9565 2234 9590 2252
rect 9536 2232 9590 2234
rect 9610 2232 9626 2252
rect 9536 2226 9626 2232
rect 9050 2203 9087 2204
rect 8258 2202 8295 2203
rect 7719 2174 7809 2180
rect 7719 2154 7735 2174
rect 7755 2172 7809 2174
rect 7755 2154 7780 2172
rect 7719 2152 7780 2154
rect 7800 2152 7809 2172
rect 7719 2146 7809 2152
rect 7732 2092 7769 2093
rect 7828 2092 7865 2093
rect 7884 2092 7920 2202
rect 8107 2181 8138 2202
rect 9049 2194 9087 2203
rect 8103 2180 8138 2181
rect 7981 2170 8138 2180
rect 7981 2150 7998 2170
rect 8018 2150 8138 2170
rect 7981 2143 8138 2150
rect 8205 2173 8354 2181
rect 8205 2153 8216 2173
rect 8236 2153 8275 2173
rect 8295 2153 8354 2173
rect 8877 2176 8917 2186
rect 8205 2146 8354 2153
rect 8420 2149 8472 2167
rect 8205 2145 8246 2146
rect 7939 2092 7976 2093
rect 7632 2083 7770 2092
rect 7104 2072 7137 2074
rect 6733 2060 7180 2072
rect 5965 1938 6133 1940
rect 5689 1912 6133 1938
rect 5199 1890 5337 1899
rect 4993 1889 5030 1890
rect 4490 1835 4527 1838
rect 4723 1836 4764 1837
rect 2846 1813 2877 1814
rect 2470 1753 2811 1754
rect 2992 1753 3029 1824
rect 4615 1829 4764 1836
rect 4059 1816 4096 1821
rect 4050 1812 4097 1816
rect 4050 1794 4069 1812
rect 4087 1794 4097 1812
rect 4615 1809 4674 1829
rect 4694 1809 4733 1829
rect 4753 1809 4764 1829
rect 4615 1801 4764 1809
rect 4831 1832 4988 1839
rect 4831 1812 4951 1832
rect 4971 1812 4988 1832
rect 4831 1802 4988 1812
rect 4831 1801 4866 1802
rect 2395 1748 2811 1753
rect 2395 1728 2398 1748
rect 2418 1728 2811 1748
rect 2842 1729 3029 1753
rect 3654 1751 3694 1756
rect 4050 1751 4097 1794
rect 4831 1780 4862 1801
rect 5049 1780 5085 1890
rect 5104 1889 5141 1890
rect 5200 1889 5237 1890
rect 5160 1830 5250 1836
rect 5160 1810 5169 1830
rect 5189 1828 5250 1830
rect 5189 1810 5214 1828
rect 5160 1808 5214 1810
rect 5234 1808 5250 1828
rect 5160 1802 5250 1808
rect 4674 1779 4711 1780
rect 3654 1712 4097 1751
rect 4487 1771 4524 1773
rect 4487 1763 4529 1771
rect 4487 1745 4497 1763
rect 4515 1745 4529 1763
rect 4487 1736 4529 1745
rect 4673 1770 4711 1779
rect 4673 1750 4682 1770
rect 4702 1750 4711 1770
rect 4673 1742 4711 1750
rect 4777 1774 4862 1780
rect 4892 1779 4929 1780
rect 4777 1754 4785 1774
rect 4805 1754 4862 1774
rect 4777 1746 4862 1754
rect 4891 1770 4929 1779
rect 4891 1750 4900 1770
rect 4920 1750 4929 1770
rect 4777 1745 4813 1746
rect 4891 1742 4929 1750
rect 4995 1778 5139 1780
rect 4995 1774 5047 1778
rect 4995 1754 5003 1774
rect 5023 1758 5047 1774
rect 5067 1774 5139 1778
rect 5067 1758 5111 1774
rect 5023 1754 5111 1758
rect 5131 1754 5139 1774
rect 4995 1746 5139 1754
rect 4995 1745 5031 1746
rect 5103 1745 5139 1746
rect 5205 1779 5242 1780
rect 5205 1778 5243 1779
rect 5205 1770 5269 1778
rect 5205 1750 5214 1770
rect 5234 1756 5269 1770
rect 5289 1756 5292 1776
rect 5234 1751 5292 1756
rect 5234 1750 5269 1751
rect 1435 1653 1443 1675
rect 1467 1653 1475 1675
rect 1435 1645 1475 1653
rect 2748 1697 2788 1705
rect 2748 1675 2756 1697
rect 2780 1675 2788 1697
rect 126 1599 569 1638
rect 126 1556 173 1599
rect 529 1594 569 1599
rect 1194 1597 1381 1621
rect 1412 1602 1805 1622
rect 1825 1602 1828 1622
rect 1412 1597 1828 1602
rect 126 1538 136 1556
rect 154 1538 173 1556
rect 126 1534 173 1538
rect 127 1529 164 1534
rect 1194 1526 1231 1597
rect 1412 1596 1753 1597
rect 1346 1536 1377 1537
rect 1194 1506 1203 1526
rect 1223 1506 1231 1526
rect 1194 1496 1231 1506
rect 1290 1526 1377 1536
rect 1290 1506 1299 1526
rect 1319 1506 1377 1526
rect 1290 1497 1377 1506
rect 1290 1496 1327 1497
rect 115 1467 167 1469
rect 113 1463 546 1467
rect 113 1457 552 1463
rect 113 1439 134 1457
rect 152 1439 552 1457
rect 1346 1446 1377 1497
rect 1412 1526 1449 1596
rect 1715 1595 1752 1596
rect 1564 1536 1600 1537
rect 1412 1506 1421 1526
rect 1441 1506 1449 1526
rect 1412 1496 1449 1506
rect 1508 1526 1656 1536
rect 1756 1533 1852 1535
rect 1508 1506 1517 1526
rect 1537 1506 1627 1526
rect 1647 1506 1656 1526
rect 1508 1497 1656 1506
rect 1714 1526 1852 1533
rect 1714 1506 1723 1526
rect 1743 1506 1852 1526
rect 1714 1497 1852 1506
rect 1508 1496 1545 1497
rect 1238 1443 1279 1444
rect 113 1421 552 1439
rect 115 1232 167 1421
rect 513 1396 552 1421
rect 1130 1436 1279 1443
rect 1130 1416 1189 1436
rect 1209 1416 1248 1436
rect 1268 1416 1279 1436
rect 1130 1408 1279 1416
rect 1346 1439 1503 1446
rect 1346 1419 1466 1439
rect 1486 1419 1503 1439
rect 1346 1409 1503 1419
rect 1346 1408 1381 1409
rect 297 1371 484 1395
rect 513 1376 908 1396
rect 928 1376 931 1396
rect 1346 1387 1377 1408
rect 1564 1387 1600 1497
rect 1619 1496 1656 1497
rect 1715 1496 1752 1497
rect 1675 1437 1765 1443
rect 1675 1417 1684 1437
rect 1704 1435 1765 1437
rect 1704 1417 1729 1435
rect 1675 1415 1729 1417
rect 1749 1415 1765 1435
rect 1675 1409 1765 1415
rect 1189 1386 1226 1387
rect 513 1371 931 1376
rect 1188 1377 1226 1386
rect 297 1300 334 1371
rect 513 1370 856 1371
rect 513 1367 552 1370
rect 818 1369 855 1370
rect 449 1310 480 1311
rect 297 1280 306 1300
rect 326 1280 334 1300
rect 297 1270 334 1280
rect 393 1300 480 1310
rect 393 1280 402 1300
rect 422 1280 480 1300
rect 393 1271 480 1280
rect 393 1270 430 1271
rect 115 1214 131 1232
rect 149 1214 167 1232
rect 449 1220 480 1271
rect 515 1300 552 1367
rect 1188 1357 1197 1377
rect 1217 1357 1226 1377
rect 1188 1349 1226 1357
rect 1292 1381 1377 1387
rect 1407 1386 1444 1387
rect 1292 1361 1300 1381
rect 1320 1361 1377 1381
rect 1292 1353 1377 1361
rect 1406 1377 1444 1386
rect 1406 1357 1415 1377
rect 1435 1357 1444 1377
rect 1292 1352 1328 1353
rect 1406 1349 1444 1357
rect 1510 1381 1654 1387
rect 1510 1361 1518 1381
rect 1538 1376 1626 1381
rect 1538 1361 1574 1376
rect 1510 1359 1574 1361
rect 1593 1361 1626 1376
rect 1646 1361 1654 1381
rect 1593 1359 1654 1361
rect 1510 1353 1654 1359
rect 1510 1352 1546 1353
rect 1618 1352 1654 1353
rect 1720 1386 1757 1387
rect 1720 1385 1758 1386
rect 1720 1377 1784 1385
rect 1720 1357 1729 1377
rect 1749 1363 1784 1377
rect 1804 1363 1807 1383
rect 1749 1358 1807 1363
rect 1749 1357 1784 1358
rect 1189 1320 1226 1349
rect 1190 1318 1226 1320
rect 667 1310 703 1311
rect 515 1280 524 1300
rect 544 1280 552 1300
rect 515 1270 552 1280
rect 611 1300 759 1310
rect 859 1307 955 1309
rect 611 1280 620 1300
rect 640 1280 730 1300
rect 750 1280 759 1300
rect 611 1271 759 1280
rect 817 1300 955 1307
rect 817 1280 826 1300
rect 846 1280 955 1300
rect 1190 1296 1381 1318
rect 1407 1317 1444 1349
rect 1720 1345 1784 1357
rect 1824 1319 1851 1497
rect 1683 1317 1851 1319
rect 1407 1303 1851 1317
rect 2454 1451 2622 1452
rect 2748 1451 2788 1675
rect 3251 1679 3419 1680
rect 3654 1679 3694 1712
rect 4050 1679 4097 1712
rect 4488 1711 4529 1736
rect 4674 1711 4711 1742
rect 4892 1711 4929 1742
rect 5205 1738 5269 1750
rect 5309 1712 5336 1890
rect 4488 1684 4537 1711
rect 4673 1685 4722 1711
rect 4891 1710 4972 1711
rect 5168 1710 5336 1712
rect 4891 1685 5336 1710
rect 4892 1684 5336 1685
rect 3251 1678 3695 1679
rect 3251 1653 3696 1678
rect 3251 1651 3419 1653
rect 3615 1652 3696 1653
rect 3865 1652 3914 1678
rect 4050 1652 4099 1679
rect 3251 1473 3278 1651
rect 3318 1613 3382 1625
rect 3658 1621 3695 1652
rect 3876 1621 3913 1652
rect 4058 1627 4099 1652
rect 4490 1651 4537 1684
rect 4893 1651 4933 1684
rect 5168 1683 5336 1684
rect 5799 1688 5839 1912
rect 5965 1911 6133 1912
rect 6736 2046 7180 2060
rect 6736 2044 6904 2046
rect 6736 1866 6763 2044
rect 6803 2006 6867 2018
rect 7143 2014 7180 2046
rect 7206 2045 7397 2067
rect 7632 2063 7741 2083
rect 7761 2063 7770 2083
rect 7632 2056 7770 2063
rect 7828 2083 7976 2092
rect 7828 2063 7837 2083
rect 7857 2063 7947 2083
rect 7967 2063 7976 2083
rect 7632 2054 7728 2056
rect 7828 2053 7976 2063
rect 8035 2083 8072 2093
rect 8035 2063 8043 2083
rect 8063 2063 8072 2083
rect 7884 2052 7920 2053
rect 7361 2043 7397 2045
rect 7361 2014 7398 2043
rect 6803 2005 6838 2006
rect 6780 2000 6838 2005
rect 6780 1980 6783 2000
rect 6803 1986 6838 2000
rect 6858 1986 6867 2006
rect 6803 1978 6867 1986
rect 6829 1977 6867 1978
rect 6830 1976 6867 1977
rect 6933 2010 6969 2011
rect 7041 2010 7077 2011
rect 6933 2002 7077 2010
rect 6933 1982 6941 2002
rect 6961 2000 7049 2002
rect 6961 1982 6994 2000
rect 6933 1981 6994 1982
rect 7015 1982 7049 2000
rect 7069 1982 7077 2002
rect 7015 1981 7077 1982
rect 6933 1976 7077 1981
rect 7143 2006 7181 2014
rect 7259 2010 7295 2011
rect 7143 1986 7152 2006
rect 7172 1986 7181 2006
rect 7143 1977 7181 1986
rect 7210 2002 7295 2010
rect 7210 1982 7267 2002
rect 7287 1982 7295 2002
rect 7143 1976 7180 1977
rect 7210 1976 7295 1982
rect 7361 2006 7399 2014
rect 7361 1986 7370 2006
rect 7390 1986 7399 2006
rect 8035 1996 8072 2063
rect 8107 2092 8138 2143
rect 8420 2131 8438 2149
rect 8456 2131 8472 2149
rect 8157 2092 8194 2093
rect 8107 2083 8194 2092
rect 8107 2063 8165 2083
rect 8185 2063 8194 2083
rect 8107 2053 8194 2063
rect 8253 2083 8290 2093
rect 8253 2063 8261 2083
rect 8281 2063 8290 2083
rect 8107 2052 8138 2053
rect 7732 1993 7769 1994
rect 8035 1993 8074 1996
rect 7731 1992 8074 1993
rect 8253 1992 8290 2063
rect 7361 1977 7399 1986
rect 7656 1987 8074 1992
rect 7361 1976 7398 1977
rect 6822 1948 6912 1954
rect 6822 1928 6838 1948
rect 6858 1946 6912 1948
rect 6858 1928 6883 1946
rect 6822 1926 6883 1928
rect 6903 1926 6912 1946
rect 6822 1920 6912 1926
rect 6835 1866 6872 1867
rect 6931 1866 6968 1867
rect 6987 1866 7023 1976
rect 7210 1955 7241 1976
rect 7656 1967 7659 1987
rect 7679 1967 8074 1987
rect 8103 1968 8290 1992
rect 7206 1954 7241 1955
rect 7084 1944 7241 1954
rect 7084 1924 7101 1944
rect 7121 1924 7241 1944
rect 7084 1917 7241 1924
rect 7308 1947 7457 1955
rect 7308 1927 7319 1947
rect 7339 1927 7378 1947
rect 7398 1927 7457 1947
rect 7308 1920 7457 1927
rect 8035 1942 8074 1967
rect 8420 1942 8472 2131
rect 8877 2158 8887 2176
rect 8905 2158 8917 2176
rect 9049 2174 9058 2194
rect 9078 2174 9087 2194
rect 9049 2166 9087 2174
rect 9153 2198 9238 2204
rect 9268 2203 9305 2204
rect 9153 2178 9161 2198
rect 9181 2178 9238 2198
rect 9153 2170 9238 2178
rect 9267 2194 9305 2203
rect 9267 2174 9276 2194
rect 9296 2174 9305 2194
rect 9153 2169 9189 2170
rect 9267 2166 9305 2174
rect 9371 2198 9515 2204
rect 9371 2178 9379 2198
rect 9399 2178 9432 2198
rect 9452 2178 9487 2198
rect 9507 2178 9515 2198
rect 9371 2170 9515 2178
rect 9371 2169 9407 2170
rect 9479 2169 9515 2170
rect 9581 2203 9618 2204
rect 9581 2202 9619 2203
rect 9581 2194 9645 2202
rect 9581 2174 9590 2194
rect 9610 2180 9645 2194
rect 9665 2180 9668 2200
rect 9610 2175 9668 2180
rect 9610 2174 9645 2175
rect 8877 2102 8917 2158
rect 9050 2137 9087 2166
rect 9051 2135 9087 2137
rect 9051 2113 9242 2135
rect 9268 2134 9305 2166
rect 9581 2162 9645 2174
rect 9685 2136 9712 2314
rect 9544 2134 9712 2136
rect 9268 2124 9712 2134
rect 9853 2230 10040 2254
rect 10071 2235 10464 2255
rect 10484 2235 10487 2255
rect 10071 2230 10487 2235
rect 9853 2159 9890 2230
rect 10071 2229 10412 2230
rect 10005 2169 10036 2170
rect 9853 2139 9862 2159
rect 9882 2139 9890 2159
rect 9853 2129 9890 2139
rect 9949 2159 10036 2169
rect 9949 2139 9958 2159
rect 9978 2139 10036 2159
rect 9949 2130 10036 2139
rect 9949 2129 9986 2130
rect 8874 2097 8917 2102
rect 9265 2108 9712 2124
rect 9265 2102 9293 2108
rect 9544 2107 9712 2108
rect 8874 2094 9024 2097
rect 9265 2094 9292 2102
rect 8874 2092 9292 2094
rect 8874 2074 8883 2092
rect 8901 2074 9292 2092
rect 10005 2079 10036 2130
rect 10071 2159 10108 2229
rect 10374 2228 10411 2229
rect 10612 2171 10645 2330
rect 10223 2169 10259 2170
rect 10071 2139 10080 2159
rect 10100 2139 10108 2159
rect 10071 2129 10108 2139
rect 10167 2159 10315 2169
rect 10415 2166 10511 2168
rect 10167 2139 10176 2159
rect 10196 2139 10286 2159
rect 10306 2139 10315 2159
rect 10167 2130 10315 2139
rect 10373 2159 10511 2166
rect 10373 2139 10382 2159
rect 10402 2139 10511 2159
rect 10612 2167 10648 2171
rect 10612 2149 10621 2167
rect 10643 2149 10648 2167
rect 10612 2143 10648 2149
rect 10373 2130 10511 2139
rect 10167 2129 10204 2130
rect 9897 2076 9938 2077
rect 8874 2071 9292 2074
rect 8874 2065 8917 2071
rect 8877 2062 8917 2065
rect 9789 2069 9938 2076
rect 9274 2053 9314 2054
rect 8985 2036 9314 2053
rect 9789 2049 9848 2069
rect 9868 2049 9907 2069
rect 9927 2049 9938 2069
rect 9789 2041 9938 2049
rect 10005 2072 10162 2079
rect 10005 2052 10125 2072
rect 10145 2052 10162 2072
rect 10005 2042 10162 2052
rect 10005 2041 10040 2042
rect 8869 1993 8912 2004
rect 8869 1975 8881 1993
rect 8899 1975 8912 1993
rect 8869 1949 8912 1975
rect 8985 1949 9012 2036
rect 9274 2027 9314 2036
rect 8035 1924 8474 1942
rect 7308 1919 7349 1920
rect 7042 1866 7079 1867
rect 6735 1857 6873 1866
rect 6735 1837 6844 1857
rect 6864 1837 6873 1857
rect 6735 1830 6873 1837
rect 6931 1857 7079 1866
rect 6931 1837 6940 1857
rect 6960 1837 7050 1857
rect 7070 1837 7079 1857
rect 6735 1828 6831 1830
rect 6931 1827 7079 1837
rect 7138 1857 7175 1867
rect 7138 1837 7146 1857
rect 7166 1837 7175 1857
rect 6987 1826 7023 1827
rect 6835 1767 6872 1768
rect 7138 1767 7175 1837
rect 7210 1866 7241 1917
rect 8035 1906 8435 1924
rect 8453 1906 8474 1924
rect 8035 1900 8474 1906
rect 8041 1896 8474 1900
rect 8869 1928 9012 1949
rect 9056 2001 9090 2017
rect 9274 2007 9667 2027
rect 9687 2007 9690 2027
rect 10005 2020 10036 2041
rect 10223 2020 10259 2130
rect 10278 2129 10315 2130
rect 10374 2129 10411 2130
rect 10334 2070 10424 2076
rect 10334 2050 10343 2070
rect 10363 2068 10424 2070
rect 10363 2050 10388 2068
rect 10334 2048 10388 2050
rect 10408 2048 10424 2068
rect 10334 2042 10424 2048
rect 9848 2019 9885 2020
rect 9274 2002 9690 2007
rect 9847 2010 9885 2019
rect 9274 2001 9615 2002
rect 9056 1931 9093 2001
rect 9208 1941 9239 1942
rect 8869 1926 9006 1928
rect 8420 1894 8472 1896
rect 8869 1884 8912 1926
rect 9056 1911 9065 1931
rect 9085 1911 9093 1931
rect 9056 1901 9093 1911
rect 9152 1931 9239 1941
rect 9152 1911 9161 1931
rect 9181 1911 9239 1931
rect 9152 1902 9239 1911
rect 9152 1901 9189 1902
rect 8867 1874 8912 1884
rect 7260 1866 7297 1867
rect 7210 1857 7297 1866
rect 7210 1837 7268 1857
rect 7288 1837 7297 1857
rect 7210 1827 7297 1837
rect 7356 1857 7393 1867
rect 7356 1837 7364 1857
rect 7384 1837 7393 1857
rect 8867 1856 8876 1874
rect 8894 1856 8912 1874
rect 8867 1850 8912 1856
rect 9208 1851 9239 1902
rect 9274 1931 9311 2001
rect 9577 2000 9614 2001
rect 9847 1990 9856 2010
rect 9876 1990 9885 2010
rect 9847 1982 9885 1990
rect 9951 2014 10036 2020
rect 10066 2019 10103 2020
rect 9951 1994 9959 2014
rect 9979 1994 10036 2014
rect 9951 1986 10036 1994
rect 10065 2010 10103 2019
rect 10065 1990 10074 2010
rect 10094 1990 10103 2010
rect 9951 1985 9987 1986
rect 10065 1982 10103 1990
rect 10169 2014 10313 2020
rect 10169 1994 10177 2014
rect 10197 1995 10229 2014
rect 10250 1995 10285 2014
rect 10197 1994 10285 1995
rect 10305 1994 10313 2014
rect 10169 1986 10313 1994
rect 10169 1985 10205 1986
rect 10277 1985 10313 1986
rect 10379 2019 10416 2020
rect 10379 2018 10417 2019
rect 10379 2010 10443 2018
rect 10379 1990 10388 2010
rect 10408 1996 10443 2010
rect 10463 1996 10466 2016
rect 10408 1991 10466 1996
rect 10408 1990 10443 1991
rect 9848 1953 9885 1982
rect 9849 1951 9885 1953
rect 9426 1941 9462 1942
rect 9274 1911 9283 1931
rect 9303 1911 9311 1931
rect 9274 1901 9311 1911
rect 9370 1931 9518 1941
rect 9618 1938 9714 1940
rect 9370 1911 9379 1931
rect 9399 1911 9489 1931
rect 9509 1911 9518 1931
rect 9370 1902 9518 1911
rect 9576 1931 9714 1938
rect 9576 1911 9585 1931
rect 9605 1911 9714 1931
rect 9849 1929 10040 1951
rect 10066 1950 10103 1982
rect 10379 1978 10443 1990
rect 10483 1952 10510 2130
rect 11115 2129 11148 2462
rect 11212 2494 11380 2495
rect 11506 2494 11546 2718
rect 12009 2722 12177 2723
rect 12413 2722 12454 2756
rect 12811 2735 12858 2756
rect 12009 2712 12454 2722
rect 12526 2720 12669 2721
rect 12009 2696 12453 2712
rect 12009 2694 12177 2696
rect 12373 2695 12453 2696
rect 12526 2695 12671 2720
rect 12813 2695 12858 2735
rect 12009 2516 12036 2694
rect 12076 2656 12140 2668
rect 12416 2664 12453 2695
rect 12634 2664 12671 2695
rect 12816 2688 12858 2695
rect 13248 2754 13290 2761
rect 13435 2754 13472 2785
rect 13653 2754 13690 2785
rect 13966 2781 14030 2793
rect 14070 2755 14097 2933
rect 13248 2714 13293 2754
rect 13435 2729 13580 2754
rect 13653 2753 13733 2754
rect 13929 2753 14097 2755
rect 13653 2737 14097 2753
rect 13437 2728 13580 2729
rect 13652 2727 14097 2737
rect 13248 2693 13295 2714
rect 13652 2693 13693 2727
rect 13929 2726 14097 2727
rect 14560 2731 14600 2955
rect 14726 2954 14894 2955
rect 14958 2987 14991 3320
rect 14958 2979 14995 2987
rect 14958 2960 14966 2979
rect 14987 2960 14995 2979
rect 14958 2954 14995 2960
rect 14560 2709 14568 2731
rect 14592 2709 14600 2731
rect 14560 2701 14600 2709
rect 12076 2655 12111 2656
rect 12053 2650 12111 2655
rect 12053 2630 12056 2650
rect 12076 2636 12111 2650
rect 12131 2636 12140 2656
rect 12076 2628 12140 2636
rect 12102 2627 12140 2628
rect 12103 2626 12140 2627
rect 12206 2660 12242 2661
rect 12314 2660 12350 2661
rect 12206 2652 12350 2660
rect 12206 2632 12214 2652
rect 12234 2648 12322 2652
rect 12234 2632 12278 2648
rect 12206 2628 12278 2632
rect 12298 2632 12322 2648
rect 12342 2632 12350 2652
rect 12298 2628 12350 2632
rect 12206 2626 12350 2628
rect 12416 2656 12454 2664
rect 12532 2660 12568 2661
rect 12416 2636 12425 2656
rect 12445 2636 12454 2656
rect 12416 2627 12454 2636
rect 12483 2652 12568 2660
rect 12483 2632 12540 2652
rect 12560 2632 12568 2652
rect 12416 2626 12453 2627
rect 12483 2626 12568 2632
rect 12634 2656 12672 2664
rect 12634 2636 12643 2656
rect 12663 2636 12672 2656
rect 12634 2627 12672 2636
rect 12816 2661 12859 2688
rect 12816 2643 12830 2661
rect 12848 2643 12859 2661
rect 12816 2635 12859 2643
rect 12821 2633 12859 2635
rect 13248 2663 13693 2693
rect 14731 2676 14796 2677
rect 13248 2660 13671 2663
rect 12634 2626 12671 2627
rect 12095 2598 12185 2604
rect 12095 2578 12111 2598
rect 12131 2596 12185 2598
rect 12131 2578 12156 2596
rect 12095 2576 12156 2578
rect 12176 2576 12185 2596
rect 12095 2570 12185 2576
rect 12108 2516 12145 2517
rect 12204 2516 12241 2517
rect 12260 2516 12296 2626
rect 12483 2605 12514 2626
rect 13248 2612 13295 2660
rect 12479 2604 12514 2605
rect 12357 2594 12514 2604
rect 12357 2574 12374 2594
rect 12394 2574 12514 2594
rect 12357 2567 12514 2574
rect 12581 2597 12730 2605
rect 12581 2577 12592 2597
rect 12612 2577 12651 2597
rect 12671 2577 12730 2597
rect 13248 2594 13258 2612
rect 13276 2594 13295 2612
rect 13248 2590 13295 2594
rect 14382 2651 14569 2675
rect 14600 2656 14993 2676
rect 15013 2656 15016 2676
rect 14600 2651 15016 2656
rect 13249 2585 13286 2590
rect 12581 2570 12730 2577
rect 14382 2580 14419 2651
rect 14600 2650 14941 2651
rect 14534 2590 14565 2591
rect 12581 2569 12622 2570
rect 12818 2568 12855 2571
rect 12315 2516 12352 2517
rect 12008 2507 12146 2516
rect 11212 2468 11656 2494
rect 11212 2466 11380 2468
rect 11212 2288 11239 2466
rect 11279 2428 11343 2440
rect 11619 2436 11656 2468
rect 11682 2467 11873 2489
rect 12008 2487 12117 2507
rect 12137 2487 12146 2507
rect 12008 2480 12146 2487
rect 12204 2507 12352 2516
rect 12204 2487 12213 2507
rect 12233 2487 12323 2507
rect 12343 2487 12352 2507
rect 12008 2478 12104 2480
rect 12204 2477 12352 2487
rect 12411 2507 12448 2517
rect 12411 2487 12419 2507
rect 12439 2487 12448 2507
rect 12260 2476 12296 2477
rect 11837 2465 11873 2467
rect 11837 2436 11874 2465
rect 11279 2427 11314 2428
rect 11256 2422 11314 2427
rect 11256 2402 11259 2422
rect 11279 2408 11314 2422
rect 11334 2408 11343 2428
rect 11279 2402 11343 2408
rect 11256 2400 11343 2402
rect 11256 2396 11283 2400
rect 11305 2399 11343 2400
rect 11306 2398 11343 2399
rect 11409 2432 11445 2433
rect 11517 2432 11553 2433
rect 11409 2425 11553 2432
rect 11409 2424 11471 2425
rect 11409 2404 11417 2424
rect 11437 2407 11471 2424
rect 11490 2424 11553 2425
rect 11490 2407 11525 2424
rect 11437 2404 11525 2407
rect 11545 2404 11553 2424
rect 11409 2398 11553 2404
rect 11619 2428 11657 2436
rect 11735 2432 11771 2433
rect 11619 2408 11628 2428
rect 11648 2408 11657 2428
rect 11619 2399 11657 2408
rect 11686 2424 11771 2432
rect 11686 2404 11743 2424
rect 11763 2404 11771 2424
rect 11619 2398 11656 2399
rect 11686 2398 11771 2404
rect 11837 2428 11875 2436
rect 11837 2408 11846 2428
rect 11866 2408 11875 2428
rect 12108 2417 12145 2418
rect 12411 2417 12448 2487
rect 12483 2516 12514 2567
rect 12810 2562 12855 2568
rect 12810 2544 12828 2562
rect 12846 2544 12855 2562
rect 14382 2560 14391 2580
rect 14411 2560 14419 2580
rect 14382 2550 14419 2560
rect 14478 2580 14565 2590
rect 14478 2560 14487 2580
rect 14507 2560 14565 2580
rect 14478 2551 14565 2560
rect 14478 2550 14515 2551
rect 12810 2534 12855 2544
rect 12533 2516 12570 2517
rect 12483 2507 12570 2516
rect 12483 2487 12541 2507
rect 12561 2487 12570 2507
rect 12483 2477 12570 2487
rect 12629 2507 12666 2517
rect 12629 2487 12637 2507
rect 12657 2487 12666 2507
rect 12810 2492 12853 2534
rect 13237 2523 13289 2525
rect 12716 2490 12853 2492
rect 12483 2476 12514 2477
rect 12629 2417 12666 2487
rect 12107 2416 12448 2417
rect 11837 2399 11875 2408
rect 12032 2411 12448 2416
rect 11837 2398 11874 2399
rect 11298 2370 11388 2376
rect 11298 2350 11314 2370
rect 11334 2368 11388 2370
rect 11334 2350 11359 2368
rect 11298 2348 11359 2350
rect 11379 2348 11388 2368
rect 11298 2342 11388 2348
rect 11311 2288 11348 2289
rect 11407 2288 11444 2289
rect 11463 2288 11499 2398
rect 11686 2377 11717 2398
rect 12032 2391 12035 2411
rect 12055 2391 12448 2411
rect 12632 2401 12666 2417
rect 12710 2469 12853 2490
rect 13235 2519 13668 2523
rect 13235 2513 13674 2519
rect 13235 2495 13256 2513
rect 13274 2495 13674 2513
rect 14534 2500 14565 2551
rect 14600 2580 14637 2650
rect 14903 2649 14940 2650
rect 14752 2590 14788 2591
rect 14600 2560 14609 2580
rect 14629 2560 14637 2580
rect 14600 2550 14637 2560
rect 14696 2580 14844 2590
rect 14944 2587 15040 2589
rect 14696 2560 14705 2580
rect 14725 2560 14815 2580
rect 14835 2560 14844 2580
rect 14696 2551 14844 2560
rect 14902 2580 15040 2587
rect 14902 2560 14911 2580
rect 14931 2560 15040 2580
rect 14902 2551 15040 2560
rect 14696 2550 14733 2551
rect 14426 2497 14467 2498
rect 13235 2477 13674 2495
rect 12408 2382 12448 2391
rect 12710 2382 12737 2469
rect 12810 2443 12853 2469
rect 12810 2425 12823 2443
rect 12841 2425 12853 2443
rect 12810 2414 12853 2425
rect 11682 2376 11717 2377
rect 11560 2366 11717 2376
rect 11560 2346 11577 2366
rect 11597 2346 11717 2366
rect 11560 2339 11717 2346
rect 11784 2369 11930 2377
rect 11784 2349 11795 2369
rect 11815 2349 11854 2369
rect 11874 2349 11930 2369
rect 12408 2365 12737 2382
rect 12408 2364 12448 2365
rect 11784 2342 11930 2349
rect 12805 2353 12845 2356
rect 12805 2347 12848 2353
rect 12430 2344 12848 2347
rect 11784 2341 11825 2342
rect 11518 2288 11555 2289
rect 11211 2279 11349 2288
rect 11211 2259 11320 2279
rect 11340 2259 11349 2279
rect 11211 2252 11349 2259
rect 11407 2279 11555 2288
rect 11407 2259 11416 2279
rect 11436 2259 11526 2279
rect 11546 2259 11555 2279
rect 11211 2250 11307 2252
rect 11407 2249 11555 2259
rect 11614 2279 11651 2289
rect 11614 2259 11622 2279
rect 11642 2259 11651 2279
rect 11463 2248 11499 2249
rect 11311 2189 11348 2190
rect 11614 2189 11651 2259
rect 11686 2288 11717 2339
rect 12430 2326 12821 2344
rect 12839 2326 12848 2344
rect 12430 2324 12848 2326
rect 12430 2316 12457 2324
rect 12698 2321 12848 2324
rect 12010 2310 12178 2311
rect 12429 2310 12457 2316
rect 12010 2294 12457 2310
rect 12805 2316 12848 2321
rect 11736 2288 11773 2289
rect 11686 2279 11773 2288
rect 11686 2259 11744 2279
rect 11764 2259 11773 2279
rect 11686 2249 11773 2259
rect 11832 2279 11869 2289
rect 11832 2259 11840 2279
rect 11860 2259 11869 2279
rect 11686 2248 11717 2249
rect 11310 2188 11651 2189
rect 11832 2188 11869 2259
rect 11235 2183 11651 2188
rect 11235 2163 11238 2183
rect 11258 2163 11651 2183
rect 11682 2164 11869 2188
rect 12010 2284 12454 2294
rect 12010 2282 12178 2284
rect 11110 2084 11152 2129
rect 12010 2104 12037 2282
rect 12077 2244 12141 2256
rect 12417 2252 12454 2284
rect 12480 2283 12671 2305
rect 12635 2281 12671 2283
rect 12635 2252 12672 2281
rect 12805 2260 12845 2316
rect 12077 2243 12112 2244
rect 12054 2238 12112 2243
rect 12054 2218 12057 2238
rect 12077 2224 12112 2238
rect 12132 2224 12141 2244
rect 12077 2216 12141 2224
rect 12103 2215 12141 2216
rect 12104 2214 12141 2215
rect 12207 2248 12243 2249
rect 12315 2248 12351 2249
rect 12207 2240 12351 2248
rect 12207 2220 12215 2240
rect 12235 2220 12270 2240
rect 12290 2220 12323 2240
rect 12343 2220 12351 2240
rect 12207 2214 12351 2220
rect 12417 2244 12455 2252
rect 12533 2248 12569 2249
rect 12417 2224 12426 2244
rect 12446 2224 12455 2244
rect 12417 2215 12455 2224
rect 12484 2240 12569 2248
rect 12484 2220 12541 2240
rect 12561 2220 12569 2240
rect 12417 2214 12454 2215
rect 12484 2214 12569 2220
rect 12635 2244 12673 2252
rect 12635 2224 12644 2244
rect 12664 2224 12673 2244
rect 12805 2242 12817 2260
rect 12835 2242 12845 2260
rect 13237 2288 13289 2477
rect 13635 2452 13674 2477
rect 14318 2490 14467 2497
rect 14318 2470 14377 2490
rect 14397 2470 14436 2490
rect 14456 2470 14467 2490
rect 14318 2462 14467 2470
rect 14534 2493 14691 2500
rect 14534 2473 14654 2493
rect 14674 2473 14691 2493
rect 14534 2463 14691 2473
rect 14534 2462 14569 2463
rect 13419 2427 13606 2451
rect 13635 2432 14030 2452
rect 14050 2432 14053 2452
rect 14534 2441 14565 2462
rect 14752 2441 14788 2551
rect 14807 2550 14844 2551
rect 14903 2550 14940 2551
rect 14863 2491 14953 2497
rect 14863 2471 14872 2491
rect 14892 2489 14953 2491
rect 14892 2471 14917 2489
rect 14863 2469 14917 2471
rect 14937 2469 14953 2489
rect 14863 2463 14953 2469
rect 14377 2440 14414 2441
rect 13635 2427 14053 2432
rect 14376 2431 14414 2440
rect 13419 2356 13456 2427
rect 13635 2426 13978 2427
rect 13635 2423 13674 2426
rect 13940 2425 13977 2426
rect 13571 2366 13602 2367
rect 13419 2336 13428 2356
rect 13448 2336 13456 2356
rect 13419 2326 13456 2336
rect 13515 2356 13602 2366
rect 13515 2336 13524 2356
rect 13544 2336 13602 2356
rect 13515 2327 13602 2336
rect 13515 2326 13552 2327
rect 13237 2270 13253 2288
rect 13271 2270 13289 2288
rect 13571 2276 13602 2327
rect 13637 2356 13674 2423
rect 14376 2411 14385 2431
rect 14405 2411 14414 2431
rect 14376 2403 14414 2411
rect 14480 2435 14565 2441
rect 14595 2440 14632 2441
rect 14480 2415 14488 2435
rect 14508 2415 14565 2435
rect 14480 2407 14565 2415
rect 14594 2431 14632 2440
rect 14594 2411 14603 2431
rect 14623 2411 14632 2431
rect 14480 2406 14516 2407
rect 14594 2403 14632 2411
rect 14698 2439 14842 2441
rect 14698 2435 14758 2439
rect 14698 2415 14706 2435
rect 14726 2417 14758 2435
rect 14781 2435 14842 2439
rect 14781 2417 14814 2435
rect 14726 2415 14814 2417
rect 14834 2415 14842 2435
rect 14698 2407 14842 2415
rect 14698 2406 14734 2407
rect 14806 2406 14842 2407
rect 14908 2440 14945 2441
rect 14908 2439 14946 2440
rect 14908 2431 14972 2439
rect 14908 2411 14917 2431
rect 14937 2417 14972 2431
rect 14992 2417 14995 2437
rect 14937 2412 14995 2417
rect 14937 2411 14972 2412
rect 14377 2374 14414 2403
rect 14378 2372 14414 2374
rect 13789 2366 13825 2367
rect 13637 2336 13646 2356
rect 13666 2336 13674 2356
rect 13637 2326 13674 2336
rect 13733 2356 13881 2366
rect 13981 2363 14077 2365
rect 13733 2336 13742 2356
rect 13762 2336 13852 2356
rect 13872 2336 13881 2356
rect 13733 2327 13881 2336
rect 13939 2356 14077 2363
rect 13939 2336 13948 2356
rect 13968 2336 14077 2356
rect 14378 2350 14569 2372
rect 14595 2371 14632 2403
rect 14908 2399 14972 2411
rect 14595 2370 14870 2371
rect 15012 2370 15039 2551
rect 14595 2345 15039 2370
rect 15175 2376 15214 4191
rect 15516 4178 15549 4511
rect 15613 4543 15781 4544
rect 15907 4543 15947 4767
rect 16410 4771 16578 4772
rect 16819 4771 16854 4788
rect 17211 4778 17258 4789
rect 16410 4745 16854 4771
rect 16410 4743 16578 4745
rect 16774 4744 16854 4745
rect 17009 4744 17076 4770
rect 17215 4744 17258 4778
rect 16410 4565 16437 4743
rect 16477 4705 16541 4717
rect 16817 4713 16854 4744
rect 17035 4713 17072 4744
rect 17217 4719 17258 4744
rect 16477 4704 16512 4705
rect 16454 4699 16512 4704
rect 16454 4679 16457 4699
rect 16477 4685 16512 4699
rect 16532 4685 16541 4705
rect 16477 4677 16541 4685
rect 16503 4676 16541 4677
rect 16504 4675 16541 4676
rect 16607 4709 16643 4710
rect 16715 4709 16751 4710
rect 16607 4701 16751 4709
rect 16607 4681 16615 4701
rect 16635 4697 16723 4701
rect 16635 4681 16679 4697
rect 16607 4677 16679 4681
rect 16699 4681 16723 4697
rect 16743 4681 16751 4701
rect 16699 4677 16751 4681
rect 16607 4675 16751 4677
rect 16817 4705 16855 4713
rect 16933 4709 16969 4710
rect 16817 4685 16826 4705
rect 16846 4685 16855 4705
rect 16817 4676 16855 4685
rect 16884 4701 16969 4709
rect 16884 4681 16941 4701
rect 16961 4681 16969 4701
rect 16817 4675 16854 4676
rect 16884 4675 16969 4681
rect 17035 4705 17073 4713
rect 17035 4685 17044 4705
rect 17064 4685 17073 4705
rect 17035 4676 17073 4685
rect 17217 4710 17259 4719
rect 17217 4692 17231 4710
rect 17249 4692 17259 4710
rect 17217 4684 17259 4692
rect 17222 4682 17259 4684
rect 17035 4675 17072 4676
rect 16496 4647 16586 4653
rect 16496 4627 16512 4647
rect 16532 4645 16586 4647
rect 16532 4627 16557 4645
rect 16496 4625 16557 4627
rect 16577 4625 16586 4645
rect 16496 4619 16586 4625
rect 16509 4565 16546 4566
rect 16605 4565 16642 4566
rect 16661 4565 16697 4675
rect 16884 4654 16915 4675
rect 16880 4653 16915 4654
rect 16758 4643 16915 4653
rect 16758 4623 16775 4643
rect 16795 4623 16915 4643
rect 16758 4616 16915 4623
rect 16982 4646 17131 4654
rect 16982 4626 16993 4646
rect 17013 4626 17052 4646
rect 17072 4626 17131 4646
rect 16982 4619 17131 4626
rect 16982 4618 17023 4619
rect 17219 4617 17256 4620
rect 16716 4565 16753 4566
rect 16409 4556 16547 4565
rect 15613 4517 16057 4543
rect 15613 4515 15781 4517
rect 15613 4337 15640 4515
rect 15680 4477 15744 4489
rect 16020 4485 16057 4517
rect 16083 4516 16274 4538
rect 16409 4536 16518 4556
rect 16538 4536 16547 4556
rect 16409 4529 16547 4536
rect 16605 4556 16753 4565
rect 16605 4536 16614 4556
rect 16634 4536 16724 4556
rect 16744 4536 16753 4556
rect 16409 4527 16505 4529
rect 16605 4526 16753 4536
rect 16812 4556 16849 4566
rect 16812 4536 16820 4556
rect 16840 4536 16849 4556
rect 16661 4525 16697 4526
rect 16238 4514 16274 4516
rect 16238 4485 16275 4514
rect 15680 4476 15715 4477
rect 15657 4471 15715 4476
rect 15657 4451 15660 4471
rect 15680 4457 15715 4471
rect 15735 4457 15744 4477
rect 15680 4451 15744 4457
rect 15657 4449 15744 4451
rect 15657 4445 15684 4449
rect 15706 4448 15744 4449
rect 15707 4447 15744 4448
rect 15810 4481 15846 4482
rect 15918 4481 15954 4482
rect 15810 4474 15954 4481
rect 15810 4473 15872 4474
rect 15810 4453 15818 4473
rect 15838 4456 15872 4473
rect 15891 4473 15954 4474
rect 15891 4456 15926 4473
rect 15838 4453 15926 4456
rect 15946 4453 15954 4473
rect 15810 4447 15954 4453
rect 16020 4477 16058 4485
rect 16136 4481 16172 4482
rect 16020 4457 16029 4477
rect 16049 4457 16058 4477
rect 16020 4448 16058 4457
rect 16087 4473 16172 4481
rect 16087 4453 16144 4473
rect 16164 4453 16172 4473
rect 16020 4447 16057 4448
rect 16087 4447 16172 4453
rect 16238 4477 16276 4485
rect 16238 4457 16247 4477
rect 16267 4457 16276 4477
rect 16509 4466 16546 4467
rect 16812 4466 16849 4536
rect 16884 4565 16915 4616
rect 17211 4611 17256 4617
rect 17211 4593 17229 4611
rect 17247 4593 17256 4611
rect 17211 4583 17256 4593
rect 16934 4565 16971 4566
rect 16884 4556 16971 4565
rect 16884 4536 16942 4556
rect 16962 4536 16971 4556
rect 16884 4526 16971 4536
rect 17030 4556 17067 4566
rect 17030 4536 17038 4556
rect 17058 4536 17067 4556
rect 17211 4541 17254 4583
rect 17117 4539 17254 4541
rect 16884 4525 16915 4526
rect 17030 4466 17067 4536
rect 16508 4465 16849 4466
rect 16238 4448 16276 4457
rect 16433 4460 16849 4465
rect 16238 4447 16275 4448
rect 15699 4419 15789 4425
rect 15699 4399 15715 4419
rect 15735 4417 15789 4419
rect 15735 4399 15760 4417
rect 15699 4397 15760 4399
rect 15780 4397 15789 4417
rect 15699 4391 15789 4397
rect 15712 4337 15749 4338
rect 15808 4337 15845 4338
rect 15864 4337 15900 4447
rect 16087 4426 16118 4447
rect 16433 4440 16436 4460
rect 16456 4440 16849 4460
rect 17033 4450 17067 4466
rect 17111 4518 17254 4539
rect 16809 4431 16849 4440
rect 17111 4431 17138 4518
rect 17211 4492 17254 4518
rect 17211 4474 17224 4492
rect 17242 4474 17254 4492
rect 17211 4463 17254 4474
rect 16083 4425 16118 4426
rect 15961 4415 16118 4425
rect 15961 4395 15978 4415
rect 15998 4395 16118 4415
rect 15961 4388 16118 4395
rect 16185 4418 16331 4426
rect 16185 4398 16196 4418
rect 16216 4398 16255 4418
rect 16275 4398 16331 4418
rect 16809 4414 17138 4431
rect 16809 4413 16849 4414
rect 16185 4391 16331 4398
rect 17206 4402 17246 4405
rect 17206 4396 17249 4402
rect 16831 4393 17249 4396
rect 16185 4390 16226 4391
rect 15919 4337 15956 4338
rect 15612 4328 15750 4337
rect 15612 4308 15721 4328
rect 15741 4308 15750 4328
rect 15612 4301 15750 4308
rect 15808 4328 15956 4337
rect 15808 4308 15817 4328
rect 15837 4308 15927 4328
rect 15947 4308 15956 4328
rect 15612 4299 15708 4301
rect 15808 4298 15956 4308
rect 16015 4328 16052 4338
rect 16015 4308 16023 4328
rect 16043 4308 16052 4328
rect 15864 4297 15900 4298
rect 15712 4238 15749 4239
rect 16015 4238 16052 4308
rect 16087 4337 16118 4388
rect 16831 4375 17222 4393
rect 17240 4375 17249 4393
rect 16831 4373 17249 4375
rect 16831 4365 16858 4373
rect 17099 4370 17249 4373
rect 16411 4359 16579 4360
rect 16830 4359 16858 4365
rect 16411 4343 16858 4359
rect 17206 4365 17249 4370
rect 16137 4337 16174 4338
rect 16087 4328 16174 4337
rect 16087 4308 16145 4328
rect 16165 4308 16174 4328
rect 16087 4298 16174 4308
rect 16233 4328 16270 4338
rect 16233 4308 16241 4328
rect 16261 4308 16270 4328
rect 16087 4297 16118 4298
rect 15711 4237 16052 4238
rect 16233 4237 16270 4308
rect 15636 4232 16052 4237
rect 15636 4212 15639 4232
rect 15659 4212 16052 4232
rect 16083 4213 16270 4237
rect 16411 4333 16855 4343
rect 16411 4331 16579 4333
rect 15445 4138 15489 4139
rect 15445 4132 15490 4138
rect 15445 4114 15457 4132
rect 15479 4114 15490 4132
rect 15511 4133 15553 4178
rect 16411 4153 16438 4331
rect 16478 4293 16542 4305
rect 16818 4301 16855 4333
rect 16881 4332 17072 4354
rect 17036 4330 17072 4332
rect 17036 4301 17073 4330
rect 17206 4309 17246 4365
rect 16478 4292 16513 4293
rect 16455 4287 16513 4292
rect 16455 4267 16458 4287
rect 16478 4273 16513 4287
rect 16533 4273 16542 4293
rect 16478 4265 16542 4273
rect 16504 4264 16542 4265
rect 16505 4263 16542 4264
rect 16608 4297 16644 4298
rect 16716 4297 16752 4298
rect 16608 4289 16752 4297
rect 16608 4269 16616 4289
rect 16636 4269 16671 4289
rect 16691 4269 16724 4289
rect 16744 4269 16752 4289
rect 16608 4263 16752 4269
rect 16818 4293 16856 4301
rect 16934 4297 16970 4298
rect 16818 4273 16827 4293
rect 16847 4273 16856 4293
rect 16818 4264 16856 4273
rect 16885 4289 16970 4297
rect 16885 4269 16942 4289
rect 16962 4269 16970 4289
rect 16818 4263 16855 4264
rect 16885 4263 16970 4269
rect 17036 4293 17074 4301
rect 17036 4273 17045 4293
rect 17065 4273 17074 4293
rect 17206 4291 17218 4309
rect 17236 4291 17246 4309
rect 17206 4281 17246 4291
rect 17036 4264 17074 4273
rect 17036 4263 17073 4264
rect 16497 4235 16587 4241
rect 16497 4215 16513 4235
rect 16533 4233 16587 4235
rect 16533 4215 16558 4233
rect 16497 4213 16558 4215
rect 16578 4213 16587 4233
rect 16497 4207 16587 4213
rect 16510 4153 16547 4154
rect 16606 4153 16643 4154
rect 16662 4153 16698 4263
rect 16885 4242 16916 4263
rect 16881 4241 16916 4242
rect 16759 4231 16916 4241
rect 16759 4211 16776 4231
rect 16796 4211 16916 4231
rect 16759 4204 16916 4211
rect 16983 4234 17132 4242
rect 16983 4214 16994 4234
rect 17014 4214 17053 4234
rect 17073 4214 17132 4234
rect 16983 4207 17132 4214
rect 17198 4210 17250 4228
rect 16983 4206 17024 4207
rect 16717 4153 16754 4154
rect 16410 4144 16548 4153
rect 15882 4133 15915 4135
rect 15511 4121 15958 4133
rect 15445 4084 15490 4114
rect 15462 3138 15490 4084
rect 15514 4107 15958 4121
rect 15514 4105 15682 4107
rect 15514 3927 15541 4105
rect 15581 4067 15645 4079
rect 15921 4075 15958 4107
rect 15984 4106 16175 4128
rect 16410 4124 16519 4144
rect 16539 4124 16548 4144
rect 16410 4117 16548 4124
rect 16606 4144 16754 4153
rect 16606 4124 16615 4144
rect 16635 4124 16725 4144
rect 16745 4124 16754 4144
rect 16410 4115 16506 4117
rect 16606 4114 16754 4124
rect 16813 4144 16850 4154
rect 16813 4124 16821 4144
rect 16841 4124 16850 4144
rect 16662 4113 16698 4114
rect 16139 4104 16175 4106
rect 16139 4075 16176 4104
rect 15581 4066 15616 4067
rect 15558 4061 15616 4066
rect 15558 4041 15561 4061
rect 15581 4047 15616 4061
rect 15636 4047 15645 4067
rect 15581 4039 15645 4047
rect 15607 4038 15645 4039
rect 15608 4037 15645 4038
rect 15711 4071 15747 4072
rect 15819 4071 15855 4072
rect 15711 4065 15855 4071
rect 15711 4063 15772 4065
rect 15711 4043 15719 4063
rect 15739 4048 15772 4063
rect 15791 4063 15855 4065
rect 15791 4048 15827 4063
rect 15739 4043 15827 4048
rect 15847 4043 15855 4063
rect 15711 4037 15855 4043
rect 15921 4067 15959 4075
rect 16037 4071 16073 4072
rect 15921 4047 15930 4067
rect 15950 4047 15959 4067
rect 15921 4038 15959 4047
rect 15988 4063 16073 4071
rect 15988 4043 16045 4063
rect 16065 4043 16073 4063
rect 15921 4037 15958 4038
rect 15988 4037 16073 4043
rect 16139 4067 16177 4075
rect 16139 4047 16148 4067
rect 16168 4047 16177 4067
rect 16813 4057 16850 4124
rect 16885 4153 16916 4204
rect 17198 4192 17216 4210
rect 17234 4192 17250 4210
rect 16935 4153 16972 4154
rect 16885 4144 16972 4153
rect 16885 4124 16943 4144
rect 16963 4124 16972 4144
rect 16885 4114 16972 4124
rect 17031 4144 17068 4154
rect 17031 4124 17039 4144
rect 17059 4124 17068 4144
rect 16885 4113 16916 4114
rect 16510 4054 16547 4055
rect 16813 4054 16852 4057
rect 16509 4053 16852 4054
rect 17031 4053 17068 4124
rect 16139 4038 16177 4047
rect 16434 4048 16852 4053
rect 16139 4037 16176 4038
rect 15600 4009 15690 4015
rect 15600 3989 15616 4009
rect 15636 4007 15690 4009
rect 15636 3989 15661 4007
rect 15600 3987 15661 3989
rect 15681 3987 15690 4007
rect 15600 3981 15690 3987
rect 15613 3927 15650 3928
rect 15709 3927 15746 3928
rect 15765 3927 15801 4037
rect 15988 4016 16019 4037
rect 16434 4028 16437 4048
rect 16457 4028 16852 4048
rect 16881 4029 17068 4053
rect 15984 4015 16019 4016
rect 15862 4005 16019 4015
rect 15862 3985 15879 4005
rect 15899 3985 16019 4005
rect 15862 3978 16019 3985
rect 16086 4008 16235 4016
rect 16086 3988 16097 4008
rect 16117 3988 16156 4008
rect 16176 3988 16235 4008
rect 16086 3981 16235 3988
rect 16813 4003 16852 4028
rect 17198 4003 17250 4192
rect 16813 3985 17252 4003
rect 16086 3980 16127 3981
rect 15820 3927 15857 3928
rect 15513 3918 15651 3927
rect 15513 3898 15622 3918
rect 15642 3898 15651 3918
rect 15513 3891 15651 3898
rect 15709 3918 15857 3927
rect 15709 3898 15718 3918
rect 15738 3898 15828 3918
rect 15848 3898 15857 3918
rect 15513 3889 15609 3891
rect 15709 3888 15857 3898
rect 15916 3918 15953 3928
rect 15916 3898 15924 3918
rect 15944 3898 15953 3918
rect 15765 3887 15801 3888
rect 15613 3828 15650 3829
rect 15916 3828 15953 3898
rect 15988 3927 16019 3978
rect 16813 3967 17213 3985
rect 17231 3967 17252 3985
rect 16813 3961 17252 3967
rect 16819 3957 17252 3961
rect 17198 3955 17250 3957
rect 16038 3927 16075 3928
rect 15988 3918 16075 3927
rect 15988 3898 16046 3918
rect 16066 3898 16075 3918
rect 15988 3888 16075 3898
rect 16134 3918 16171 3928
rect 16134 3898 16142 3918
rect 16162 3898 16171 3918
rect 15988 3887 16019 3888
rect 15612 3827 15953 3828
rect 16134 3827 16171 3898
rect 17201 3890 17238 3895
rect 17192 3886 17239 3890
rect 17192 3868 17211 3886
rect 17229 3868 17239 3886
rect 15537 3822 15953 3827
rect 15537 3802 15540 3822
rect 15560 3802 15953 3822
rect 15984 3803 16171 3827
rect 16796 3825 16836 3830
rect 17192 3825 17239 3868
rect 16796 3786 17239 3825
rect 15890 3771 15930 3779
rect 15890 3749 15898 3771
rect 15922 3749 15930 3771
rect 15596 3525 15764 3526
rect 15890 3525 15930 3749
rect 16393 3753 16561 3754
rect 16796 3753 16836 3786
rect 17192 3753 17239 3786
rect 16393 3752 16837 3753
rect 16393 3727 16838 3752
rect 16393 3725 16561 3727
rect 16757 3726 16838 3727
rect 17007 3726 17056 3752
rect 17192 3726 17241 3753
rect 16393 3547 16420 3725
rect 16460 3687 16524 3699
rect 16800 3695 16837 3726
rect 17018 3695 17055 3726
rect 17200 3701 17241 3726
rect 16460 3686 16495 3687
rect 16437 3681 16495 3686
rect 16437 3661 16440 3681
rect 16460 3667 16495 3681
rect 16515 3667 16524 3687
rect 16460 3659 16524 3667
rect 16486 3658 16524 3659
rect 16487 3657 16524 3658
rect 16590 3691 16626 3692
rect 16698 3691 16734 3692
rect 16590 3683 16734 3691
rect 16590 3663 16598 3683
rect 16618 3679 16706 3683
rect 16618 3663 16662 3679
rect 16590 3659 16662 3663
rect 16682 3663 16706 3679
rect 16726 3663 16734 3683
rect 16682 3659 16734 3663
rect 16590 3657 16734 3659
rect 16800 3687 16838 3695
rect 16916 3691 16952 3692
rect 16800 3667 16809 3687
rect 16829 3667 16838 3687
rect 16800 3658 16838 3667
rect 16867 3683 16952 3691
rect 16867 3663 16924 3683
rect 16944 3663 16952 3683
rect 16800 3657 16837 3658
rect 16867 3657 16952 3663
rect 17018 3687 17056 3695
rect 17018 3667 17027 3687
rect 17047 3667 17056 3687
rect 17018 3658 17056 3667
rect 17200 3692 17242 3701
rect 17200 3674 17214 3692
rect 17232 3674 17242 3692
rect 17200 3666 17242 3674
rect 17205 3664 17242 3666
rect 17018 3657 17055 3658
rect 16479 3629 16569 3635
rect 16479 3609 16495 3629
rect 16515 3627 16569 3629
rect 16515 3609 16540 3627
rect 16479 3607 16540 3609
rect 16560 3607 16569 3627
rect 16479 3601 16569 3607
rect 16492 3547 16529 3548
rect 16588 3547 16625 3548
rect 16644 3547 16680 3657
rect 16867 3636 16898 3657
rect 16863 3635 16898 3636
rect 16741 3625 16898 3635
rect 16741 3605 16758 3625
rect 16778 3605 16898 3625
rect 16741 3598 16898 3605
rect 16965 3628 17114 3636
rect 16965 3608 16976 3628
rect 16996 3608 17035 3628
rect 17055 3608 17114 3628
rect 16965 3601 17114 3608
rect 16965 3600 17006 3601
rect 17202 3599 17239 3602
rect 16699 3547 16736 3548
rect 16392 3538 16530 3547
rect 15596 3499 16040 3525
rect 15596 3497 15764 3499
rect 15596 3319 15623 3497
rect 15663 3459 15727 3471
rect 16003 3467 16040 3499
rect 16066 3498 16257 3520
rect 16392 3518 16501 3538
rect 16521 3518 16530 3538
rect 16392 3511 16530 3518
rect 16588 3538 16736 3547
rect 16588 3518 16597 3538
rect 16617 3518 16707 3538
rect 16727 3518 16736 3538
rect 16392 3509 16488 3511
rect 16588 3508 16736 3518
rect 16795 3538 16832 3548
rect 16795 3518 16803 3538
rect 16823 3518 16832 3538
rect 16644 3507 16680 3508
rect 16221 3496 16257 3498
rect 16221 3467 16258 3496
rect 15663 3458 15698 3459
rect 15640 3453 15698 3458
rect 15640 3433 15643 3453
rect 15663 3439 15698 3453
rect 15718 3439 15727 3459
rect 15663 3431 15727 3439
rect 15689 3430 15727 3431
rect 15690 3429 15727 3430
rect 15793 3463 15829 3464
rect 15901 3463 15937 3464
rect 15793 3455 15937 3463
rect 15793 3435 15801 3455
rect 15821 3454 15909 3455
rect 15821 3435 15856 3454
rect 15877 3435 15909 3454
rect 15929 3435 15937 3455
rect 15793 3429 15937 3435
rect 16003 3459 16041 3467
rect 16119 3463 16155 3464
rect 16003 3439 16012 3459
rect 16032 3439 16041 3459
rect 16003 3430 16041 3439
rect 16070 3455 16155 3463
rect 16070 3435 16127 3455
rect 16147 3435 16155 3455
rect 16003 3429 16040 3430
rect 16070 3429 16155 3435
rect 16221 3459 16259 3467
rect 16221 3439 16230 3459
rect 16250 3439 16259 3459
rect 16492 3448 16529 3449
rect 16795 3448 16832 3518
rect 16867 3547 16898 3598
rect 17194 3593 17239 3599
rect 17194 3575 17212 3593
rect 17230 3575 17239 3593
rect 17194 3565 17239 3575
rect 16917 3547 16954 3548
rect 16867 3538 16954 3547
rect 16867 3518 16925 3538
rect 16945 3518 16954 3538
rect 16867 3508 16954 3518
rect 17013 3538 17050 3548
rect 17013 3518 17021 3538
rect 17041 3518 17050 3538
rect 17194 3523 17237 3565
rect 17100 3521 17237 3523
rect 16867 3507 16898 3508
rect 17013 3448 17050 3518
rect 16491 3447 16832 3448
rect 16221 3430 16259 3439
rect 16416 3442 16832 3447
rect 16221 3429 16258 3430
rect 15682 3401 15772 3407
rect 15682 3381 15698 3401
rect 15718 3399 15772 3401
rect 15718 3381 15743 3399
rect 15682 3379 15743 3381
rect 15763 3379 15772 3399
rect 15682 3373 15772 3379
rect 15695 3319 15732 3320
rect 15791 3319 15828 3320
rect 15847 3319 15883 3429
rect 16070 3408 16101 3429
rect 16416 3422 16419 3442
rect 16439 3422 16832 3442
rect 17016 3432 17050 3448
rect 17094 3500 17237 3521
rect 16792 3413 16832 3422
rect 17094 3413 17121 3500
rect 17194 3474 17237 3500
rect 17194 3456 17207 3474
rect 17225 3456 17237 3474
rect 17194 3445 17237 3456
rect 16066 3407 16101 3408
rect 15944 3397 16101 3407
rect 15944 3377 15961 3397
rect 15981 3377 16101 3397
rect 15944 3370 16101 3377
rect 16168 3400 16317 3408
rect 16168 3380 16179 3400
rect 16199 3380 16238 3400
rect 16258 3380 16317 3400
rect 16792 3396 17121 3413
rect 16792 3395 16832 3396
rect 16168 3373 16317 3380
rect 17189 3384 17229 3387
rect 17189 3378 17232 3384
rect 16814 3375 17232 3378
rect 16168 3372 16209 3373
rect 15902 3319 15939 3320
rect 15595 3310 15733 3319
rect 15595 3290 15704 3310
rect 15724 3290 15733 3310
rect 15595 3283 15733 3290
rect 15791 3310 15939 3319
rect 15791 3290 15800 3310
rect 15820 3290 15910 3310
rect 15930 3290 15939 3310
rect 15595 3281 15691 3283
rect 15791 3280 15939 3290
rect 15998 3310 16035 3320
rect 15998 3290 16006 3310
rect 16026 3290 16035 3310
rect 15847 3279 15883 3280
rect 15695 3220 15732 3221
rect 15998 3220 16035 3290
rect 16070 3319 16101 3370
rect 16814 3357 17205 3375
rect 17223 3357 17232 3375
rect 16814 3355 17232 3357
rect 16814 3347 16841 3355
rect 17082 3352 17232 3355
rect 16394 3341 16562 3342
rect 16813 3341 16841 3347
rect 16394 3325 16841 3341
rect 17189 3347 17232 3352
rect 16120 3319 16157 3320
rect 16070 3310 16157 3319
rect 16070 3290 16128 3310
rect 16148 3290 16157 3310
rect 16070 3280 16157 3290
rect 16216 3310 16253 3320
rect 16216 3290 16224 3310
rect 16244 3290 16253 3310
rect 16070 3279 16101 3280
rect 15694 3219 16035 3220
rect 16216 3219 16253 3290
rect 15619 3214 16035 3219
rect 15619 3194 15622 3214
rect 15642 3194 16035 3214
rect 16066 3195 16253 3219
rect 16394 3315 16838 3325
rect 16394 3313 16562 3315
rect 15461 3120 15490 3138
rect 16394 3135 16421 3313
rect 16461 3275 16525 3287
rect 16801 3283 16838 3315
rect 16864 3314 17055 3336
rect 17019 3312 17055 3314
rect 17019 3283 17056 3312
rect 17189 3291 17229 3347
rect 16461 3274 16496 3275
rect 16438 3269 16496 3274
rect 16438 3249 16441 3269
rect 16461 3255 16496 3269
rect 16516 3255 16525 3275
rect 16461 3247 16525 3255
rect 16487 3246 16525 3247
rect 16488 3245 16525 3246
rect 16591 3279 16627 3280
rect 16699 3279 16735 3280
rect 16591 3271 16735 3279
rect 16591 3251 16599 3271
rect 16619 3251 16654 3271
rect 16674 3251 16707 3271
rect 16727 3251 16735 3271
rect 16591 3245 16735 3251
rect 16801 3275 16839 3283
rect 16917 3279 16953 3280
rect 16801 3255 16810 3275
rect 16830 3255 16839 3275
rect 16801 3246 16839 3255
rect 16868 3271 16953 3279
rect 16868 3251 16925 3271
rect 16945 3251 16953 3271
rect 16801 3245 16838 3246
rect 16868 3245 16953 3251
rect 17019 3275 17057 3283
rect 17019 3255 17028 3275
rect 17048 3255 17057 3275
rect 17189 3273 17201 3291
rect 17219 3273 17229 3291
rect 17189 3263 17229 3273
rect 17019 3246 17057 3255
rect 17019 3245 17056 3246
rect 16480 3217 16570 3223
rect 16480 3197 16496 3217
rect 16516 3215 16570 3217
rect 16516 3197 16541 3215
rect 16480 3195 16541 3197
rect 16561 3195 16570 3215
rect 16480 3189 16570 3195
rect 16493 3135 16530 3136
rect 16589 3135 16626 3136
rect 16645 3135 16681 3245
rect 16868 3224 16899 3245
rect 16864 3223 16899 3224
rect 16742 3213 16899 3223
rect 16742 3193 16759 3213
rect 16779 3193 16899 3213
rect 16742 3186 16899 3193
rect 16966 3216 17115 3224
rect 16966 3196 16977 3216
rect 16997 3196 17036 3216
rect 17056 3196 17115 3216
rect 16966 3189 17115 3196
rect 17181 3192 17233 3210
rect 16966 3188 17007 3189
rect 16700 3135 16737 3136
rect 15431 3118 15490 3120
rect 16393 3126 16531 3135
rect 15431 3117 15599 3118
rect 15725 3117 15765 3119
rect 15431 3091 15875 3117
rect 15431 3089 15599 3091
rect 15431 3087 15512 3089
rect 15431 2911 15458 3087
rect 15498 3051 15562 3063
rect 15838 3059 15875 3091
rect 15901 3090 16092 3112
rect 16393 3106 16502 3126
rect 16522 3106 16531 3126
rect 16393 3099 16531 3106
rect 16589 3126 16737 3135
rect 16589 3106 16598 3126
rect 16618 3106 16708 3126
rect 16728 3106 16737 3126
rect 16393 3097 16489 3099
rect 16589 3096 16737 3106
rect 16796 3126 16833 3136
rect 16796 3106 16804 3126
rect 16824 3106 16833 3126
rect 16645 3095 16681 3096
rect 16056 3088 16092 3090
rect 16056 3059 16093 3088
rect 15498 3050 15533 3051
rect 15475 3045 15533 3050
rect 15475 3025 15478 3045
rect 15498 3031 15533 3045
rect 15553 3031 15562 3051
rect 15498 3023 15562 3031
rect 15524 3022 15562 3023
rect 15525 3021 15562 3022
rect 15628 3055 15664 3056
rect 15736 3055 15772 3056
rect 15628 3047 15772 3055
rect 15628 3027 15636 3047
rect 15656 3046 15744 3047
rect 15656 3028 15691 3046
rect 15709 3028 15744 3046
rect 15656 3027 15744 3028
rect 15764 3027 15772 3047
rect 15628 3021 15772 3027
rect 15838 3051 15876 3059
rect 15954 3055 15990 3056
rect 15838 3031 15847 3051
rect 15867 3031 15876 3051
rect 15838 3022 15876 3031
rect 15905 3047 15990 3055
rect 15905 3027 15962 3047
rect 15982 3027 15990 3047
rect 15838 3021 15875 3022
rect 15905 3021 15990 3027
rect 16056 3051 16094 3059
rect 16056 3031 16065 3051
rect 16085 3031 16094 3051
rect 16796 3039 16833 3106
rect 16868 3135 16899 3186
rect 17181 3174 17199 3192
rect 17217 3174 17233 3192
rect 16918 3135 16955 3136
rect 16868 3126 16955 3135
rect 16868 3106 16926 3126
rect 16946 3106 16955 3126
rect 16868 3096 16955 3106
rect 17014 3126 17051 3136
rect 17014 3106 17022 3126
rect 17042 3106 17051 3126
rect 16868 3095 16899 3096
rect 16493 3036 16530 3037
rect 16796 3036 16835 3039
rect 16492 3035 16835 3036
rect 17014 3035 17051 3106
rect 16056 3022 16094 3031
rect 16417 3030 16835 3035
rect 16056 3021 16093 3022
rect 15517 2993 15607 2999
rect 15517 2973 15533 2993
rect 15553 2991 15607 2993
rect 15553 2973 15578 2991
rect 15517 2971 15578 2973
rect 15598 2971 15607 2991
rect 15517 2965 15607 2971
rect 15530 2911 15567 2912
rect 15626 2911 15663 2912
rect 15682 2911 15718 3021
rect 15905 3000 15936 3021
rect 16417 3010 16420 3030
rect 16440 3010 16835 3030
rect 16864 3011 17051 3035
rect 15901 2999 15936 3000
rect 15779 2989 15936 2999
rect 15779 2969 15796 2989
rect 15816 2969 15936 2989
rect 15779 2962 15936 2969
rect 16003 2992 16152 3000
rect 16003 2972 16014 2992
rect 16034 2972 16073 2992
rect 16093 2972 16152 2992
rect 16003 2965 16152 2972
rect 16796 2985 16835 3010
rect 17181 2985 17233 3174
rect 16796 2967 17235 2985
rect 16003 2964 16044 2965
rect 15737 2911 15774 2912
rect 15430 2902 15568 2911
rect 15430 2882 15539 2902
rect 15559 2882 15568 2902
rect 15430 2875 15568 2882
rect 15626 2902 15774 2911
rect 15626 2882 15635 2902
rect 15655 2882 15745 2902
rect 15765 2882 15774 2902
rect 15430 2873 15526 2875
rect 15626 2872 15774 2882
rect 15833 2902 15870 2912
rect 15833 2882 15841 2902
rect 15861 2882 15870 2902
rect 15682 2871 15718 2872
rect 15530 2812 15567 2813
rect 15833 2812 15870 2882
rect 15905 2911 15936 2962
rect 16796 2949 17196 2967
rect 17214 2949 17235 2967
rect 16796 2943 17235 2949
rect 16802 2939 17235 2943
rect 17181 2937 17233 2939
rect 15955 2911 15992 2912
rect 15905 2902 15992 2911
rect 15905 2882 15963 2902
rect 15983 2882 15992 2902
rect 15905 2872 15992 2882
rect 16051 2902 16088 2912
rect 16051 2882 16059 2902
rect 16079 2882 16088 2902
rect 15905 2871 15936 2872
rect 15529 2811 15870 2812
rect 16051 2811 16088 2882
rect 17184 2872 17221 2877
rect 15454 2806 15870 2811
rect 15454 2786 15457 2806
rect 15477 2786 15870 2806
rect 15901 2787 16088 2811
rect 17175 2868 17222 2872
rect 17175 2850 17194 2868
rect 17212 2850 17222 2868
rect 17175 2802 17222 2850
rect 16799 2799 17222 2802
rect 15674 2785 15739 2786
rect 16777 2769 17222 2799
rect 15870 2753 15910 2761
rect 15870 2731 15878 2753
rect 15902 2731 15910 2753
rect 15475 2502 15512 2508
rect 15475 2483 15483 2502
rect 15504 2483 15512 2502
rect 15475 2475 15512 2483
rect 15175 2354 15182 2376
rect 15206 2354 15214 2376
rect 15175 2348 15214 2354
rect 14705 2343 14745 2345
rect 14871 2344 15039 2345
rect 14973 2343 15010 2344
rect 13939 2327 14077 2336
rect 13733 2326 13770 2327
rect 13463 2273 13504 2274
rect 13237 2252 13289 2270
rect 13355 2266 13504 2273
rect 12805 2232 12845 2242
rect 13355 2246 13414 2266
rect 13434 2246 13473 2266
rect 13493 2246 13504 2266
rect 13355 2238 13504 2246
rect 13571 2269 13728 2276
rect 13571 2249 13691 2269
rect 13711 2249 13728 2269
rect 13571 2239 13728 2249
rect 13571 2238 13606 2239
rect 12635 2215 12673 2224
rect 13571 2217 13602 2238
rect 13789 2217 13825 2327
rect 13844 2326 13881 2327
rect 13940 2326 13977 2327
rect 13900 2267 13990 2273
rect 13900 2247 13909 2267
rect 13929 2265 13990 2267
rect 13929 2247 13954 2265
rect 13900 2245 13954 2247
rect 13974 2245 13990 2265
rect 13900 2239 13990 2245
rect 13414 2216 13451 2217
rect 12635 2214 12672 2215
rect 12096 2186 12186 2192
rect 12096 2166 12112 2186
rect 12132 2184 12186 2186
rect 12132 2166 12157 2184
rect 12096 2164 12157 2166
rect 12177 2164 12186 2184
rect 12096 2158 12186 2164
rect 12109 2104 12146 2105
rect 12205 2104 12242 2105
rect 12261 2104 12297 2214
rect 12484 2193 12515 2214
rect 13413 2207 13451 2216
rect 12480 2192 12515 2193
rect 12358 2182 12515 2192
rect 12358 2162 12375 2182
rect 12395 2162 12515 2182
rect 12358 2155 12515 2162
rect 12582 2185 12731 2193
rect 12582 2165 12593 2185
rect 12613 2165 12652 2185
rect 12672 2165 12731 2185
rect 13241 2189 13281 2199
rect 12582 2158 12731 2165
rect 12797 2161 12849 2179
rect 12582 2157 12623 2158
rect 12316 2104 12353 2105
rect 12009 2095 12147 2104
rect 11481 2084 11514 2086
rect 11110 2072 11557 2084
rect 10342 1950 10510 1952
rect 10066 1924 10510 1950
rect 9576 1902 9714 1911
rect 9370 1901 9407 1902
rect 8867 1847 8904 1850
rect 9100 1848 9141 1849
rect 7210 1826 7241 1827
rect 6834 1766 7175 1767
rect 7356 1766 7393 1837
rect 8992 1841 9141 1848
rect 8423 1829 8460 1834
rect 8414 1825 8461 1829
rect 8414 1807 8433 1825
rect 8451 1807 8461 1825
rect 8992 1821 9051 1841
rect 9071 1821 9110 1841
rect 9130 1821 9141 1841
rect 8992 1813 9141 1821
rect 9208 1844 9365 1851
rect 9208 1824 9328 1844
rect 9348 1824 9365 1844
rect 9208 1814 9365 1824
rect 9208 1813 9243 1814
rect 6759 1761 7175 1766
rect 6759 1741 6762 1761
rect 6782 1741 7175 1761
rect 7206 1742 7393 1766
rect 8018 1764 8058 1769
rect 8414 1764 8461 1807
rect 9208 1792 9239 1813
rect 9426 1792 9462 1902
rect 9481 1901 9518 1902
rect 9577 1901 9614 1902
rect 9537 1842 9627 1848
rect 9537 1822 9546 1842
rect 9566 1840 9627 1842
rect 9566 1822 9591 1840
rect 9537 1820 9591 1822
rect 9611 1820 9627 1840
rect 9537 1814 9627 1820
rect 9051 1791 9088 1792
rect 8018 1725 8461 1764
rect 8864 1783 8901 1785
rect 8864 1775 8906 1783
rect 8864 1757 8874 1775
rect 8892 1757 8906 1775
rect 8864 1748 8906 1757
rect 9050 1782 9088 1791
rect 9050 1762 9059 1782
rect 9079 1762 9088 1782
rect 9050 1754 9088 1762
rect 9154 1786 9239 1792
rect 9269 1791 9306 1792
rect 9154 1766 9162 1786
rect 9182 1766 9239 1786
rect 9154 1758 9239 1766
rect 9268 1782 9306 1791
rect 9268 1762 9277 1782
rect 9297 1762 9306 1782
rect 9154 1757 9190 1758
rect 9268 1754 9306 1762
rect 9372 1790 9516 1792
rect 9372 1786 9424 1790
rect 9372 1766 9380 1786
rect 9400 1770 9424 1786
rect 9444 1786 9516 1790
rect 9444 1770 9488 1786
rect 9400 1766 9488 1770
rect 9508 1766 9516 1786
rect 9372 1758 9516 1766
rect 9372 1757 9408 1758
rect 9480 1757 9516 1758
rect 9582 1791 9619 1792
rect 9582 1790 9620 1791
rect 9582 1782 9646 1790
rect 9582 1762 9591 1782
rect 9611 1768 9646 1782
rect 9666 1768 9669 1788
rect 9611 1763 9669 1768
rect 9611 1762 9646 1763
rect 5799 1666 5807 1688
rect 5831 1666 5839 1688
rect 5799 1658 5839 1666
rect 7112 1710 7152 1718
rect 7112 1688 7120 1710
rect 7144 1688 7152 1710
rect 3318 1612 3353 1613
rect 3295 1607 3353 1612
rect 3295 1587 3298 1607
rect 3318 1593 3353 1607
rect 3373 1593 3382 1613
rect 3318 1585 3382 1593
rect 3344 1584 3382 1585
rect 3345 1583 3382 1584
rect 3448 1617 3484 1618
rect 3556 1617 3592 1618
rect 3448 1609 3592 1617
rect 3448 1589 3456 1609
rect 3476 1605 3564 1609
rect 3476 1589 3520 1605
rect 3448 1585 3520 1589
rect 3540 1589 3564 1605
rect 3584 1589 3592 1609
rect 3540 1585 3592 1589
rect 3448 1583 3592 1585
rect 3658 1613 3696 1621
rect 3774 1617 3810 1618
rect 3658 1593 3667 1613
rect 3687 1593 3696 1613
rect 3658 1584 3696 1593
rect 3725 1609 3810 1617
rect 3725 1589 3782 1609
rect 3802 1589 3810 1609
rect 3658 1583 3695 1584
rect 3725 1583 3810 1589
rect 3876 1613 3914 1621
rect 3876 1593 3885 1613
rect 3905 1593 3914 1613
rect 3876 1584 3914 1593
rect 4058 1618 4100 1627
rect 4058 1600 4072 1618
rect 4090 1600 4100 1618
rect 4058 1592 4100 1600
rect 4063 1590 4100 1592
rect 4490 1612 4933 1651
rect 3876 1583 3913 1584
rect 3337 1555 3427 1561
rect 3337 1535 3353 1555
rect 3373 1553 3427 1555
rect 3373 1535 3398 1553
rect 3337 1533 3398 1535
rect 3418 1533 3427 1553
rect 3337 1527 3427 1533
rect 3350 1473 3387 1474
rect 3446 1473 3483 1474
rect 3502 1473 3538 1583
rect 3725 1562 3756 1583
rect 4490 1569 4537 1612
rect 4893 1607 4933 1612
rect 5558 1610 5745 1634
rect 5776 1615 6169 1635
rect 6189 1615 6192 1635
rect 5776 1610 6192 1615
rect 3721 1561 3756 1562
rect 3599 1551 3756 1561
rect 3599 1531 3616 1551
rect 3636 1531 3756 1551
rect 3599 1524 3756 1531
rect 3823 1554 3972 1562
rect 3823 1534 3834 1554
rect 3854 1534 3893 1554
rect 3913 1534 3972 1554
rect 4490 1551 4500 1569
rect 4518 1551 4537 1569
rect 4490 1547 4537 1551
rect 4491 1542 4528 1547
rect 3823 1527 3972 1534
rect 5558 1539 5595 1610
rect 5776 1609 6117 1610
rect 5710 1549 5741 1550
rect 3823 1526 3864 1527
rect 4060 1525 4097 1528
rect 3557 1473 3594 1474
rect 3250 1464 3388 1473
rect 2454 1425 2898 1451
rect 2454 1423 2622 1425
rect 1407 1291 1854 1303
rect 1450 1289 1483 1291
rect 817 1271 955 1280
rect 611 1270 648 1271
rect 341 1217 382 1218
rect 115 1196 167 1214
rect 233 1210 382 1217
rect 233 1190 292 1210
rect 312 1190 351 1210
rect 371 1190 382 1210
rect 233 1182 382 1190
rect 449 1213 606 1220
rect 449 1193 569 1213
rect 589 1193 606 1213
rect 449 1183 606 1193
rect 449 1182 484 1183
rect 449 1161 480 1182
rect 667 1161 703 1271
rect 722 1270 759 1271
rect 818 1270 855 1271
rect 778 1211 868 1217
rect 778 1191 787 1211
rect 807 1209 868 1211
rect 807 1191 832 1209
rect 778 1189 832 1191
rect 852 1189 868 1209
rect 778 1183 868 1189
rect 292 1160 329 1161
rect 291 1151 329 1160
rect 119 1133 159 1143
rect 119 1115 129 1133
rect 147 1115 159 1133
rect 291 1131 300 1151
rect 320 1131 329 1151
rect 291 1123 329 1131
rect 395 1155 480 1161
rect 510 1160 547 1161
rect 395 1135 403 1155
rect 423 1135 480 1155
rect 395 1127 480 1135
rect 509 1151 547 1160
rect 509 1131 518 1151
rect 538 1131 547 1151
rect 395 1126 431 1127
rect 509 1123 547 1131
rect 613 1155 757 1161
rect 613 1135 621 1155
rect 641 1135 674 1155
rect 694 1135 729 1155
rect 749 1135 757 1155
rect 613 1127 757 1135
rect 613 1126 649 1127
rect 721 1126 757 1127
rect 823 1160 860 1161
rect 823 1159 861 1160
rect 823 1151 887 1159
rect 823 1131 832 1151
rect 852 1137 887 1151
rect 907 1137 910 1157
rect 852 1132 910 1137
rect 852 1131 887 1132
rect 119 1059 159 1115
rect 292 1094 329 1123
rect 293 1092 329 1094
rect 293 1070 484 1092
rect 510 1091 547 1123
rect 823 1119 887 1131
rect 927 1093 954 1271
rect 1812 1246 1854 1291
rect 786 1091 954 1093
rect 510 1081 954 1091
rect 1095 1187 1282 1211
rect 1313 1192 1706 1212
rect 1726 1192 1729 1212
rect 1313 1187 1729 1192
rect 1095 1116 1132 1187
rect 1313 1186 1654 1187
rect 1247 1126 1278 1127
rect 1095 1096 1104 1116
rect 1124 1096 1132 1116
rect 1095 1086 1132 1096
rect 1191 1116 1278 1126
rect 1191 1096 1200 1116
rect 1220 1096 1278 1116
rect 1191 1087 1278 1096
rect 1191 1086 1228 1087
rect 116 1054 159 1059
rect 507 1065 954 1081
rect 507 1059 535 1065
rect 786 1064 954 1065
rect 116 1051 266 1054
rect 507 1051 534 1059
rect 116 1049 534 1051
rect 116 1031 125 1049
rect 143 1031 534 1049
rect 1247 1036 1278 1087
rect 1313 1116 1350 1186
rect 1616 1185 1653 1186
rect 1465 1126 1501 1127
rect 1313 1096 1322 1116
rect 1342 1096 1350 1116
rect 1313 1086 1350 1096
rect 1409 1116 1557 1126
rect 1657 1123 1753 1125
rect 1409 1096 1418 1116
rect 1438 1096 1528 1116
rect 1548 1096 1557 1116
rect 1409 1087 1557 1096
rect 1615 1116 1753 1123
rect 1615 1096 1624 1116
rect 1644 1096 1753 1116
rect 1615 1087 1753 1096
rect 1409 1086 1446 1087
rect 1139 1033 1180 1034
rect 116 1028 534 1031
rect 116 1022 159 1028
rect 119 1019 159 1022
rect 1034 1026 1180 1033
rect 516 1010 556 1011
rect 227 993 556 1010
rect 1034 1006 1090 1026
rect 1110 1006 1149 1026
rect 1169 1006 1180 1026
rect 1034 998 1180 1006
rect 1247 1029 1404 1036
rect 1247 1009 1367 1029
rect 1387 1009 1404 1029
rect 1247 999 1404 1009
rect 1247 998 1282 999
rect 111 950 154 961
rect 111 932 123 950
rect 141 932 154 950
rect 111 906 154 932
rect 227 906 254 993
rect 516 984 556 993
rect 111 885 254 906
rect 298 958 332 974
rect 516 964 909 984
rect 929 964 932 984
rect 1247 977 1278 998
rect 1465 977 1501 1087
rect 1520 1086 1557 1087
rect 1616 1086 1653 1087
rect 1576 1027 1666 1033
rect 1576 1007 1585 1027
rect 1605 1025 1666 1027
rect 1605 1007 1630 1025
rect 1576 1005 1630 1007
rect 1650 1005 1666 1025
rect 1576 999 1666 1005
rect 1090 976 1127 977
rect 516 959 932 964
rect 1089 967 1127 976
rect 516 958 857 959
rect 298 888 335 958
rect 450 898 481 899
rect 111 883 248 885
rect 111 841 154 883
rect 298 868 307 888
rect 327 868 335 888
rect 298 858 335 868
rect 394 888 481 898
rect 394 868 403 888
rect 423 868 481 888
rect 394 859 481 868
rect 394 858 431 859
rect 109 831 154 841
rect 109 813 118 831
rect 136 813 154 831
rect 109 807 154 813
rect 450 808 481 859
rect 516 888 553 958
rect 819 957 856 958
rect 1089 947 1098 967
rect 1118 947 1127 967
rect 1089 939 1127 947
rect 1193 971 1278 977
rect 1308 976 1345 977
rect 1193 951 1201 971
rect 1221 951 1278 971
rect 1193 943 1278 951
rect 1307 967 1345 976
rect 1307 947 1316 967
rect 1336 947 1345 967
rect 1193 942 1229 943
rect 1307 939 1345 947
rect 1411 971 1555 977
rect 1411 951 1419 971
rect 1439 968 1527 971
rect 1439 951 1474 968
rect 1411 950 1474 951
rect 1493 951 1527 968
rect 1547 951 1555 971
rect 1493 950 1555 951
rect 1411 943 1555 950
rect 1411 942 1447 943
rect 1519 942 1555 943
rect 1621 976 1658 977
rect 1621 975 1659 976
rect 1681 975 1708 979
rect 1621 973 1708 975
rect 1621 967 1685 973
rect 1621 947 1630 967
rect 1650 953 1685 967
rect 1705 953 1708 973
rect 1650 948 1708 953
rect 1650 947 1685 948
rect 1090 910 1127 939
rect 1091 908 1127 910
rect 668 898 704 899
rect 516 868 525 888
rect 545 868 553 888
rect 516 858 553 868
rect 612 888 760 898
rect 860 895 956 897
rect 612 868 621 888
rect 641 868 731 888
rect 751 868 760 888
rect 612 859 760 868
rect 818 888 956 895
rect 818 868 827 888
rect 847 868 956 888
rect 1091 886 1282 908
rect 1308 907 1345 939
rect 1621 935 1685 947
rect 1725 909 1752 1087
rect 1584 907 1752 909
rect 1308 881 1752 907
rect 818 859 956 868
rect 612 858 649 859
rect 109 804 146 807
rect 342 805 383 806
rect 234 798 383 805
rect 234 778 293 798
rect 313 778 352 798
rect 372 778 383 798
rect 234 770 383 778
rect 450 801 607 808
rect 450 781 570 801
rect 590 781 607 801
rect 450 771 607 781
rect 450 770 485 771
rect 450 749 481 770
rect 668 749 704 859
rect 723 858 760 859
rect 819 858 856 859
rect 779 799 869 805
rect 779 779 788 799
rect 808 797 869 799
rect 808 779 833 797
rect 779 777 833 779
rect 853 777 869 797
rect 779 771 869 777
rect 293 748 330 749
rect 106 740 143 742
rect 106 732 148 740
rect 106 714 116 732
rect 134 714 148 732
rect 106 705 148 714
rect 292 739 330 748
rect 292 719 301 739
rect 321 719 330 739
rect 292 711 330 719
rect 396 743 481 749
rect 511 748 548 749
rect 396 723 404 743
rect 424 723 481 743
rect 396 715 481 723
rect 510 739 548 748
rect 510 719 519 739
rect 539 719 548 739
rect 396 714 432 715
rect 510 711 548 719
rect 614 747 758 749
rect 614 743 666 747
rect 614 723 622 743
rect 642 727 666 743
rect 686 743 758 747
rect 686 727 730 743
rect 642 723 730 727
rect 750 723 758 743
rect 614 715 758 723
rect 614 714 650 715
rect 722 714 758 715
rect 824 748 861 749
rect 824 747 862 748
rect 824 739 888 747
rect 824 719 833 739
rect 853 725 888 739
rect 908 725 911 745
rect 853 720 911 725
rect 853 719 888 720
rect 107 680 148 705
rect 293 680 330 711
rect 511 689 548 711
rect 824 707 888 719
rect 506 680 548 689
rect 928 681 955 859
rect 107 668 152 680
rect 103 610 152 668
rect 293 654 355 680
rect 506 679 591 680
rect 787 679 955 681
rect 506 653 955 679
rect 506 610 545 653
rect 787 652 955 653
rect 1418 657 1458 881
rect 1584 880 1752 881
rect 1816 913 1849 1246
rect 2454 1245 2481 1423
rect 2521 1385 2585 1397
rect 2861 1393 2898 1425
rect 2924 1424 3115 1446
rect 3250 1444 3359 1464
rect 3379 1444 3388 1464
rect 3250 1437 3388 1444
rect 3446 1464 3594 1473
rect 3446 1444 3455 1464
rect 3475 1444 3565 1464
rect 3585 1444 3594 1464
rect 3250 1435 3346 1437
rect 3446 1434 3594 1444
rect 3653 1464 3690 1474
rect 3653 1444 3661 1464
rect 3681 1444 3690 1464
rect 3502 1433 3538 1434
rect 3079 1422 3115 1424
rect 3079 1393 3116 1422
rect 2521 1384 2556 1385
rect 2498 1379 2556 1384
rect 2498 1359 2501 1379
rect 2521 1365 2556 1379
rect 2576 1365 2585 1385
rect 2521 1357 2585 1365
rect 2547 1356 2585 1357
rect 2548 1355 2585 1356
rect 2651 1389 2687 1390
rect 2759 1389 2795 1390
rect 2651 1381 2795 1389
rect 2651 1361 2659 1381
rect 2679 1380 2767 1381
rect 2679 1361 2714 1380
rect 2735 1361 2767 1380
rect 2787 1361 2795 1381
rect 2651 1355 2795 1361
rect 2861 1385 2899 1393
rect 2977 1389 3013 1390
rect 2861 1365 2870 1385
rect 2890 1365 2899 1385
rect 2861 1356 2899 1365
rect 2928 1381 3013 1389
rect 2928 1361 2985 1381
rect 3005 1361 3013 1381
rect 2861 1355 2898 1356
rect 2928 1355 3013 1361
rect 3079 1385 3117 1393
rect 3079 1365 3088 1385
rect 3108 1365 3117 1385
rect 3350 1374 3387 1375
rect 3653 1374 3690 1444
rect 3725 1473 3756 1524
rect 4052 1519 4097 1525
rect 4052 1501 4070 1519
rect 4088 1501 4097 1519
rect 5558 1519 5567 1539
rect 5587 1519 5595 1539
rect 5558 1509 5595 1519
rect 5654 1539 5741 1549
rect 5654 1519 5663 1539
rect 5683 1519 5741 1539
rect 5654 1510 5741 1519
rect 5654 1509 5691 1510
rect 4052 1491 4097 1501
rect 3775 1473 3812 1474
rect 3725 1464 3812 1473
rect 3725 1444 3783 1464
rect 3803 1444 3812 1464
rect 3725 1434 3812 1444
rect 3871 1464 3908 1474
rect 3871 1444 3879 1464
rect 3899 1444 3908 1464
rect 4052 1449 4095 1491
rect 4479 1480 4531 1482
rect 3958 1447 4095 1449
rect 3725 1433 3756 1434
rect 3871 1374 3908 1444
rect 3349 1373 3690 1374
rect 3079 1356 3117 1365
rect 3274 1368 3690 1373
rect 3079 1355 3116 1356
rect 2540 1327 2630 1333
rect 2540 1307 2556 1327
rect 2576 1325 2630 1327
rect 2576 1307 2601 1325
rect 2540 1305 2601 1307
rect 2621 1305 2630 1325
rect 2540 1299 2630 1305
rect 2553 1245 2590 1246
rect 2649 1245 2686 1246
rect 2705 1245 2741 1355
rect 2928 1334 2959 1355
rect 3274 1348 3277 1368
rect 3297 1348 3690 1368
rect 3874 1358 3908 1374
rect 3952 1426 4095 1447
rect 4477 1476 4910 1480
rect 4477 1470 4916 1476
rect 4477 1452 4498 1470
rect 4516 1452 4916 1470
rect 5710 1459 5741 1510
rect 5776 1539 5813 1609
rect 6079 1608 6116 1609
rect 5928 1549 5964 1550
rect 5776 1519 5785 1539
rect 5805 1519 5813 1539
rect 5776 1509 5813 1519
rect 5872 1539 6020 1549
rect 6120 1546 6216 1548
rect 5872 1519 5881 1539
rect 5901 1519 5991 1539
rect 6011 1519 6020 1539
rect 5872 1510 6020 1519
rect 6078 1539 6216 1546
rect 6078 1519 6087 1539
rect 6107 1519 6216 1539
rect 6078 1510 6216 1519
rect 5872 1509 5909 1510
rect 5602 1456 5643 1457
rect 4477 1434 4916 1452
rect 3650 1339 3690 1348
rect 3952 1339 3979 1426
rect 4052 1400 4095 1426
rect 4052 1382 4065 1400
rect 4083 1382 4095 1400
rect 4052 1371 4095 1382
rect 2924 1333 2959 1334
rect 2802 1323 2959 1333
rect 2802 1303 2819 1323
rect 2839 1303 2959 1323
rect 2802 1296 2959 1303
rect 3026 1326 3175 1334
rect 3026 1306 3037 1326
rect 3057 1306 3096 1326
rect 3116 1306 3175 1326
rect 3650 1322 3979 1339
rect 3650 1321 3690 1322
rect 3026 1299 3175 1306
rect 4047 1310 4087 1313
rect 4047 1304 4090 1310
rect 3672 1301 4090 1304
rect 3026 1298 3067 1299
rect 2760 1245 2797 1246
rect 2453 1236 2591 1245
rect 2453 1216 2562 1236
rect 2582 1216 2591 1236
rect 2453 1209 2591 1216
rect 2649 1236 2797 1245
rect 2649 1216 2658 1236
rect 2678 1216 2768 1236
rect 2788 1216 2797 1236
rect 2453 1207 2549 1209
rect 2649 1206 2797 1216
rect 2856 1236 2893 1246
rect 2856 1216 2864 1236
rect 2884 1216 2893 1236
rect 2705 1205 2741 1206
rect 2553 1146 2590 1147
rect 2856 1146 2893 1216
rect 2928 1245 2959 1296
rect 3672 1283 4063 1301
rect 4081 1283 4090 1301
rect 3672 1281 4090 1283
rect 3672 1273 3699 1281
rect 3940 1278 4090 1281
rect 3252 1267 3420 1268
rect 3671 1267 3699 1273
rect 3252 1251 3699 1267
rect 4047 1273 4090 1278
rect 2978 1245 3015 1246
rect 2928 1236 3015 1245
rect 2928 1216 2986 1236
rect 3006 1216 3015 1236
rect 2928 1206 3015 1216
rect 3074 1236 3111 1246
rect 3074 1216 3082 1236
rect 3102 1216 3111 1236
rect 2928 1205 2959 1206
rect 2552 1145 2893 1146
rect 3074 1145 3111 1216
rect 2477 1140 2893 1145
rect 2477 1120 2480 1140
rect 2500 1120 2893 1140
rect 2924 1121 3111 1145
rect 3252 1241 3696 1251
rect 3252 1239 3420 1241
rect 3252 1061 3279 1239
rect 3319 1201 3383 1213
rect 3659 1209 3696 1241
rect 3722 1240 3913 1262
rect 3877 1238 3913 1240
rect 3877 1209 3914 1238
rect 4047 1217 4087 1273
rect 3319 1200 3354 1201
rect 3296 1195 3354 1200
rect 3296 1175 3299 1195
rect 3319 1181 3354 1195
rect 3374 1181 3383 1201
rect 3319 1173 3383 1181
rect 3345 1172 3383 1173
rect 3346 1171 3383 1172
rect 3449 1205 3485 1206
rect 3557 1205 3593 1206
rect 3449 1197 3593 1205
rect 3449 1177 3457 1197
rect 3477 1177 3512 1197
rect 3532 1177 3565 1197
rect 3585 1177 3593 1197
rect 3449 1171 3593 1177
rect 3659 1201 3697 1209
rect 3775 1205 3811 1206
rect 3659 1181 3668 1201
rect 3688 1181 3697 1201
rect 3659 1172 3697 1181
rect 3726 1197 3811 1205
rect 3726 1177 3783 1197
rect 3803 1177 3811 1197
rect 3659 1171 3696 1172
rect 3726 1171 3811 1177
rect 3877 1201 3915 1209
rect 3877 1181 3886 1201
rect 3906 1181 3915 1201
rect 4047 1199 4059 1217
rect 4077 1199 4087 1217
rect 4479 1245 4531 1434
rect 4877 1409 4916 1434
rect 5494 1449 5643 1456
rect 5494 1429 5553 1449
rect 5573 1429 5612 1449
rect 5632 1429 5643 1449
rect 5494 1421 5643 1429
rect 5710 1452 5867 1459
rect 5710 1432 5830 1452
rect 5850 1432 5867 1452
rect 5710 1422 5867 1432
rect 5710 1421 5745 1422
rect 4661 1384 4848 1408
rect 4877 1389 5272 1409
rect 5292 1389 5295 1409
rect 5710 1400 5741 1421
rect 5928 1400 5964 1510
rect 5983 1509 6020 1510
rect 6079 1509 6116 1510
rect 6039 1450 6129 1456
rect 6039 1430 6048 1450
rect 6068 1448 6129 1450
rect 6068 1430 6093 1448
rect 6039 1428 6093 1430
rect 6113 1428 6129 1448
rect 6039 1422 6129 1428
rect 5553 1399 5590 1400
rect 4877 1384 5295 1389
rect 5552 1390 5590 1399
rect 4661 1313 4698 1384
rect 4877 1383 5220 1384
rect 4877 1380 4916 1383
rect 5182 1382 5219 1383
rect 4813 1323 4844 1324
rect 4661 1293 4670 1313
rect 4690 1293 4698 1313
rect 4661 1283 4698 1293
rect 4757 1313 4844 1323
rect 4757 1293 4766 1313
rect 4786 1293 4844 1313
rect 4757 1284 4844 1293
rect 4757 1283 4794 1284
rect 4479 1227 4495 1245
rect 4513 1227 4531 1245
rect 4813 1233 4844 1284
rect 4879 1313 4916 1380
rect 5552 1370 5561 1390
rect 5581 1370 5590 1390
rect 5552 1362 5590 1370
rect 5656 1394 5741 1400
rect 5771 1399 5808 1400
rect 5656 1374 5664 1394
rect 5684 1374 5741 1394
rect 5656 1366 5741 1374
rect 5770 1390 5808 1399
rect 5770 1370 5779 1390
rect 5799 1370 5808 1390
rect 5656 1365 5692 1366
rect 5770 1362 5808 1370
rect 5874 1394 6018 1400
rect 5874 1374 5882 1394
rect 5902 1389 5990 1394
rect 5902 1374 5938 1389
rect 5874 1372 5938 1374
rect 5957 1374 5990 1389
rect 6010 1374 6018 1394
rect 5957 1372 6018 1374
rect 5874 1366 6018 1372
rect 5874 1365 5910 1366
rect 5982 1365 6018 1366
rect 6084 1399 6121 1400
rect 6084 1398 6122 1399
rect 6084 1390 6148 1398
rect 6084 1370 6093 1390
rect 6113 1376 6148 1390
rect 6168 1376 6171 1396
rect 6113 1371 6171 1376
rect 6113 1370 6148 1371
rect 5553 1333 5590 1362
rect 5554 1331 5590 1333
rect 5031 1323 5067 1324
rect 4879 1293 4888 1313
rect 4908 1293 4916 1313
rect 4879 1283 4916 1293
rect 4975 1313 5123 1323
rect 5223 1320 5319 1322
rect 4975 1293 4984 1313
rect 5004 1293 5094 1313
rect 5114 1293 5123 1313
rect 4975 1284 5123 1293
rect 5181 1313 5319 1320
rect 5181 1293 5190 1313
rect 5210 1293 5319 1313
rect 5554 1309 5745 1331
rect 5771 1330 5808 1362
rect 6084 1358 6148 1370
rect 6188 1332 6215 1510
rect 6047 1330 6215 1332
rect 5771 1316 6215 1330
rect 6818 1464 6986 1465
rect 7112 1464 7152 1688
rect 7615 1692 7783 1693
rect 8018 1692 8058 1725
rect 8414 1692 8461 1725
rect 8865 1723 8906 1748
rect 9051 1723 9088 1754
rect 9269 1723 9306 1754
rect 9582 1750 9646 1762
rect 9686 1724 9713 1902
rect 8865 1696 8914 1723
rect 9050 1697 9099 1723
rect 9268 1722 9349 1723
rect 9545 1722 9713 1724
rect 9268 1697 9713 1722
rect 9269 1696 9713 1697
rect 7615 1691 8059 1692
rect 7615 1666 8060 1691
rect 7615 1664 7783 1666
rect 7979 1665 8060 1666
rect 8229 1665 8278 1691
rect 8414 1665 8463 1692
rect 7615 1486 7642 1664
rect 7682 1626 7746 1638
rect 8022 1634 8059 1665
rect 8240 1634 8277 1665
rect 8422 1640 8463 1665
rect 8867 1663 8914 1696
rect 9270 1663 9310 1696
rect 9545 1695 9713 1696
rect 10176 1700 10216 1924
rect 10342 1923 10510 1924
rect 11113 2058 11557 2072
rect 11113 2056 11281 2058
rect 11113 1878 11140 2056
rect 11180 2018 11244 2030
rect 11520 2026 11557 2058
rect 11583 2057 11774 2079
rect 12009 2075 12118 2095
rect 12138 2075 12147 2095
rect 12009 2068 12147 2075
rect 12205 2095 12353 2104
rect 12205 2075 12214 2095
rect 12234 2075 12324 2095
rect 12344 2075 12353 2095
rect 12009 2066 12105 2068
rect 12205 2065 12353 2075
rect 12412 2095 12449 2105
rect 12412 2075 12420 2095
rect 12440 2075 12449 2095
rect 12261 2064 12297 2065
rect 11738 2055 11774 2057
rect 11738 2026 11775 2055
rect 11180 2017 11215 2018
rect 11157 2012 11215 2017
rect 11157 1992 11160 2012
rect 11180 1998 11215 2012
rect 11235 1998 11244 2018
rect 11180 1990 11244 1998
rect 11206 1989 11244 1990
rect 11207 1988 11244 1989
rect 11310 2022 11346 2023
rect 11418 2022 11454 2023
rect 11310 2014 11454 2022
rect 11310 1994 11318 2014
rect 11338 2012 11426 2014
rect 11338 1994 11371 2012
rect 11310 1993 11371 1994
rect 11392 1994 11426 2012
rect 11446 1994 11454 2014
rect 11392 1993 11454 1994
rect 11310 1988 11454 1993
rect 11520 2018 11558 2026
rect 11636 2022 11672 2023
rect 11520 1998 11529 2018
rect 11549 1998 11558 2018
rect 11520 1989 11558 1998
rect 11587 2014 11672 2022
rect 11587 1994 11644 2014
rect 11664 1994 11672 2014
rect 11520 1988 11557 1989
rect 11587 1988 11672 1994
rect 11738 2018 11776 2026
rect 11738 1998 11747 2018
rect 11767 1998 11776 2018
rect 12412 2008 12449 2075
rect 12484 2104 12515 2155
rect 12797 2143 12815 2161
rect 12833 2143 12849 2161
rect 12534 2104 12571 2105
rect 12484 2095 12571 2104
rect 12484 2075 12542 2095
rect 12562 2075 12571 2095
rect 12484 2065 12571 2075
rect 12630 2095 12667 2105
rect 12630 2075 12638 2095
rect 12658 2075 12667 2095
rect 12484 2064 12515 2065
rect 12109 2005 12146 2006
rect 12412 2005 12451 2008
rect 12108 2004 12451 2005
rect 12630 2004 12667 2075
rect 11738 1989 11776 1998
rect 12033 1999 12451 2004
rect 11738 1988 11775 1989
rect 11199 1960 11289 1966
rect 11199 1940 11215 1960
rect 11235 1958 11289 1960
rect 11235 1940 11260 1958
rect 11199 1938 11260 1940
rect 11280 1938 11289 1958
rect 11199 1932 11289 1938
rect 11212 1878 11249 1879
rect 11308 1878 11345 1879
rect 11364 1878 11400 1988
rect 11587 1967 11618 1988
rect 12033 1979 12036 1999
rect 12056 1979 12451 1999
rect 12480 1980 12667 2004
rect 11583 1966 11618 1967
rect 11461 1956 11618 1966
rect 11461 1936 11478 1956
rect 11498 1936 11618 1956
rect 11461 1929 11618 1936
rect 11685 1959 11834 1967
rect 11685 1939 11696 1959
rect 11716 1939 11755 1959
rect 11775 1939 11834 1959
rect 11685 1932 11834 1939
rect 12412 1954 12451 1979
rect 12797 1954 12849 2143
rect 13241 2171 13251 2189
rect 13269 2171 13281 2189
rect 13413 2187 13422 2207
rect 13442 2187 13451 2207
rect 13413 2179 13451 2187
rect 13517 2211 13602 2217
rect 13632 2216 13669 2217
rect 13517 2191 13525 2211
rect 13545 2191 13602 2211
rect 13517 2183 13602 2191
rect 13631 2207 13669 2216
rect 13631 2187 13640 2207
rect 13660 2187 13669 2207
rect 13517 2182 13553 2183
rect 13631 2179 13669 2187
rect 13735 2211 13879 2217
rect 13735 2191 13743 2211
rect 13763 2191 13796 2211
rect 13816 2191 13851 2211
rect 13871 2191 13879 2211
rect 13735 2183 13879 2191
rect 13735 2182 13771 2183
rect 13843 2182 13879 2183
rect 13945 2216 13982 2217
rect 13945 2215 13983 2216
rect 13945 2207 14009 2215
rect 13945 2187 13954 2207
rect 13974 2193 14009 2207
rect 14029 2193 14032 2213
rect 13974 2188 14032 2193
rect 13974 2187 14009 2188
rect 13241 2115 13281 2171
rect 13414 2150 13451 2179
rect 13415 2148 13451 2150
rect 13415 2126 13606 2148
rect 13632 2147 13669 2179
rect 13945 2175 14009 2187
rect 14049 2149 14076 2327
rect 13908 2147 14076 2149
rect 13632 2137 14076 2147
rect 14217 2243 14404 2267
rect 14435 2248 14828 2268
rect 14848 2248 14851 2268
rect 14435 2243 14851 2248
rect 14217 2172 14254 2243
rect 14435 2242 14776 2243
rect 14369 2182 14400 2183
rect 14217 2152 14226 2172
rect 14246 2152 14254 2172
rect 14217 2142 14254 2152
rect 14313 2172 14400 2182
rect 14313 2152 14322 2172
rect 14342 2152 14400 2172
rect 14313 2143 14400 2152
rect 14313 2142 14350 2143
rect 13238 2110 13281 2115
rect 13629 2121 14076 2137
rect 13629 2115 13657 2121
rect 13908 2120 14076 2121
rect 13238 2107 13388 2110
rect 13629 2107 13656 2115
rect 13238 2105 13656 2107
rect 13238 2087 13247 2105
rect 13265 2087 13656 2105
rect 14369 2092 14400 2143
rect 14435 2172 14472 2242
rect 14738 2241 14775 2242
rect 14976 2184 15009 2343
rect 14587 2182 14623 2183
rect 14435 2152 14444 2172
rect 14464 2152 14472 2172
rect 14435 2142 14472 2152
rect 14531 2172 14679 2182
rect 14779 2179 14875 2181
rect 14531 2152 14540 2172
rect 14560 2152 14650 2172
rect 14670 2152 14679 2172
rect 14531 2143 14679 2152
rect 14737 2172 14875 2179
rect 14737 2152 14746 2172
rect 14766 2152 14875 2172
rect 14976 2180 15012 2184
rect 14976 2162 14985 2180
rect 15007 2162 15012 2180
rect 14976 2156 15012 2162
rect 14737 2143 14875 2152
rect 14531 2142 14568 2143
rect 14261 2089 14302 2090
rect 13238 2084 13656 2087
rect 13238 2078 13281 2084
rect 13241 2075 13281 2078
rect 14153 2082 14302 2089
rect 13638 2066 13678 2067
rect 13349 2049 13678 2066
rect 14153 2062 14212 2082
rect 14232 2062 14271 2082
rect 14291 2062 14302 2082
rect 14153 2054 14302 2062
rect 14369 2085 14526 2092
rect 14369 2065 14489 2085
rect 14509 2065 14526 2085
rect 14369 2055 14526 2065
rect 14369 2054 14404 2055
rect 13233 2006 13276 2017
rect 13233 1988 13245 2006
rect 13263 1988 13276 2006
rect 13233 1962 13276 1988
rect 13349 1962 13376 2049
rect 13638 2040 13678 2049
rect 12412 1936 12851 1954
rect 11685 1931 11726 1932
rect 11419 1878 11456 1879
rect 11112 1869 11250 1878
rect 11112 1849 11221 1869
rect 11241 1849 11250 1869
rect 11112 1842 11250 1849
rect 11308 1869 11456 1878
rect 11308 1849 11317 1869
rect 11337 1849 11427 1869
rect 11447 1849 11456 1869
rect 11112 1840 11208 1842
rect 11308 1839 11456 1849
rect 11515 1869 11552 1879
rect 11515 1849 11523 1869
rect 11543 1849 11552 1869
rect 11364 1838 11400 1839
rect 11212 1779 11249 1780
rect 11515 1779 11552 1849
rect 11587 1878 11618 1929
rect 12412 1918 12812 1936
rect 12830 1918 12851 1936
rect 12412 1912 12851 1918
rect 12418 1908 12851 1912
rect 13233 1941 13376 1962
rect 13420 2014 13454 2030
rect 13638 2020 14031 2040
rect 14051 2020 14054 2040
rect 14369 2033 14400 2054
rect 14587 2033 14623 2143
rect 14642 2142 14679 2143
rect 14738 2142 14775 2143
rect 14698 2083 14788 2089
rect 14698 2063 14707 2083
rect 14727 2081 14788 2083
rect 14727 2063 14752 2081
rect 14698 2061 14752 2063
rect 14772 2061 14788 2081
rect 14698 2055 14788 2061
rect 14212 2032 14249 2033
rect 13638 2015 14054 2020
rect 14211 2023 14249 2032
rect 13638 2014 13979 2015
rect 13420 1944 13457 2014
rect 13572 1954 13603 1955
rect 13233 1939 13370 1941
rect 12797 1906 12849 1908
rect 13233 1897 13276 1939
rect 13420 1924 13429 1944
rect 13449 1924 13457 1944
rect 13420 1914 13457 1924
rect 13516 1944 13603 1954
rect 13516 1924 13525 1944
rect 13545 1924 13603 1944
rect 13516 1915 13603 1924
rect 13516 1914 13553 1915
rect 13231 1887 13276 1897
rect 11637 1878 11674 1879
rect 11587 1869 11674 1878
rect 11587 1849 11645 1869
rect 11665 1849 11674 1869
rect 11587 1839 11674 1849
rect 11733 1869 11770 1879
rect 11733 1849 11741 1869
rect 11761 1849 11770 1869
rect 13231 1869 13240 1887
rect 13258 1869 13276 1887
rect 13231 1863 13276 1869
rect 13572 1864 13603 1915
rect 13638 1944 13675 2014
rect 13941 2013 13978 2014
rect 14211 2003 14220 2023
rect 14240 2003 14249 2023
rect 14211 1995 14249 2003
rect 14315 2027 14400 2033
rect 14430 2032 14467 2033
rect 14315 2007 14323 2027
rect 14343 2007 14400 2027
rect 14315 1999 14400 2007
rect 14429 2023 14467 2032
rect 14429 2003 14438 2023
rect 14458 2003 14467 2023
rect 14315 1998 14351 1999
rect 14429 1995 14467 2003
rect 14533 2027 14677 2033
rect 14533 2007 14541 2027
rect 14561 2008 14593 2027
rect 14614 2008 14649 2027
rect 14561 2007 14649 2008
rect 14669 2007 14677 2027
rect 14533 1999 14677 2007
rect 14533 1998 14569 1999
rect 14641 1998 14677 1999
rect 14743 2032 14780 2033
rect 14743 2031 14781 2032
rect 14743 2023 14807 2031
rect 14743 2003 14752 2023
rect 14772 2009 14807 2023
rect 14827 2009 14830 2029
rect 14772 2004 14830 2009
rect 14772 2003 14807 2004
rect 14212 1966 14249 1995
rect 14213 1964 14249 1966
rect 13790 1954 13826 1955
rect 13638 1924 13647 1944
rect 13667 1924 13675 1944
rect 13638 1914 13675 1924
rect 13734 1944 13882 1954
rect 13982 1951 14078 1953
rect 13734 1924 13743 1944
rect 13763 1924 13853 1944
rect 13873 1924 13882 1944
rect 13734 1915 13882 1924
rect 13940 1944 14078 1951
rect 13940 1924 13949 1944
rect 13969 1924 14078 1944
rect 14213 1942 14404 1964
rect 14430 1963 14467 1995
rect 14743 1991 14807 2003
rect 14847 1965 14874 2143
rect 15479 2142 15512 2475
rect 15576 2507 15744 2508
rect 15870 2507 15910 2731
rect 16373 2735 16541 2736
rect 16777 2735 16818 2769
rect 17175 2748 17222 2769
rect 16373 2725 16818 2735
rect 16890 2733 17033 2734
rect 16373 2709 16817 2725
rect 16373 2707 16541 2709
rect 16737 2708 16817 2709
rect 16890 2708 17035 2733
rect 17177 2708 17222 2748
rect 16373 2529 16400 2707
rect 16440 2669 16504 2681
rect 16780 2677 16817 2708
rect 16998 2677 17035 2708
rect 17180 2701 17222 2708
rect 16440 2668 16475 2669
rect 16417 2663 16475 2668
rect 16417 2643 16420 2663
rect 16440 2649 16475 2663
rect 16495 2649 16504 2669
rect 16440 2641 16504 2649
rect 16466 2640 16504 2641
rect 16467 2639 16504 2640
rect 16570 2673 16606 2674
rect 16678 2673 16714 2674
rect 16570 2665 16714 2673
rect 16570 2645 16578 2665
rect 16598 2661 16686 2665
rect 16598 2645 16642 2661
rect 16570 2641 16642 2645
rect 16662 2645 16686 2661
rect 16706 2645 16714 2665
rect 16662 2641 16714 2645
rect 16570 2639 16714 2641
rect 16780 2669 16818 2677
rect 16896 2673 16932 2674
rect 16780 2649 16789 2669
rect 16809 2649 16818 2669
rect 16780 2640 16818 2649
rect 16847 2665 16932 2673
rect 16847 2645 16904 2665
rect 16924 2645 16932 2665
rect 16780 2639 16817 2640
rect 16847 2639 16932 2645
rect 16998 2669 17036 2677
rect 16998 2649 17007 2669
rect 17027 2649 17036 2669
rect 16998 2640 17036 2649
rect 17180 2674 17223 2701
rect 17180 2656 17194 2674
rect 17212 2656 17223 2674
rect 17180 2648 17223 2656
rect 17185 2646 17223 2648
rect 16998 2639 17035 2640
rect 16459 2611 16549 2617
rect 16459 2591 16475 2611
rect 16495 2609 16549 2611
rect 16495 2591 16520 2609
rect 16459 2589 16520 2591
rect 16540 2589 16549 2609
rect 16459 2583 16549 2589
rect 16472 2529 16509 2530
rect 16568 2529 16605 2530
rect 16624 2529 16660 2639
rect 16847 2618 16878 2639
rect 16843 2617 16878 2618
rect 16721 2607 16878 2617
rect 16721 2587 16738 2607
rect 16758 2587 16878 2607
rect 16721 2580 16878 2587
rect 16945 2610 17094 2618
rect 16945 2590 16956 2610
rect 16976 2590 17015 2610
rect 17035 2590 17094 2610
rect 16945 2583 17094 2590
rect 16945 2582 16986 2583
rect 17182 2581 17219 2584
rect 16679 2529 16716 2530
rect 16372 2520 16510 2529
rect 15576 2481 16020 2507
rect 15576 2479 15744 2481
rect 15576 2301 15603 2479
rect 15643 2441 15707 2453
rect 15983 2449 16020 2481
rect 16046 2480 16237 2502
rect 16372 2500 16481 2520
rect 16501 2500 16510 2520
rect 16372 2493 16510 2500
rect 16568 2520 16716 2529
rect 16568 2500 16577 2520
rect 16597 2500 16687 2520
rect 16707 2500 16716 2520
rect 16372 2491 16468 2493
rect 16568 2490 16716 2500
rect 16775 2520 16812 2530
rect 16775 2500 16783 2520
rect 16803 2500 16812 2520
rect 16624 2489 16660 2490
rect 16201 2478 16237 2480
rect 16201 2449 16238 2478
rect 15643 2440 15678 2441
rect 15620 2435 15678 2440
rect 15620 2415 15623 2435
rect 15643 2421 15678 2435
rect 15698 2421 15707 2441
rect 15643 2415 15707 2421
rect 15620 2413 15707 2415
rect 15620 2409 15647 2413
rect 15669 2412 15707 2413
rect 15670 2411 15707 2412
rect 15773 2445 15809 2446
rect 15881 2445 15917 2446
rect 15773 2438 15917 2445
rect 15773 2437 15835 2438
rect 15773 2417 15781 2437
rect 15801 2420 15835 2437
rect 15854 2437 15917 2438
rect 15854 2420 15889 2437
rect 15801 2417 15889 2420
rect 15909 2417 15917 2437
rect 15773 2411 15917 2417
rect 15983 2441 16021 2449
rect 16099 2445 16135 2446
rect 15983 2421 15992 2441
rect 16012 2421 16021 2441
rect 15983 2412 16021 2421
rect 16050 2437 16135 2445
rect 16050 2417 16107 2437
rect 16127 2417 16135 2437
rect 15983 2411 16020 2412
rect 16050 2411 16135 2417
rect 16201 2441 16239 2449
rect 16201 2421 16210 2441
rect 16230 2421 16239 2441
rect 16472 2430 16509 2431
rect 16775 2430 16812 2500
rect 16847 2529 16878 2580
rect 17174 2575 17219 2581
rect 17174 2557 17192 2575
rect 17210 2557 17219 2575
rect 17174 2547 17219 2557
rect 16897 2529 16934 2530
rect 16847 2520 16934 2529
rect 16847 2500 16905 2520
rect 16925 2500 16934 2520
rect 16847 2490 16934 2500
rect 16993 2520 17030 2530
rect 16993 2500 17001 2520
rect 17021 2500 17030 2520
rect 17174 2505 17217 2547
rect 17080 2503 17217 2505
rect 16847 2489 16878 2490
rect 16993 2430 17030 2500
rect 16471 2429 16812 2430
rect 16201 2412 16239 2421
rect 16396 2424 16812 2429
rect 16201 2411 16238 2412
rect 15662 2383 15752 2389
rect 15662 2363 15678 2383
rect 15698 2381 15752 2383
rect 15698 2363 15723 2381
rect 15662 2361 15723 2363
rect 15743 2361 15752 2381
rect 15662 2355 15752 2361
rect 15675 2301 15712 2302
rect 15771 2301 15808 2302
rect 15827 2301 15863 2411
rect 16050 2390 16081 2411
rect 16396 2404 16399 2424
rect 16419 2404 16812 2424
rect 16996 2414 17030 2430
rect 17074 2482 17217 2503
rect 16772 2395 16812 2404
rect 17074 2395 17101 2482
rect 17174 2456 17217 2482
rect 17174 2438 17187 2456
rect 17205 2438 17217 2456
rect 17174 2427 17217 2438
rect 16046 2389 16081 2390
rect 15924 2379 16081 2389
rect 15924 2359 15941 2379
rect 15961 2359 16081 2379
rect 15924 2352 16081 2359
rect 16148 2382 16294 2390
rect 16148 2362 16159 2382
rect 16179 2362 16218 2382
rect 16238 2362 16294 2382
rect 16772 2378 17101 2395
rect 16772 2377 16812 2378
rect 16148 2355 16294 2362
rect 17169 2366 17209 2369
rect 17169 2360 17212 2366
rect 16794 2357 17212 2360
rect 16148 2354 16189 2355
rect 15882 2301 15919 2302
rect 15575 2292 15713 2301
rect 15575 2272 15684 2292
rect 15704 2272 15713 2292
rect 15575 2265 15713 2272
rect 15771 2292 15919 2301
rect 15771 2272 15780 2292
rect 15800 2272 15890 2292
rect 15910 2272 15919 2292
rect 15575 2263 15671 2265
rect 15771 2262 15919 2272
rect 15978 2292 16015 2302
rect 15978 2272 15986 2292
rect 16006 2272 16015 2292
rect 15827 2261 15863 2262
rect 15675 2202 15712 2203
rect 15978 2202 16015 2272
rect 16050 2301 16081 2352
rect 16794 2339 17185 2357
rect 17203 2339 17212 2357
rect 16794 2337 17212 2339
rect 16794 2329 16821 2337
rect 17062 2334 17212 2337
rect 16374 2323 16542 2324
rect 16793 2323 16821 2329
rect 16374 2307 16821 2323
rect 17169 2329 17212 2334
rect 16100 2301 16137 2302
rect 16050 2292 16137 2301
rect 16050 2272 16108 2292
rect 16128 2272 16137 2292
rect 16050 2262 16137 2272
rect 16196 2292 16233 2302
rect 16196 2272 16204 2292
rect 16224 2272 16233 2292
rect 16050 2261 16081 2262
rect 15674 2201 16015 2202
rect 16196 2201 16233 2272
rect 15599 2196 16015 2201
rect 15599 2176 15602 2196
rect 15622 2176 16015 2196
rect 16046 2177 16233 2201
rect 16374 2297 16818 2307
rect 16374 2295 16542 2297
rect 15474 2097 15516 2142
rect 16374 2117 16401 2295
rect 16441 2257 16505 2269
rect 16781 2265 16818 2297
rect 16844 2296 17035 2318
rect 16999 2294 17035 2296
rect 16999 2265 17036 2294
rect 17169 2273 17209 2329
rect 16441 2256 16476 2257
rect 16418 2251 16476 2256
rect 16418 2231 16421 2251
rect 16441 2237 16476 2251
rect 16496 2237 16505 2257
rect 16441 2229 16505 2237
rect 16467 2228 16505 2229
rect 16468 2227 16505 2228
rect 16571 2261 16607 2262
rect 16679 2261 16715 2262
rect 16571 2253 16715 2261
rect 16571 2233 16579 2253
rect 16599 2233 16634 2253
rect 16654 2233 16687 2253
rect 16707 2233 16715 2253
rect 16571 2227 16715 2233
rect 16781 2257 16819 2265
rect 16897 2261 16933 2262
rect 16781 2237 16790 2257
rect 16810 2237 16819 2257
rect 16781 2228 16819 2237
rect 16848 2253 16933 2261
rect 16848 2233 16905 2253
rect 16925 2233 16933 2253
rect 16781 2227 16818 2228
rect 16848 2227 16933 2233
rect 16999 2257 17037 2265
rect 16999 2237 17008 2257
rect 17028 2237 17037 2257
rect 17169 2255 17181 2273
rect 17199 2255 17209 2273
rect 17169 2245 17209 2255
rect 16999 2228 17037 2237
rect 16999 2227 17036 2228
rect 16460 2199 16550 2205
rect 16460 2179 16476 2199
rect 16496 2197 16550 2199
rect 16496 2179 16521 2197
rect 16460 2177 16521 2179
rect 16541 2177 16550 2197
rect 16460 2171 16550 2177
rect 16473 2117 16510 2118
rect 16569 2117 16606 2118
rect 16625 2117 16661 2227
rect 16848 2206 16879 2227
rect 16844 2205 16879 2206
rect 16722 2195 16879 2205
rect 16722 2175 16739 2195
rect 16759 2175 16879 2195
rect 16722 2168 16879 2175
rect 16946 2198 17095 2206
rect 16946 2178 16957 2198
rect 16977 2178 17016 2198
rect 17036 2178 17095 2198
rect 16946 2171 17095 2178
rect 17161 2174 17213 2192
rect 16946 2170 16987 2171
rect 16680 2117 16717 2118
rect 16373 2108 16511 2117
rect 15845 2097 15878 2099
rect 15474 2085 15921 2097
rect 14706 1963 14874 1965
rect 14430 1937 14874 1963
rect 13940 1915 14078 1924
rect 13734 1914 13771 1915
rect 13231 1860 13268 1863
rect 13464 1861 13505 1862
rect 11587 1838 11618 1839
rect 11211 1778 11552 1779
rect 11733 1778 11770 1849
rect 13356 1854 13505 1861
rect 12800 1841 12837 1846
rect 12791 1837 12838 1841
rect 12791 1819 12810 1837
rect 12828 1819 12838 1837
rect 13356 1834 13415 1854
rect 13435 1834 13474 1854
rect 13494 1834 13505 1854
rect 13356 1826 13505 1834
rect 13572 1857 13729 1864
rect 13572 1837 13692 1857
rect 13712 1837 13729 1857
rect 13572 1827 13729 1837
rect 13572 1826 13607 1827
rect 11136 1773 11552 1778
rect 11136 1753 11139 1773
rect 11159 1753 11552 1773
rect 11583 1754 11770 1778
rect 12395 1776 12435 1781
rect 12791 1776 12838 1819
rect 13572 1805 13603 1826
rect 13790 1805 13826 1915
rect 13845 1914 13882 1915
rect 13941 1914 13978 1915
rect 13901 1855 13991 1861
rect 13901 1835 13910 1855
rect 13930 1853 13991 1855
rect 13930 1835 13955 1853
rect 13901 1833 13955 1835
rect 13975 1833 13991 1853
rect 13901 1827 13991 1833
rect 13415 1804 13452 1805
rect 12395 1737 12838 1776
rect 13228 1796 13265 1798
rect 13228 1788 13270 1796
rect 13228 1770 13238 1788
rect 13256 1770 13270 1788
rect 13228 1761 13270 1770
rect 13414 1795 13452 1804
rect 13414 1775 13423 1795
rect 13443 1775 13452 1795
rect 13414 1767 13452 1775
rect 13518 1799 13603 1805
rect 13633 1804 13670 1805
rect 13518 1779 13526 1799
rect 13546 1779 13603 1799
rect 13518 1771 13603 1779
rect 13632 1795 13670 1804
rect 13632 1775 13641 1795
rect 13661 1775 13670 1795
rect 13518 1770 13554 1771
rect 13632 1767 13670 1775
rect 13736 1803 13880 1805
rect 13736 1799 13788 1803
rect 13736 1779 13744 1799
rect 13764 1783 13788 1799
rect 13808 1799 13880 1803
rect 13808 1783 13852 1799
rect 13764 1779 13852 1783
rect 13872 1779 13880 1799
rect 13736 1771 13880 1779
rect 13736 1770 13772 1771
rect 13844 1770 13880 1771
rect 13946 1804 13983 1805
rect 13946 1803 13984 1804
rect 13946 1795 14010 1803
rect 13946 1775 13955 1795
rect 13975 1781 14010 1795
rect 14030 1781 14033 1801
rect 13975 1776 14033 1781
rect 13975 1775 14010 1776
rect 10176 1678 10184 1700
rect 10208 1678 10216 1700
rect 10176 1670 10216 1678
rect 11489 1722 11529 1730
rect 11489 1700 11497 1722
rect 11521 1700 11529 1722
rect 7682 1625 7717 1626
rect 7659 1620 7717 1625
rect 7659 1600 7662 1620
rect 7682 1606 7717 1620
rect 7737 1606 7746 1626
rect 7682 1598 7746 1606
rect 7708 1597 7746 1598
rect 7709 1596 7746 1597
rect 7812 1630 7848 1631
rect 7920 1630 7956 1631
rect 7812 1622 7956 1630
rect 7812 1602 7820 1622
rect 7840 1618 7928 1622
rect 7840 1602 7884 1618
rect 7812 1598 7884 1602
rect 7904 1602 7928 1618
rect 7948 1602 7956 1622
rect 7904 1598 7956 1602
rect 7812 1596 7956 1598
rect 8022 1626 8060 1634
rect 8138 1630 8174 1631
rect 8022 1606 8031 1626
rect 8051 1606 8060 1626
rect 8022 1597 8060 1606
rect 8089 1622 8174 1630
rect 8089 1602 8146 1622
rect 8166 1602 8174 1622
rect 8022 1596 8059 1597
rect 8089 1596 8174 1602
rect 8240 1626 8278 1634
rect 8240 1606 8249 1626
rect 8269 1606 8278 1626
rect 8240 1597 8278 1606
rect 8422 1631 8464 1640
rect 8422 1613 8436 1631
rect 8454 1613 8464 1631
rect 8422 1605 8464 1613
rect 8427 1603 8464 1605
rect 8867 1624 9310 1663
rect 8240 1596 8277 1597
rect 7701 1568 7791 1574
rect 7701 1548 7717 1568
rect 7737 1566 7791 1568
rect 7737 1548 7762 1566
rect 7701 1546 7762 1548
rect 7782 1546 7791 1566
rect 7701 1540 7791 1546
rect 7714 1486 7751 1487
rect 7810 1486 7847 1487
rect 7866 1486 7902 1596
rect 8089 1575 8120 1596
rect 8867 1581 8914 1624
rect 9270 1619 9310 1624
rect 9935 1622 10122 1646
rect 10153 1627 10546 1647
rect 10566 1627 10569 1647
rect 10153 1622 10569 1627
rect 8085 1574 8120 1575
rect 7963 1564 8120 1574
rect 7963 1544 7980 1564
rect 8000 1544 8120 1564
rect 7963 1537 8120 1544
rect 8187 1567 8336 1575
rect 8187 1547 8198 1567
rect 8218 1547 8257 1567
rect 8277 1547 8336 1567
rect 8867 1563 8877 1581
rect 8895 1563 8914 1581
rect 8867 1559 8914 1563
rect 8868 1554 8905 1559
rect 8187 1540 8336 1547
rect 9935 1551 9972 1622
rect 10153 1621 10494 1622
rect 10087 1561 10118 1562
rect 8187 1539 8228 1540
rect 8424 1538 8461 1541
rect 7921 1486 7958 1487
rect 7614 1477 7752 1486
rect 6818 1438 7262 1464
rect 6818 1436 6986 1438
rect 5771 1304 6218 1316
rect 5814 1302 5847 1304
rect 5181 1284 5319 1293
rect 4975 1283 5012 1284
rect 4705 1230 4746 1231
rect 4479 1209 4531 1227
rect 4597 1223 4746 1230
rect 4047 1189 4087 1199
rect 4597 1203 4656 1223
rect 4676 1203 4715 1223
rect 4735 1203 4746 1223
rect 4597 1195 4746 1203
rect 4813 1226 4970 1233
rect 4813 1206 4933 1226
rect 4953 1206 4970 1226
rect 4813 1196 4970 1206
rect 4813 1195 4848 1196
rect 3877 1172 3915 1181
rect 4813 1174 4844 1195
rect 5031 1174 5067 1284
rect 5086 1283 5123 1284
rect 5182 1283 5219 1284
rect 5142 1224 5232 1230
rect 5142 1204 5151 1224
rect 5171 1222 5232 1224
rect 5171 1204 5196 1222
rect 5142 1202 5196 1204
rect 5216 1202 5232 1222
rect 5142 1196 5232 1202
rect 4656 1173 4693 1174
rect 3877 1171 3914 1172
rect 3338 1143 3428 1149
rect 3338 1123 3354 1143
rect 3374 1141 3428 1143
rect 3374 1123 3399 1141
rect 3338 1121 3399 1123
rect 3419 1121 3428 1141
rect 3338 1115 3428 1121
rect 3351 1061 3388 1062
rect 3447 1061 3484 1062
rect 3503 1061 3539 1171
rect 3726 1150 3757 1171
rect 4655 1164 4693 1173
rect 3722 1149 3757 1150
rect 3600 1139 3757 1149
rect 3600 1119 3617 1139
rect 3637 1119 3757 1139
rect 3600 1112 3757 1119
rect 3824 1142 3973 1150
rect 3824 1122 3835 1142
rect 3855 1122 3894 1142
rect 3914 1122 3973 1142
rect 4483 1146 4523 1156
rect 3824 1115 3973 1122
rect 4039 1118 4091 1136
rect 3824 1114 3865 1115
rect 3558 1061 3595 1062
rect 3251 1052 3389 1061
rect 3251 1032 3360 1052
rect 3380 1032 3389 1052
rect 3251 1025 3389 1032
rect 3447 1052 3595 1061
rect 3447 1032 3456 1052
rect 3476 1032 3566 1052
rect 3586 1032 3595 1052
rect 3251 1023 3347 1025
rect 3447 1022 3595 1032
rect 3654 1052 3691 1062
rect 3654 1032 3662 1052
rect 3682 1032 3691 1052
rect 3503 1021 3539 1022
rect 3654 965 3691 1032
rect 3726 1061 3757 1112
rect 4039 1100 4057 1118
rect 4075 1100 4091 1118
rect 3776 1061 3813 1062
rect 3726 1052 3813 1061
rect 3726 1032 3784 1052
rect 3804 1032 3813 1052
rect 3726 1022 3813 1032
rect 3872 1052 3909 1062
rect 3872 1032 3880 1052
rect 3900 1032 3909 1052
rect 3726 1021 3757 1022
rect 3351 962 3388 963
rect 3654 962 3693 965
rect 3350 961 3693 962
rect 3872 961 3909 1032
rect 3275 956 3693 961
rect 3275 936 3278 956
rect 3298 936 3693 956
rect 3722 937 3909 961
rect 1816 905 1853 913
rect 1816 886 1824 905
rect 1845 886 1853 905
rect 1816 880 1853 886
rect 3654 911 3693 936
rect 4039 911 4091 1100
rect 4483 1128 4493 1146
rect 4511 1128 4523 1146
rect 4655 1144 4664 1164
rect 4684 1144 4693 1164
rect 4655 1136 4693 1144
rect 4759 1168 4844 1174
rect 4874 1173 4911 1174
rect 4759 1148 4767 1168
rect 4787 1148 4844 1168
rect 4759 1140 4844 1148
rect 4873 1164 4911 1173
rect 4873 1144 4882 1164
rect 4902 1144 4911 1164
rect 4759 1139 4795 1140
rect 4873 1136 4911 1144
rect 4977 1168 5121 1174
rect 4977 1148 4985 1168
rect 5005 1148 5038 1168
rect 5058 1148 5093 1168
rect 5113 1148 5121 1168
rect 4977 1140 5121 1148
rect 4977 1139 5013 1140
rect 5085 1139 5121 1140
rect 5187 1173 5224 1174
rect 5187 1172 5225 1173
rect 5187 1164 5251 1172
rect 5187 1144 5196 1164
rect 5216 1150 5251 1164
rect 5271 1150 5274 1170
rect 5216 1145 5274 1150
rect 5216 1144 5251 1145
rect 4483 1072 4523 1128
rect 4656 1107 4693 1136
rect 4657 1105 4693 1107
rect 4657 1083 4848 1105
rect 4874 1104 4911 1136
rect 5187 1132 5251 1144
rect 5291 1106 5318 1284
rect 6176 1259 6218 1304
rect 5150 1104 5318 1106
rect 4874 1094 5318 1104
rect 5459 1200 5646 1224
rect 5677 1205 6070 1225
rect 6090 1205 6093 1225
rect 5677 1200 6093 1205
rect 5459 1129 5496 1200
rect 5677 1199 6018 1200
rect 5611 1139 5642 1140
rect 5459 1109 5468 1129
rect 5488 1109 5496 1129
rect 5459 1099 5496 1109
rect 5555 1129 5642 1139
rect 5555 1109 5564 1129
rect 5584 1109 5642 1129
rect 5555 1100 5642 1109
rect 5555 1099 5592 1100
rect 4480 1067 4523 1072
rect 4871 1078 5318 1094
rect 4871 1072 4899 1078
rect 5150 1077 5318 1078
rect 4480 1064 4630 1067
rect 4871 1064 4898 1072
rect 4480 1062 4898 1064
rect 4480 1044 4489 1062
rect 4507 1044 4898 1062
rect 5611 1049 5642 1100
rect 5677 1129 5714 1199
rect 5980 1198 6017 1199
rect 5829 1139 5865 1140
rect 5677 1109 5686 1129
rect 5706 1109 5714 1129
rect 5677 1099 5714 1109
rect 5773 1129 5921 1139
rect 6021 1136 6117 1138
rect 5773 1109 5782 1129
rect 5802 1109 5892 1129
rect 5912 1109 5921 1129
rect 5773 1100 5921 1109
rect 5979 1129 6117 1136
rect 5979 1109 5988 1129
rect 6008 1109 6117 1129
rect 5979 1100 6117 1109
rect 5773 1099 5810 1100
rect 5503 1046 5544 1047
rect 4480 1041 4898 1044
rect 4480 1035 4523 1041
rect 4483 1032 4523 1035
rect 5398 1039 5544 1046
rect 4880 1023 4920 1024
rect 4591 1006 4920 1023
rect 5398 1019 5454 1039
rect 5474 1019 5513 1039
rect 5533 1019 5544 1039
rect 5398 1011 5544 1019
rect 5611 1042 5768 1049
rect 5611 1022 5731 1042
rect 5751 1022 5768 1042
rect 5611 1012 5768 1022
rect 5611 1011 5646 1012
rect 4475 963 4518 974
rect 4475 945 4487 963
rect 4505 945 4518 963
rect 4475 919 4518 945
rect 4591 919 4618 1006
rect 4880 997 4920 1006
rect 3654 893 4093 911
rect 3654 875 4054 893
rect 4072 875 4093 893
rect 3654 869 4093 875
rect 3660 865 4093 869
rect 4475 898 4618 919
rect 4662 971 4696 987
rect 4880 977 5273 997
rect 5293 977 5296 997
rect 5611 990 5642 1011
rect 5829 990 5865 1100
rect 5884 1099 5921 1100
rect 5980 1099 6017 1100
rect 5940 1040 6030 1046
rect 5940 1020 5949 1040
rect 5969 1038 6030 1040
rect 5969 1020 5994 1038
rect 5940 1018 5994 1020
rect 6014 1018 6030 1038
rect 5940 1012 6030 1018
rect 5454 989 5491 990
rect 4880 972 5296 977
rect 5453 980 5491 989
rect 4880 971 5221 972
rect 4662 901 4699 971
rect 4814 911 4845 912
rect 4475 896 4612 898
rect 4039 863 4091 865
rect 4475 854 4518 896
rect 4662 881 4671 901
rect 4691 881 4699 901
rect 4662 871 4699 881
rect 4758 901 4845 911
rect 4758 881 4767 901
rect 4787 881 4845 901
rect 4758 872 4845 881
rect 4758 871 4795 872
rect 4473 844 4518 854
rect 4473 826 4482 844
rect 4500 826 4518 844
rect 4473 820 4518 826
rect 4814 821 4845 872
rect 4880 901 4917 971
rect 5183 970 5220 971
rect 5453 960 5462 980
rect 5482 960 5491 980
rect 5453 952 5491 960
rect 5557 984 5642 990
rect 5672 989 5709 990
rect 5557 964 5565 984
rect 5585 964 5642 984
rect 5557 956 5642 964
rect 5671 980 5709 989
rect 5671 960 5680 980
rect 5700 960 5709 980
rect 5557 955 5593 956
rect 5671 952 5709 960
rect 5775 984 5919 990
rect 5775 964 5783 984
rect 5803 981 5891 984
rect 5803 964 5838 981
rect 5775 963 5838 964
rect 5857 964 5891 981
rect 5911 964 5919 984
rect 5857 963 5919 964
rect 5775 956 5919 963
rect 5775 955 5811 956
rect 5883 955 5919 956
rect 5985 989 6022 990
rect 5985 988 6023 989
rect 6045 988 6072 992
rect 5985 986 6072 988
rect 5985 980 6049 986
rect 5985 960 5994 980
rect 6014 966 6049 980
rect 6069 966 6072 986
rect 6014 961 6072 966
rect 6014 960 6049 961
rect 5454 923 5491 952
rect 5455 921 5491 923
rect 5032 911 5068 912
rect 4880 881 4889 901
rect 4909 881 4917 901
rect 4880 871 4917 881
rect 4976 901 5124 911
rect 5224 908 5320 910
rect 4976 881 4985 901
rect 5005 881 5095 901
rect 5115 881 5124 901
rect 4976 872 5124 881
rect 5182 901 5320 908
rect 5182 881 5191 901
rect 5211 881 5320 901
rect 5455 899 5646 921
rect 5672 920 5709 952
rect 5985 948 6049 960
rect 6089 922 6116 1100
rect 5948 920 6116 922
rect 5672 894 6116 920
rect 5182 872 5320 881
rect 4976 871 5013 872
rect 4473 817 4510 820
rect 4706 818 4747 819
rect 4598 811 4747 818
rect 4042 798 4079 803
rect 4033 794 4080 798
rect 4033 776 4052 794
rect 4070 776 4080 794
rect 4598 791 4657 811
rect 4677 791 4716 811
rect 4736 791 4747 811
rect 4598 783 4747 791
rect 4814 814 4971 821
rect 4814 794 4934 814
rect 4954 794 4971 814
rect 4814 784 4971 794
rect 4814 783 4849 784
rect 4033 713 4080 776
rect 4814 762 4845 783
rect 5032 762 5068 872
rect 5087 871 5124 872
rect 5183 871 5220 872
rect 5143 812 5233 818
rect 5143 792 5152 812
rect 5172 810 5233 812
rect 5172 792 5197 810
rect 5143 790 5197 792
rect 5217 790 5233 810
rect 5143 784 5233 790
rect 4657 761 4694 762
rect 4470 753 4507 755
rect 4470 745 4512 753
rect 4470 727 4480 745
rect 4498 727 4512 745
rect 4470 718 4512 727
rect 4656 752 4694 761
rect 4656 732 4665 752
rect 4685 732 4694 752
rect 4656 724 4694 732
rect 4760 756 4845 762
rect 4875 761 4912 762
rect 4760 736 4768 756
rect 4788 736 4845 756
rect 4760 728 4845 736
rect 4874 752 4912 761
rect 4874 732 4883 752
rect 4903 732 4912 752
rect 4760 727 4796 728
rect 4874 724 4912 732
rect 4978 760 5122 762
rect 4978 756 5030 760
rect 4978 736 4986 756
rect 5006 740 5030 756
rect 5050 756 5122 760
rect 5050 740 5094 756
rect 5006 736 5094 740
rect 5114 736 5122 756
rect 4978 728 5122 736
rect 4978 727 5014 728
rect 5086 727 5122 728
rect 5188 761 5225 762
rect 5188 760 5226 761
rect 5188 752 5252 760
rect 5188 732 5197 752
rect 5217 738 5252 752
rect 5272 738 5275 758
rect 5217 733 5275 738
rect 5217 732 5252 733
rect 4033 698 4083 713
rect 4033 673 4047 698
rect 4079 673 4083 698
rect 4471 693 4512 718
rect 4657 693 4694 724
rect 4875 702 4912 724
rect 5188 720 5252 732
rect 4870 693 4912 702
rect 5292 694 5319 872
rect 4471 681 4516 693
rect 4033 660 4080 673
rect 1418 635 1426 657
rect 1450 635 1458 657
rect 1418 627 1458 635
rect 4467 623 4516 681
rect 4657 667 4719 693
rect 4870 692 4955 693
rect 5151 692 5319 694
rect 4870 666 5319 692
rect 4870 623 4909 666
rect 5151 665 5319 666
rect 5782 670 5822 894
rect 5948 893 6116 894
rect 6180 926 6213 1259
rect 6818 1258 6845 1436
rect 6885 1398 6949 1410
rect 7225 1406 7262 1438
rect 7288 1437 7479 1459
rect 7614 1457 7723 1477
rect 7743 1457 7752 1477
rect 7614 1450 7752 1457
rect 7810 1477 7958 1486
rect 7810 1457 7819 1477
rect 7839 1457 7929 1477
rect 7949 1457 7958 1477
rect 7614 1448 7710 1450
rect 7810 1447 7958 1457
rect 8017 1477 8054 1487
rect 8017 1457 8025 1477
rect 8045 1457 8054 1477
rect 7866 1446 7902 1447
rect 7443 1435 7479 1437
rect 7443 1406 7480 1435
rect 6885 1397 6920 1398
rect 6862 1392 6920 1397
rect 6862 1372 6865 1392
rect 6885 1378 6920 1392
rect 6940 1378 6949 1398
rect 6885 1370 6949 1378
rect 6911 1369 6949 1370
rect 6912 1368 6949 1369
rect 7015 1402 7051 1403
rect 7123 1402 7159 1403
rect 7015 1394 7159 1402
rect 7015 1374 7023 1394
rect 7043 1393 7131 1394
rect 7043 1374 7078 1393
rect 7099 1374 7131 1393
rect 7151 1374 7159 1394
rect 7015 1368 7159 1374
rect 7225 1398 7263 1406
rect 7341 1402 7377 1403
rect 7225 1378 7234 1398
rect 7254 1378 7263 1398
rect 7225 1369 7263 1378
rect 7292 1394 7377 1402
rect 7292 1374 7349 1394
rect 7369 1374 7377 1394
rect 7225 1368 7262 1369
rect 7292 1368 7377 1374
rect 7443 1398 7481 1406
rect 7443 1378 7452 1398
rect 7472 1378 7481 1398
rect 7714 1387 7751 1388
rect 8017 1387 8054 1457
rect 8089 1486 8120 1537
rect 8416 1532 8461 1538
rect 8416 1514 8434 1532
rect 8452 1514 8461 1532
rect 9935 1531 9944 1551
rect 9964 1531 9972 1551
rect 9935 1521 9972 1531
rect 10031 1551 10118 1561
rect 10031 1531 10040 1551
rect 10060 1531 10118 1551
rect 10031 1522 10118 1531
rect 10031 1521 10068 1522
rect 8416 1504 8461 1514
rect 8139 1486 8176 1487
rect 8089 1477 8176 1486
rect 8089 1457 8147 1477
rect 8167 1457 8176 1477
rect 8089 1447 8176 1457
rect 8235 1477 8272 1487
rect 8235 1457 8243 1477
rect 8263 1457 8272 1477
rect 8416 1462 8459 1504
rect 8856 1492 8908 1494
rect 8322 1460 8459 1462
rect 8089 1446 8120 1447
rect 8235 1387 8272 1457
rect 7713 1386 8054 1387
rect 7443 1369 7481 1378
rect 7638 1381 8054 1386
rect 7443 1368 7480 1369
rect 6904 1340 6994 1346
rect 6904 1320 6920 1340
rect 6940 1338 6994 1340
rect 6940 1320 6965 1338
rect 6904 1318 6965 1320
rect 6985 1318 6994 1338
rect 6904 1312 6994 1318
rect 6917 1258 6954 1259
rect 7013 1258 7050 1259
rect 7069 1258 7105 1368
rect 7292 1347 7323 1368
rect 7638 1361 7641 1381
rect 7661 1361 8054 1381
rect 8238 1371 8272 1387
rect 8316 1439 8459 1460
rect 8854 1488 9287 1492
rect 8854 1482 9293 1488
rect 8854 1464 8875 1482
rect 8893 1464 9293 1482
rect 10087 1471 10118 1522
rect 10153 1551 10190 1621
rect 10456 1620 10493 1621
rect 10305 1561 10341 1562
rect 10153 1531 10162 1551
rect 10182 1531 10190 1551
rect 10153 1521 10190 1531
rect 10249 1551 10397 1561
rect 10497 1558 10593 1560
rect 10249 1531 10258 1551
rect 10278 1531 10368 1551
rect 10388 1531 10397 1551
rect 10249 1522 10397 1531
rect 10455 1551 10593 1558
rect 10455 1531 10464 1551
rect 10484 1531 10593 1551
rect 10455 1522 10593 1531
rect 10249 1521 10286 1522
rect 9979 1468 10020 1469
rect 8854 1446 9293 1464
rect 8014 1352 8054 1361
rect 8316 1352 8343 1439
rect 8416 1413 8459 1439
rect 8416 1395 8429 1413
rect 8447 1395 8459 1413
rect 8416 1384 8459 1395
rect 7288 1346 7323 1347
rect 7166 1336 7323 1346
rect 7166 1316 7183 1336
rect 7203 1316 7323 1336
rect 7166 1309 7323 1316
rect 7390 1339 7539 1347
rect 7390 1319 7401 1339
rect 7421 1319 7460 1339
rect 7480 1319 7539 1339
rect 8014 1335 8343 1352
rect 8014 1334 8054 1335
rect 7390 1312 7539 1319
rect 8411 1323 8451 1326
rect 8411 1317 8454 1323
rect 8036 1314 8454 1317
rect 7390 1311 7431 1312
rect 7124 1258 7161 1259
rect 6817 1249 6955 1258
rect 6817 1229 6926 1249
rect 6946 1229 6955 1249
rect 6817 1222 6955 1229
rect 7013 1249 7161 1258
rect 7013 1229 7022 1249
rect 7042 1229 7132 1249
rect 7152 1229 7161 1249
rect 6817 1220 6913 1222
rect 7013 1219 7161 1229
rect 7220 1249 7257 1259
rect 7220 1229 7228 1249
rect 7248 1229 7257 1249
rect 7069 1218 7105 1219
rect 6917 1159 6954 1160
rect 7220 1159 7257 1229
rect 7292 1258 7323 1309
rect 8036 1296 8427 1314
rect 8445 1296 8454 1314
rect 8036 1294 8454 1296
rect 8036 1286 8063 1294
rect 8304 1291 8454 1294
rect 7616 1280 7784 1281
rect 8035 1280 8063 1286
rect 7616 1264 8063 1280
rect 8411 1286 8454 1291
rect 7342 1258 7379 1259
rect 7292 1249 7379 1258
rect 7292 1229 7350 1249
rect 7370 1229 7379 1249
rect 7292 1219 7379 1229
rect 7438 1249 7475 1259
rect 7438 1229 7446 1249
rect 7466 1229 7475 1249
rect 7292 1218 7323 1219
rect 6916 1158 7257 1159
rect 7438 1158 7475 1229
rect 6841 1153 7257 1158
rect 6841 1133 6844 1153
rect 6864 1133 7257 1153
rect 7288 1134 7475 1158
rect 7616 1254 8060 1264
rect 7616 1252 7784 1254
rect 7616 1074 7643 1252
rect 7683 1214 7747 1226
rect 8023 1222 8060 1254
rect 8086 1253 8277 1275
rect 8241 1251 8277 1253
rect 8241 1222 8278 1251
rect 8411 1230 8451 1286
rect 7683 1213 7718 1214
rect 7660 1208 7718 1213
rect 7660 1188 7663 1208
rect 7683 1194 7718 1208
rect 7738 1194 7747 1214
rect 7683 1186 7747 1194
rect 7709 1185 7747 1186
rect 7710 1184 7747 1185
rect 7813 1218 7849 1219
rect 7921 1218 7957 1219
rect 7813 1210 7957 1218
rect 7813 1190 7821 1210
rect 7841 1190 7876 1210
rect 7896 1190 7929 1210
rect 7949 1190 7957 1210
rect 7813 1184 7957 1190
rect 8023 1214 8061 1222
rect 8139 1218 8175 1219
rect 8023 1194 8032 1214
rect 8052 1194 8061 1214
rect 8023 1185 8061 1194
rect 8090 1210 8175 1218
rect 8090 1190 8147 1210
rect 8167 1190 8175 1210
rect 8023 1184 8060 1185
rect 8090 1184 8175 1190
rect 8241 1214 8279 1222
rect 8241 1194 8250 1214
rect 8270 1194 8279 1214
rect 8411 1212 8423 1230
rect 8441 1212 8451 1230
rect 8856 1257 8908 1446
rect 9254 1421 9293 1446
rect 9871 1461 10020 1468
rect 9871 1441 9930 1461
rect 9950 1441 9989 1461
rect 10009 1441 10020 1461
rect 9871 1433 10020 1441
rect 10087 1464 10244 1471
rect 10087 1444 10207 1464
rect 10227 1444 10244 1464
rect 10087 1434 10244 1444
rect 10087 1433 10122 1434
rect 9038 1396 9225 1420
rect 9254 1401 9649 1421
rect 9669 1401 9672 1421
rect 10087 1412 10118 1433
rect 10305 1412 10341 1522
rect 10360 1521 10397 1522
rect 10456 1521 10493 1522
rect 10416 1462 10506 1468
rect 10416 1442 10425 1462
rect 10445 1460 10506 1462
rect 10445 1442 10470 1460
rect 10416 1440 10470 1442
rect 10490 1440 10506 1460
rect 10416 1434 10506 1440
rect 9930 1411 9967 1412
rect 9254 1396 9672 1401
rect 9929 1402 9967 1411
rect 9038 1325 9075 1396
rect 9254 1395 9597 1396
rect 9254 1392 9293 1395
rect 9559 1394 9596 1395
rect 9190 1335 9221 1336
rect 9038 1305 9047 1325
rect 9067 1305 9075 1325
rect 9038 1295 9075 1305
rect 9134 1325 9221 1335
rect 9134 1305 9143 1325
rect 9163 1305 9221 1325
rect 9134 1296 9221 1305
rect 9134 1295 9171 1296
rect 8856 1239 8872 1257
rect 8890 1239 8908 1257
rect 9190 1245 9221 1296
rect 9256 1325 9293 1392
rect 9929 1382 9938 1402
rect 9958 1382 9967 1402
rect 9929 1374 9967 1382
rect 10033 1406 10118 1412
rect 10148 1411 10185 1412
rect 10033 1386 10041 1406
rect 10061 1386 10118 1406
rect 10033 1378 10118 1386
rect 10147 1402 10185 1411
rect 10147 1382 10156 1402
rect 10176 1382 10185 1402
rect 10033 1377 10069 1378
rect 10147 1374 10185 1382
rect 10251 1406 10395 1412
rect 10251 1386 10259 1406
rect 10279 1401 10367 1406
rect 10279 1386 10315 1401
rect 10251 1384 10315 1386
rect 10334 1386 10367 1401
rect 10387 1386 10395 1406
rect 10334 1384 10395 1386
rect 10251 1378 10395 1384
rect 10251 1377 10287 1378
rect 10359 1377 10395 1378
rect 10461 1411 10498 1412
rect 10461 1410 10499 1411
rect 10461 1402 10525 1410
rect 10461 1382 10470 1402
rect 10490 1388 10525 1402
rect 10545 1388 10548 1408
rect 10490 1383 10548 1388
rect 10490 1382 10525 1383
rect 9930 1345 9967 1374
rect 9931 1343 9967 1345
rect 9408 1335 9444 1336
rect 9256 1305 9265 1325
rect 9285 1305 9293 1325
rect 9256 1295 9293 1305
rect 9352 1325 9500 1335
rect 9600 1332 9696 1334
rect 9352 1305 9361 1325
rect 9381 1305 9471 1325
rect 9491 1305 9500 1325
rect 9352 1296 9500 1305
rect 9558 1325 9696 1332
rect 9558 1305 9567 1325
rect 9587 1305 9696 1325
rect 9931 1321 10122 1343
rect 10148 1342 10185 1374
rect 10461 1370 10525 1382
rect 10565 1344 10592 1522
rect 10424 1342 10592 1344
rect 10148 1328 10592 1342
rect 11195 1476 11363 1477
rect 11489 1476 11529 1700
rect 11992 1704 12160 1705
rect 12395 1704 12435 1737
rect 12791 1704 12838 1737
rect 13229 1736 13270 1761
rect 13415 1736 13452 1767
rect 13633 1736 13670 1767
rect 13946 1763 14010 1775
rect 14050 1737 14077 1915
rect 13229 1709 13278 1736
rect 13414 1710 13463 1736
rect 13632 1735 13713 1736
rect 13909 1735 14077 1737
rect 13632 1710 14077 1735
rect 13633 1709 14077 1710
rect 11992 1703 12436 1704
rect 11992 1678 12437 1703
rect 11992 1676 12160 1678
rect 12356 1677 12437 1678
rect 12606 1677 12655 1703
rect 12791 1677 12840 1704
rect 11992 1498 12019 1676
rect 12059 1638 12123 1650
rect 12399 1646 12436 1677
rect 12617 1646 12654 1677
rect 12799 1652 12840 1677
rect 13231 1676 13278 1709
rect 13634 1676 13674 1709
rect 13909 1708 14077 1709
rect 14540 1713 14580 1937
rect 14706 1936 14874 1937
rect 15477 2071 15921 2085
rect 15477 2069 15645 2071
rect 15477 1891 15504 2069
rect 15544 2031 15608 2043
rect 15884 2039 15921 2071
rect 15947 2070 16138 2092
rect 16373 2088 16482 2108
rect 16502 2088 16511 2108
rect 16373 2081 16511 2088
rect 16569 2108 16717 2117
rect 16569 2088 16578 2108
rect 16598 2088 16688 2108
rect 16708 2088 16717 2108
rect 16373 2079 16469 2081
rect 16569 2078 16717 2088
rect 16776 2108 16813 2118
rect 16776 2088 16784 2108
rect 16804 2088 16813 2108
rect 16625 2077 16661 2078
rect 16102 2068 16138 2070
rect 16102 2039 16139 2068
rect 15544 2030 15579 2031
rect 15521 2025 15579 2030
rect 15521 2005 15524 2025
rect 15544 2011 15579 2025
rect 15599 2011 15608 2031
rect 15544 2003 15608 2011
rect 15570 2002 15608 2003
rect 15571 2001 15608 2002
rect 15674 2035 15710 2036
rect 15782 2035 15818 2036
rect 15674 2027 15818 2035
rect 15674 2007 15682 2027
rect 15702 2025 15790 2027
rect 15702 2007 15735 2025
rect 15674 2006 15735 2007
rect 15756 2007 15790 2025
rect 15810 2007 15818 2027
rect 15756 2006 15818 2007
rect 15674 2001 15818 2006
rect 15884 2031 15922 2039
rect 16000 2035 16036 2036
rect 15884 2011 15893 2031
rect 15913 2011 15922 2031
rect 15884 2002 15922 2011
rect 15951 2027 16036 2035
rect 15951 2007 16008 2027
rect 16028 2007 16036 2027
rect 15884 2001 15921 2002
rect 15951 2001 16036 2007
rect 16102 2031 16140 2039
rect 16102 2011 16111 2031
rect 16131 2011 16140 2031
rect 16776 2021 16813 2088
rect 16848 2117 16879 2168
rect 17161 2156 17179 2174
rect 17197 2156 17213 2174
rect 16898 2117 16935 2118
rect 16848 2108 16935 2117
rect 16848 2088 16906 2108
rect 16926 2088 16935 2108
rect 16848 2078 16935 2088
rect 16994 2108 17031 2118
rect 16994 2088 17002 2108
rect 17022 2088 17031 2108
rect 16848 2077 16879 2078
rect 16473 2018 16510 2019
rect 16776 2018 16815 2021
rect 16472 2017 16815 2018
rect 16994 2017 17031 2088
rect 16102 2002 16140 2011
rect 16397 2012 16815 2017
rect 16102 2001 16139 2002
rect 15563 1973 15653 1979
rect 15563 1953 15579 1973
rect 15599 1971 15653 1973
rect 15599 1953 15624 1971
rect 15563 1951 15624 1953
rect 15644 1951 15653 1971
rect 15563 1945 15653 1951
rect 15576 1891 15613 1892
rect 15672 1891 15709 1892
rect 15728 1891 15764 2001
rect 15951 1980 15982 2001
rect 16397 1992 16400 2012
rect 16420 1992 16815 2012
rect 16844 1993 17031 2017
rect 15947 1979 15982 1980
rect 15825 1969 15982 1979
rect 15825 1949 15842 1969
rect 15862 1949 15982 1969
rect 15825 1942 15982 1949
rect 16049 1972 16198 1980
rect 16049 1952 16060 1972
rect 16080 1952 16119 1972
rect 16139 1952 16198 1972
rect 16049 1945 16198 1952
rect 16776 1967 16815 1992
rect 17161 1967 17213 2156
rect 16776 1949 17215 1967
rect 16049 1944 16090 1945
rect 15783 1891 15820 1892
rect 15476 1882 15614 1891
rect 15476 1862 15585 1882
rect 15605 1862 15614 1882
rect 15476 1855 15614 1862
rect 15672 1882 15820 1891
rect 15672 1862 15681 1882
rect 15701 1862 15791 1882
rect 15811 1862 15820 1882
rect 15476 1853 15572 1855
rect 15672 1852 15820 1862
rect 15879 1882 15916 1892
rect 15879 1862 15887 1882
rect 15907 1862 15916 1882
rect 15728 1851 15764 1852
rect 15576 1792 15613 1793
rect 15879 1792 15916 1862
rect 15951 1891 15982 1942
rect 16776 1931 17176 1949
rect 17194 1931 17215 1949
rect 16776 1925 17215 1931
rect 16782 1921 17215 1925
rect 17161 1919 17213 1921
rect 16001 1891 16038 1892
rect 15951 1882 16038 1891
rect 15951 1862 16009 1882
rect 16029 1862 16038 1882
rect 15951 1852 16038 1862
rect 16097 1882 16134 1892
rect 16097 1862 16105 1882
rect 16125 1862 16134 1882
rect 15951 1851 15982 1852
rect 15575 1791 15916 1792
rect 16097 1791 16134 1862
rect 17164 1854 17201 1859
rect 17155 1850 17202 1854
rect 17155 1832 17174 1850
rect 17192 1832 17202 1850
rect 15500 1786 15916 1791
rect 15500 1766 15503 1786
rect 15523 1766 15916 1786
rect 15947 1767 16134 1791
rect 16759 1789 16799 1794
rect 17155 1789 17202 1832
rect 16759 1750 17202 1789
rect 14540 1691 14548 1713
rect 14572 1691 14580 1713
rect 14540 1683 14580 1691
rect 15853 1735 15893 1743
rect 15853 1713 15861 1735
rect 15885 1713 15893 1735
rect 12059 1637 12094 1638
rect 12036 1632 12094 1637
rect 12036 1612 12039 1632
rect 12059 1618 12094 1632
rect 12114 1618 12123 1638
rect 12059 1610 12123 1618
rect 12085 1609 12123 1610
rect 12086 1608 12123 1609
rect 12189 1642 12225 1643
rect 12297 1642 12333 1643
rect 12189 1634 12333 1642
rect 12189 1614 12197 1634
rect 12217 1630 12305 1634
rect 12217 1614 12261 1630
rect 12189 1610 12261 1614
rect 12281 1614 12305 1630
rect 12325 1614 12333 1634
rect 12281 1610 12333 1614
rect 12189 1608 12333 1610
rect 12399 1638 12437 1646
rect 12515 1642 12551 1643
rect 12399 1618 12408 1638
rect 12428 1618 12437 1638
rect 12399 1609 12437 1618
rect 12466 1634 12551 1642
rect 12466 1614 12523 1634
rect 12543 1614 12551 1634
rect 12399 1608 12436 1609
rect 12466 1608 12551 1614
rect 12617 1638 12655 1646
rect 12617 1618 12626 1638
rect 12646 1618 12655 1638
rect 12617 1609 12655 1618
rect 12799 1643 12841 1652
rect 12799 1625 12813 1643
rect 12831 1625 12841 1643
rect 12799 1617 12841 1625
rect 12804 1615 12841 1617
rect 13231 1637 13674 1676
rect 12617 1608 12654 1609
rect 12078 1580 12168 1586
rect 12078 1560 12094 1580
rect 12114 1578 12168 1580
rect 12114 1560 12139 1578
rect 12078 1558 12139 1560
rect 12159 1558 12168 1578
rect 12078 1552 12168 1558
rect 12091 1498 12128 1499
rect 12187 1498 12224 1499
rect 12243 1498 12279 1608
rect 12466 1587 12497 1608
rect 13231 1594 13278 1637
rect 13634 1632 13674 1637
rect 14299 1635 14486 1659
rect 14517 1640 14910 1660
rect 14930 1640 14933 1660
rect 14517 1635 14933 1640
rect 12462 1586 12497 1587
rect 12340 1576 12497 1586
rect 12340 1556 12357 1576
rect 12377 1556 12497 1576
rect 12340 1549 12497 1556
rect 12564 1579 12713 1587
rect 12564 1559 12575 1579
rect 12595 1559 12634 1579
rect 12654 1559 12713 1579
rect 13231 1576 13241 1594
rect 13259 1576 13278 1594
rect 13231 1572 13278 1576
rect 13232 1567 13269 1572
rect 12564 1552 12713 1559
rect 14299 1564 14336 1635
rect 14517 1634 14858 1635
rect 14451 1574 14482 1575
rect 12564 1551 12605 1552
rect 12801 1550 12838 1553
rect 12298 1498 12335 1499
rect 11991 1489 12129 1498
rect 11195 1450 11639 1476
rect 11195 1448 11363 1450
rect 10148 1316 10595 1328
rect 10191 1314 10224 1316
rect 9558 1296 9696 1305
rect 9352 1295 9389 1296
rect 9082 1242 9123 1243
rect 8856 1221 8908 1239
rect 8974 1235 9123 1242
rect 8411 1202 8451 1212
rect 8974 1215 9033 1235
rect 9053 1215 9092 1235
rect 9112 1215 9123 1235
rect 8974 1207 9123 1215
rect 9190 1238 9347 1245
rect 9190 1218 9310 1238
rect 9330 1218 9347 1238
rect 9190 1208 9347 1218
rect 9190 1207 9225 1208
rect 8241 1185 8279 1194
rect 9190 1186 9221 1207
rect 9408 1186 9444 1296
rect 9463 1295 9500 1296
rect 9559 1295 9596 1296
rect 9519 1236 9609 1242
rect 9519 1216 9528 1236
rect 9548 1234 9609 1236
rect 9548 1216 9573 1234
rect 9519 1214 9573 1216
rect 9593 1214 9609 1234
rect 9519 1208 9609 1214
rect 9033 1185 9070 1186
rect 8241 1184 8278 1185
rect 7702 1156 7792 1162
rect 7702 1136 7718 1156
rect 7738 1154 7792 1156
rect 7738 1136 7763 1154
rect 7702 1134 7763 1136
rect 7783 1134 7792 1154
rect 7702 1128 7792 1134
rect 7715 1074 7752 1075
rect 7811 1074 7848 1075
rect 7867 1074 7903 1184
rect 8090 1163 8121 1184
rect 9032 1176 9070 1185
rect 8086 1162 8121 1163
rect 7964 1152 8121 1162
rect 7964 1132 7981 1152
rect 8001 1132 8121 1152
rect 7964 1125 8121 1132
rect 8188 1155 8337 1163
rect 8188 1135 8199 1155
rect 8219 1135 8258 1155
rect 8278 1135 8337 1155
rect 8860 1158 8900 1168
rect 8188 1128 8337 1135
rect 8403 1131 8455 1149
rect 8188 1127 8229 1128
rect 7922 1074 7959 1075
rect 7615 1065 7753 1074
rect 7615 1045 7724 1065
rect 7744 1045 7753 1065
rect 7615 1038 7753 1045
rect 7811 1065 7959 1074
rect 7811 1045 7820 1065
rect 7840 1045 7930 1065
rect 7950 1045 7959 1065
rect 7615 1036 7711 1038
rect 7811 1035 7959 1045
rect 8018 1065 8055 1075
rect 8018 1045 8026 1065
rect 8046 1045 8055 1065
rect 7867 1034 7903 1035
rect 8018 978 8055 1045
rect 8090 1074 8121 1125
rect 8403 1113 8421 1131
rect 8439 1113 8455 1131
rect 8140 1074 8177 1075
rect 8090 1065 8177 1074
rect 8090 1045 8148 1065
rect 8168 1045 8177 1065
rect 8090 1035 8177 1045
rect 8236 1065 8273 1075
rect 8236 1045 8244 1065
rect 8264 1045 8273 1065
rect 8090 1034 8121 1035
rect 7715 975 7752 976
rect 8018 975 8057 978
rect 7714 974 8057 975
rect 8236 974 8273 1045
rect 7639 969 8057 974
rect 7639 949 7642 969
rect 7662 949 8057 969
rect 8086 950 8273 974
rect 6180 918 6217 926
rect 6180 899 6188 918
rect 6209 899 6217 918
rect 6180 893 6217 899
rect 8018 924 8057 949
rect 8403 924 8455 1113
rect 8860 1140 8870 1158
rect 8888 1140 8900 1158
rect 9032 1156 9041 1176
rect 9061 1156 9070 1176
rect 9032 1148 9070 1156
rect 9136 1180 9221 1186
rect 9251 1185 9288 1186
rect 9136 1160 9144 1180
rect 9164 1160 9221 1180
rect 9136 1152 9221 1160
rect 9250 1176 9288 1185
rect 9250 1156 9259 1176
rect 9279 1156 9288 1176
rect 9136 1151 9172 1152
rect 9250 1148 9288 1156
rect 9354 1180 9498 1186
rect 9354 1160 9362 1180
rect 9382 1160 9415 1180
rect 9435 1160 9470 1180
rect 9490 1160 9498 1180
rect 9354 1152 9498 1160
rect 9354 1151 9390 1152
rect 9462 1151 9498 1152
rect 9564 1185 9601 1186
rect 9564 1184 9602 1185
rect 9564 1176 9628 1184
rect 9564 1156 9573 1176
rect 9593 1162 9628 1176
rect 9648 1162 9651 1182
rect 9593 1157 9651 1162
rect 9593 1156 9628 1157
rect 8860 1084 8900 1140
rect 9033 1119 9070 1148
rect 9034 1117 9070 1119
rect 9034 1095 9225 1117
rect 9251 1116 9288 1148
rect 9564 1144 9628 1156
rect 9668 1118 9695 1296
rect 10553 1271 10595 1316
rect 9527 1116 9695 1118
rect 9251 1106 9695 1116
rect 9836 1212 10023 1236
rect 10054 1217 10447 1237
rect 10467 1217 10470 1237
rect 10054 1212 10470 1217
rect 9836 1141 9873 1212
rect 10054 1211 10395 1212
rect 9988 1151 10019 1152
rect 9836 1121 9845 1141
rect 9865 1121 9873 1141
rect 9836 1111 9873 1121
rect 9932 1141 10019 1151
rect 9932 1121 9941 1141
rect 9961 1121 10019 1141
rect 9932 1112 10019 1121
rect 9932 1111 9969 1112
rect 8857 1079 8900 1084
rect 9248 1090 9695 1106
rect 9248 1084 9276 1090
rect 9527 1089 9695 1090
rect 8857 1076 9007 1079
rect 9248 1076 9275 1084
rect 8857 1074 9275 1076
rect 8857 1056 8866 1074
rect 8884 1056 9275 1074
rect 9988 1061 10019 1112
rect 10054 1141 10091 1211
rect 10357 1210 10394 1211
rect 10206 1151 10242 1152
rect 10054 1121 10063 1141
rect 10083 1121 10091 1141
rect 10054 1111 10091 1121
rect 10150 1141 10298 1151
rect 10398 1148 10494 1150
rect 10150 1121 10159 1141
rect 10179 1121 10269 1141
rect 10289 1121 10298 1141
rect 10150 1112 10298 1121
rect 10356 1141 10494 1148
rect 10356 1121 10365 1141
rect 10385 1121 10494 1141
rect 10356 1112 10494 1121
rect 10150 1111 10187 1112
rect 9880 1058 9921 1059
rect 8857 1053 9275 1056
rect 8857 1047 8900 1053
rect 8860 1044 8900 1047
rect 9775 1051 9921 1058
rect 9257 1035 9297 1036
rect 8968 1018 9297 1035
rect 9775 1031 9831 1051
rect 9851 1031 9890 1051
rect 9910 1031 9921 1051
rect 9775 1023 9921 1031
rect 9988 1054 10145 1061
rect 9988 1034 10108 1054
rect 10128 1034 10145 1054
rect 9988 1024 10145 1034
rect 9988 1023 10023 1024
rect 8852 975 8895 986
rect 8852 957 8864 975
rect 8882 957 8895 975
rect 8852 931 8895 957
rect 8968 931 8995 1018
rect 9257 1009 9297 1018
rect 8018 906 8457 924
rect 8018 888 8418 906
rect 8436 888 8457 906
rect 8018 882 8457 888
rect 8024 878 8457 882
rect 8852 910 8995 931
rect 9039 983 9073 999
rect 9257 989 9650 1009
rect 9670 989 9673 1009
rect 9988 1002 10019 1023
rect 10206 1002 10242 1112
rect 10261 1111 10298 1112
rect 10357 1111 10394 1112
rect 10317 1052 10407 1058
rect 10317 1032 10326 1052
rect 10346 1050 10407 1052
rect 10346 1032 10371 1050
rect 10317 1030 10371 1032
rect 10391 1030 10407 1050
rect 10317 1024 10407 1030
rect 9831 1001 9868 1002
rect 9257 984 9673 989
rect 9830 992 9868 1001
rect 9257 983 9598 984
rect 9039 913 9076 983
rect 9191 923 9222 924
rect 8852 908 8989 910
rect 8403 876 8455 878
rect 8852 866 8895 908
rect 9039 893 9048 913
rect 9068 893 9076 913
rect 9039 883 9076 893
rect 9135 913 9222 923
rect 9135 893 9144 913
rect 9164 893 9222 913
rect 9135 884 9222 893
rect 9135 883 9172 884
rect 8850 856 8895 866
rect 8850 838 8859 856
rect 8877 838 8895 856
rect 8850 832 8895 838
rect 9191 833 9222 884
rect 9257 913 9294 983
rect 9560 982 9597 983
rect 9830 972 9839 992
rect 9859 972 9868 992
rect 9830 964 9868 972
rect 9934 996 10019 1002
rect 10049 1001 10086 1002
rect 9934 976 9942 996
rect 9962 976 10019 996
rect 9934 968 10019 976
rect 10048 992 10086 1001
rect 10048 972 10057 992
rect 10077 972 10086 992
rect 9934 967 9970 968
rect 10048 964 10086 972
rect 10152 996 10296 1002
rect 10152 976 10160 996
rect 10180 993 10268 996
rect 10180 976 10215 993
rect 10152 975 10215 976
rect 10234 976 10268 993
rect 10288 976 10296 996
rect 10234 975 10296 976
rect 10152 968 10296 975
rect 10152 967 10188 968
rect 10260 967 10296 968
rect 10362 1001 10399 1002
rect 10362 1000 10400 1001
rect 10422 1000 10449 1004
rect 10362 998 10449 1000
rect 10362 992 10426 998
rect 10362 972 10371 992
rect 10391 978 10426 992
rect 10446 978 10449 998
rect 10391 973 10449 978
rect 10391 972 10426 973
rect 9831 935 9868 964
rect 9832 933 9868 935
rect 9409 923 9445 924
rect 9257 893 9266 913
rect 9286 893 9294 913
rect 9257 883 9294 893
rect 9353 913 9501 923
rect 9601 920 9697 922
rect 9353 893 9362 913
rect 9382 893 9472 913
rect 9492 893 9501 913
rect 9353 884 9501 893
rect 9559 913 9697 920
rect 9559 893 9568 913
rect 9588 893 9697 913
rect 9832 911 10023 933
rect 10049 932 10086 964
rect 10362 960 10426 972
rect 10466 934 10493 1112
rect 10325 932 10493 934
rect 10049 906 10493 932
rect 9559 884 9697 893
rect 9353 883 9390 884
rect 8850 829 8887 832
rect 9083 830 9124 831
rect 8975 823 9124 830
rect 8406 811 8443 816
rect 8397 807 8444 811
rect 8397 789 8416 807
rect 8434 789 8444 807
rect 8975 803 9034 823
rect 9054 803 9093 823
rect 9113 803 9124 823
rect 8975 795 9124 803
rect 9191 826 9348 833
rect 9191 806 9311 826
rect 9331 806 9348 826
rect 9191 796 9348 806
rect 9191 795 9226 796
rect 8397 726 8444 789
rect 9191 774 9222 795
rect 9409 774 9445 884
rect 9464 883 9501 884
rect 9560 883 9597 884
rect 9520 824 9610 830
rect 9520 804 9529 824
rect 9549 822 9610 824
rect 9549 804 9574 822
rect 9520 802 9574 804
rect 9594 802 9610 822
rect 9520 796 9610 802
rect 9034 773 9071 774
rect 8847 765 8884 767
rect 8847 757 8889 765
rect 8847 739 8857 757
rect 8875 739 8889 757
rect 8847 730 8889 739
rect 9033 764 9071 773
rect 9033 744 9042 764
rect 9062 744 9071 764
rect 9033 736 9071 744
rect 9137 768 9222 774
rect 9252 773 9289 774
rect 9137 748 9145 768
rect 9165 748 9222 768
rect 9137 740 9222 748
rect 9251 764 9289 773
rect 9251 744 9260 764
rect 9280 744 9289 764
rect 9137 739 9173 740
rect 9251 736 9289 744
rect 9355 772 9499 774
rect 9355 768 9407 772
rect 9355 748 9363 768
rect 9383 752 9407 768
rect 9427 768 9499 772
rect 9427 752 9471 768
rect 9383 748 9471 752
rect 9491 748 9499 768
rect 9355 740 9499 748
rect 9355 739 9391 740
rect 9463 739 9499 740
rect 9565 773 9602 774
rect 9565 772 9603 773
rect 9565 764 9629 772
rect 9565 744 9574 764
rect 9594 750 9629 764
rect 9649 750 9652 770
rect 9594 745 9652 750
rect 9594 744 9629 745
rect 8397 711 8447 726
rect 8397 686 8411 711
rect 8443 686 8447 711
rect 8848 705 8889 730
rect 9034 705 9071 736
rect 9252 714 9289 736
rect 9565 732 9629 744
rect 9247 705 9289 714
rect 9669 706 9696 884
rect 8848 693 8893 705
rect 8397 673 8444 686
rect 5782 648 5790 670
rect 5814 648 5822 670
rect 5782 640 5822 648
rect 8844 635 8893 693
rect 9034 679 9096 705
rect 9247 704 9332 705
rect 9528 704 9696 706
rect 9247 678 9696 704
rect 9247 635 9286 678
rect 9528 677 9696 678
rect 10159 682 10199 906
rect 10325 905 10493 906
rect 10557 938 10590 1271
rect 11195 1270 11222 1448
rect 11262 1410 11326 1422
rect 11602 1418 11639 1450
rect 11665 1449 11856 1471
rect 11991 1469 12100 1489
rect 12120 1469 12129 1489
rect 11991 1462 12129 1469
rect 12187 1489 12335 1498
rect 12187 1469 12196 1489
rect 12216 1469 12306 1489
rect 12326 1469 12335 1489
rect 11991 1460 12087 1462
rect 12187 1459 12335 1469
rect 12394 1489 12431 1499
rect 12394 1469 12402 1489
rect 12422 1469 12431 1489
rect 12243 1458 12279 1459
rect 11820 1447 11856 1449
rect 11820 1418 11857 1447
rect 11262 1409 11297 1410
rect 11239 1404 11297 1409
rect 11239 1384 11242 1404
rect 11262 1390 11297 1404
rect 11317 1390 11326 1410
rect 11262 1382 11326 1390
rect 11288 1381 11326 1382
rect 11289 1380 11326 1381
rect 11392 1414 11428 1415
rect 11500 1414 11536 1415
rect 11392 1406 11536 1414
rect 11392 1386 11400 1406
rect 11420 1405 11508 1406
rect 11420 1386 11455 1405
rect 11476 1386 11508 1405
rect 11528 1386 11536 1406
rect 11392 1380 11536 1386
rect 11602 1410 11640 1418
rect 11718 1414 11754 1415
rect 11602 1390 11611 1410
rect 11631 1390 11640 1410
rect 11602 1381 11640 1390
rect 11669 1406 11754 1414
rect 11669 1386 11726 1406
rect 11746 1386 11754 1406
rect 11602 1380 11639 1381
rect 11669 1380 11754 1386
rect 11820 1410 11858 1418
rect 11820 1390 11829 1410
rect 11849 1390 11858 1410
rect 12091 1399 12128 1400
rect 12394 1399 12431 1469
rect 12466 1498 12497 1549
rect 12793 1544 12838 1550
rect 12793 1526 12811 1544
rect 12829 1526 12838 1544
rect 14299 1544 14308 1564
rect 14328 1544 14336 1564
rect 14299 1534 14336 1544
rect 14395 1564 14482 1574
rect 14395 1544 14404 1564
rect 14424 1544 14482 1564
rect 14395 1535 14482 1544
rect 14395 1534 14432 1535
rect 12793 1516 12838 1526
rect 12516 1498 12553 1499
rect 12466 1489 12553 1498
rect 12466 1469 12524 1489
rect 12544 1469 12553 1489
rect 12466 1459 12553 1469
rect 12612 1489 12649 1499
rect 12612 1469 12620 1489
rect 12640 1469 12649 1489
rect 12793 1474 12836 1516
rect 13220 1505 13272 1507
rect 12699 1472 12836 1474
rect 12466 1458 12497 1459
rect 12612 1399 12649 1469
rect 12090 1398 12431 1399
rect 11820 1381 11858 1390
rect 12015 1393 12431 1398
rect 11820 1380 11857 1381
rect 11281 1352 11371 1358
rect 11281 1332 11297 1352
rect 11317 1350 11371 1352
rect 11317 1332 11342 1350
rect 11281 1330 11342 1332
rect 11362 1330 11371 1350
rect 11281 1324 11371 1330
rect 11294 1270 11331 1271
rect 11390 1270 11427 1271
rect 11446 1270 11482 1380
rect 11669 1359 11700 1380
rect 12015 1373 12018 1393
rect 12038 1373 12431 1393
rect 12615 1383 12649 1399
rect 12693 1451 12836 1472
rect 13218 1501 13651 1505
rect 13218 1495 13657 1501
rect 13218 1477 13239 1495
rect 13257 1477 13657 1495
rect 14451 1484 14482 1535
rect 14517 1564 14554 1634
rect 14820 1633 14857 1634
rect 14669 1574 14705 1575
rect 14517 1544 14526 1564
rect 14546 1544 14554 1564
rect 14517 1534 14554 1544
rect 14613 1564 14761 1574
rect 14861 1571 14957 1573
rect 14613 1544 14622 1564
rect 14642 1544 14732 1564
rect 14752 1544 14761 1564
rect 14613 1535 14761 1544
rect 14819 1564 14957 1571
rect 14819 1544 14828 1564
rect 14848 1544 14957 1564
rect 14819 1535 14957 1544
rect 14613 1534 14650 1535
rect 14343 1481 14384 1482
rect 13218 1459 13657 1477
rect 12391 1364 12431 1373
rect 12693 1364 12720 1451
rect 12793 1425 12836 1451
rect 12793 1407 12806 1425
rect 12824 1407 12836 1425
rect 12793 1396 12836 1407
rect 11665 1358 11700 1359
rect 11543 1348 11700 1358
rect 11543 1328 11560 1348
rect 11580 1328 11700 1348
rect 11543 1321 11700 1328
rect 11767 1351 11916 1359
rect 11767 1331 11778 1351
rect 11798 1331 11837 1351
rect 11857 1331 11916 1351
rect 12391 1347 12720 1364
rect 12391 1346 12431 1347
rect 11767 1324 11916 1331
rect 12788 1335 12828 1338
rect 12788 1329 12831 1335
rect 12413 1326 12831 1329
rect 11767 1323 11808 1324
rect 11501 1270 11538 1271
rect 11194 1261 11332 1270
rect 11194 1241 11303 1261
rect 11323 1241 11332 1261
rect 11194 1234 11332 1241
rect 11390 1261 11538 1270
rect 11390 1241 11399 1261
rect 11419 1241 11509 1261
rect 11529 1241 11538 1261
rect 11194 1232 11290 1234
rect 11390 1231 11538 1241
rect 11597 1261 11634 1271
rect 11597 1241 11605 1261
rect 11625 1241 11634 1261
rect 11446 1230 11482 1231
rect 11294 1171 11331 1172
rect 11597 1171 11634 1241
rect 11669 1270 11700 1321
rect 12413 1308 12804 1326
rect 12822 1308 12831 1326
rect 12413 1306 12831 1308
rect 12413 1298 12440 1306
rect 12681 1303 12831 1306
rect 11993 1292 12161 1293
rect 12412 1292 12440 1298
rect 11993 1276 12440 1292
rect 12788 1298 12831 1303
rect 11719 1270 11756 1271
rect 11669 1261 11756 1270
rect 11669 1241 11727 1261
rect 11747 1241 11756 1261
rect 11669 1231 11756 1241
rect 11815 1261 11852 1271
rect 11815 1241 11823 1261
rect 11843 1241 11852 1261
rect 11669 1230 11700 1231
rect 11293 1170 11634 1171
rect 11815 1170 11852 1241
rect 11218 1165 11634 1170
rect 11218 1145 11221 1165
rect 11241 1145 11634 1165
rect 11665 1146 11852 1170
rect 11993 1266 12437 1276
rect 11993 1264 12161 1266
rect 11993 1086 12020 1264
rect 12060 1226 12124 1238
rect 12400 1234 12437 1266
rect 12463 1265 12654 1287
rect 12618 1263 12654 1265
rect 12618 1234 12655 1263
rect 12788 1242 12828 1298
rect 12060 1225 12095 1226
rect 12037 1220 12095 1225
rect 12037 1200 12040 1220
rect 12060 1206 12095 1220
rect 12115 1206 12124 1226
rect 12060 1198 12124 1206
rect 12086 1197 12124 1198
rect 12087 1196 12124 1197
rect 12190 1230 12226 1231
rect 12298 1230 12334 1231
rect 12190 1222 12334 1230
rect 12190 1202 12198 1222
rect 12218 1202 12253 1222
rect 12273 1202 12306 1222
rect 12326 1202 12334 1222
rect 12190 1196 12334 1202
rect 12400 1226 12438 1234
rect 12516 1230 12552 1231
rect 12400 1206 12409 1226
rect 12429 1206 12438 1226
rect 12400 1197 12438 1206
rect 12467 1222 12552 1230
rect 12467 1202 12524 1222
rect 12544 1202 12552 1222
rect 12400 1196 12437 1197
rect 12467 1196 12552 1202
rect 12618 1226 12656 1234
rect 12618 1206 12627 1226
rect 12647 1206 12656 1226
rect 12788 1224 12800 1242
rect 12818 1224 12828 1242
rect 13220 1270 13272 1459
rect 13618 1434 13657 1459
rect 14235 1474 14384 1481
rect 14235 1454 14294 1474
rect 14314 1454 14353 1474
rect 14373 1454 14384 1474
rect 14235 1446 14384 1454
rect 14451 1477 14608 1484
rect 14451 1457 14571 1477
rect 14591 1457 14608 1477
rect 14451 1447 14608 1457
rect 14451 1446 14486 1447
rect 13402 1409 13589 1433
rect 13618 1414 14013 1434
rect 14033 1414 14036 1434
rect 14451 1425 14482 1446
rect 14669 1425 14705 1535
rect 14724 1534 14761 1535
rect 14820 1534 14857 1535
rect 14780 1475 14870 1481
rect 14780 1455 14789 1475
rect 14809 1473 14870 1475
rect 14809 1455 14834 1473
rect 14780 1453 14834 1455
rect 14854 1453 14870 1473
rect 14780 1447 14870 1453
rect 14294 1424 14331 1425
rect 13618 1409 14036 1414
rect 14293 1415 14331 1424
rect 13402 1338 13439 1409
rect 13618 1408 13961 1409
rect 13618 1405 13657 1408
rect 13923 1407 13960 1408
rect 13554 1348 13585 1349
rect 13402 1318 13411 1338
rect 13431 1318 13439 1338
rect 13402 1308 13439 1318
rect 13498 1338 13585 1348
rect 13498 1318 13507 1338
rect 13527 1318 13585 1338
rect 13498 1309 13585 1318
rect 13498 1308 13535 1309
rect 13220 1252 13236 1270
rect 13254 1252 13272 1270
rect 13554 1258 13585 1309
rect 13620 1338 13657 1405
rect 14293 1395 14302 1415
rect 14322 1395 14331 1415
rect 14293 1387 14331 1395
rect 14397 1419 14482 1425
rect 14512 1424 14549 1425
rect 14397 1399 14405 1419
rect 14425 1399 14482 1419
rect 14397 1391 14482 1399
rect 14511 1415 14549 1424
rect 14511 1395 14520 1415
rect 14540 1395 14549 1415
rect 14397 1390 14433 1391
rect 14511 1387 14549 1395
rect 14615 1419 14759 1425
rect 14615 1399 14623 1419
rect 14643 1414 14731 1419
rect 14643 1399 14679 1414
rect 14615 1397 14679 1399
rect 14698 1399 14731 1414
rect 14751 1399 14759 1419
rect 14698 1397 14759 1399
rect 14615 1391 14759 1397
rect 14615 1390 14651 1391
rect 14723 1390 14759 1391
rect 14825 1424 14862 1425
rect 14825 1423 14863 1424
rect 14825 1415 14889 1423
rect 14825 1395 14834 1415
rect 14854 1401 14889 1415
rect 14909 1401 14912 1421
rect 14854 1396 14912 1401
rect 14854 1395 14889 1396
rect 14294 1358 14331 1387
rect 14295 1356 14331 1358
rect 13772 1348 13808 1349
rect 13620 1318 13629 1338
rect 13649 1318 13657 1338
rect 13620 1308 13657 1318
rect 13716 1338 13864 1348
rect 13964 1345 14060 1347
rect 13716 1318 13725 1338
rect 13745 1318 13835 1338
rect 13855 1318 13864 1338
rect 13716 1309 13864 1318
rect 13922 1338 14060 1345
rect 13922 1318 13931 1338
rect 13951 1318 14060 1338
rect 14295 1334 14486 1356
rect 14512 1355 14549 1387
rect 14825 1383 14889 1395
rect 14929 1357 14956 1535
rect 14788 1355 14956 1357
rect 14512 1341 14956 1355
rect 15559 1489 15727 1490
rect 15853 1489 15893 1713
rect 16356 1717 16524 1718
rect 16759 1717 16799 1750
rect 17155 1717 17202 1750
rect 16356 1716 16800 1717
rect 16356 1691 16801 1716
rect 16356 1689 16524 1691
rect 16720 1690 16801 1691
rect 16970 1690 17019 1716
rect 17155 1690 17204 1717
rect 16356 1511 16383 1689
rect 16423 1651 16487 1663
rect 16763 1659 16800 1690
rect 16981 1659 17018 1690
rect 17163 1665 17204 1690
rect 16423 1650 16458 1651
rect 16400 1645 16458 1650
rect 16400 1625 16403 1645
rect 16423 1631 16458 1645
rect 16478 1631 16487 1651
rect 16423 1623 16487 1631
rect 16449 1622 16487 1623
rect 16450 1621 16487 1622
rect 16553 1655 16589 1656
rect 16661 1655 16697 1656
rect 16553 1647 16697 1655
rect 16553 1627 16561 1647
rect 16581 1643 16669 1647
rect 16581 1627 16625 1643
rect 16553 1623 16625 1627
rect 16645 1627 16669 1643
rect 16689 1627 16697 1647
rect 16645 1623 16697 1627
rect 16553 1621 16697 1623
rect 16763 1651 16801 1659
rect 16879 1655 16915 1656
rect 16763 1631 16772 1651
rect 16792 1631 16801 1651
rect 16763 1622 16801 1631
rect 16830 1647 16915 1655
rect 16830 1627 16887 1647
rect 16907 1627 16915 1647
rect 16763 1621 16800 1622
rect 16830 1621 16915 1627
rect 16981 1651 17019 1659
rect 16981 1631 16990 1651
rect 17010 1631 17019 1651
rect 16981 1622 17019 1631
rect 17163 1656 17205 1665
rect 17163 1638 17177 1656
rect 17195 1638 17205 1656
rect 17163 1630 17205 1638
rect 17168 1628 17205 1630
rect 16981 1621 17018 1622
rect 16442 1593 16532 1599
rect 16442 1573 16458 1593
rect 16478 1591 16532 1593
rect 16478 1573 16503 1591
rect 16442 1571 16503 1573
rect 16523 1571 16532 1591
rect 16442 1565 16532 1571
rect 16455 1511 16492 1512
rect 16551 1511 16588 1512
rect 16607 1511 16643 1621
rect 16830 1600 16861 1621
rect 16826 1599 16861 1600
rect 16704 1589 16861 1599
rect 16704 1569 16721 1589
rect 16741 1569 16861 1589
rect 16704 1562 16861 1569
rect 16928 1592 17077 1600
rect 16928 1572 16939 1592
rect 16959 1572 16998 1592
rect 17018 1572 17077 1592
rect 16928 1565 17077 1572
rect 16928 1564 16969 1565
rect 17165 1563 17202 1566
rect 16662 1511 16699 1512
rect 16355 1502 16493 1511
rect 15559 1463 16003 1489
rect 15559 1461 15727 1463
rect 14512 1329 14959 1341
rect 14555 1327 14588 1329
rect 13922 1309 14060 1318
rect 13716 1308 13753 1309
rect 13446 1255 13487 1256
rect 13220 1234 13272 1252
rect 13338 1248 13487 1255
rect 12788 1214 12828 1224
rect 13338 1228 13397 1248
rect 13417 1228 13456 1248
rect 13476 1228 13487 1248
rect 13338 1220 13487 1228
rect 13554 1251 13711 1258
rect 13554 1231 13674 1251
rect 13694 1231 13711 1251
rect 13554 1221 13711 1231
rect 13554 1220 13589 1221
rect 12618 1197 12656 1206
rect 13554 1199 13585 1220
rect 13772 1199 13808 1309
rect 13827 1308 13864 1309
rect 13923 1308 13960 1309
rect 13883 1249 13973 1255
rect 13883 1229 13892 1249
rect 13912 1247 13973 1249
rect 13912 1229 13937 1247
rect 13883 1227 13937 1229
rect 13957 1227 13973 1247
rect 13883 1221 13973 1227
rect 13397 1198 13434 1199
rect 12618 1196 12655 1197
rect 12079 1168 12169 1174
rect 12079 1148 12095 1168
rect 12115 1166 12169 1168
rect 12115 1148 12140 1166
rect 12079 1146 12140 1148
rect 12160 1146 12169 1166
rect 12079 1140 12169 1146
rect 12092 1086 12129 1087
rect 12188 1086 12225 1087
rect 12244 1086 12280 1196
rect 12467 1175 12498 1196
rect 13396 1189 13434 1198
rect 12463 1174 12498 1175
rect 12341 1164 12498 1174
rect 12341 1144 12358 1164
rect 12378 1144 12498 1164
rect 12341 1137 12498 1144
rect 12565 1167 12714 1175
rect 12565 1147 12576 1167
rect 12596 1147 12635 1167
rect 12655 1147 12714 1167
rect 13224 1171 13264 1181
rect 12565 1140 12714 1147
rect 12780 1143 12832 1161
rect 12565 1139 12606 1140
rect 12299 1086 12336 1087
rect 11992 1077 12130 1086
rect 11992 1057 12101 1077
rect 12121 1057 12130 1077
rect 11992 1050 12130 1057
rect 12188 1077 12336 1086
rect 12188 1057 12197 1077
rect 12217 1057 12307 1077
rect 12327 1057 12336 1077
rect 11992 1048 12088 1050
rect 12188 1047 12336 1057
rect 12395 1077 12432 1087
rect 12395 1057 12403 1077
rect 12423 1057 12432 1077
rect 12244 1046 12280 1047
rect 12395 990 12432 1057
rect 12467 1086 12498 1137
rect 12780 1125 12798 1143
rect 12816 1125 12832 1143
rect 12517 1086 12554 1087
rect 12467 1077 12554 1086
rect 12467 1057 12525 1077
rect 12545 1057 12554 1077
rect 12467 1047 12554 1057
rect 12613 1077 12650 1087
rect 12613 1057 12621 1077
rect 12641 1057 12650 1077
rect 12467 1046 12498 1047
rect 12092 987 12129 988
rect 12395 987 12434 990
rect 12091 986 12434 987
rect 12613 986 12650 1057
rect 12016 981 12434 986
rect 12016 961 12019 981
rect 12039 961 12434 981
rect 12463 962 12650 986
rect 10557 930 10594 938
rect 10557 911 10565 930
rect 10586 911 10594 930
rect 10557 905 10594 911
rect 12395 936 12434 961
rect 12780 936 12832 1125
rect 13224 1153 13234 1171
rect 13252 1153 13264 1171
rect 13396 1169 13405 1189
rect 13425 1169 13434 1189
rect 13396 1161 13434 1169
rect 13500 1193 13585 1199
rect 13615 1198 13652 1199
rect 13500 1173 13508 1193
rect 13528 1173 13585 1193
rect 13500 1165 13585 1173
rect 13614 1189 13652 1198
rect 13614 1169 13623 1189
rect 13643 1169 13652 1189
rect 13500 1164 13536 1165
rect 13614 1161 13652 1169
rect 13718 1193 13862 1199
rect 13718 1173 13726 1193
rect 13746 1173 13779 1193
rect 13799 1173 13834 1193
rect 13854 1173 13862 1193
rect 13718 1165 13862 1173
rect 13718 1164 13754 1165
rect 13826 1164 13862 1165
rect 13928 1198 13965 1199
rect 13928 1197 13966 1198
rect 13928 1189 13992 1197
rect 13928 1169 13937 1189
rect 13957 1175 13992 1189
rect 14012 1175 14015 1195
rect 13957 1170 14015 1175
rect 13957 1169 13992 1170
rect 13224 1097 13264 1153
rect 13397 1132 13434 1161
rect 13398 1130 13434 1132
rect 13398 1108 13589 1130
rect 13615 1129 13652 1161
rect 13928 1157 13992 1169
rect 14032 1131 14059 1309
rect 14917 1284 14959 1329
rect 13891 1129 14059 1131
rect 13615 1119 14059 1129
rect 14200 1225 14387 1249
rect 14418 1230 14811 1250
rect 14831 1230 14834 1250
rect 14418 1225 14834 1230
rect 14200 1154 14237 1225
rect 14418 1224 14759 1225
rect 14352 1164 14383 1165
rect 14200 1134 14209 1154
rect 14229 1134 14237 1154
rect 14200 1124 14237 1134
rect 14296 1154 14383 1164
rect 14296 1134 14305 1154
rect 14325 1134 14383 1154
rect 14296 1125 14383 1134
rect 14296 1124 14333 1125
rect 13221 1092 13264 1097
rect 13612 1103 14059 1119
rect 13612 1097 13640 1103
rect 13891 1102 14059 1103
rect 13221 1089 13371 1092
rect 13612 1089 13639 1097
rect 13221 1087 13639 1089
rect 13221 1069 13230 1087
rect 13248 1069 13639 1087
rect 14352 1074 14383 1125
rect 14418 1154 14455 1224
rect 14721 1223 14758 1224
rect 14570 1164 14606 1165
rect 14418 1134 14427 1154
rect 14447 1134 14455 1154
rect 14418 1124 14455 1134
rect 14514 1154 14662 1164
rect 14762 1161 14858 1163
rect 14514 1134 14523 1154
rect 14543 1134 14633 1154
rect 14653 1134 14662 1154
rect 14514 1125 14662 1134
rect 14720 1154 14858 1161
rect 14720 1134 14729 1154
rect 14749 1134 14858 1154
rect 14720 1125 14858 1134
rect 14514 1124 14551 1125
rect 14244 1071 14285 1072
rect 13221 1066 13639 1069
rect 13221 1060 13264 1066
rect 13224 1057 13264 1060
rect 14139 1064 14285 1071
rect 13621 1048 13661 1049
rect 13332 1031 13661 1048
rect 14139 1044 14195 1064
rect 14215 1044 14254 1064
rect 14274 1044 14285 1064
rect 14139 1036 14285 1044
rect 14352 1067 14509 1074
rect 14352 1047 14472 1067
rect 14492 1047 14509 1067
rect 14352 1037 14509 1047
rect 14352 1036 14387 1037
rect 13216 988 13259 999
rect 13216 970 13228 988
rect 13246 970 13259 988
rect 13216 944 13259 970
rect 13332 944 13359 1031
rect 13621 1022 13661 1031
rect 12395 918 12834 936
rect 12395 900 12795 918
rect 12813 900 12834 918
rect 12395 894 12834 900
rect 12401 890 12834 894
rect 13216 923 13359 944
rect 13403 996 13437 1012
rect 13621 1002 14014 1022
rect 14034 1002 14037 1022
rect 14352 1015 14383 1036
rect 14570 1015 14606 1125
rect 14625 1124 14662 1125
rect 14721 1124 14758 1125
rect 14681 1065 14771 1071
rect 14681 1045 14690 1065
rect 14710 1063 14771 1065
rect 14710 1045 14735 1063
rect 14681 1043 14735 1045
rect 14755 1043 14771 1063
rect 14681 1037 14771 1043
rect 14195 1014 14232 1015
rect 13621 997 14037 1002
rect 14194 1005 14232 1014
rect 13621 996 13962 997
rect 13403 926 13440 996
rect 13555 936 13586 937
rect 13216 921 13353 923
rect 12780 888 12832 890
rect 13216 879 13259 921
rect 13403 906 13412 926
rect 13432 906 13440 926
rect 13403 896 13440 906
rect 13499 926 13586 936
rect 13499 906 13508 926
rect 13528 906 13586 926
rect 13499 897 13586 906
rect 13499 896 13536 897
rect 13214 869 13259 879
rect 13214 851 13223 869
rect 13241 851 13259 869
rect 13214 845 13259 851
rect 13555 846 13586 897
rect 13621 926 13658 996
rect 13924 995 13961 996
rect 14194 985 14203 1005
rect 14223 985 14232 1005
rect 14194 977 14232 985
rect 14298 1009 14383 1015
rect 14413 1014 14450 1015
rect 14298 989 14306 1009
rect 14326 989 14383 1009
rect 14298 981 14383 989
rect 14412 1005 14450 1014
rect 14412 985 14421 1005
rect 14441 985 14450 1005
rect 14298 980 14334 981
rect 14412 977 14450 985
rect 14516 1009 14660 1015
rect 14516 989 14524 1009
rect 14544 1006 14632 1009
rect 14544 989 14579 1006
rect 14516 988 14579 989
rect 14598 989 14632 1006
rect 14652 989 14660 1009
rect 14598 988 14660 989
rect 14516 981 14660 988
rect 14516 980 14552 981
rect 14624 980 14660 981
rect 14726 1014 14763 1015
rect 14726 1013 14764 1014
rect 14786 1013 14813 1017
rect 14726 1011 14813 1013
rect 14726 1005 14790 1011
rect 14726 985 14735 1005
rect 14755 991 14790 1005
rect 14810 991 14813 1011
rect 14755 986 14813 991
rect 14755 985 14790 986
rect 14195 948 14232 977
rect 14196 946 14232 948
rect 13773 936 13809 937
rect 13621 906 13630 926
rect 13650 906 13658 926
rect 13621 896 13658 906
rect 13717 926 13865 936
rect 13965 933 14061 935
rect 13717 906 13726 926
rect 13746 906 13836 926
rect 13856 906 13865 926
rect 13717 897 13865 906
rect 13923 926 14061 933
rect 13923 906 13932 926
rect 13952 906 14061 926
rect 14196 924 14387 946
rect 14413 945 14450 977
rect 14726 973 14790 985
rect 14830 947 14857 1125
rect 14689 945 14857 947
rect 14413 919 14857 945
rect 13923 897 14061 906
rect 13717 896 13754 897
rect 13214 842 13251 845
rect 13447 843 13488 844
rect 13339 836 13488 843
rect 12783 823 12820 828
rect 12774 819 12821 823
rect 12774 801 12793 819
rect 12811 801 12821 819
rect 13339 816 13398 836
rect 13418 816 13457 836
rect 13477 816 13488 836
rect 13339 808 13488 816
rect 13555 839 13712 846
rect 13555 819 13675 839
rect 13695 819 13712 839
rect 13555 809 13712 819
rect 13555 808 13590 809
rect 12774 738 12821 801
rect 13555 787 13586 808
rect 13773 787 13809 897
rect 13828 896 13865 897
rect 13924 896 13961 897
rect 13884 837 13974 843
rect 13884 817 13893 837
rect 13913 835 13974 837
rect 13913 817 13938 835
rect 13884 815 13938 817
rect 13958 815 13974 835
rect 13884 809 13974 815
rect 13398 786 13435 787
rect 13211 778 13248 780
rect 13211 770 13253 778
rect 13211 752 13221 770
rect 13239 752 13253 770
rect 13211 743 13253 752
rect 13397 777 13435 786
rect 13397 757 13406 777
rect 13426 757 13435 777
rect 13397 749 13435 757
rect 13501 781 13586 787
rect 13616 786 13653 787
rect 13501 761 13509 781
rect 13529 761 13586 781
rect 13501 753 13586 761
rect 13615 777 13653 786
rect 13615 757 13624 777
rect 13644 757 13653 777
rect 13501 752 13537 753
rect 13615 749 13653 757
rect 13719 785 13863 787
rect 13719 781 13771 785
rect 13719 761 13727 781
rect 13747 765 13771 781
rect 13791 781 13863 785
rect 13791 765 13835 781
rect 13747 761 13835 765
rect 13855 761 13863 781
rect 13719 753 13863 761
rect 13719 752 13755 753
rect 13827 752 13863 753
rect 13929 786 13966 787
rect 13929 785 13967 786
rect 13929 777 13993 785
rect 13929 757 13938 777
rect 13958 763 13993 777
rect 14013 763 14016 783
rect 13958 758 14016 763
rect 13958 757 13993 758
rect 12774 723 12824 738
rect 12774 698 12788 723
rect 12820 698 12824 723
rect 13212 718 13253 743
rect 13398 718 13435 749
rect 13616 727 13653 749
rect 13929 745 13993 757
rect 13611 718 13653 727
rect 14033 719 14060 897
rect 13212 706 13257 718
rect 12774 685 12821 698
rect 10159 660 10167 682
rect 10191 660 10199 682
rect 10159 652 10199 660
rect 13208 648 13257 706
rect 13398 692 13460 718
rect 13611 717 13696 718
rect 13892 717 14060 719
rect 13611 691 14060 717
rect 13611 648 13650 691
rect 13892 690 14060 691
rect 14523 695 14563 919
rect 14689 918 14857 919
rect 14921 951 14954 1284
rect 15559 1283 15586 1461
rect 15626 1423 15690 1435
rect 15966 1431 16003 1463
rect 16029 1462 16220 1484
rect 16355 1482 16464 1502
rect 16484 1482 16493 1502
rect 16355 1475 16493 1482
rect 16551 1502 16699 1511
rect 16551 1482 16560 1502
rect 16580 1482 16670 1502
rect 16690 1482 16699 1502
rect 16355 1473 16451 1475
rect 16551 1472 16699 1482
rect 16758 1502 16795 1512
rect 16758 1482 16766 1502
rect 16786 1482 16795 1502
rect 16607 1471 16643 1472
rect 16184 1460 16220 1462
rect 16184 1431 16221 1460
rect 15626 1422 15661 1423
rect 15603 1417 15661 1422
rect 15603 1397 15606 1417
rect 15626 1403 15661 1417
rect 15681 1403 15690 1423
rect 15626 1395 15690 1403
rect 15652 1394 15690 1395
rect 15653 1393 15690 1394
rect 15756 1427 15792 1428
rect 15864 1427 15900 1428
rect 15756 1419 15900 1427
rect 15756 1399 15764 1419
rect 15784 1418 15872 1419
rect 15784 1399 15819 1418
rect 15840 1399 15872 1418
rect 15892 1399 15900 1419
rect 15756 1393 15900 1399
rect 15966 1423 16004 1431
rect 16082 1427 16118 1428
rect 15966 1403 15975 1423
rect 15995 1403 16004 1423
rect 15966 1394 16004 1403
rect 16033 1419 16118 1427
rect 16033 1399 16090 1419
rect 16110 1399 16118 1419
rect 15966 1393 16003 1394
rect 16033 1393 16118 1399
rect 16184 1423 16222 1431
rect 16184 1403 16193 1423
rect 16213 1403 16222 1423
rect 16455 1412 16492 1413
rect 16758 1412 16795 1482
rect 16830 1511 16861 1562
rect 17157 1557 17202 1563
rect 17157 1539 17175 1557
rect 17193 1539 17202 1557
rect 17157 1529 17202 1539
rect 16880 1511 16917 1512
rect 16830 1502 16917 1511
rect 16830 1482 16888 1502
rect 16908 1482 16917 1502
rect 16830 1472 16917 1482
rect 16976 1502 17013 1512
rect 16976 1482 16984 1502
rect 17004 1482 17013 1502
rect 17157 1487 17200 1529
rect 17063 1485 17200 1487
rect 16830 1471 16861 1472
rect 16976 1412 17013 1482
rect 16454 1411 16795 1412
rect 16184 1394 16222 1403
rect 16379 1406 16795 1411
rect 16184 1393 16221 1394
rect 15645 1365 15735 1371
rect 15645 1345 15661 1365
rect 15681 1363 15735 1365
rect 15681 1345 15706 1363
rect 15645 1343 15706 1345
rect 15726 1343 15735 1363
rect 15645 1337 15735 1343
rect 15658 1283 15695 1284
rect 15754 1283 15791 1284
rect 15810 1283 15846 1393
rect 16033 1372 16064 1393
rect 16379 1386 16382 1406
rect 16402 1386 16795 1406
rect 16979 1396 17013 1412
rect 17057 1464 17200 1485
rect 16755 1377 16795 1386
rect 17057 1377 17084 1464
rect 17157 1438 17200 1464
rect 17157 1420 17170 1438
rect 17188 1420 17200 1438
rect 17157 1409 17200 1420
rect 16029 1371 16064 1372
rect 15907 1361 16064 1371
rect 15907 1341 15924 1361
rect 15944 1341 16064 1361
rect 15907 1334 16064 1341
rect 16131 1364 16280 1372
rect 16131 1344 16142 1364
rect 16162 1344 16201 1364
rect 16221 1344 16280 1364
rect 16755 1360 17084 1377
rect 16755 1359 16795 1360
rect 16131 1337 16280 1344
rect 17152 1348 17192 1351
rect 17152 1342 17195 1348
rect 16777 1339 17195 1342
rect 16131 1336 16172 1337
rect 15865 1283 15902 1284
rect 15558 1274 15696 1283
rect 15558 1254 15667 1274
rect 15687 1254 15696 1274
rect 15558 1247 15696 1254
rect 15754 1274 15902 1283
rect 15754 1254 15763 1274
rect 15783 1254 15873 1274
rect 15893 1254 15902 1274
rect 15558 1245 15654 1247
rect 15754 1244 15902 1254
rect 15961 1274 15998 1284
rect 15961 1254 15969 1274
rect 15989 1254 15998 1274
rect 15810 1243 15846 1244
rect 15658 1184 15695 1185
rect 15961 1184 15998 1254
rect 16033 1283 16064 1334
rect 16777 1321 17168 1339
rect 17186 1321 17195 1339
rect 16777 1319 17195 1321
rect 16777 1311 16804 1319
rect 17045 1316 17195 1319
rect 16357 1305 16525 1306
rect 16776 1305 16804 1311
rect 16357 1289 16804 1305
rect 17152 1311 17195 1316
rect 16083 1283 16120 1284
rect 16033 1274 16120 1283
rect 16033 1254 16091 1274
rect 16111 1254 16120 1274
rect 16033 1244 16120 1254
rect 16179 1274 16216 1284
rect 16179 1254 16187 1274
rect 16207 1254 16216 1274
rect 16033 1243 16064 1244
rect 15657 1183 15998 1184
rect 16179 1183 16216 1254
rect 15582 1178 15998 1183
rect 15582 1158 15585 1178
rect 15605 1158 15998 1178
rect 16029 1159 16216 1183
rect 16357 1279 16801 1289
rect 16357 1277 16525 1279
rect 16357 1099 16384 1277
rect 16424 1239 16488 1251
rect 16764 1247 16801 1279
rect 16827 1278 17018 1300
rect 16982 1276 17018 1278
rect 16982 1247 17019 1276
rect 17152 1255 17192 1311
rect 16424 1238 16459 1239
rect 16401 1233 16459 1238
rect 16401 1213 16404 1233
rect 16424 1219 16459 1233
rect 16479 1219 16488 1239
rect 16424 1211 16488 1219
rect 16450 1210 16488 1211
rect 16451 1209 16488 1210
rect 16554 1243 16590 1244
rect 16662 1243 16698 1244
rect 16554 1235 16698 1243
rect 16554 1215 16562 1235
rect 16582 1215 16617 1235
rect 16637 1215 16670 1235
rect 16690 1215 16698 1235
rect 16554 1209 16698 1215
rect 16764 1239 16802 1247
rect 16880 1243 16916 1244
rect 16764 1219 16773 1239
rect 16793 1219 16802 1239
rect 16764 1210 16802 1219
rect 16831 1235 16916 1243
rect 16831 1215 16888 1235
rect 16908 1215 16916 1235
rect 16764 1209 16801 1210
rect 16831 1209 16916 1215
rect 16982 1239 17020 1247
rect 16982 1219 16991 1239
rect 17011 1219 17020 1239
rect 17152 1237 17164 1255
rect 17182 1237 17192 1255
rect 17152 1227 17192 1237
rect 16982 1210 17020 1219
rect 16982 1209 17019 1210
rect 16443 1181 16533 1187
rect 16443 1161 16459 1181
rect 16479 1179 16533 1181
rect 16479 1161 16504 1179
rect 16443 1159 16504 1161
rect 16524 1159 16533 1179
rect 16443 1153 16533 1159
rect 16456 1099 16493 1100
rect 16552 1099 16589 1100
rect 16608 1099 16644 1209
rect 16831 1188 16862 1209
rect 16827 1187 16862 1188
rect 16705 1177 16862 1187
rect 16705 1157 16722 1177
rect 16742 1157 16862 1177
rect 16705 1150 16862 1157
rect 16929 1180 17078 1188
rect 16929 1160 16940 1180
rect 16960 1160 16999 1180
rect 17019 1160 17078 1180
rect 16929 1153 17078 1160
rect 17144 1156 17196 1174
rect 16929 1152 16970 1153
rect 16663 1099 16700 1100
rect 16356 1090 16494 1099
rect 16356 1070 16465 1090
rect 16485 1070 16494 1090
rect 16356 1063 16494 1070
rect 16552 1090 16700 1099
rect 16552 1070 16561 1090
rect 16581 1070 16671 1090
rect 16691 1070 16700 1090
rect 16356 1061 16452 1063
rect 16552 1060 16700 1070
rect 16759 1090 16796 1100
rect 16759 1070 16767 1090
rect 16787 1070 16796 1090
rect 16608 1059 16644 1060
rect 16759 1003 16796 1070
rect 16831 1099 16862 1150
rect 17144 1138 17162 1156
rect 17180 1138 17196 1156
rect 16881 1099 16918 1100
rect 16831 1090 16918 1099
rect 16831 1070 16889 1090
rect 16909 1070 16918 1090
rect 16831 1060 16918 1070
rect 16977 1090 17014 1100
rect 16977 1070 16985 1090
rect 17005 1070 17014 1090
rect 16831 1059 16862 1060
rect 16456 1000 16493 1001
rect 16759 1000 16798 1003
rect 16455 999 16798 1000
rect 16977 999 17014 1070
rect 16380 994 16798 999
rect 16380 974 16383 994
rect 16403 974 16798 994
rect 16827 975 17014 999
rect 14921 943 14958 951
rect 14921 924 14929 943
rect 14950 924 14958 943
rect 14921 918 14958 924
rect 16759 949 16798 974
rect 17144 949 17196 1138
rect 16759 931 17198 949
rect 16759 913 17159 931
rect 17177 913 17198 931
rect 16759 907 17198 913
rect 16765 903 17198 907
rect 17144 901 17196 903
rect 17147 836 17184 841
rect 17138 832 17185 836
rect 17138 814 17157 832
rect 17175 814 17185 832
rect 17138 751 17185 814
rect 17138 736 17188 751
rect 17138 711 17152 736
rect 17184 711 17188 736
rect 17138 698 17185 711
rect 14523 673 14531 695
rect 14555 673 14563 695
rect 14523 665 14563 673
rect 101 583 506 610
rect 542 583 545 610
rect 4465 596 4870 623
rect 4906 596 4909 623
rect 8842 608 9247 635
rect 9283 608 9286 635
rect 13206 621 13611 648
rect 13647 621 13650 648
rect 13206 617 13650 621
rect 13206 616 13632 617
rect 8842 604 9286 608
rect 8842 603 9268 604
rect 4465 592 4909 596
rect 4465 591 4891 592
rect 101 579 545 583
rect 101 578 527 579
rect 14965 446 15030 447
rect 10601 433 10666 434
rect 6224 421 6289 422
rect 1860 408 1925 409
rect 1511 383 1698 407
rect 1729 387 2122 408
rect 2143 387 2145 408
rect 1729 383 2145 387
rect 5875 396 6062 420
rect 6093 400 6486 421
rect 6507 400 6509 421
rect 6093 396 6509 400
rect 10252 408 10439 432
rect 10470 412 10863 433
rect 10884 412 10886 433
rect 10470 408 10886 412
rect 14616 421 14803 445
rect 14834 425 15227 446
rect 15248 425 15250 446
rect 14834 421 15250 425
rect 1511 312 1548 383
rect 1729 382 2070 383
rect 1663 322 1694 323
rect 1511 292 1520 312
rect 1540 292 1548 312
rect 1511 282 1548 292
rect 1607 312 1694 322
rect 1607 292 1616 312
rect 1636 292 1694 312
rect 1607 283 1694 292
rect 1607 282 1644 283
rect 1663 232 1694 283
rect 1729 312 1766 382
rect 2032 381 2069 382
rect 4349 334 4414 335
rect 1881 322 1917 323
rect 1729 292 1738 312
rect 1758 292 1766 312
rect 1729 282 1766 292
rect 1825 312 1973 322
rect 2073 319 2234 321
rect 1825 292 1834 312
rect 1854 292 1944 312
rect 1964 292 1973 312
rect 1825 283 1973 292
rect 2031 314 2234 319
rect 2031 312 2204 314
rect 2031 292 2040 312
rect 2060 294 2204 312
rect 2224 294 2234 314
rect 2060 292 2234 294
rect 2031 285 2234 292
rect 4000 309 4187 333
rect 4218 313 4611 334
rect 4632 313 4634 334
rect 4218 309 4634 313
rect 5875 325 5912 396
rect 6093 395 6434 396
rect 6027 335 6058 336
rect 2031 283 2169 285
rect 1825 282 1862 283
rect 1555 229 1596 230
rect 1447 222 1596 229
rect 1447 202 1506 222
rect 1526 202 1565 222
rect 1585 202 1596 222
rect 1447 194 1596 202
rect 1663 225 1820 232
rect 1663 205 1783 225
rect 1803 205 1820 225
rect 1663 195 1820 205
rect 1663 194 1698 195
rect 1663 173 1694 194
rect 1881 173 1917 283
rect 1936 282 1973 283
rect 2032 282 2069 283
rect 1992 223 2082 229
rect 1992 203 2001 223
rect 2021 221 2082 223
rect 2021 203 2046 221
rect 1992 201 2046 203
rect 2066 201 2082 221
rect 1992 195 2082 201
rect 1506 172 1543 173
rect 1505 163 1543 172
rect 1505 143 1514 163
rect 1534 143 1543 163
rect 1505 135 1543 143
rect 1609 167 1694 173
rect 1724 172 1761 173
rect 1609 147 1617 167
rect 1637 147 1694 167
rect 1609 139 1694 147
rect 1723 163 1761 172
rect 1723 143 1732 163
rect 1752 143 1761 163
rect 1609 138 1645 139
rect 1723 135 1761 143
rect 1827 168 1971 173
rect 1827 167 1888 168
rect 1827 147 1835 167
rect 1855 147 1888 167
rect 1827 144 1888 147
rect 1911 167 1971 168
rect 1911 147 1943 167
rect 1963 147 1971 167
rect 1911 144 1971 147
rect 1827 139 1971 144
rect 1827 138 1863 139
rect 1935 138 1971 139
rect 2037 172 2074 173
rect 2037 171 2075 172
rect 2037 163 2101 171
rect 2037 143 2046 163
rect 2066 149 2101 163
rect 2121 149 2124 169
rect 2066 144 2124 149
rect 2066 143 2101 144
rect 1506 106 1543 135
rect 1507 104 1543 106
rect 1507 82 1698 104
rect 1724 103 1761 135
rect 2037 131 2101 143
rect 2141 105 2168 283
rect 4000 238 4037 309
rect 4218 308 4559 309
rect 4152 248 4183 249
rect 4000 218 4009 238
rect 4029 218 4037 238
rect 4000 208 4037 218
rect 4096 238 4183 248
rect 4096 218 4105 238
rect 4125 218 4183 238
rect 4096 209 4183 218
rect 4096 208 4133 209
rect 4152 158 4183 209
rect 4218 238 4255 308
rect 4521 307 4558 308
rect 5875 305 5884 325
rect 5904 305 5912 325
rect 5875 295 5912 305
rect 5971 325 6058 335
rect 5971 305 5980 325
rect 6000 305 6058 325
rect 5971 296 6058 305
rect 5971 295 6008 296
rect 4370 248 4406 249
rect 4218 218 4227 238
rect 4247 218 4255 238
rect 4218 208 4255 218
rect 4314 238 4462 248
rect 4562 245 4684 247
rect 4314 218 4323 238
rect 4343 218 4433 238
rect 4453 218 4462 238
rect 4314 209 4462 218
rect 4520 243 4684 245
rect 6027 245 6058 296
rect 6093 325 6130 395
rect 6396 394 6433 395
rect 8797 358 8862 359
rect 6245 335 6281 336
rect 6093 305 6102 325
rect 6122 305 6130 325
rect 6093 295 6130 305
rect 6189 325 6337 335
rect 6437 332 6598 334
rect 6189 305 6198 325
rect 6218 305 6308 325
rect 6328 305 6337 325
rect 6189 296 6337 305
rect 6395 327 6598 332
rect 6395 325 6568 327
rect 6395 305 6404 325
rect 6424 307 6568 325
rect 6588 307 6598 327
rect 6424 305 6598 307
rect 6395 298 6598 305
rect 8448 333 8635 357
rect 8666 337 9059 358
rect 9080 337 9082 358
rect 8666 333 9082 337
rect 10252 337 10289 408
rect 10470 407 10811 408
rect 10404 347 10435 348
rect 6395 296 6533 298
rect 6189 295 6226 296
rect 4520 240 4723 243
rect 5919 242 5960 243
rect 4520 238 4693 240
rect 4520 218 4529 238
rect 4549 220 4693 238
rect 4713 220 4723 240
rect 4549 218 4723 220
rect 4520 211 4723 218
rect 5811 235 5960 242
rect 5811 215 5870 235
rect 5890 215 5929 235
rect 5949 215 5960 235
rect 4520 209 4658 211
rect 4314 208 4351 209
rect 4044 155 4085 156
rect 3936 148 4085 155
rect 3936 128 3995 148
rect 4015 128 4054 148
rect 4074 128 4085 148
rect 3936 120 4085 128
rect 4152 151 4309 158
rect 4152 131 4272 151
rect 4292 131 4309 151
rect 4152 121 4309 131
rect 4152 120 4187 121
rect 2000 103 2168 105
rect 1724 77 2168 103
rect 4152 99 4183 120
rect 4370 99 4406 209
rect 4425 208 4462 209
rect 4521 208 4558 209
rect 4481 149 4571 155
rect 4481 129 4490 149
rect 4510 147 4571 149
rect 4510 129 4535 147
rect 4481 127 4535 129
rect 4555 127 4571 147
rect 4481 121 4571 127
rect 3995 98 4032 99
rect 1834 74 1874 77
rect 2000 76 2168 77
rect 3994 89 4032 98
rect 3994 69 4003 89
rect 4023 69 4032 89
rect 3994 61 4032 69
rect 4098 93 4183 99
rect 4213 98 4250 99
rect 4098 73 4106 93
rect 4126 73 4183 93
rect 4098 65 4183 73
rect 4212 89 4250 98
rect 4212 69 4221 89
rect 4241 69 4250 89
rect 4098 64 4134 65
rect 4212 61 4250 69
rect 4316 93 4460 99
rect 4316 73 4324 93
rect 4344 90 4432 93
rect 4344 73 4380 90
rect 4316 69 4380 73
rect 4397 73 4432 90
rect 4452 73 4460 93
rect 4397 69 4460 73
rect 4316 65 4460 69
rect 4316 64 4352 65
rect 4424 64 4460 65
rect 4526 98 4563 99
rect 4526 97 4564 98
rect 4526 89 4590 97
rect 4526 69 4535 89
rect 4555 75 4590 89
rect 4610 75 4613 95
rect 4555 70 4613 75
rect 4555 69 4590 70
rect 3995 32 4032 61
rect 3996 30 4032 32
rect 3996 8 4187 30
rect 4213 29 4250 61
rect 4526 57 4590 69
rect 4630 31 4657 209
rect 5811 207 5960 215
rect 6027 238 6184 245
rect 6027 218 6147 238
rect 6167 218 6184 238
rect 6027 208 6184 218
rect 6027 207 6062 208
rect 6027 186 6058 207
rect 6245 186 6281 296
rect 6300 295 6337 296
rect 6396 295 6433 296
rect 6356 236 6446 242
rect 6356 216 6365 236
rect 6385 234 6446 236
rect 6385 216 6410 234
rect 6356 214 6410 216
rect 6430 214 6446 234
rect 6356 208 6446 214
rect 5870 185 5907 186
rect 5869 176 5907 185
rect 5869 156 5878 176
rect 5898 156 5907 176
rect 5869 148 5907 156
rect 5973 180 6058 186
rect 6088 185 6125 186
rect 5973 160 5981 180
rect 6001 160 6058 180
rect 5973 152 6058 160
rect 6087 176 6125 185
rect 6087 156 6096 176
rect 6116 156 6125 176
rect 5973 151 6009 152
rect 6087 148 6125 156
rect 6191 182 6335 186
rect 6191 180 6255 182
rect 6191 160 6199 180
rect 6219 160 6255 180
rect 6191 158 6255 160
rect 6278 180 6335 182
rect 6278 160 6307 180
rect 6327 160 6335 180
rect 6278 158 6335 160
rect 6191 152 6335 158
rect 6191 151 6227 152
rect 6299 151 6335 152
rect 6401 185 6438 186
rect 6401 184 6439 185
rect 6401 176 6465 184
rect 6401 156 6410 176
rect 6430 162 6465 176
rect 6485 162 6488 182
rect 6430 157 6488 162
rect 6430 156 6465 157
rect 5870 119 5907 148
rect 5871 117 5907 119
rect 5871 95 6062 117
rect 6088 116 6125 148
rect 6401 144 6465 156
rect 6505 118 6532 296
rect 8448 262 8485 333
rect 8666 332 9007 333
rect 8600 272 8631 273
rect 8448 242 8457 262
rect 8477 242 8485 262
rect 8448 232 8485 242
rect 8544 262 8631 272
rect 8544 242 8553 262
rect 8573 242 8631 262
rect 8544 233 8631 242
rect 8544 232 8581 233
rect 8600 182 8631 233
rect 8666 262 8703 332
rect 8969 331 9006 332
rect 10252 317 10261 337
rect 10281 317 10289 337
rect 10252 307 10289 317
rect 10348 337 10435 347
rect 10348 317 10357 337
rect 10377 317 10435 337
rect 10348 308 10435 317
rect 10348 307 10385 308
rect 8818 272 8854 273
rect 8666 242 8675 262
rect 8695 242 8703 262
rect 8666 232 8703 242
rect 8762 262 8910 272
rect 9010 269 9132 271
rect 8762 242 8771 262
rect 8791 242 8881 262
rect 8901 242 8910 262
rect 8762 233 8910 242
rect 8968 267 9132 269
rect 8968 264 9171 267
rect 8968 262 9141 264
rect 8968 242 8977 262
rect 8997 244 9141 262
rect 9161 244 9171 264
rect 10404 257 10435 308
rect 10470 337 10507 407
rect 10773 406 10810 407
rect 13090 359 13155 360
rect 10622 347 10658 348
rect 10470 317 10479 337
rect 10499 317 10507 337
rect 10470 307 10507 317
rect 10566 337 10714 347
rect 10814 344 10975 346
rect 10566 317 10575 337
rect 10595 317 10685 337
rect 10705 317 10714 337
rect 10566 308 10714 317
rect 10772 339 10975 344
rect 10772 337 10945 339
rect 10772 317 10781 337
rect 10801 319 10945 337
rect 10965 319 10975 339
rect 10801 317 10975 319
rect 10772 310 10975 317
rect 12741 334 12928 358
rect 12959 338 13352 359
rect 13373 338 13375 359
rect 12959 334 13375 338
rect 14616 350 14653 421
rect 14834 420 15175 421
rect 14768 360 14799 361
rect 10772 308 10910 310
rect 10566 307 10603 308
rect 10296 254 10337 255
rect 8997 242 9171 244
rect 8968 235 9171 242
rect 10188 247 10337 254
rect 8968 233 9106 235
rect 8762 232 8799 233
rect 8492 179 8533 180
rect 8379 172 8533 179
rect 8379 152 8443 172
rect 8463 152 8502 172
rect 8522 152 8533 172
rect 8379 145 8533 152
rect 8384 144 8533 145
rect 8600 175 8757 182
rect 8600 155 8720 175
rect 8740 155 8757 175
rect 8600 145 8757 155
rect 8600 144 8635 145
rect 8600 123 8631 144
rect 8818 123 8854 233
rect 8873 232 8910 233
rect 8969 232 9006 233
rect 8929 173 9019 179
rect 8929 153 8938 173
rect 8958 171 9019 173
rect 8958 153 8983 171
rect 8929 151 8983 153
rect 9003 151 9019 171
rect 8929 145 9019 151
rect 8443 122 8480 123
rect 6364 116 6532 118
rect 6088 90 6532 116
rect 6198 87 6238 90
rect 6364 89 6532 90
rect 8442 113 8480 122
rect 8442 93 8451 113
rect 8471 93 8480 113
rect 8442 85 8480 93
rect 8546 117 8631 123
rect 8661 122 8698 123
rect 8546 97 8554 117
rect 8574 97 8631 117
rect 8546 89 8631 97
rect 8660 113 8698 122
rect 8660 93 8669 113
rect 8689 93 8698 113
rect 8546 88 8582 89
rect 8660 85 8698 93
rect 8764 117 8908 123
rect 8764 97 8772 117
rect 8792 97 8880 117
rect 8900 97 8908 117
rect 8764 89 8908 97
rect 8764 88 8800 89
rect 8872 88 8908 89
rect 8974 122 9011 123
rect 8974 121 9012 122
rect 8974 113 9038 121
rect 8974 93 8983 113
rect 9003 99 9038 113
rect 9058 99 9061 119
rect 9003 94 9061 99
rect 9003 93 9038 94
rect 8443 56 8480 85
rect 8444 54 8480 56
rect 8444 32 8635 54
rect 8661 53 8698 85
rect 8974 81 9038 93
rect 9078 55 9105 233
rect 10188 227 10247 247
rect 10267 227 10306 247
rect 10326 227 10337 247
rect 10188 219 10337 227
rect 10404 250 10561 257
rect 10404 230 10524 250
rect 10544 230 10561 250
rect 10404 220 10561 230
rect 10404 219 10439 220
rect 10404 198 10435 219
rect 10622 198 10658 308
rect 10677 307 10714 308
rect 10773 307 10810 308
rect 10733 248 10823 254
rect 10733 228 10742 248
rect 10762 246 10823 248
rect 10762 228 10787 246
rect 10733 226 10787 228
rect 10807 226 10823 246
rect 10733 220 10823 226
rect 10247 197 10284 198
rect 10246 188 10284 197
rect 10246 168 10255 188
rect 10275 168 10284 188
rect 10246 160 10284 168
rect 10350 192 10435 198
rect 10465 197 10502 198
rect 10350 172 10358 192
rect 10378 172 10435 192
rect 10350 164 10435 172
rect 10464 188 10502 197
rect 10464 168 10473 188
rect 10493 168 10502 188
rect 10350 163 10386 164
rect 10464 160 10502 168
rect 10568 193 10712 198
rect 10568 192 10629 193
rect 10568 172 10576 192
rect 10596 172 10629 192
rect 10568 169 10629 172
rect 10652 192 10712 193
rect 10652 172 10684 192
rect 10704 172 10712 192
rect 10652 169 10712 172
rect 10568 164 10712 169
rect 10568 163 10604 164
rect 10676 163 10712 164
rect 10778 197 10815 198
rect 10778 196 10816 197
rect 10778 188 10842 196
rect 10778 168 10787 188
rect 10807 174 10842 188
rect 10862 174 10865 194
rect 10807 169 10865 174
rect 10807 168 10842 169
rect 10247 131 10284 160
rect 10248 129 10284 131
rect 10248 107 10439 129
rect 10465 128 10502 160
rect 10778 156 10842 168
rect 10882 130 10909 308
rect 12741 263 12778 334
rect 12959 333 13300 334
rect 12893 273 12924 274
rect 12741 243 12750 263
rect 12770 243 12778 263
rect 12741 233 12778 243
rect 12837 263 12924 273
rect 12837 243 12846 263
rect 12866 243 12924 263
rect 12837 234 12924 243
rect 12837 233 12874 234
rect 12893 183 12924 234
rect 12959 263 12996 333
rect 13262 332 13299 333
rect 14616 330 14625 350
rect 14645 330 14653 350
rect 14616 320 14653 330
rect 14712 350 14799 360
rect 14712 330 14721 350
rect 14741 330 14799 350
rect 14712 321 14799 330
rect 14712 320 14749 321
rect 13111 273 13147 274
rect 12959 243 12968 263
rect 12988 243 12996 263
rect 12959 233 12996 243
rect 13055 263 13203 273
rect 13303 270 13425 272
rect 13055 243 13064 263
rect 13084 243 13174 263
rect 13194 243 13203 263
rect 13055 234 13203 243
rect 13261 268 13425 270
rect 14768 270 14799 321
rect 14834 350 14871 420
rect 15137 419 15174 420
rect 14986 360 15022 361
rect 14834 330 14843 350
rect 14863 330 14871 350
rect 14834 320 14871 330
rect 14930 350 15078 360
rect 15178 357 15339 359
rect 14930 330 14939 350
rect 14959 330 15049 350
rect 15069 330 15078 350
rect 14930 321 15078 330
rect 15136 352 15339 357
rect 15136 350 15309 352
rect 15136 330 15145 350
rect 15165 332 15309 350
rect 15329 332 15339 352
rect 15165 330 15339 332
rect 15136 323 15339 330
rect 15136 321 15274 323
rect 14930 320 14967 321
rect 13261 265 13464 268
rect 14660 267 14701 268
rect 13261 263 13434 265
rect 13261 243 13270 263
rect 13290 245 13434 263
rect 13454 245 13464 265
rect 13290 243 13464 245
rect 13261 236 13464 243
rect 14552 260 14701 267
rect 14552 240 14611 260
rect 14631 240 14670 260
rect 14690 240 14701 260
rect 13261 234 13399 236
rect 13055 233 13092 234
rect 12785 180 12826 181
rect 12677 173 12826 180
rect 12677 153 12736 173
rect 12756 153 12795 173
rect 12815 153 12826 173
rect 12677 145 12826 153
rect 12893 176 13050 183
rect 12893 156 13013 176
rect 13033 156 13050 176
rect 12893 146 13050 156
rect 12893 145 12928 146
rect 10741 128 10909 130
rect 10465 102 10909 128
rect 12893 124 12924 145
rect 13111 124 13147 234
rect 13166 233 13203 234
rect 13262 233 13299 234
rect 13222 174 13312 180
rect 13222 154 13231 174
rect 13251 172 13312 174
rect 13251 154 13276 172
rect 13222 152 13276 154
rect 13296 152 13312 172
rect 13222 146 13312 152
rect 12736 123 12773 124
rect 10575 99 10615 102
rect 10741 101 10909 102
rect 12735 114 12773 123
rect 12735 94 12744 114
rect 12764 94 12773 114
rect 12735 86 12773 94
rect 12839 118 12924 124
rect 12954 123 12991 124
rect 12839 98 12847 118
rect 12867 98 12924 118
rect 12839 90 12924 98
rect 12953 114 12991 123
rect 12953 94 12962 114
rect 12982 94 12991 114
rect 12839 89 12875 90
rect 12953 86 12991 94
rect 13057 118 13201 124
rect 13057 98 13065 118
rect 13085 98 13117 118
rect 13057 96 13117 98
rect 13138 98 13173 118
rect 13193 98 13201 118
rect 13138 96 13201 98
rect 13057 90 13201 96
rect 13057 89 13093 90
rect 13165 89 13201 90
rect 13267 123 13304 124
rect 13267 122 13305 123
rect 13267 114 13331 122
rect 13267 94 13276 114
rect 13296 100 13331 114
rect 13351 100 13354 120
rect 13296 95 13354 100
rect 13296 94 13331 95
rect 12736 57 12773 86
rect 8937 53 9105 55
rect 4489 29 4657 31
rect 4213 3 4657 29
rect 8661 27 9105 53
rect 12737 55 12773 57
rect 12737 33 12928 55
rect 12954 54 12991 86
rect 13267 82 13331 94
rect 13371 56 13398 234
rect 14552 232 14701 240
rect 14768 263 14925 270
rect 14768 243 14888 263
rect 14908 243 14925 263
rect 14768 233 14925 243
rect 14768 232 14803 233
rect 14768 211 14799 232
rect 14986 211 15022 321
rect 15041 320 15078 321
rect 15137 320 15174 321
rect 15097 261 15187 267
rect 15097 241 15106 261
rect 15126 259 15187 261
rect 15126 241 15151 259
rect 15097 239 15151 241
rect 15171 239 15187 259
rect 15097 233 15187 239
rect 14611 210 14648 211
rect 14610 201 14648 210
rect 14610 181 14619 201
rect 14639 181 14648 201
rect 14610 173 14648 181
rect 14714 205 14799 211
rect 14829 210 14866 211
rect 14714 185 14722 205
rect 14742 185 14799 205
rect 14714 177 14799 185
rect 14828 201 14866 210
rect 14828 181 14837 201
rect 14857 181 14866 201
rect 14714 176 14750 177
rect 14828 173 14866 181
rect 14932 207 15076 211
rect 14932 205 14996 207
rect 14932 185 14940 205
rect 14960 185 14996 205
rect 14932 183 14996 185
rect 15019 205 15076 207
rect 15019 185 15048 205
rect 15068 185 15076 205
rect 15019 183 15076 185
rect 14932 177 15076 183
rect 14932 176 14968 177
rect 15040 176 15076 177
rect 15142 210 15179 211
rect 15142 209 15180 210
rect 15142 201 15206 209
rect 15142 181 15151 201
rect 15171 187 15206 201
rect 15226 187 15229 207
rect 15171 182 15229 187
rect 15171 181 15206 182
rect 14611 144 14648 173
rect 14612 142 14648 144
rect 14612 120 14803 142
rect 14829 141 14866 173
rect 15142 169 15206 181
rect 15246 143 15273 321
rect 15105 141 15273 143
rect 14829 115 15273 141
rect 14939 112 14979 115
rect 15105 114 15273 115
rect 13230 54 13398 56
rect 12954 28 13398 54
rect 8771 24 8811 27
rect 8937 26 9105 27
rect 13064 25 13104 28
rect 13230 27 13398 28
rect 4323 0 4363 3
rect 4489 2 4657 3
<< viali >>
rect 2883 8801 2907 8823
rect 2488 8553 2509 8572
rect 1035 8502 1055 8522
rect 419 8316 439 8336
rect 959 8315 979 8335
rect 801 8261 821 8281
rect 1014 8263 1034 8283
rect 1833 8318 1853 8338
rect 1217 8132 1237 8152
rect 1036 8090 1056 8110
rect 1757 8131 1777 8151
rect 1598 8078 1619 8097
rect 1812 8079 1832 8099
rect 7247 8814 7271 8836
rect 3425 8713 3445 8733
rect 3647 8711 3667 8731
rect 3480 8661 3500 8681
rect 4020 8660 4040 8680
rect 2628 8485 2648 8505
rect 2840 8490 2859 8508
rect 2683 8433 2703 8453
rect 3404 8474 3424 8494
rect 3223 8432 3243 8452
rect 2607 8246 2627 8266
rect 3426 8301 3446 8321
rect 3639 8303 3659 8323
rect 6852 8566 6873 8585
rect 5399 8515 5419 8535
rect 4783 8329 4803 8349
rect 5323 8328 5343 8348
rect 3481 8249 3501 8269
rect 4021 8248 4041 8268
rect 420 7904 440 7924
rect 960 7903 980 7923
rect 793 7853 813 7873
rect 1015 7851 1035 7871
rect 2529 8075 2549 8095
rect 2740 8082 2759 8099
rect 2584 8023 2604 8043
rect 3405 8062 3425 8082
rect 3124 8022 3144 8042
rect 5165 8274 5185 8294
rect 5378 8276 5398 8296
rect 6197 8331 6217 8351
rect 5581 8145 5601 8165
rect 5400 8103 5420 8123
rect 6121 8144 6141 8164
rect 5962 8091 5983 8110
rect 6176 8092 6196 8112
rect 7789 8726 7809 8746
rect 8011 8724 8031 8744
rect 11624 8826 11648 8848
rect 7844 8674 7864 8694
rect 8384 8673 8404 8693
rect 6992 8498 7012 8518
rect 7204 8503 7223 8521
rect 7047 8446 7067 8466
rect 7768 8487 7788 8507
rect 7587 8445 7607 8465
rect 6971 8259 6991 8279
rect 7790 8314 7810 8334
rect 8003 8316 8023 8336
rect 11229 8578 11250 8597
rect 9776 8527 9796 8547
rect 9160 8341 9180 8361
rect 9700 8340 9720 8360
rect 7845 8262 7865 8282
rect 8385 8261 8405 8281
rect 4784 7917 4804 7937
rect 2508 7836 2528 7856
rect 5324 7916 5344 7936
rect 5157 7866 5177 7886
rect 5379 7864 5399 7884
rect 1553 7761 1577 7783
rect 2866 7783 2890 7805
rect 1915 7710 1935 7730
rect 1299 7524 1319 7544
rect 1018 7484 1038 7504
rect 1839 7523 1859 7543
rect 1682 7471 1703 7490
rect 1894 7471 1914 7491
rect 6893 8088 6913 8108
rect 7104 8095 7123 8112
rect 6948 8036 6968 8056
rect 7769 8075 7789 8095
rect 7488 8035 7508 8055
rect 9542 8286 9562 8306
rect 9755 8288 9775 8308
rect 10574 8343 10594 8363
rect 9958 8157 9978 8177
rect 9777 8115 9797 8135
rect 10498 8156 10518 8176
rect 10339 8103 10360 8122
rect 10553 8104 10573 8124
rect 15988 8839 16012 8861
rect 12166 8738 12186 8758
rect 12388 8736 12408 8756
rect 12221 8686 12241 8706
rect 12761 8685 12781 8705
rect 11369 8510 11389 8530
rect 11581 8515 11600 8533
rect 11424 8458 11444 8478
rect 12145 8499 12165 8519
rect 11964 8457 11984 8477
rect 11348 8271 11368 8291
rect 12167 8326 12187 8346
rect 12380 8328 12400 8348
rect 15593 8591 15614 8610
rect 14140 8540 14160 8560
rect 13524 8354 13544 8374
rect 14064 8353 14084 8373
rect 12222 8274 12242 8294
rect 12762 8273 12782 8293
rect 9161 7929 9181 7949
rect 6872 7849 6892 7869
rect 9701 7928 9721 7948
rect 9534 7878 9554 7898
rect 9756 7876 9776 7896
rect 5917 7774 5941 7796
rect 7230 7796 7254 7818
rect 3408 7695 3428 7715
rect 3630 7693 3650 7713
rect 3463 7643 3483 7663
rect 6279 7723 6299 7743
rect 4003 7642 4023 7662
rect 402 7298 422 7318
rect 942 7297 962 7317
rect 784 7243 804 7263
rect 997 7245 1017 7265
rect 1816 7300 1836 7320
rect 1200 7114 1220 7134
rect 1019 7072 1039 7092
rect 1740 7113 1760 7133
rect 1584 7058 1603 7076
rect 1795 7061 1815 7081
rect 403 6886 423 6906
rect 943 6885 963 6905
rect 776 6835 796 6855
rect 998 6833 1018 6853
rect 2611 7467 2631 7487
rect 2824 7469 2845 7488
rect 2666 7415 2686 7435
rect 3387 7456 3407 7476
rect 3206 7414 3226 7434
rect 2431 7316 2453 7334
rect 2590 7228 2610 7248
rect 3409 7283 3429 7303
rect 3622 7285 3642 7305
rect 5663 7537 5683 7557
rect 5382 7497 5402 7517
rect 6203 7536 6223 7556
rect 6046 7484 6067 7503
rect 6258 7484 6278 7504
rect 11270 8100 11290 8120
rect 11481 8107 11500 8124
rect 11325 8048 11345 8068
rect 12146 8087 12166 8107
rect 11865 8047 11885 8067
rect 13906 8299 13926 8319
rect 14119 8301 14139 8321
rect 14938 8356 14958 8376
rect 14322 8170 14342 8190
rect 14141 8128 14161 8148
rect 14862 8169 14882 8189
rect 14703 8116 14724 8135
rect 14917 8117 14937 8137
rect 16530 8751 16550 8771
rect 16752 8749 16772 8769
rect 16585 8699 16605 8719
rect 17125 8698 17145 8718
rect 15733 8523 15753 8543
rect 15945 8528 15964 8546
rect 15788 8471 15808 8491
rect 16509 8512 16529 8532
rect 16328 8470 16348 8490
rect 15712 8284 15732 8304
rect 16531 8339 16551 8359
rect 16744 8341 16764 8361
rect 16586 8287 16606 8307
rect 17126 8286 17146 8306
rect 13525 7942 13545 7962
rect 11249 7861 11269 7881
rect 14065 7941 14085 7961
rect 13898 7891 13918 7911
rect 14120 7889 14140 7909
rect 10294 7786 10318 7808
rect 11607 7808 11631 7830
rect 7772 7708 7792 7728
rect 7994 7706 8014 7726
rect 7827 7656 7847 7676
rect 10656 7735 10676 7755
rect 8367 7655 8387 7675
rect 4766 7311 4786 7331
rect 5306 7310 5326 7330
rect 3464 7231 3484 7251
rect 4004 7230 4024 7250
rect 2232 7120 2256 7142
rect 1934 6994 1955 7013
rect 1536 6743 1560 6765
rect 1961 6690 1981 6710
rect 1345 6504 1365 6524
rect 998 6466 1018 6486
rect 1885 6503 1905 6523
rect 1729 6450 1747 6468
rect 1940 6451 1960 6471
rect 382 6280 402 6300
rect 922 6279 942 6299
rect 764 6225 784 6245
rect 977 6227 997 6247
rect 1796 6282 1816 6302
rect 1180 6096 1200 6116
rect 999 6054 1019 6074
rect 1720 6095 1740 6115
rect 1561 6042 1582 6061
rect 1775 6043 1795 6063
rect 383 5868 403 5888
rect 923 5867 943 5887
rect 756 5817 776 5837
rect 978 5815 998 5835
rect 1516 5725 1540 5747
rect 1878 5674 1898 5694
rect 1262 5488 1282 5508
rect 981 5448 1001 5468
rect 1802 5487 1822 5507
rect 1647 5431 1666 5448
rect 1857 5435 1877 5455
rect 365 5262 385 5282
rect 905 5261 925 5281
rect 747 5207 767 5227
rect 960 5209 980 5229
rect 1959 5364 1981 5382
rect 1779 5264 1799 5284
rect 1163 5078 1183 5098
rect 982 5036 1002 5056
rect 1703 5077 1723 5097
rect 1547 5022 1566 5040
rect 1758 5025 1778 5045
rect 366 4850 386 4870
rect 906 4849 926 4869
rect 739 4799 759 4819
rect 961 4797 981 4817
rect 2446 7059 2466 7079
rect 2657 7057 2680 7079
rect 2501 7007 2521 7027
rect 3388 7044 3408 7064
rect 3041 7006 3061 7026
rect 5148 7256 5168 7276
rect 5361 7258 5381 7278
rect 6180 7313 6200 7333
rect 5564 7127 5584 7147
rect 5383 7085 5403 7105
rect 6104 7126 6124 7146
rect 5948 7071 5967 7089
rect 6159 7074 6179 7094
rect 2425 6820 2445 6840
rect 4767 6899 4787 6919
rect 5307 6898 5327 6918
rect 5140 6848 5160 6868
rect 5362 6846 5382 6866
rect 2846 6765 2870 6787
rect 2451 6517 2472 6536
rect 6975 7480 6995 7500
rect 7188 7482 7209 7501
rect 7030 7428 7050 7448
rect 7751 7469 7771 7489
rect 7570 7427 7590 7447
rect 6795 7329 6817 7347
rect 6954 7241 6974 7261
rect 7773 7296 7793 7316
rect 7986 7298 8006 7318
rect 10040 7549 10060 7569
rect 9759 7509 9779 7529
rect 10580 7548 10600 7568
rect 10423 7496 10444 7515
rect 10635 7496 10655 7516
rect 15634 8113 15654 8133
rect 15845 8120 15864 8137
rect 15689 8061 15709 8081
rect 16510 8100 16530 8120
rect 16229 8060 16249 8080
rect 15613 7874 15633 7894
rect 14658 7799 14682 7821
rect 15971 7821 15995 7843
rect 12149 7720 12169 7740
rect 12371 7718 12391 7738
rect 12204 7668 12224 7688
rect 15020 7748 15040 7768
rect 12744 7667 12764 7687
rect 9143 7323 9163 7343
rect 9683 7322 9703 7342
rect 7828 7244 7848 7264
rect 8368 7243 8388 7263
rect 6596 7133 6620 7155
rect 6298 7007 6319 7026
rect 5900 6756 5924 6778
rect 3388 6677 3408 6697
rect 3610 6675 3630 6695
rect 3443 6625 3463 6645
rect 3983 6624 4003 6644
rect 6325 6703 6345 6723
rect 2591 6449 2611 6469
rect 2803 6454 2822 6472
rect 2646 6397 2666 6417
rect 3367 6438 3387 6458
rect 3186 6396 3206 6416
rect 2570 6210 2590 6230
rect 3389 6265 3409 6285
rect 3602 6267 3622 6287
rect 5709 6517 5729 6537
rect 5362 6479 5382 6499
rect 6249 6516 6269 6536
rect 6093 6463 6111 6481
rect 6304 6464 6324 6484
rect 4746 6293 4766 6313
rect 5286 6292 5306 6312
rect 3444 6213 3464 6233
rect 3984 6212 4004 6232
rect 2492 6039 2512 6059
rect 2703 6040 2724 6059
rect 2547 5987 2567 6007
rect 3368 6026 3388 6046
rect 3087 5986 3107 6006
rect 5128 6238 5148 6258
rect 5341 6240 5361 6260
rect 6160 6295 6180 6315
rect 5544 6109 5564 6129
rect 5363 6067 5383 6087
rect 6084 6108 6104 6128
rect 5925 6055 5946 6074
rect 6139 6056 6159 6076
rect 4747 5881 4767 5901
rect 2471 5800 2491 5820
rect 5287 5880 5307 5900
rect 5120 5830 5140 5850
rect 5342 5828 5362 5848
rect 2829 5747 2853 5769
rect 5880 5738 5904 5760
rect 3371 5659 3391 5679
rect 3593 5657 3613 5677
rect 3426 5607 3446 5627
rect 6242 5687 6262 5707
rect 3966 5606 3986 5626
rect 2574 5431 2594 5451
rect 2787 5433 2808 5452
rect 2629 5379 2649 5399
rect 3350 5420 3370 5440
rect 3169 5378 3189 5398
rect 2553 5192 2573 5212
rect 3372 5247 3392 5267
rect 3585 5249 3605 5269
rect 5626 5501 5646 5521
rect 5345 5461 5365 5481
rect 6166 5500 6186 5520
rect 6011 5444 6030 5461
rect 6221 5448 6241 5468
rect 4729 5275 4749 5295
rect 5269 5274 5289 5294
rect 3427 5195 3447 5215
rect 3967 5194 3987 5214
rect 1897 4958 1918 4977
rect 2270 5025 2290 5045
rect 2482 5024 2508 5050
rect 2325 4973 2345 4993
rect 3351 5008 3371 5028
rect 2865 4972 2885 4992
rect 5111 5220 5131 5240
rect 5324 5222 5344 5242
rect 6323 5377 6345 5395
rect 6143 5277 6163 5297
rect 5527 5091 5547 5111
rect 5346 5049 5366 5069
rect 6067 5090 6087 5110
rect 5911 5035 5930 5053
rect 6122 5038 6142 5058
rect 2249 4786 2269 4806
rect 4730 4863 4750 4883
rect 5270 4862 5290 4882
rect 5103 4812 5123 4832
rect 5325 4810 5345 4830
rect 1499 4707 1523 4729
rect 2810 4729 2834 4751
rect 2064 4652 2084 4672
rect 1448 4466 1468 4486
rect 962 4430 982 4450
rect 1988 4465 2008 4485
rect 1826 4402 1849 4425
rect 2043 4413 2063 4433
rect 2415 4481 2436 4500
rect 346 4244 366 4264
rect 886 4243 906 4263
rect 728 4189 748 4209
rect 941 4191 961 4211
rect 1760 4246 1780 4266
rect 1144 4060 1164 4080
rect 963 4018 983 4038
rect 1684 4059 1704 4079
rect 1525 4006 1546 4025
rect 1739 4007 1759 4027
rect 347 3832 367 3852
rect 887 3831 907 3851
rect 720 3781 740 3801
rect 942 3779 962 3799
rect 1480 3689 1504 3711
rect 1842 3638 1862 3658
rect 1226 3452 1246 3472
rect 945 3412 965 3432
rect 1766 3451 1786 3471
rect 1609 3399 1630 3418
rect 1821 3399 1841 3419
rect 329 3226 349 3246
rect 869 3225 889 3245
rect 711 3171 731 3191
rect 924 3173 944 3193
rect 1743 3228 1763 3248
rect 1127 3042 1147 3062
rect 946 3000 966 3020
rect 1667 3041 1687 3061
rect 1511 2986 1530 3004
rect 1722 2989 1742 3009
rect 330 2814 350 2834
rect 870 2813 890 2833
rect 703 2763 723 2783
rect 925 2761 945 2781
rect 1861 2922 1882 2941
rect 1463 2671 1487 2693
rect 1888 2618 1908 2638
rect 1272 2432 1292 2452
rect 925 2394 945 2414
rect 1812 2431 1832 2451
rect 1653 2379 1676 2401
rect 1867 2379 1887 2399
rect 6810 7072 6830 7092
rect 7021 7070 7044 7092
rect 6865 7020 6885 7040
rect 7752 7057 7772 7077
rect 7405 7019 7425 7039
rect 9525 7268 9545 7288
rect 9738 7270 9758 7290
rect 10557 7325 10577 7345
rect 9941 7139 9961 7159
rect 9760 7097 9780 7117
rect 10481 7138 10501 7158
rect 10325 7083 10344 7101
rect 10536 7086 10556 7106
rect 6789 6833 6809 6853
rect 9144 6911 9164 6931
rect 9684 6910 9704 6930
rect 9517 6860 9537 6880
rect 9739 6858 9759 6878
rect 7210 6778 7234 6800
rect 6815 6530 6836 6549
rect 11352 7492 11372 7512
rect 11565 7494 11586 7513
rect 11407 7440 11427 7460
rect 12128 7481 12148 7501
rect 11947 7439 11967 7459
rect 11172 7341 11194 7359
rect 11331 7253 11351 7273
rect 12150 7308 12170 7328
rect 12363 7310 12383 7330
rect 14404 7562 14424 7582
rect 14123 7522 14143 7542
rect 14944 7561 14964 7581
rect 14787 7509 14808 7528
rect 14999 7509 15019 7529
rect 16513 7733 16533 7753
rect 16735 7731 16755 7751
rect 16568 7681 16588 7701
rect 17108 7680 17128 7700
rect 13507 7336 13527 7356
rect 14047 7335 14067 7355
rect 12205 7256 12225 7276
rect 12745 7255 12765 7275
rect 10973 7145 10997 7167
rect 10675 7019 10696 7038
rect 10277 6768 10301 6790
rect 7752 6690 7772 6710
rect 7974 6688 7994 6708
rect 7807 6638 7827 6658
rect 8347 6637 8367 6657
rect 10702 6715 10722 6735
rect 6955 6462 6975 6482
rect 7167 6467 7186 6485
rect 7010 6410 7030 6430
rect 7731 6451 7751 6471
rect 7550 6409 7570 6429
rect 6934 6223 6954 6243
rect 7753 6278 7773 6298
rect 7966 6280 7986 6300
rect 10086 6529 10106 6549
rect 9739 6491 9759 6511
rect 10626 6528 10646 6548
rect 10470 6475 10488 6493
rect 10681 6476 10701 6496
rect 9123 6305 9143 6325
rect 9663 6304 9683 6324
rect 7808 6226 7828 6246
rect 8348 6225 8368 6245
rect 6856 6052 6876 6072
rect 7067 6053 7088 6072
rect 6911 6000 6931 6020
rect 7732 6039 7752 6059
rect 7451 5999 7471 6019
rect 9505 6250 9525 6270
rect 9718 6252 9738 6272
rect 10537 6307 10557 6327
rect 9921 6121 9941 6141
rect 9740 6079 9760 6099
rect 10461 6120 10481 6140
rect 10302 6067 10323 6086
rect 10516 6068 10536 6088
rect 9124 5893 9144 5913
rect 6835 5813 6855 5833
rect 9664 5892 9684 5912
rect 9497 5842 9517 5862
rect 9719 5840 9739 5860
rect 7193 5760 7217 5782
rect 10257 5750 10281 5772
rect 7735 5672 7755 5692
rect 7957 5670 7977 5690
rect 7790 5620 7810 5640
rect 10619 5699 10639 5719
rect 8330 5619 8350 5639
rect 6938 5444 6958 5464
rect 7151 5446 7172 5465
rect 6993 5392 7013 5412
rect 7714 5433 7734 5453
rect 7533 5391 7553 5411
rect 6917 5205 6937 5225
rect 7736 5260 7756 5280
rect 7949 5262 7969 5282
rect 10003 5513 10023 5533
rect 9722 5473 9742 5493
rect 10543 5512 10563 5532
rect 10388 5456 10407 5473
rect 10598 5460 10618 5480
rect 9106 5287 9126 5307
rect 9646 5286 9666 5306
rect 7791 5208 7811 5228
rect 8331 5207 8351 5227
rect 6261 4971 6282 4990
rect 6634 5038 6654 5058
rect 6846 5037 6872 5063
rect 6689 4986 6709 5006
rect 7715 5021 7735 5041
rect 7229 4985 7249 5005
rect 9488 5232 9508 5252
rect 9701 5234 9721 5254
rect 10700 5389 10722 5407
rect 10520 5289 10540 5309
rect 9904 5103 9924 5123
rect 9723 5061 9743 5081
rect 10444 5102 10464 5122
rect 10288 5047 10307 5065
rect 10499 5050 10519 5070
rect 6613 4799 6633 4819
rect 9107 4875 9127 4895
rect 9647 4874 9667 4894
rect 9480 4824 9500 4844
rect 9702 4822 9722 4842
rect 5863 4720 5887 4742
rect 7174 4742 7198 4764
rect 3352 4641 3372 4661
rect 3574 4639 3594 4659
rect 3407 4589 3427 4609
rect 3947 4588 3967 4608
rect 6428 4665 6448 4685
rect 2555 4413 2575 4433
rect 2767 4418 2786 4436
rect 2610 4361 2630 4381
rect 3331 4402 3351 4422
rect 3150 4360 3170 4380
rect 2534 4174 2554 4194
rect 2352 4076 2374 4094
rect 3353 4229 3373 4249
rect 3566 4231 3586 4251
rect 5812 4479 5832 4499
rect 5326 4443 5346 4463
rect 6352 4478 6372 4498
rect 6190 4415 6213 4438
rect 6407 4426 6427 4446
rect 6779 4494 6800 4513
rect 4710 4257 4730 4277
rect 5250 4256 5270 4276
rect 3408 4177 3428 4197
rect 3948 4176 3968 4196
rect 2456 4003 2476 4023
rect 2667 4010 2686 4027
rect 2511 3951 2531 3971
rect 3332 3990 3352 4010
rect 3051 3950 3071 3970
rect 5092 4202 5112 4222
rect 5305 4204 5325 4224
rect 6124 4259 6144 4279
rect 5508 4073 5528 4093
rect 5327 4031 5347 4051
rect 6048 4072 6068 4092
rect 5889 4019 5910 4038
rect 6103 4020 6123 4040
rect 4711 3845 4731 3865
rect 2435 3764 2455 3784
rect 5251 3844 5271 3864
rect 5084 3794 5104 3814
rect 5306 3792 5326 3812
rect 2793 3711 2817 3733
rect 5844 3702 5868 3724
rect 3335 3623 3355 3643
rect 3557 3621 3577 3641
rect 3390 3571 3410 3591
rect 6206 3651 6226 3671
rect 3930 3570 3950 3590
rect 2538 3395 2558 3415
rect 2751 3397 2772 3416
rect 2593 3343 2613 3363
rect 3314 3384 3334 3404
rect 3133 3342 3153 3362
rect 2517 3156 2537 3176
rect 3336 3211 3356 3231
rect 3549 3213 3569 3233
rect 5590 3465 5610 3485
rect 5309 3425 5329 3445
rect 6130 3464 6150 3484
rect 5973 3412 5994 3431
rect 6185 3412 6205 3432
rect 4693 3239 4713 3259
rect 5233 3238 5253 3258
rect 3391 3159 3411 3179
rect 3931 3158 3951 3178
rect 2373 2987 2393 3007
rect 2586 2990 2604 3008
rect 2428 2935 2448 2955
rect 3315 2972 3335 2992
rect 2968 2934 2988 2954
rect 5075 3184 5095 3204
rect 5288 3186 5308 3206
rect 6107 3241 6127 3261
rect 5491 3055 5511 3075
rect 5310 3013 5330 3033
rect 6031 3054 6051 3074
rect 5875 2999 5894 3017
rect 6086 3002 6106 3022
rect 2352 2748 2372 2768
rect 4694 2827 4714 2847
rect 5234 2826 5254 2846
rect 5067 2776 5087 2796
rect 5289 2774 5309 2794
rect 2773 2693 2797 2715
rect 2378 2445 2399 2464
rect 2077 2316 2101 2338
rect 309 2208 329 2228
rect 849 2207 869 2227
rect 691 2153 711 2173
rect 904 2155 924 2175
rect 1723 2210 1743 2230
rect 1880 2124 1902 2142
rect 1107 2024 1127 2044
rect 926 1982 946 2002
rect 1647 2023 1667 2043
rect 1488 1970 1509 1989
rect 1702 1971 1722 1991
rect 6225 2935 6246 2954
rect 5827 2684 5851 2706
rect 3315 2605 3335 2625
rect 3537 2603 3557 2623
rect 3370 2553 3390 2573
rect 3910 2552 3930 2572
rect 6252 2631 6272 2651
rect 2518 2377 2538 2397
rect 2730 2382 2749 2400
rect 2573 2325 2593 2345
rect 3294 2366 3314 2386
rect 3113 2324 3133 2344
rect 2497 2138 2517 2158
rect 3316 2193 3336 2213
rect 3529 2195 3549 2215
rect 5636 2445 5656 2465
rect 5289 2407 5309 2427
rect 6176 2444 6196 2464
rect 6017 2392 6040 2414
rect 6231 2392 6251 2412
rect 11187 7084 11207 7104
rect 11398 7082 11421 7104
rect 11242 7032 11262 7052
rect 12129 7069 12149 7089
rect 11782 7031 11802 7051
rect 13889 7281 13909 7301
rect 14102 7283 14122 7303
rect 14921 7338 14941 7358
rect 14305 7152 14325 7172
rect 14124 7110 14144 7130
rect 14845 7151 14865 7171
rect 14689 7096 14708 7114
rect 14900 7099 14920 7119
rect 11166 6845 11186 6865
rect 13508 6924 13528 6944
rect 14048 6923 14068 6943
rect 13881 6873 13901 6893
rect 14103 6871 14123 6891
rect 11587 6790 11611 6812
rect 11192 6542 11213 6561
rect 15716 7505 15736 7525
rect 15929 7507 15950 7526
rect 15771 7453 15791 7473
rect 16492 7494 16512 7514
rect 16311 7452 16331 7472
rect 15536 7354 15558 7372
rect 15695 7266 15715 7286
rect 16514 7321 16534 7341
rect 16727 7323 16747 7343
rect 16569 7269 16589 7289
rect 17109 7268 17129 7288
rect 15337 7158 15361 7180
rect 15039 7032 15060 7051
rect 14641 6781 14665 6803
rect 12129 6702 12149 6722
rect 12351 6700 12371 6720
rect 12184 6650 12204 6670
rect 12724 6649 12744 6669
rect 15066 6728 15086 6748
rect 11332 6474 11352 6494
rect 11544 6479 11563 6497
rect 11387 6422 11407 6442
rect 12108 6463 12128 6483
rect 11927 6421 11947 6441
rect 11311 6235 11331 6255
rect 12130 6290 12150 6310
rect 12343 6292 12363 6312
rect 14450 6542 14470 6562
rect 14103 6504 14123 6524
rect 14990 6541 15010 6561
rect 14834 6488 14852 6506
rect 15045 6489 15065 6509
rect 13487 6318 13507 6338
rect 14027 6317 14047 6337
rect 12185 6238 12205 6258
rect 12725 6237 12745 6257
rect 11233 6064 11253 6084
rect 11444 6065 11465 6084
rect 11288 6012 11308 6032
rect 12109 6051 12129 6071
rect 11828 6011 11848 6031
rect 13869 6263 13889 6283
rect 14082 6265 14102 6285
rect 14901 6320 14921 6340
rect 14285 6134 14305 6154
rect 14104 6092 14124 6112
rect 14825 6133 14845 6153
rect 14666 6080 14687 6099
rect 14880 6081 14900 6101
rect 13488 5906 13508 5926
rect 11212 5825 11232 5845
rect 14028 5905 14048 5925
rect 13861 5855 13881 5875
rect 14083 5853 14103 5873
rect 11570 5772 11594 5794
rect 14621 5763 14645 5785
rect 12112 5684 12132 5704
rect 12334 5682 12354 5702
rect 12167 5632 12187 5652
rect 14983 5712 15003 5732
rect 12707 5631 12727 5651
rect 11315 5456 11335 5476
rect 11528 5458 11549 5477
rect 11370 5404 11390 5424
rect 12091 5445 12111 5465
rect 11910 5403 11930 5423
rect 11294 5217 11314 5237
rect 12113 5272 12133 5292
rect 12326 5274 12346 5294
rect 14367 5526 14387 5546
rect 14086 5486 14106 5506
rect 14907 5525 14927 5545
rect 14752 5469 14771 5486
rect 14962 5473 14982 5493
rect 13470 5300 13490 5320
rect 14010 5299 14030 5319
rect 12168 5220 12188 5240
rect 12708 5219 12728 5239
rect 10638 4983 10659 5002
rect 11011 5050 11031 5070
rect 11223 5049 11249 5075
rect 11066 4998 11086 5018
rect 12092 5033 12112 5053
rect 11606 4997 11626 5017
rect 13852 5245 13872 5265
rect 14065 5247 14085 5267
rect 15064 5402 15086 5420
rect 14884 5302 14904 5322
rect 14268 5116 14288 5136
rect 14087 5074 14107 5094
rect 14808 5115 14828 5135
rect 14652 5060 14671 5078
rect 14863 5063 14883 5083
rect 10990 4811 11010 4831
rect 13471 4888 13491 4908
rect 14011 4887 14031 4907
rect 13844 4837 13864 4857
rect 14066 4835 14086 4855
rect 10240 4732 10264 4754
rect 11551 4754 11575 4776
rect 7716 4654 7736 4674
rect 7938 4652 7958 4672
rect 7771 4602 7791 4622
rect 8311 4601 8331 4621
rect 10805 4677 10825 4697
rect 6919 4426 6939 4446
rect 7131 4431 7150 4449
rect 6974 4374 6994 4394
rect 7695 4415 7715 4435
rect 7514 4373 7534 4393
rect 6898 4187 6918 4207
rect 6716 4089 6738 4107
rect 7717 4242 7737 4262
rect 7930 4244 7950 4264
rect 10189 4491 10209 4511
rect 9703 4455 9723 4475
rect 10729 4490 10749 4510
rect 10567 4427 10590 4450
rect 10784 4438 10804 4458
rect 11156 4506 11177 4525
rect 9087 4269 9107 4289
rect 9627 4268 9647 4288
rect 7772 4190 7792 4210
rect 8312 4189 8332 4209
rect 6820 4016 6840 4036
rect 7031 4023 7050 4040
rect 6875 3964 6895 3984
rect 7696 4003 7716 4023
rect 7415 3963 7435 3983
rect 9469 4214 9489 4234
rect 9682 4216 9702 4236
rect 10501 4271 10521 4291
rect 9885 4085 9905 4105
rect 9704 4043 9724 4063
rect 10425 4084 10445 4104
rect 10266 4031 10287 4050
rect 10480 4032 10500 4052
rect 9088 3857 9108 3877
rect 6799 3777 6819 3797
rect 9628 3856 9648 3876
rect 9461 3806 9481 3826
rect 9683 3804 9703 3824
rect 7157 3724 7181 3746
rect 10221 3714 10245 3736
rect 7699 3636 7719 3656
rect 7921 3634 7941 3654
rect 7754 3584 7774 3604
rect 10583 3663 10603 3683
rect 8294 3583 8314 3603
rect 6902 3408 6922 3428
rect 7115 3410 7136 3429
rect 6957 3356 6977 3376
rect 7678 3397 7698 3417
rect 7497 3355 7517 3375
rect 6881 3169 6901 3189
rect 7700 3224 7720 3244
rect 7913 3226 7933 3246
rect 9967 3477 9987 3497
rect 9686 3437 9706 3457
rect 10507 3476 10527 3496
rect 10350 3424 10371 3443
rect 10562 3424 10582 3444
rect 9070 3251 9090 3271
rect 9610 3250 9630 3270
rect 7755 3172 7775 3192
rect 8295 3171 8315 3191
rect 6737 3000 6757 3020
rect 6950 3003 6968 3021
rect 6792 2948 6812 2968
rect 7679 2985 7699 3005
rect 7332 2947 7352 2967
rect 9452 3196 9472 3216
rect 9665 3198 9685 3218
rect 10484 3253 10504 3273
rect 9868 3067 9888 3087
rect 9687 3025 9707 3045
rect 10408 3066 10428 3086
rect 10252 3011 10271 3029
rect 10463 3014 10483 3034
rect 6716 2761 6736 2781
rect 9071 2839 9091 2859
rect 9611 2838 9631 2858
rect 9444 2788 9464 2808
rect 9666 2786 9686 2806
rect 7137 2706 7161 2728
rect 6742 2458 6763 2477
rect 6441 2329 6465 2351
rect 4673 2221 4693 2241
rect 5213 2220 5233 2240
rect 3371 2141 3391 2161
rect 3911 2140 3931 2160
rect 310 1796 330 1816
rect 850 1795 870 1815
rect 683 1745 703 1765
rect 905 1743 925 1763
rect 2419 1967 2439 1987
rect 2630 1968 2651 1987
rect 2474 1915 2494 1935
rect 3295 1954 3315 1974
rect 3014 1914 3034 1934
rect 5055 2166 5075 2186
rect 5268 2168 5288 2188
rect 6087 2223 6107 2243
rect 6244 2137 6266 2155
rect 5471 2037 5491 2057
rect 5290 1995 5310 2015
rect 6011 2036 6031 2056
rect 5852 1983 5873 2002
rect 6066 1984 6086 2004
rect 10602 2947 10623 2966
rect 10204 2696 10228 2718
rect 7679 2618 7699 2638
rect 7901 2616 7921 2636
rect 7734 2566 7754 2586
rect 8274 2565 8294 2585
rect 10629 2643 10649 2663
rect 6882 2390 6902 2410
rect 7094 2395 7113 2413
rect 6937 2338 6957 2358
rect 7658 2379 7678 2399
rect 7477 2337 7497 2357
rect 6861 2151 6881 2171
rect 7680 2206 7700 2226
rect 7893 2208 7913 2228
rect 10013 2457 10033 2477
rect 9666 2419 9686 2439
rect 10553 2456 10573 2476
rect 10394 2404 10417 2426
rect 10608 2404 10628 2424
rect 15551 7097 15571 7117
rect 15762 7095 15785 7117
rect 15606 7045 15626 7065
rect 16493 7082 16513 7102
rect 16146 7044 16166 7064
rect 15530 6858 15550 6878
rect 15951 6803 15975 6825
rect 15556 6555 15577 6574
rect 16493 6715 16513 6735
rect 16715 6713 16735 6733
rect 16548 6663 16568 6683
rect 17088 6662 17108 6682
rect 15696 6487 15716 6507
rect 15908 6492 15927 6510
rect 15751 6435 15771 6455
rect 16472 6476 16492 6496
rect 16291 6434 16311 6454
rect 15675 6248 15695 6268
rect 16494 6303 16514 6323
rect 16707 6305 16727 6325
rect 16549 6251 16569 6271
rect 17089 6250 17109 6270
rect 15597 6077 15617 6097
rect 15808 6078 15829 6097
rect 15652 6025 15672 6045
rect 16473 6064 16493 6084
rect 16192 6024 16212 6044
rect 15576 5838 15596 5858
rect 15934 5785 15958 5807
rect 16476 5697 16496 5717
rect 16698 5695 16718 5715
rect 16531 5645 16551 5665
rect 17071 5644 17091 5664
rect 15679 5469 15699 5489
rect 15892 5471 15913 5490
rect 15734 5417 15754 5437
rect 16455 5458 16475 5478
rect 16274 5416 16294 5436
rect 15658 5230 15678 5250
rect 16477 5285 16497 5305
rect 16690 5287 16710 5307
rect 16532 5233 16552 5253
rect 17072 5232 17092 5252
rect 15002 4996 15023 5015
rect 15375 5063 15395 5083
rect 15587 5062 15613 5088
rect 15430 5011 15450 5031
rect 16456 5046 16476 5066
rect 15970 5010 15990 5030
rect 15354 4824 15374 4844
rect 14604 4745 14628 4767
rect 15915 4767 15939 4789
rect 12093 4666 12113 4686
rect 12315 4664 12335 4684
rect 12148 4614 12168 4634
rect 12688 4613 12708 4633
rect 15169 4690 15189 4710
rect 11296 4438 11316 4458
rect 11508 4443 11527 4461
rect 11351 4386 11371 4406
rect 12072 4427 12092 4447
rect 11891 4385 11911 4405
rect 11275 4199 11295 4219
rect 11093 4101 11115 4119
rect 12094 4254 12114 4274
rect 12307 4256 12327 4276
rect 14553 4504 14573 4524
rect 14067 4468 14087 4488
rect 15093 4503 15113 4523
rect 14931 4440 14954 4463
rect 15148 4451 15168 4471
rect 15520 4519 15541 4538
rect 13451 4282 13471 4302
rect 13991 4281 14011 4301
rect 12149 4202 12169 4222
rect 12689 4201 12709 4221
rect 11197 4028 11217 4048
rect 11408 4035 11427 4052
rect 11252 3976 11272 3996
rect 12073 4015 12093 4035
rect 11792 3975 11812 3995
rect 13833 4227 13853 4247
rect 14046 4229 14066 4249
rect 14865 4284 14885 4304
rect 14249 4098 14269 4118
rect 14068 4056 14088 4076
rect 14789 4097 14809 4117
rect 14630 4044 14651 4063
rect 14844 4045 14864 4065
rect 13452 3870 13472 3890
rect 11176 3789 11196 3809
rect 13992 3869 14012 3889
rect 13825 3819 13845 3839
rect 14047 3817 14067 3837
rect 11534 3736 11558 3758
rect 14585 3727 14609 3749
rect 12076 3648 12096 3668
rect 12298 3646 12318 3666
rect 12131 3596 12151 3616
rect 14947 3676 14967 3696
rect 12671 3595 12691 3615
rect 11279 3420 11299 3440
rect 11492 3422 11513 3441
rect 11334 3368 11354 3388
rect 12055 3409 12075 3429
rect 11874 3367 11894 3387
rect 11258 3181 11278 3201
rect 12077 3236 12097 3256
rect 12290 3238 12310 3258
rect 14331 3490 14351 3510
rect 14050 3450 14070 3470
rect 14871 3489 14891 3509
rect 14714 3437 14735 3456
rect 14926 3437 14946 3457
rect 13434 3264 13454 3284
rect 13974 3263 13994 3283
rect 12132 3184 12152 3204
rect 12672 3183 12692 3203
rect 11114 3012 11134 3032
rect 11327 3015 11345 3033
rect 11169 2960 11189 2980
rect 12056 2997 12076 3017
rect 11709 2959 11729 2979
rect 13816 3209 13836 3229
rect 14029 3211 14049 3231
rect 14848 3266 14868 3286
rect 14232 3080 14252 3100
rect 14051 3038 14071 3058
rect 14772 3079 14792 3099
rect 14616 3024 14635 3042
rect 14827 3027 14847 3047
rect 11093 2773 11113 2793
rect 13435 2852 13455 2872
rect 13975 2851 13995 2871
rect 13808 2801 13828 2821
rect 14030 2799 14050 2819
rect 11514 2718 11538 2740
rect 11119 2470 11140 2489
rect 10818 2341 10842 2363
rect 9050 2233 9070 2253
rect 9590 2232 9610 2252
rect 7735 2154 7755 2174
rect 8275 2153 8295 2173
rect 4674 1809 4694 1829
rect 2398 1728 2418 1748
rect 5214 1808 5234 1828
rect 5047 1758 5067 1778
rect 5269 1756 5289 1776
rect 1443 1653 1467 1675
rect 2756 1675 2780 1697
rect 1805 1602 1825 1622
rect 1189 1416 1209 1436
rect 908 1376 928 1396
rect 1729 1415 1749 1435
rect 1574 1359 1593 1376
rect 1784 1363 1804 1383
rect 6783 1980 6803 2000
rect 6994 1981 7015 2000
rect 6838 1928 6858 1948
rect 7659 1967 7679 1987
rect 7378 1927 7398 1947
rect 9432 2178 9452 2198
rect 9645 2180 9665 2200
rect 10464 2235 10484 2255
rect 10621 2149 10643 2167
rect 9848 2049 9868 2069
rect 9667 2007 9687 2027
rect 10388 2048 10408 2068
rect 10229 1995 10250 2014
rect 10443 1996 10463 2016
rect 14966 2960 14987 2979
rect 14568 2709 14592 2731
rect 12056 2630 12076 2650
rect 12278 2628 12298 2648
rect 12111 2578 12131 2598
rect 12651 2577 12671 2597
rect 14993 2656 15013 2676
rect 11259 2402 11279 2422
rect 11471 2407 11490 2425
rect 11314 2350 11334 2370
rect 12035 2391 12055 2411
rect 11854 2349 11874 2369
rect 11238 2163 11258 2183
rect 12057 2218 12077 2238
rect 12270 2220 12290 2240
rect 14377 2470 14397 2490
rect 14030 2432 14050 2452
rect 14917 2469 14937 2489
rect 14758 2417 14781 2439
rect 14972 2417 14992 2437
rect 16457 4679 16477 4699
rect 16679 4677 16699 4697
rect 16512 4627 16532 4647
rect 17052 4626 17072 4646
rect 15660 4451 15680 4471
rect 15872 4456 15891 4474
rect 15715 4399 15735 4419
rect 16436 4440 16456 4460
rect 16255 4398 16275 4418
rect 15639 4212 15659 4232
rect 15457 4114 15479 4132
rect 16458 4267 16478 4287
rect 16671 4269 16691 4289
rect 16513 4215 16533 4235
rect 17053 4214 17073 4234
rect 15561 4041 15581 4061
rect 15772 4048 15791 4065
rect 15616 3989 15636 4009
rect 16437 4028 16457 4048
rect 16156 3988 16176 4008
rect 15540 3802 15560 3822
rect 15898 3749 15922 3771
rect 16440 3661 16460 3681
rect 16662 3659 16682 3679
rect 16495 3609 16515 3629
rect 17035 3608 17055 3628
rect 15643 3433 15663 3453
rect 15856 3435 15877 3454
rect 15698 3381 15718 3401
rect 16419 3422 16439 3442
rect 16238 3380 16258 3400
rect 15622 3194 15642 3214
rect 16441 3249 16461 3269
rect 16654 3251 16674 3271
rect 16496 3197 16516 3217
rect 17036 3196 17056 3216
rect 15478 3025 15498 3045
rect 15691 3028 15709 3046
rect 15533 2973 15553 2993
rect 16420 3010 16440 3030
rect 16073 2972 16093 2992
rect 15457 2786 15477 2806
rect 15878 2731 15902 2753
rect 15483 2483 15504 2502
rect 15182 2354 15206 2376
rect 13414 2246 13434 2266
rect 13954 2245 13974 2265
rect 12112 2166 12132 2186
rect 12652 2165 12672 2185
rect 9051 1821 9071 1841
rect 6762 1741 6782 1761
rect 9591 1820 9611 1840
rect 9424 1770 9444 1790
rect 9646 1768 9666 1788
rect 5807 1666 5831 1688
rect 7120 1688 7144 1710
rect 3298 1587 3318 1607
rect 3520 1585 3540 1605
rect 3353 1535 3373 1555
rect 6169 1615 6189 1635
rect 3893 1534 3913 1554
rect 292 1190 312 1210
rect 832 1189 852 1209
rect 674 1135 694 1155
rect 887 1137 907 1157
rect 1706 1192 1726 1212
rect 1090 1006 1110 1026
rect 909 964 929 984
rect 1630 1005 1650 1025
rect 1474 950 1493 968
rect 1685 953 1705 973
rect 293 778 313 798
rect 833 777 853 797
rect 666 727 686 747
rect 888 725 908 745
rect 2501 1359 2521 1379
rect 2714 1361 2735 1380
rect 2556 1307 2576 1327
rect 3277 1348 3297 1368
rect 3096 1306 3116 1326
rect 2480 1120 2500 1140
rect 3299 1175 3319 1195
rect 3512 1177 3532 1197
rect 5553 1429 5573 1449
rect 5272 1389 5292 1409
rect 6093 1428 6113 1448
rect 5938 1372 5957 1389
rect 6148 1376 6168 1396
rect 11160 1992 11180 2012
rect 11371 1993 11392 2012
rect 11215 1940 11235 1960
rect 12036 1979 12056 1999
rect 11755 1939 11775 1959
rect 13796 2191 13816 2211
rect 14009 2193 14029 2213
rect 14828 2248 14848 2268
rect 14985 2162 15007 2180
rect 14212 2062 14232 2082
rect 14031 2020 14051 2040
rect 14752 2061 14772 2081
rect 14593 2008 14614 2027
rect 14807 2009 14827 2029
rect 16420 2643 16440 2663
rect 16642 2641 16662 2661
rect 16475 2591 16495 2611
rect 17015 2590 17035 2610
rect 15623 2415 15643 2435
rect 15835 2420 15854 2438
rect 15678 2363 15698 2383
rect 16399 2404 16419 2424
rect 16218 2362 16238 2382
rect 15602 2176 15622 2196
rect 16421 2231 16441 2251
rect 16634 2233 16654 2253
rect 16476 2179 16496 2199
rect 17016 2178 17036 2198
rect 13415 1834 13435 1854
rect 11139 1753 11159 1773
rect 13955 1833 13975 1853
rect 13788 1783 13808 1803
rect 14010 1781 14030 1801
rect 10184 1678 10208 1700
rect 11497 1700 11521 1722
rect 7662 1600 7682 1620
rect 7884 1598 7904 1618
rect 7717 1548 7737 1568
rect 10546 1627 10566 1647
rect 8257 1547 8277 1567
rect 4656 1203 4676 1223
rect 5196 1202 5216 1222
rect 3354 1123 3374 1143
rect 3894 1122 3914 1142
rect 3278 936 3298 956
rect 1824 886 1845 905
rect 5038 1148 5058 1168
rect 5251 1150 5271 1170
rect 6070 1205 6090 1225
rect 5454 1019 5474 1039
rect 5273 977 5293 997
rect 5994 1018 6014 1038
rect 5838 963 5857 981
rect 6049 966 6069 986
rect 4657 791 4677 811
rect 5197 790 5217 810
rect 5030 740 5050 760
rect 5252 738 5272 758
rect 4047 673 4079 698
rect 1426 635 1450 657
rect 6865 1372 6885 1392
rect 7078 1374 7099 1393
rect 6920 1320 6940 1340
rect 7641 1361 7661 1381
rect 7460 1319 7480 1339
rect 6844 1133 6864 1153
rect 7663 1188 7683 1208
rect 7876 1190 7896 1210
rect 9930 1441 9950 1461
rect 9649 1401 9669 1421
rect 10470 1440 10490 1460
rect 10315 1384 10334 1401
rect 10525 1388 10545 1408
rect 15524 2005 15544 2025
rect 15735 2006 15756 2025
rect 15579 1953 15599 1973
rect 16400 1992 16420 2012
rect 16119 1952 16139 1972
rect 15503 1766 15523 1786
rect 14548 1691 14572 1713
rect 15861 1713 15885 1735
rect 12039 1612 12059 1632
rect 12261 1610 12281 1630
rect 12094 1560 12114 1580
rect 14910 1640 14930 1660
rect 12634 1559 12654 1579
rect 9033 1215 9053 1235
rect 9573 1214 9593 1234
rect 7718 1136 7738 1156
rect 8258 1135 8278 1155
rect 7642 949 7662 969
rect 6188 899 6209 918
rect 9415 1160 9435 1180
rect 9628 1162 9648 1182
rect 10447 1217 10467 1237
rect 9831 1031 9851 1051
rect 9650 989 9670 1009
rect 10371 1030 10391 1050
rect 10215 975 10234 993
rect 10426 978 10446 998
rect 9034 803 9054 823
rect 9574 802 9594 822
rect 9407 752 9427 772
rect 9629 750 9649 770
rect 8411 686 8443 711
rect 5790 648 5814 670
rect 11242 1384 11262 1404
rect 11455 1386 11476 1405
rect 11297 1332 11317 1352
rect 12018 1373 12038 1393
rect 11837 1331 11857 1351
rect 11221 1145 11241 1165
rect 12040 1200 12060 1220
rect 12253 1202 12273 1222
rect 14294 1454 14314 1474
rect 14013 1414 14033 1434
rect 14834 1453 14854 1473
rect 14679 1397 14698 1414
rect 14889 1401 14909 1421
rect 16403 1625 16423 1645
rect 16625 1623 16645 1643
rect 16458 1573 16478 1593
rect 16998 1572 17018 1592
rect 13397 1228 13417 1248
rect 13937 1227 13957 1247
rect 12095 1148 12115 1168
rect 12635 1147 12655 1167
rect 12019 961 12039 981
rect 10565 911 10586 930
rect 13779 1173 13799 1193
rect 13992 1175 14012 1195
rect 14811 1230 14831 1250
rect 14195 1044 14215 1064
rect 14014 1002 14034 1022
rect 14735 1043 14755 1063
rect 14579 988 14598 1006
rect 14790 991 14810 1011
rect 13398 816 13418 836
rect 13938 815 13958 835
rect 13771 765 13791 785
rect 13993 763 14013 783
rect 12788 698 12820 723
rect 10167 660 10191 682
rect 15606 1397 15626 1417
rect 15819 1399 15840 1418
rect 15661 1345 15681 1365
rect 16382 1386 16402 1406
rect 16201 1344 16221 1364
rect 15585 1158 15605 1178
rect 16404 1213 16424 1233
rect 16617 1215 16637 1235
rect 16459 1161 16479 1181
rect 16999 1160 17019 1180
rect 16383 974 16403 994
rect 14929 924 14950 943
rect 17152 711 17184 736
rect 14531 673 14555 695
rect 506 583 542 610
rect 4870 596 4906 623
rect 9247 608 9283 635
rect 13611 621 13647 648
rect 2122 387 2143 408
rect 6486 400 6507 421
rect 10863 412 10884 433
rect 15227 425 15248 446
rect 2204 294 2224 314
rect 4611 313 4632 334
rect 1506 202 1526 222
rect 2046 201 2066 221
rect 1888 144 1911 168
rect 2101 149 2121 169
rect 6568 307 6588 327
rect 9059 337 9080 358
rect 4693 220 4713 240
rect 5870 215 5890 235
rect 3995 128 4015 148
rect 4535 127 4555 147
rect 4380 69 4397 90
rect 4590 75 4610 95
rect 6410 214 6430 234
rect 6255 158 6278 182
rect 6465 162 6485 182
rect 9141 244 9161 264
rect 10945 319 10965 339
rect 13352 338 13373 359
rect 8443 152 8463 172
rect 8983 151 9003 171
rect 9038 99 9058 119
rect 10247 227 10267 247
rect 10787 226 10807 246
rect 10629 169 10652 193
rect 10842 174 10862 194
rect 15309 332 15329 352
rect 13434 245 13454 265
rect 14611 240 14631 260
rect 12736 153 12756 173
rect 13276 152 13296 172
rect 13117 96 13138 118
rect 13331 100 13351 120
rect 15151 239 15171 259
rect 14996 183 15019 207
rect 15206 187 15226 207
<< metal1 >>
rect 16492 8869 16778 8870
rect 15977 8861 16780 8869
rect 12128 8856 12414 8857
rect 11613 8848 12416 8856
rect 7751 8844 8037 8845
rect 7236 8836 8039 8844
rect 3387 8831 3673 8832
rect 2872 8823 3675 8831
rect 2872 8806 2883 8823
rect 2873 8801 2883 8806
rect 2907 8806 3675 8823
rect 7236 8819 7247 8836
rect 2907 8801 2912 8806
rect 2873 8788 2912 8801
rect 3417 8740 3452 8741
rect 3396 8733 3452 8740
rect 3396 8713 3425 8733
rect 3445 8713 3452 8733
rect 3396 8708 3452 8713
rect 3636 8731 3675 8806
rect 7237 8814 7247 8819
rect 7271 8819 8039 8836
rect 11613 8831 11624 8848
rect 7271 8814 7276 8819
rect 7237 8801 7276 8814
rect 7781 8753 7816 8754
rect 3636 8711 3647 8731
rect 3667 8711 3675 8731
rect 2480 8572 2862 8577
rect 2480 8553 2488 8572
rect 2509 8553 2862 8572
rect 2480 8545 2862 8553
rect 1031 8527 1063 8528
rect 1028 8522 1063 8527
rect 1028 8502 1035 8522
rect 1055 8502 1063 8522
rect 2833 8515 2862 8545
rect 2620 8512 2655 8513
rect 1028 8494 1063 8502
rect 410 8336 995 8344
rect 410 8316 419 8336
rect 439 8335 995 8336
rect 439 8316 959 8335
rect 410 8315 959 8316
rect 979 8315 995 8335
rect 410 8309 995 8315
rect 1029 8288 1063 8494
rect 2599 8505 2655 8512
rect 2599 8485 2628 8505
rect 2648 8485 2655 8505
rect 2599 8480 2655 8485
rect 2832 8508 2866 8515
rect 2832 8490 2840 8508
rect 2859 8490 2866 8508
rect 2832 8482 2866 8490
rect 3396 8502 3430 8708
rect 3636 8707 3675 8711
rect 7760 8746 7816 8753
rect 7760 8726 7789 8746
rect 7809 8726 7816 8746
rect 7760 8721 7816 8726
rect 8000 8744 8039 8819
rect 11614 8826 11624 8831
rect 11648 8831 12416 8848
rect 15977 8844 15988 8861
rect 11648 8826 11653 8831
rect 11614 8813 11653 8826
rect 12158 8765 12193 8766
rect 8000 8724 8011 8744
rect 8031 8724 8039 8744
rect 3464 8681 4049 8687
rect 3464 8661 3480 8681
rect 3500 8680 4049 8681
rect 3500 8661 4020 8680
rect 3464 8660 4020 8661
rect 4040 8660 4049 8680
rect 3464 8652 4049 8660
rect 6844 8585 7226 8590
rect 6844 8566 6852 8585
rect 6873 8566 7226 8585
rect 6844 8558 7226 8566
rect 5395 8540 5427 8541
rect 5392 8535 5427 8540
rect 5392 8515 5399 8535
rect 5419 8515 5427 8535
rect 7197 8528 7226 8558
rect 6984 8525 7019 8526
rect 5392 8507 5427 8515
rect 3396 8494 3431 8502
rect 793 8281 828 8288
rect 793 8261 801 8281
rect 821 8261 828 8281
rect 793 8188 828 8261
rect 1007 8283 1063 8288
rect 1007 8263 1014 8283
rect 1034 8263 1063 8283
rect 1007 8256 1063 8263
rect 1098 8390 1128 8392
rect 1827 8390 1860 8391
rect 1098 8364 1861 8390
rect 1007 8255 1042 8256
rect 1098 8189 1128 8364
rect 1827 8343 1861 8364
rect 1826 8338 1861 8343
rect 1826 8318 1833 8338
rect 1853 8318 1861 8338
rect 1826 8310 1861 8318
rect 1093 8188 1128 8189
rect 792 8161 1128 8188
rect 1098 8160 1128 8161
rect 1208 8152 1793 8160
rect 1208 8132 1217 8152
rect 1237 8151 1793 8152
rect 1237 8132 1757 8151
rect 1208 8131 1757 8132
rect 1777 8131 1793 8151
rect 1208 8125 1793 8131
rect 1032 8115 1064 8116
rect 1029 8110 1064 8115
rect 1029 8090 1036 8110
rect 1056 8090 1064 8110
rect 1827 8104 1861 8310
rect 2599 8274 2633 8480
rect 3396 8474 3404 8494
rect 3424 8474 3431 8494
rect 3396 8469 3431 8474
rect 3396 8468 3428 8469
rect 2667 8453 3252 8459
rect 2667 8433 2683 8453
rect 2703 8452 3252 8453
rect 2703 8433 3223 8452
rect 2667 8432 3223 8433
rect 3243 8432 3252 8452
rect 2667 8424 3252 8432
rect 3332 8423 3362 8424
rect 3332 8396 3668 8423
rect 3332 8395 3367 8396
rect 2599 8266 2634 8274
rect 2599 8246 2607 8266
rect 2627 8246 2634 8266
rect 2599 8241 2634 8246
rect 2599 8220 2633 8241
rect 3332 8220 3362 8395
rect 3418 8328 3453 8329
rect 2599 8194 3362 8220
rect 2600 8193 2633 8194
rect 3332 8192 3362 8194
rect 3397 8321 3453 8328
rect 3397 8301 3426 8321
rect 3446 8301 3453 8321
rect 3397 8296 3453 8301
rect 3632 8323 3667 8396
rect 3632 8303 3639 8323
rect 3659 8303 3667 8323
rect 4774 8349 5359 8357
rect 4774 8329 4783 8349
rect 4803 8348 5359 8349
rect 4803 8329 5323 8348
rect 4774 8328 5323 8329
rect 5343 8328 5359 8348
rect 4774 8322 5359 8328
rect 3632 8296 3667 8303
rect 5393 8301 5427 8507
rect 6963 8518 7019 8525
rect 6963 8498 6992 8518
rect 7012 8498 7019 8518
rect 6963 8493 7019 8498
rect 7196 8521 7230 8528
rect 7196 8503 7204 8521
rect 7223 8503 7230 8521
rect 7196 8495 7230 8503
rect 7760 8515 7794 8721
rect 8000 8720 8039 8724
rect 12137 8758 12193 8765
rect 12137 8738 12166 8758
rect 12186 8738 12193 8758
rect 12137 8733 12193 8738
rect 12377 8756 12416 8831
rect 15978 8839 15988 8844
rect 16012 8844 16780 8861
rect 16012 8839 16017 8844
rect 15978 8826 16017 8839
rect 16522 8778 16557 8779
rect 12377 8736 12388 8756
rect 12408 8736 12416 8756
rect 7828 8694 8413 8700
rect 7828 8674 7844 8694
rect 7864 8693 8413 8694
rect 7864 8674 8384 8693
rect 7828 8673 8384 8674
rect 8404 8673 8413 8693
rect 7828 8665 8413 8673
rect 11221 8597 11603 8602
rect 11221 8578 11229 8597
rect 11250 8578 11603 8597
rect 11221 8570 11603 8578
rect 9772 8552 9804 8553
rect 9769 8547 9804 8552
rect 9769 8527 9776 8547
rect 9796 8527 9804 8547
rect 11574 8540 11603 8570
rect 11361 8537 11396 8538
rect 9769 8519 9804 8527
rect 7760 8507 7795 8515
rect 1029 8082 1064 8090
rect 411 7924 996 7932
rect 411 7904 420 7924
rect 440 7923 996 7924
rect 440 7904 960 7923
rect 411 7903 960 7904
rect 980 7903 996 7923
rect 411 7897 996 7903
rect 785 7873 824 7877
rect 1030 7876 1064 8082
rect 1593 8097 1628 8103
rect 1593 8078 1598 8097
rect 1619 8078 1628 8097
rect 1593 8069 1628 8078
rect 1805 8099 1861 8104
rect 1805 8079 1812 8099
rect 1832 8079 1861 8099
rect 1805 8072 1861 8079
rect 2428 8143 2762 8171
rect 1805 8071 1840 8072
rect 1597 8001 1626 8069
rect 1597 7967 1943 8001
rect 785 7853 793 7873
rect 813 7853 824 7873
rect 785 7778 824 7853
rect 1008 7871 1064 7876
rect 1008 7851 1015 7871
rect 1035 7851 1064 7871
rect 1008 7844 1064 7851
rect 1008 7843 1043 7844
rect 1548 7783 1587 7796
rect 1548 7778 1553 7783
rect 785 7761 1553 7778
rect 1577 7778 1587 7783
rect 1577 7761 1588 7778
rect 785 7753 1588 7761
rect 787 7752 1073 7753
rect 1904 7730 1943 7967
rect 1904 7718 1915 7730
rect 1908 7710 1915 7718
rect 1935 7710 1943 7730
rect 1908 7702 1943 7710
rect 1290 7544 1875 7552
rect 1290 7524 1299 7544
rect 1319 7543 1875 7544
rect 1319 7524 1839 7543
rect 1290 7523 1839 7524
rect 1859 7523 1875 7543
rect 1290 7517 1875 7523
rect 1014 7509 1046 7510
rect 1011 7504 1046 7509
rect 1011 7484 1018 7504
rect 1038 7484 1046 7504
rect 1909 7496 1943 7702
rect 1011 7476 1046 7484
rect 393 7318 978 7326
rect 393 7298 402 7318
rect 422 7317 978 7318
rect 422 7298 942 7317
rect 393 7297 942 7298
rect 962 7297 978 7317
rect 393 7291 978 7297
rect 1012 7270 1046 7476
rect 1677 7490 1708 7496
rect 1677 7471 1682 7490
rect 1703 7471 1708 7490
rect 1677 7429 1708 7471
rect 1887 7491 1943 7496
rect 1887 7471 1894 7491
rect 1914 7471 1943 7491
rect 1887 7464 1943 7471
rect 1887 7463 1922 7464
rect 1677 7401 2016 7429
rect 776 7263 811 7270
rect 776 7243 784 7263
rect 804 7243 811 7263
rect 776 7170 811 7243
rect 990 7265 1046 7270
rect 990 7245 997 7265
rect 1017 7245 1046 7265
rect 990 7238 1046 7245
rect 1081 7372 1111 7374
rect 1810 7372 1843 7373
rect 1081 7346 1844 7372
rect 990 7237 1025 7238
rect 1081 7171 1111 7346
rect 1810 7325 1844 7346
rect 1809 7320 1844 7325
rect 1809 7300 1816 7320
rect 1836 7300 1844 7320
rect 1809 7292 1844 7300
rect 1076 7170 1111 7171
rect 775 7143 1111 7170
rect 1081 7142 1111 7143
rect 1191 7134 1776 7142
rect 1191 7114 1200 7134
rect 1220 7133 1776 7134
rect 1220 7114 1740 7133
rect 1191 7113 1740 7114
rect 1760 7113 1776 7133
rect 1191 7107 1776 7113
rect 1015 7097 1047 7098
rect 1012 7092 1047 7097
rect 1012 7072 1019 7092
rect 1039 7072 1047 7092
rect 1810 7086 1844 7292
rect 1012 7064 1047 7072
rect 394 6906 979 6914
rect 394 6886 403 6906
rect 423 6905 979 6906
rect 423 6886 943 6905
rect 394 6885 943 6886
rect 963 6885 979 6905
rect 394 6879 979 6885
rect 768 6855 807 6859
rect 1013 6858 1047 7064
rect 1577 7076 1611 7084
rect 1577 7058 1584 7076
rect 1603 7058 1611 7076
rect 1577 7051 1611 7058
rect 1788 7081 1844 7086
rect 1788 7061 1795 7081
rect 1815 7061 1844 7081
rect 1788 7054 1844 7061
rect 1788 7053 1823 7054
rect 1581 7021 1610 7051
rect 1581 7013 1963 7021
rect 1581 6994 1934 7013
rect 1955 6994 1963 7013
rect 1581 6989 1963 6994
rect 768 6835 776 6855
rect 796 6835 807 6855
rect 768 6760 807 6835
rect 991 6853 1047 6858
rect 991 6833 998 6853
rect 1018 6833 1047 6853
rect 991 6826 1047 6833
rect 991 6825 1026 6826
rect 1531 6765 1570 6778
rect 1531 6760 1536 6765
rect 768 6743 1536 6760
rect 1560 6760 1570 6765
rect 1560 6743 1571 6760
rect 768 6735 1571 6743
rect 770 6734 1056 6735
rect 1987 6716 2016 7401
rect 2428 7334 2460 8143
rect 2736 8108 2762 8143
rect 2521 8102 2556 8103
rect 2500 8095 2556 8102
rect 2500 8075 2529 8095
rect 2549 8075 2556 8095
rect 2500 8070 2556 8075
rect 2732 8099 2768 8108
rect 2732 8082 2740 8099
rect 2759 8082 2768 8099
rect 2732 8073 2768 8082
rect 3397 8090 3431 8296
rect 5157 8294 5192 8301
rect 3465 8269 4050 8275
rect 3465 8249 3481 8269
rect 3501 8268 4050 8269
rect 3501 8249 4021 8268
rect 3465 8248 4021 8249
rect 4041 8248 4050 8268
rect 3465 8240 4050 8248
rect 5157 8274 5165 8294
rect 5185 8274 5192 8294
rect 5157 8201 5192 8274
rect 5371 8296 5427 8301
rect 5371 8276 5378 8296
rect 5398 8276 5427 8296
rect 5371 8269 5427 8276
rect 5462 8403 5492 8405
rect 6191 8403 6224 8404
rect 5462 8377 6225 8403
rect 5371 8268 5406 8269
rect 5462 8202 5492 8377
rect 6191 8356 6225 8377
rect 6190 8351 6225 8356
rect 6190 8331 6197 8351
rect 6217 8331 6225 8351
rect 6190 8323 6225 8331
rect 5457 8201 5492 8202
rect 5156 8174 5492 8201
rect 5462 8173 5492 8174
rect 5572 8165 6157 8173
rect 5572 8145 5581 8165
rect 5601 8164 6157 8165
rect 5601 8145 6121 8164
rect 5572 8144 6121 8145
rect 6141 8144 6157 8164
rect 5572 8138 6157 8144
rect 5396 8128 5428 8129
rect 5393 8123 5428 8128
rect 5393 8103 5400 8123
rect 5420 8103 5428 8123
rect 6191 8117 6225 8323
rect 6963 8287 6997 8493
rect 7760 8487 7768 8507
rect 7788 8487 7795 8507
rect 7760 8482 7795 8487
rect 7760 8481 7792 8482
rect 7031 8466 7616 8472
rect 7031 8446 7047 8466
rect 7067 8465 7616 8466
rect 7067 8446 7587 8465
rect 7031 8445 7587 8446
rect 7607 8445 7616 8465
rect 7031 8437 7616 8445
rect 7696 8436 7726 8437
rect 7696 8409 8032 8436
rect 7696 8408 7731 8409
rect 6963 8279 6998 8287
rect 6963 8259 6971 8279
rect 6991 8259 6998 8279
rect 6963 8254 6998 8259
rect 6963 8233 6997 8254
rect 7696 8233 7726 8408
rect 7782 8341 7817 8342
rect 6963 8207 7726 8233
rect 6964 8206 6997 8207
rect 7696 8205 7726 8207
rect 7761 8334 7817 8341
rect 7761 8314 7790 8334
rect 7810 8314 7817 8334
rect 7761 8309 7817 8314
rect 7996 8336 8031 8409
rect 7996 8316 8003 8336
rect 8023 8316 8031 8336
rect 9151 8361 9736 8369
rect 9151 8341 9160 8361
rect 9180 8360 9736 8361
rect 9180 8341 9700 8360
rect 9151 8340 9700 8341
rect 9720 8340 9736 8360
rect 9151 8334 9736 8340
rect 7996 8309 8031 8316
rect 9770 8313 9804 8519
rect 11340 8530 11396 8537
rect 11340 8510 11369 8530
rect 11389 8510 11396 8530
rect 11340 8505 11396 8510
rect 11573 8533 11607 8540
rect 11573 8515 11581 8533
rect 11600 8515 11607 8533
rect 11573 8507 11607 8515
rect 12137 8527 12171 8733
rect 12377 8732 12416 8736
rect 16501 8771 16557 8778
rect 16501 8751 16530 8771
rect 16550 8751 16557 8771
rect 16501 8746 16557 8751
rect 16741 8769 16780 8844
rect 16741 8749 16752 8769
rect 16772 8749 16780 8769
rect 12205 8706 12790 8712
rect 12205 8686 12221 8706
rect 12241 8705 12790 8706
rect 12241 8686 12761 8705
rect 12205 8685 12761 8686
rect 12781 8685 12790 8705
rect 12205 8677 12790 8685
rect 15585 8610 15967 8615
rect 15585 8591 15593 8610
rect 15614 8591 15967 8610
rect 15585 8583 15967 8591
rect 14136 8565 14168 8566
rect 14133 8560 14168 8565
rect 14133 8540 14140 8560
rect 14160 8540 14168 8560
rect 15938 8553 15967 8583
rect 15725 8550 15760 8551
rect 14133 8532 14168 8540
rect 12137 8519 12172 8527
rect 5393 8095 5428 8103
rect 3397 8082 3432 8090
rect 2500 7864 2534 8070
rect 3397 8062 3405 8082
rect 3425 8062 3432 8082
rect 3397 8057 3432 8062
rect 3397 8056 3429 8057
rect 2568 8043 3153 8049
rect 2568 8023 2584 8043
rect 2604 8042 3153 8043
rect 2604 8023 3124 8042
rect 2568 8022 3124 8023
rect 3144 8022 3153 8042
rect 2568 8014 3153 8022
rect 4775 7937 5360 7945
rect 4775 7917 4784 7937
rect 4804 7936 5360 7937
rect 4804 7917 5324 7936
rect 4775 7916 5324 7917
rect 5344 7916 5360 7936
rect 4775 7910 5360 7916
rect 5149 7886 5188 7890
rect 5394 7889 5428 8095
rect 5957 8110 5992 8116
rect 5957 8091 5962 8110
rect 5983 8091 5992 8110
rect 5957 8082 5992 8091
rect 6169 8112 6225 8117
rect 6169 8092 6176 8112
rect 6196 8092 6225 8112
rect 6169 8085 6225 8092
rect 6792 8156 7126 8184
rect 6169 8084 6204 8085
rect 5961 8014 5990 8082
rect 5961 7980 6307 8014
rect 5149 7866 5157 7886
rect 5177 7866 5188 7886
rect 2500 7856 2535 7864
rect 2500 7836 2508 7856
rect 2528 7848 2535 7856
rect 2528 7836 2539 7848
rect 2500 7599 2539 7836
rect 3370 7813 3656 7814
rect 2855 7805 3658 7813
rect 2855 7788 2866 7805
rect 2856 7783 2866 7788
rect 2890 7788 3658 7805
rect 2890 7783 2895 7788
rect 2856 7770 2895 7783
rect 3400 7722 3435 7723
rect 3379 7715 3435 7722
rect 3379 7695 3408 7715
rect 3428 7695 3435 7715
rect 3379 7690 3435 7695
rect 3619 7713 3658 7788
rect 5149 7791 5188 7866
rect 5372 7884 5428 7889
rect 5372 7864 5379 7884
rect 5399 7864 5428 7884
rect 5372 7857 5428 7864
rect 5372 7856 5407 7857
rect 5912 7796 5951 7809
rect 5912 7791 5917 7796
rect 5149 7774 5917 7791
rect 5941 7791 5951 7796
rect 5941 7774 5952 7791
rect 5149 7766 5952 7774
rect 5151 7765 5437 7766
rect 6268 7743 6307 7980
rect 6268 7731 6279 7743
rect 6272 7723 6279 7731
rect 6299 7723 6307 7743
rect 6272 7715 6307 7723
rect 3619 7693 3630 7713
rect 3650 7693 3658 7713
rect 2500 7565 2846 7599
rect 2817 7497 2846 7565
rect 2603 7494 2638 7495
rect 2428 7316 2431 7334
rect 2453 7316 2460 7334
rect 2428 7304 2460 7316
rect 2582 7487 2638 7494
rect 2582 7467 2611 7487
rect 2631 7467 2638 7487
rect 2582 7462 2638 7467
rect 2815 7488 2850 7497
rect 2815 7469 2824 7488
rect 2845 7469 2850 7488
rect 2815 7463 2850 7469
rect 3379 7484 3413 7690
rect 3619 7689 3658 7693
rect 3447 7663 4032 7669
rect 3447 7643 3463 7663
rect 3483 7662 4032 7663
rect 3483 7643 4003 7662
rect 3447 7642 4003 7643
rect 4023 7642 4032 7662
rect 3447 7634 4032 7642
rect 5654 7557 6239 7565
rect 5654 7537 5663 7557
rect 5683 7556 6239 7557
rect 5683 7537 6203 7556
rect 5654 7536 6203 7537
rect 6223 7536 6239 7556
rect 5654 7530 6239 7536
rect 5378 7522 5410 7523
rect 5375 7517 5410 7522
rect 5375 7497 5382 7517
rect 5402 7497 5410 7517
rect 6273 7509 6307 7715
rect 5375 7489 5410 7497
rect 3379 7476 3414 7484
rect 2582 7256 2616 7462
rect 3379 7456 3387 7476
rect 3407 7456 3414 7476
rect 3379 7451 3414 7456
rect 3379 7450 3411 7451
rect 2650 7435 3235 7441
rect 2650 7415 2666 7435
rect 2686 7434 3235 7435
rect 2686 7415 3206 7434
rect 2650 7414 3206 7415
rect 3226 7414 3235 7434
rect 2650 7406 3235 7414
rect 3315 7405 3345 7406
rect 3315 7378 3651 7405
rect 3315 7377 3350 7378
rect 2582 7248 2617 7256
rect 2582 7228 2590 7248
rect 2610 7228 2617 7248
rect 2582 7223 2617 7228
rect 2582 7202 2616 7223
rect 3315 7202 3345 7377
rect 3401 7310 3436 7311
rect 2582 7176 3345 7202
rect 2583 7175 2616 7176
rect 3315 7174 3345 7176
rect 3380 7303 3436 7310
rect 3380 7283 3409 7303
rect 3429 7283 3436 7303
rect 3380 7278 3436 7283
rect 3615 7305 3650 7378
rect 3615 7285 3622 7305
rect 3642 7285 3650 7305
rect 4757 7331 5342 7339
rect 4757 7311 4766 7331
rect 4786 7330 5342 7331
rect 4786 7311 5306 7330
rect 4757 7310 5306 7311
rect 5326 7310 5342 7330
rect 4757 7304 5342 7310
rect 3615 7278 3650 7285
rect 5376 7283 5410 7489
rect 6041 7503 6072 7509
rect 6041 7484 6046 7503
rect 6067 7484 6072 7503
rect 6041 7442 6072 7484
rect 6251 7504 6307 7509
rect 6251 7484 6258 7504
rect 6278 7484 6307 7504
rect 6251 7477 6307 7484
rect 6251 7476 6286 7477
rect 6041 7414 6380 7442
rect 2220 7142 2683 7150
rect 2220 7120 2232 7142
rect 2256 7120 2683 7142
rect 2220 7119 2683 7120
rect 2222 7107 2261 7119
rect 2656 7088 2683 7119
rect 2438 7086 2473 7087
rect 2417 7079 2473 7086
rect 2417 7059 2446 7079
rect 2466 7059 2473 7079
rect 2417 7054 2473 7059
rect 2652 7079 2685 7088
rect 2652 7057 2657 7079
rect 2680 7057 2685 7079
rect 2417 6848 2451 7054
rect 2652 7051 2685 7057
rect 3380 7072 3414 7278
rect 5140 7276 5175 7283
rect 3448 7251 4033 7257
rect 3448 7231 3464 7251
rect 3484 7250 4033 7251
rect 3484 7231 4004 7250
rect 3448 7230 4004 7231
rect 4024 7230 4033 7250
rect 3448 7222 4033 7230
rect 5140 7256 5148 7276
rect 5168 7256 5175 7276
rect 5140 7183 5175 7256
rect 5354 7278 5410 7283
rect 5354 7258 5361 7278
rect 5381 7258 5410 7278
rect 5354 7251 5410 7258
rect 5445 7385 5475 7387
rect 6174 7385 6207 7386
rect 5445 7359 6208 7385
rect 5354 7250 5389 7251
rect 5445 7184 5475 7359
rect 6174 7338 6208 7359
rect 6173 7333 6208 7338
rect 6173 7313 6180 7333
rect 6200 7313 6208 7333
rect 6173 7305 6208 7313
rect 5440 7183 5475 7184
rect 5139 7156 5475 7183
rect 5445 7155 5475 7156
rect 5555 7147 6140 7155
rect 5555 7127 5564 7147
rect 5584 7146 6140 7147
rect 5584 7127 6104 7146
rect 5555 7126 6104 7127
rect 6124 7126 6140 7146
rect 5555 7120 6140 7126
rect 5379 7110 5411 7111
rect 5376 7105 5411 7110
rect 5376 7085 5383 7105
rect 5403 7085 5411 7105
rect 6174 7099 6208 7305
rect 5376 7077 5411 7085
rect 3380 7064 3415 7072
rect 3380 7044 3388 7064
rect 3408 7044 3415 7064
rect 3380 7039 3415 7044
rect 3380 7038 3412 7039
rect 2485 7027 3070 7033
rect 2485 7007 2501 7027
rect 2521 7026 3070 7027
rect 2521 7007 3041 7026
rect 2485 7006 3041 7007
rect 3061 7006 3070 7026
rect 2485 6998 3070 7006
rect 4758 6919 5343 6927
rect 4758 6899 4767 6919
rect 4787 6918 5343 6919
rect 4787 6899 5307 6918
rect 4758 6898 5307 6899
rect 5327 6898 5343 6918
rect 4758 6892 5343 6898
rect 5132 6868 5171 6872
rect 5377 6871 5411 7077
rect 5941 7089 5975 7097
rect 5941 7071 5948 7089
rect 5967 7071 5975 7089
rect 5941 7064 5975 7071
rect 6152 7094 6208 7099
rect 6152 7074 6159 7094
rect 6179 7074 6208 7094
rect 6152 7067 6208 7074
rect 6152 7066 6187 7067
rect 5945 7034 5974 7064
rect 5945 7026 6327 7034
rect 5945 7007 6298 7026
rect 6319 7007 6327 7026
rect 5945 7002 6327 7007
rect 5132 6848 5140 6868
rect 5160 6848 5171 6868
rect 2417 6847 2452 6848
rect 2385 6840 2452 6847
rect 2385 6820 2425 6840
rect 2445 6820 2452 6840
rect 2385 6817 2452 6820
rect 2385 6814 2450 6817
rect 1956 6713 2021 6716
rect 1954 6710 2021 6713
rect 1954 6690 1961 6710
rect 1981 6690 2021 6710
rect 1954 6683 2021 6690
rect 1954 6682 1989 6683
rect 1336 6524 1921 6532
rect 1336 6504 1345 6524
rect 1365 6523 1921 6524
rect 1365 6504 1885 6523
rect 1336 6503 1885 6504
rect 1905 6503 1921 6523
rect 1336 6497 1921 6503
rect 994 6491 1026 6492
rect 991 6486 1026 6491
rect 991 6466 998 6486
rect 1018 6466 1026 6486
rect 991 6458 1026 6466
rect 373 6300 958 6308
rect 373 6280 382 6300
rect 402 6299 958 6300
rect 402 6280 922 6299
rect 373 6279 922 6280
rect 942 6279 958 6299
rect 373 6273 958 6279
rect 992 6252 1026 6458
rect 1719 6468 1760 6479
rect 1955 6476 1989 6682
rect 1719 6450 1729 6468
rect 1747 6450 1760 6468
rect 1719 6442 1760 6450
rect 1933 6471 1989 6476
rect 1933 6451 1940 6471
rect 1960 6451 1989 6471
rect 1933 6444 1989 6451
rect 1933 6443 1968 6444
rect 1728 6412 1754 6442
rect 1728 6411 2066 6412
rect 1728 6375 2082 6411
rect 756 6245 791 6252
rect 756 6225 764 6245
rect 784 6225 791 6245
rect 756 6152 791 6225
rect 970 6247 1026 6252
rect 970 6227 977 6247
rect 997 6227 1026 6247
rect 970 6220 1026 6227
rect 1061 6354 1091 6356
rect 1790 6354 1823 6355
rect 1061 6328 1824 6354
rect 970 6219 1005 6220
rect 1061 6153 1091 6328
rect 1790 6307 1824 6328
rect 1789 6302 1824 6307
rect 1789 6282 1796 6302
rect 1816 6282 1824 6302
rect 1789 6274 1824 6282
rect 1056 6152 1091 6153
rect 755 6125 1091 6152
rect 1061 6124 1091 6125
rect 1171 6116 1756 6124
rect 1171 6096 1180 6116
rect 1200 6115 1756 6116
rect 1200 6096 1720 6115
rect 1171 6095 1720 6096
rect 1740 6095 1756 6115
rect 1171 6089 1756 6095
rect 995 6079 1027 6080
rect 992 6074 1027 6079
rect 992 6054 999 6074
rect 1019 6054 1027 6074
rect 1790 6068 1824 6274
rect 992 6046 1027 6054
rect 374 5888 959 5896
rect 374 5868 383 5888
rect 403 5887 959 5888
rect 403 5868 923 5887
rect 374 5867 923 5868
rect 943 5867 959 5887
rect 374 5861 959 5867
rect 748 5837 787 5841
rect 993 5840 1027 6046
rect 1556 6061 1591 6067
rect 1556 6042 1561 6061
rect 1582 6042 1591 6061
rect 1556 6033 1591 6042
rect 1768 6063 1824 6068
rect 1768 6043 1775 6063
rect 1795 6043 1824 6063
rect 1768 6036 1824 6043
rect 1768 6035 1803 6036
rect 1560 5965 1589 6033
rect 1560 5931 1906 5965
rect 748 5817 756 5837
rect 776 5817 787 5837
rect 748 5742 787 5817
rect 971 5835 1027 5840
rect 971 5815 978 5835
rect 998 5815 1027 5835
rect 971 5808 1027 5815
rect 971 5807 1006 5808
rect 1511 5747 1550 5760
rect 1511 5742 1516 5747
rect 748 5725 1516 5742
rect 1540 5742 1550 5747
rect 1540 5725 1551 5742
rect 748 5717 1551 5725
rect 750 5716 1036 5717
rect 1867 5694 1906 5931
rect 1867 5682 1878 5694
rect 1871 5674 1878 5682
rect 1898 5674 1906 5694
rect 1871 5666 1906 5674
rect 1253 5508 1838 5516
rect 1253 5488 1262 5508
rect 1282 5507 1838 5508
rect 1282 5488 1802 5507
rect 1253 5487 1802 5488
rect 1822 5487 1838 5507
rect 1253 5481 1838 5487
rect 977 5473 1009 5474
rect 974 5468 1009 5473
rect 974 5448 981 5468
rect 1001 5448 1009 5468
rect 1872 5460 1906 5666
rect 974 5440 1009 5448
rect 356 5282 941 5290
rect 356 5262 365 5282
rect 385 5281 941 5282
rect 385 5262 905 5281
rect 356 5261 905 5262
rect 925 5261 941 5281
rect 356 5255 941 5261
rect 975 5234 1009 5440
rect 1638 5448 1674 5457
rect 1638 5431 1647 5448
rect 1666 5431 1674 5448
rect 1638 5422 1674 5431
rect 1850 5455 1906 5460
rect 1850 5435 1857 5455
rect 1877 5435 1906 5455
rect 1850 5428 1906 5435
rect 1850 5427 1885 5428
rect 1644 5387 1670 5422
rect 1952 5387 1984 5388
rect 1644 5382 1984 5387
rect 1644 5364 1959 5382
rect 1981 5364 1984 5382
rect 1644 5359 1984 5364
rect 1952 5358 1984 5359
rect 739 5227 774 5234
rect 739 5207 747 5227
rect 767 5207 774 5227
rect 739 5134 774 5207
rect 953 5229 1009 5234
rect 953 5209 960 5229
rect 980 5209 1009 5229
rect 953 5202 1009 5209
rect 1044 5336 1074 5338
rect 1773 5336 1806 5337
rect 1044 5310 1807 5336
rect 953 5201 988 5202
rect 1044 5135 1074 5310
rect 1773 5289 1807 5310
rect 1772 5284 1807 5289
rect 1772 5264 1779 5284
rect 1799 5264 1807 5284
rect 1772 5256 1807 5264
rect 1039 5134 1074 5135
rect 738 5107 1074 5134
rect 1044 5106 1074 5107
rect 1154 5098 1739 5106
rect 1154 5078 1163 5098
rect 1183 5097 1739 5098
rect 1183 5078 1703 5097
rect 1154 5077 1703 5078
rect 1723 5077 1739 5097
rect 1154 5071 1739 5077
rect 978 5061 1010 5062
rect 975 5056 1010 5061
rect 975 5036 982 5056
rect 1002 5036 1010 5056
rect 1773 5050 1807 5256
rect 975 5028 1010 5036
rect 357 4870 942 4878
rect 357 4850 366 4870
rect 386 4869 942 4870
rect 386 4850 906 4869
rect 357 4849 906 4850
rect 926 4849 942 4869
rect 357 4843 942 4849
rect 731 4819 770 4823
rect 976 4822 1010 5028
rect 1540 5040 1574 5048
rect 1540 5022 1547 5040
rect 1566 5022 1574 5040
rect 1540 5015 1574 5022
rect 1751 5045 1807 5050
rect 1751 5025 1758 5045
rect 1778 5025 1807 5045
rect 1751 5018 1807 5025
rect 1751 5017 1786 5018
rect 1544 4985 1573 5015
rect 1544 4977 1926 4985
rect 1544 4958 1897 4977
rect 1918 4958 1926 4977
rect 1544 4953 1926 4958
rect 731 4799 739 4819
rect 759 4799 770 4819
rect 731 4724 770 4799
rect 954 4817 1010 4822
rect 954 4797 961 4817
rect 981 4797 1010 4817
rect 954 4790 1010 4797
rect 954 4789 989 4790
rect 1494 4729 1533 4742
rect 1494 4724 1499 4729
rect 731 4707 1499 4724
rect 1523 4724 1533 4729
rect 1523 4707 1534 4724
rect 731 4699 1534 4707
rect 733 4698 1019 4699
rect 2055 4675 2082 6375
rect 2390 6129 2419 6814
rect 3350 6795 3636 6796
rect 2835 6787 3638 6795
rect 2835 6770 2846 6787
rect 2836 6765 2846 6770
rect 2870 6770 3638 6787
rect 2870 6765 2875 6770
rect 2836 6752 2875 6765
rect 3380 6704 3415 6705
rect 3359 6697 3415 6704
rect 3359 6677 3388 6697
rect 3408 6677 3415 6697
rect 3359 6672 3415 6677
rect 3599 6695 3638 6770
rect 5132 6773 5171 6848
rect 5355 6866 5411 6871
rect 5355 6846 5362 6866
rect 5382 6846 5411 6866
rect 5355 6839 5411 6846
rect 5355 6838 5390 6839
rect 5895 6778 5934 6791
rect 5895 6773 5900 6778
rect 5132 6756 5900 6773
rect 5924 6773 5934 6778
rect 5924 6756 5935 6773
rect 5132 6748 5935 6756
rect 5134 6747 5420 6748
rect 6351 6729 6380 7414
rect 6792 7347 6824 8156
rect 7100 8121 7126 8156
rect 6885 8115 6920 8116
rect 6864 8108 6920 8115
rect 6864 8088 6893 8108
rect 6913 8088 6920 8108
rect 6864 8083 6920 8088
rect 7096 8112 7132 8121
rect 7096 8095 7104 8112
rect 7123 8095 7132 8112
rect 7096 8086 7132 8095
rect 7761 8103 7795 8309
rect 9534 8306 9569 8313
rect 7829 8282 8414 8288
rect 7829 8262 7845 8282
rect 7865 8281 8414 8282
rect 7865 8262 8385 8281
rect 7829 8261 8385 8262
rect 8405 8261 8414 8281
rect 7829 8253 8414 8261
rect 9534 8286 9542 8306
rect 9562 8286 9569 8306
rect 9534 8213 9569 8286
rect 9748 8308 9804 8313
rect 9748 8288 9755 8308
rect 9775 8288 9804 8308
rect 9748 8281 9804 8288
rect 9839 8415 9869 8417
rect 10568 8415 10601 8416
rect 9839 8389 10602 8415
rect 9748 8280 9783 8281
rect 9839 8214 9869 8389
rect 10568 8368 10602 8389
rect 10567 8363 10602 8368
rect 10567 8343 10574 8363
rect 10594 8343 10602 8363
rect 10567 8335 10602 8343
rect 9834 8213 9869 8214
rect 9533 8186 9869 8213
rect 9839 8185 9869 8186
rect 9949 8177 10534 8185
rect 9949 8157 9958 8177
rect 9978 8176 10534 8177
rect 9978 8157 10498 8176
rect 9949 8156 10498 8157
rect 10518 8156 10534 8176
rect 9949 8150 10534 8156
rect 9773 8140 9805 8141
rect 9770 8135 9805 8140
rect 9770 8115 9777 8135
rect 9797 8115 9805 8135
rect 10568 8129 10602 8335
rect 11340 8299 11374 8505
rect 12137 8499 12145 8519
rect 12165 8499 12172 8519
rect 12137 8494 12172 8499
rect 12137 8493 12169 8494
rect 11408 8478 11993 8484
rect 11408 8458 11424 8478
rect 11444 8477 11993 8478
rect 11444 8458 11964 8477
rect 11408 8457 11964 8458
rect 11984 8457 11993 8477
rect 11408 8449 11993 8457
rect 12073 8448 12103 8449
rect 12073 8421 12409 8448
rect 12073 8420 12108 8421
rect 11340 8291 11375 8299
rect 11340 8271 11348 8291
rect 11368 8271 11375 8291
rect 11340 8266 11375 8271
rect 11340 8245 11374 8266
rect 12073 8245 12103 8420
rect 12159 8353 12194 8354
rect 11340 8219 12103 8245
rect 11341 8218 11374 8219
rect 12073 8217 12103 8219
rect 12138 8346 12194 8353
rect 12138 8326 12167 8346
rect 12187 8326 12194 8346
rect 12138 8321 12194 8326
rect 12373 8348 12408 8421
rect 12373 8328 12380 8348
rect 12400 8328 12408 8348
rect 13515 8374 14100 8382
rect 13515 8354 13524 8374
rect 13544 8373 14100 8374
rect 13544 8354 14064 8373
rect 13515 8353 14064 8354
rect 14084 8353 14100 8373
rect 13515 8347 14100 8353
rect 12373 8321 12408 8328
rect 14134 8326 14168 8532
rect 15704 8543 15760 8550
rect 15704 8523 15733 8543
rect 15753 8523 15760 8543
rect 15704 8518 15760 8523
rect 15937 8546 15971 8553
rect 15937 8528 15945 8546
rect 15964 8528 15971 8546
rect 15937 8520 15971 8528
rect 16501 8540 16535 8746
rect 16741 8745 16780 8749
rect 16569 8719 17154 8725
rect 16569 8699 16585 8719
rect 16605 8718 17154 8719
rect 16605 8699 17125 8718
rect 16569 8698 17125 8699
rect 17145 8698 17154 8718
rect 16569 8690 17154 8698
rect 16501 8532 16536 8540
rect 9770 8107 9805 8115
rect 7761 8095 7796 8103
rect 6864 7877 6898 8083
rect 7761 8075 7769 8095
rect 7789 8075 7796 8095
rect 7761 8070 7796 8075
rect 7761 8069 7793 8070
rect 6932 8056 7517 8062
rect 6932 8036 6948 8056
rect 6968 8055 7517 8056
rect 6968 8036 7488 8055
rect 6932 8035 7488 8036
rect 7508 8035 7517 8055
rect 6932 8027 7517 8035
rect 9152 7949 9737 7957
rect 9152 7929 9161 7949
rect 9181 7948 9737 7949
rect 9181 7929 9701 7948
rect 9152 7928 9701 7929
rect 9721 7928 9737 7948
rect 9152 7922 9737 7928
rect 9526 7898 9565 7902
rect 9771 7901 9805 8107
rect 10334 8122 10369 8128
rect 10334 8103 10339 8122
rect 10360 8103 10369 8122
rect 10334 8094 10369 8103
rect 10546 8124 10602 8129
rect 10546 8104 10553 8124
rect 10573 8104 10602 8124
rect 10546 8097 10602 8104
rect 11169 8168 11503 8196
rect 10546 8096 10581 8097
rect 10338 8026 10367 8094
rect 10338 7992 10684 8026
rect 9526 7878 9534 7898
rect 9554 7878 9565 7898
rect 6864 7869 6899 7877
rect 6864 7849 6872 7869
rect 6892 7861 6899 7869
rect 6892 7849 6903 7861
rect 6864 7612 6903 7849
rect 7734 7826 8020 7827
rect 7219 7818 8022 7826
rect 7219 7801 7230 7818
rect 7220 7796 7230 7801
rect 7254 7801 8022 7818
rect 7254 7796 7259 7801
rect 7220 7783 7259 7796
rect 7764 7735 7799 7736
rect 7743 7728 7799 7735
rect 7743 7708 7772 7728
rect 7792 7708 7799 7728
rect 7743 7703 7799 7708
rect 7983 7726 8022 7801
rect 9526 7803 9565 7878
rect 9749 7896 9805 7901
rect 9749 7876 9756 7896
rect 9776 7876 9805 7896
rect 9749 7869 9805 7876
rect 9749 7868 9784 7869
rect 10289 7808 10328 7821
rect 10289 7803 10294 7808
rect 9526 7786 10294 7803
rect 10318 7803 10328 7808
rect 10318 7786 10329 7803
rect 9526 7778 10329 7786
rect 9528 7777 9814 7778
rect 10645 7755 10684 7992
rect 10645 7743 10656 7755
rect 10649 7735 10656 7743
rect 10676 7735 10684 7755
rect 10649 7727 10684 7735
rect 7983 7706 7994 7726
rect 8014 7706 8022 7726
rect 6864 7578 7210 7612
rect 7181 7510 7210 7578
rect 6967 7507 7002 7508
rect 6792 7329 6795 7347
rect 6817 7329 6824 7347
rect 6792 7317 6824 7329
rect 6946 7500 7002 7507
rect 6946 7480 6975 7500
rect 6995 7480 7002 7500
rect 6946 7475 7002 7480
rect 7179 7501 7214 7510
rect 7179 7482 7188 7501
rect 7209 7482 7214 7501
rect 7179 7476 7214 7482
rect 7743 7497 7777 7703
rect 7983 7702 8022 7706
rect 7811 7676 8396 7682
rect 7811 7656 7827 7676
rect 7847 7675 8396 7676
rect 7847 7656 8367 7675
rect 7811 7655 8367 7656
rect 8387 7655 8396 7675
rect 7811 7647 8396 7655
rect 10031 7569 10616 7577
rect 10031 7549 10040 7569
rect 10060 7568 10616 7569
rect 10060 7549 10580 7568
rect 10031 7548 10580 7549
rect 10600 7548 10616 7568
rect 10031 7542 10616 7548
rect 9755 7534 9787 7535
rect 9752 7529 9787 7534
rect 9752 7509 9759 7529
rect 9779 7509 9787 7529
rect 10650 7521 10684 7727
rect 9752 7501 9787 7509
rect 7743 7489 7778 7497
rect 6946 7269 6980 7475
rect 7743 7469 7751 7489
rect 7771 7469 7778 7489
rect 7743 7464 7778 7469
rect 7743 7463 7775 7464
rect 7014 7448 7599 7454
rect 7014 7428 7030 7448
rect 7050 7447 7599 7448
rect 7050 7428 7570 7447
rect 7014 7427 7570 7428
rect 7590 7427 7599 7447
rect 7014 7419 7599 7427
rect 7679 7418 7709 7419
rect 7679 7391 8015 7418
rect 7679 7390 7714 7391
rect 6946 7261 6981 7269
rect 6946 7241 6954 7261
rect 6974 7241 6981 7261
rect 6946 7236 6981 7241
rect 6946 7215 6980 7236
rect 7679 7215 7709 7390
rect 7765 7323 7800 7324
rect 6946 7189 7709 7215
rect 6947 7188 6980 7189
rect 7679 7187 7709 7189
rect 7744 7316 7800 7323
rect 7744 7296 7773 7316
rect 7793 7296 7800 7316
rect 7744 7291 7800 7296
rect 7979 7318 8014 7391
rect 7979 7298 7986 7318
rect 8006 7298 8014 7318
rect 9134 7343 9719 7351
rect 9134 7323 9143 7343
rect 9163 7342 9719 7343
rect 9163 7323 9683 7342
rect 9134 7322 9683 7323
rect 9703 7322 9719 7342
rect 9134 7316 9719 7322
rect 7979 7291 8014 7298
rect 9753 7295 9787 7501
rect 10418 7515 10449 7521
rect 10418 7496 10423 7515
rect 10444 7496 10449 7515
rect 10418 7454 10449 7496
rect 10628 7516 10684 7521
rect 10628 7496 10635 7516
rect 10655 7496 10684 7516
rect 10628 7489 10684 7496
rect 10628 7488 10663 7489
rect 10418 7426 10757 7454
rect 6584 7155 7047 7163
rect 6584 7133 6596 7155
rect 6620 7133 7047 7155
rect 6584 7132 7047 7133
rect 6586 7120 6625 7132
rect 7020 7101 7047 7132
rect 6802 7099 6837 7100
rect 6781 7092 6837 7099
rect 6781 7072 6810 7092
rect 6830 7072 6837 7092
rect 6781 7067 6837 7072
rect 7016 7092 7049 7101
rect 7016 7070 7021 7092
rect 7044 7070 7049 7092
rect 6781 6861 6815 7067
rect 7016 7064 7049 7070
rect 7744 7085 7778 7291
rect 9517 7288 9552 7295
rect 7812 7264 8397 7270
rect 7812 7244 7828 7264
rect 7848 7263 8397 7264
rect 7848 7244 8368 7263
rect 7812 7243 8368 7244
rect 8388 7243 8397 7263
rect 7812 7235 8397 7243
rect 9517 7268 9525 7288
rect 9545 7268 9552 7288
rect 9517 7195 9552 7268
rect 9731 7290 9787 7295
rect 9731 7270 9738 7290
rect 9758 7270 9787 7290
rect 9731 7263 9787 7270
rect 9822 7397 9852 7399
rect 10551 7397 10584 7398
rect 9822 7371 10585 7397
rect 9731 7262 9766 7263
rect 9822 7196 9852 7371
rect 10551 7350 10585 7371
rect 10550 7345 10585 7350
rect 10550 7325 10557 7345
rect 10577 7325 10585 7345
rect 10550 7317 10585 7325
rect 9817 7195 9852 7196
rect 9516 7168 9852 7195
rect 9822 7167 9852 7168
rect 9932 7159 10517 7167
rect 9932 7139 9941 7159
rect 9961 7158 10517 7159
rect 9961 7139 10481 7158
rect 9932 7138 10481 7139
rect 10501 7138 10517 7158
rect 9932 7132 10517 7138
rect 9756 7122 9788 7123
rect 9753 7117 9788 7122
rect 9753 7097 9760 7117
rect 9780 7097 9788 7117
rect 10551 7111 10585 7317
rect 9753 7089 9788 7097
rect 7744 7077 7779 7085
rect 7744 7057 7752 7077
rect 7772 7057 7779 7077
rect 7744 7052 7779 7057
rect 7744 7051 7776 7052
rect 6849 7040 7434 7046
rect 6849 7020 6865 7040
rect 6885 7039 7434 7040
rect 6885 7020 7405 7039
rect 6849 7019 7405 7020
rect 7425 7019 7434 7039
rect 6849 7011 7434 7019
rect 9135 6931 9720 6939
rect 9135 6911 9144 6931
rect 9164 6930 9720 6931
rect 9164 6911 9684 6930
rect 9135 6910 9684 6911
rect 9704 6910 9720 6930
rect 9135 6904 9720 6910
rect 9509 6880 9548 6884
rect 9754 6883 9788 7089
rect 10318 7101 10352 7109
rect 10318 7083 10325 7101
rect 10344 7083 10352 7101
rect 10318 7076 10352 7083
rect 10529 7106 10585 7111
rect 10529 7086 10536 7106
rect 10556 7086 10585 7106
rect 10529 7079 10585 7086
rect 10529 7078 10564 7079
rect 10322 7046 10351 7076
rect 10322 7038 10704 7046
rect 10322 7019 10675 7038
rect 10696 7019 10704 7038
rect 10322 7014 10704 7019
rect 6781 6860 6816 6861
rect 6749 6853 6816 6860
rect 6749 6833 6789 6853
rect 6809 6833 6816 6853
rect 6749 6830 6816 6833
rect 9509 6860 9517 6880
rect 9537 6860 9548 6880
rect 6749 6827 6814 6830
rect 6320 6726 6385 6729
rect 6318 6723 6385 6726
rect 6318 6703 6325 6723
rect 6345 6703 6385 6723
rect 6318 6696 6385 6703
rect 6318 6695 6353 6696
rect 3599 6675 3610 6695
rect 3630 6675 3638 6695
rect 2443 6536 2825 6541
rect 2443 6517 2451 6536
rect 2472 6517 2825 6536
rect 2443 6509 2825 6517
rect 2796 6479 2825 6509
rect 2583 6476 2618 6477
rect 2562 6469 2618 6476
rect 2562 6449 2591 6469
rect 2611 6449 2618 6469
rect 2562 6444 2618 6449
rect 2795 6472 2829 6479
rect 2795 6454 2803 6472
rect 2822 6454 2829 6472
rect 2795 6446 2829 6454
rect 3359 6466 3393 6672
rect 3599 6671 3638 6675
rect 3427 6645 4012 6651
rect 3427 6625 3443 6645
rect 3463 6644 4012 6645
rect 3463 6625 3983 6644
rect 3427 6624 3983 6625
rect 4003 6624 4012 6644
rect 3427 6616 4012 6624
rect 5700 6537 6285 6545
rect 5700 6517 5709 6537
rect 5729 6536 6285 6537
rect 5729 6517 6249 6536
rect 5700 6516 6249 6517
rect 6269 6516 6285 6536
rect 5700 6510 6285 6516
rect 5358 6504 5390 6505
rect 5355 6499 5390 6504
rect 5355 6479 5362 6499
rect 5382 6479 5390 6499
rect 5355 6471 5390 6479
rect 3359 6458 3394 6466
rect 2562 6238 2596 6444
rect 3359 6438 3367 6458
rect 3387 6438 3394 6458
rect 3359 6433 3394 6438
rect 3359 6432 3391 6433
rect 2630 6417 3215 6423
rect 2630 6397 2646 6417
rect 2666 6416 3215 6417
rect 2666 6397 3186 6416
rect 2630 6396 3186 6397
rect 3206 6396 3215 6416
rect 2630 6388 3215 6396
rect 3295 6387 3325 6388
rect 3295 6360 3631 6387
rect 3295 6359 3330 6360
rect 2562 6230 2597 6238
rect 2562 6210 2570 6230
rect 2590 6210 2597 6230
rect 2562 6205 2597 6210
rect 2562 6184 2596 6205
rect 3295 6184 3325 6359
rect 3381 6292 3416 6293
rect 2562 6158 3325 6184
rect 2563 6157 2596 6158
rect 3295 6156 3325 6158
rect 3360 6285 3416 6292
rect 3360 6265 3389 6285
rect 3409 6265 3416 6285
rect 3360 6260 3416 6265
rect 3595 6287 3630 6360
rect 3595 6267 3602 6287
rect 3622 6267 3630 6287
rect 4737 6313 5322 6321
rect 4737 6293 4746 6313
rect 4766 6312 5322 6313
rect 4766 6293 5286 6312
rect 4737 6292 5286 6293
rect 5306 6292 5322 6312
rect 4737 6286 5322 6292
rect 3595 6260 3630 6267
rect 5356 6265 5390 6471
rect 6083 6481 6124 6492
rect 6319 6489 6353 6695
rect 6083 6463 6093 6481
rect 6111 6463 6124 6481
rect 6083 6455 6124 6463
rect 6297 6484 6353 6489
rect 6297 6464 6304 6484
rect 6324 6464 6353 6484
rect 6297 6457 6353 6464
rect 6297 6456 6332 6457
rect 6092 6425 6118 6455
rect 6092 6424 6430 6425
rect 6092 6388 6446 6424
rect 2390 6101 2729 6129
rect 2484 6066 2519 6067
rect 2463 6059 2519 6066
rect 2463 6039 2492 6059
rect 2512 6039 2519 6059
rect 2463 6034 2519 6039
rect 2698 6059 2729 6101
rect 2698 6040 2703 6059
rect 2724 6040 2729 6059
rect 2698 6034 2729 6040
rect 3360 6054 3394 6260
rect 5120 6258 5155 6265
rect 3428 6233 4013 6239
rect 3428 6213 3444 6233
rect 3464 6232 4013 6233
rect 3464 6213 3984 6232
rect 3428 6212 3984 6213
rect 4004 6212 4013 6232
rect 3428 6204 4013 6212
rect 5120 6238 5128 6258
rect 5148 6238 5155 6258
rect 5120 6165 5155 6238
rect 5334 6260 5390 6265
rect 5334 6240 5341 6260
rect 5361 6240 5390 6260
rect 5334 6233 5390 6240
rect 5425 6367 5455 6369
rect 6154 6367 6187 6368
rect 5425 6341 6188 6367
rect 5334 6232 5369 6233
rect 5425 6166 5455 6341
rect 6154 6320 6188 6341
rect 6153 6315 6188 6320
rect 6153 6295 6160 6315
rect 6180 6295 6188 6315
rect 6153 6287 6188 6295
rect 5420 6165 5455 6166
rect 5119 6138 5455 6165
rect 5425 6137 5455 6138
rect 5535 6129 6120 6137
rect 5535 6109 5544 6129
rect 5564 6128 6120 6129
rect 5564 6109 6084 6128
rect 5535 6108 6084 6109
rect 6104 6108 6120 6128
rect 5535 6102 6120 6108
rect 5359 6092 5391 6093
rect 5356 6087 5391 6092
rect 5356 6067 5363 6087
rect 5383 6067 5391 6087
rect 6154 6081 6188 6287
rect 5356 6059 5391 6067
rect 3360 6046 3395 6054
rect 2463 5828 2497 6034
rect 3360 6026 3368 6046
rect 3388 6026 3395 6046
rect 3360 6021 3395 6026
rect 3360 6020 3392 6021
rect 2531 6007 3116 6013
rect 2531 5987 2547 6007
rect 2567 6006 3116 6007
rect 2567 5987 3087 6006
rect 2531 5986 3087 5987
rect 3107 5986 3116 6006
rect 2531 5978 3116 5986
rect 4738 5901 5323 5909
rect 4738 5881 4747 5901
rect 4767 5900 5323 5901
rect 4767 5881 5287 5900
rect 4738 5880 5287 5881
rect 5307 5880 5323 5900
rect 4738 5874 5323 5880
rect 5112 5850 5151 5854
rect 5357 5853 5391 6059
rect 5920 6074 5955 6080
rect 5920 6055 5925 6074
rect 5946 6055 5955 6074
rect 5920 6046 5955 6055
rect 6132 6076 6188 6081
rect 6132 6056 6139 6076
rect 6159 6056 6188 6076
rect 6132 6049 6188 6056
rect 6132 6048 6167 6049
rect 5924 5978 5953 6046
rect 5924 5944 6270 5978
rect 5112 5830 5120 5850
rect 5140 5830 5151 5850
rect 2463 5820 2498 5828
rect 2463 5800 2471 5820
rect 2491 5812 2498 5820
rect 2491 5800 2502 5812
rect 2463 5563 2502 5800
rect 3333 5777 3619 5778
rect 2818 5769 3621 5777
rect 2818 5752 2829 5769
rect 2819 5747 2829 5752
rect 2853 5752 3621 5769
rect 2853 5747 2858 5752
rect 2819 5734 2858 5747
rect 3363 5686 3398 5687
rect 3342 5679 3398 5686
rect 3342 5659 3371 5679
rect 3391 5659 3398 5679
rect 3342 5654 3398 5659
rect 3582 5677 3621 5752
rect 5112 5755 5151 5830
rect 5335 5848 5391 5853
rect 5335 5828 5342 5848
rect 5362 5828 5391 5848
rect 5335 5821 5391 5828
rect 5335 5820 5370 5821
rect 5875 5760 5914 5773
rect 5875 5755 5880 5760
rect 5112 5738 5880 5755
rect 5904 5755 5914 5760
rect 5904 5738 5915 5755
rect 5112 5730 5915 5738
rect 5114 5729 5400 5730
rect 6231 5707 6270 5944
rect 6231 5695 6242 5707
rect 6235 5687 6242 5695
rect 6262 5687 6270 5707
rect 6235 5679 6270 5687
rect 3582 5657 3593 5677
rect 3613 5657 3621 5677
rect 2463 5529 2809 5563
rect 2780 5461 2809 5529
rect 2566 5458 2601 5459
rect 2545 5451 2601 5458
rect 2545 5431 2574 5451
rect 2594 5431 2601 5451
rect 2545 5426 2601 5431
rect 2778 5452 2813 5461
rect 2778 5433 2787 5452
rect 2808 5433 2813 5452
rect 2778 5427 2813 5433
rect 3342 5448 3376 5654
rect 3582 5653 3621 5657
rect 3410 5627 3995 5633
rect 3410 5607 3426 5627
rect 3446 5626 3995 5627
rect 3446 5607 3966 5626
rect 3410 5606 3966 5607
rect 3986 5606 3995 5626
rect 3410 5598 3995 5606
rect 5617 5521 6202 5529
rect 5617 5501 5626 5521
rect 5646 5520 6202 5521
rect 5646 5501 6166 5520
rect 5617 5500 6166 5501
rect 6186 5500 6202 5520
rect 5617 5494 6202 5500
rect 5341 5486 5373 5487
rect 5338 5481 5373 5486
rect 5338 5461 5345 5481
rect 5365 5461 5373 5481
rect 6236 5473 6270 5679
rect 5338 5453 5373 5461
rect 3342 5440 3377 5448
rect 2545 5220 2579 5426
rect 3342 5420 3350 5440
rect 3370 5420 3377 5440
rect 3342 5415 3377 5420
rect 3342 5414 3374 5415
rect 2613 5399 3198 5405
rect 2613 5379 2629 5399
rect 2649 5398 3198 5399
rect 2649 5379 3169 5398
rect 2613 5378 3169 5379
rect 3189 5378 3198 5398
rect 2613 5370 3198 5378
rect 3278 5369 3308 5370
rect 3278 5342 3614 5369
rect 3278 5341 3313 5342
rect 2545 5212 2580 5220
rect 2545 5192 2553 5212
rect 2573 5192 2580 5212
rect 2545 5187 2580 5192
rect 2545 5166 2579 5187
rect 3278 5166 3308 5341
rect 3364 5274 3399 5275
rect 2545 5140 3308 5166
rect 2546 5139 2579 5140
rect 3278 5138 3308 5140
rect 3343 5267 3399 5274
rect 3343 5247 3372 5267
rect 3392 5247 3399 5267
rect 3343 5242 3399 5247
rect 3578 5269 3613 5342
rect 3578 5249 3585 5269
rect 3605 5249 3613 5269
rect 4720 5295 5305 5303
rect 4720 5275 4729 5295
rect 4749 5294 5305 5295
rect 4749 5275 5269 5294
rect 4720 5274 5269 5275
rect 5289 5274 5305 5294
rect 4720 5268 5305 5274
rect 3578 5242 3613 5249
rect 5339 5247 5373 5453
rect 6002 5461 6038 5470
rect 6002 5444 6011 5461
rect 6030 5444 6038 5461
rect 6002 5435 6038 5444
rect 6214 5468 6270 5473
rect 6214 5448 6221 5468
rect 6241 5448 6270 5468
rect 6214 5441 6270 5448
rect 6214 5440 6249 5441
rect 6008 5400 6034 5435
rect 6316 5400 6348 5401
rect 6008 5395 6348 5400
rect 6008 5377 6323 5395
rect 6345 5377 6348 5395
rect 6008 5372 6348 5377
rect 6316 5371 6348 5372
rect 2197 5119 2514 5122
rect 2197 5092 2200 5119
rect 2227 5092 2514 5119
rect 2197 5086 2514 5092
rect 2197 5083 2233 5086
rect 2478 5056 2514 5086
rect 2262 5052 2297 5053
rect 2241 5045 2297 5052
rect 2241 5025 2270 5045
rect 2290 5025 2297 5045
rect 2241 5020 2297 5025
rect 2476 5050 2514 5056
rect 2476 5024 2482 5050
rect 2508 5024 2514 5050
rect 2241 4821 2275 5020
rect 2476 5016 2514 5024
rect 3343 5036 3377 5242
rect 5103 5240 5138 5247
rect 3411 5215 3996 5221
rect 3411 5195 3427 5215
rect 3447 5214 3996 5215
rect 3447 5195 3967 5214
rect 3411 5194 3967 5195
rect 3987 5194 3996 5214
rect 3411 5186 3996 5194
rect 5103 5220 5111 5240
rect 5131 5220 5138 5240
rect 5103 5147 5138 5220
rect 5317 5242 5373 5247
rect 5317 5222 5324 5242
rect 5344 5222 5373 5242
rect 5317 5215 5373 5222
rect 5408 5349 5438 5351
rect 6137 5349 6170 5350
rect 5408 5323 6171 5349
rect 5317 5214 5352 5215
rect 5408 5148 5438 5323
rect 6137 5302 6171 5323
rect 6136 5297 6171 5302
rect 6136 5277 6143 5297
rect 6163 5277 6171 5297
rect 6136 5269 6171 5277
rect 5403 5147 5438 5148
rect 5102 5120 5438 5147
rect 5408 5119 5438 5120
rect 5518 5111 6103 5119
rect 5518 5091 5527 5111
rect 5547 5110 6103 5111
rect 5547 5091 6067 5110
rect 5518 5090 6067 5091
rect 6087 5090 6103 5110
rect 5518 5084 6103 5090
rect 5342 5074 5374 5075
rect 5339 5069 5374 5074
rect 5339 5049 5346 5069
rect 5366 5049 5374 5069
rect 6137 5063 6171 5269
rect 5339 5041 5374 5049
rect 3343 5028 3378 5036
rect 3343 5008 3351 5028
rect 3371 5008 3378 5028
rect 3343 5003 3378 5008
rect 3343 5002 3375 5003
rect 2309 4993 2894 4999
rect 2309 4973 2325 4993
rect 2345 4992 2894 4993
rect 2345 4973 2865 4992
rect 2309 4972 2865 4973
rect 2885 4972 2894 4992
rect 2309 4964 2894 4972
rect 4721 4883 5306 4891
rect 4721 4863 4730 4883
rect 4750 4882 5306 4883
rect 4750 4863 5270 4882
rect 4721 4862 5270 4863
rect 5290 4862 5306 4882
rect 4721 4856 5306 4862
rect 5095 4832 5134 4836
rect 5340 4835 5374 5041
rect 5904 5053 5938 5061
rect 5904 5035 5911 5053
rect 5930 5035 5938 5053
rect 5904 5028 5938 5035
rect 6115 5058 6171 5063
rect 6115 5038 6122 5058
rect 6142 5038 6171 5058
rect 6115 5031 6171 5038
rect 6115 5030 6150 5031
rect 5908 4998 5937 5028
rect 5908 4990 6290 4998
rect 5908 4971 6261 4990
rect 6282 4971 6290 4990
rect 5908 4966 6290 4971
rect 2241 4806 2278 4821
rect 2241 4786 2249 4806
rect 2269 4786 2278 4806
rect 2241 4783 2278 4786
rect 2055 4672 2092 4675
rect 2055 4652 2064 4672
rect 2084 4652 2092 4672
rect 2055 4637 2092 4652
rect 1439 4486 2024 4494
rect 1439 4466 1448 4486
rect 1468 4485 2024 4486
rect 1468 4466 1988 4485
rect 1439 4465 1988 4466
rect 2008 4465 2024 4485
rect 1439 4459 2024 4465
rect 958 4455 990 4456
rect 955 4450 990 4455
rect 955 4430 962 4450
rect 982 4430 990 4450
rect 2058 4438 2092 4637
rect 2036 4433 2092 4438
rect 955 4422 990 4430
rect 337 4264 922 4272
rect 337 4244 346 4264
rect 366 4263 922 4264
rect 366 4244 886 4263
rect 337 4243 886 4244
rect 906 4243 922 4263
rect 337 4237 922 4243
rect 956 4216 990 4422
rect 1818 4431 1853 4433
rect 1818 4425 1856 4431
rect 1818 4402 1826 4425
rect 1849 4402 1856 4425
rect 2036 4413 2043 4433
rect 2063 4413 2092 4433
rect 2036 4406 2092 4413
rect 2036 4405 2071 4406
rect 1818 4396 1856 4402
rect 1818 4383 1853 4396
rect 1816 4325 1853 4383
rect 720 4209 755 4216
rect 720 4189 728 4209
rect 748 4189 755 4209
rect 720 4116 755 4189
rect 934 4211 990 4216
rect 934 4191 941 4211
rect 961 4191 990 4211
rect 934 4184 990 4191
rect 1025 4318 1055 4320
rect 1754 4318 1787 4319
rect 1025 4292 1788 4318
rect 934 4183 969 4184
rect 1025 4117 1055 4292
rect 1754 4271 1788 4292
rect 1816 4308 1851 4325
rect 1816 4307 2110 4308
rect 1816 4306 2153 4307
rect 1816 4299 2158 4306
rect 1816 4273 2118 4299
rect 2149 4273 2158 4299
rect 1753 4266 1788 4271
rect 2109 4270 2158 4273
rect 1753 4246 1760 4266
rect 1780 4246 1788 4266
rect 2115 4265 2158 4270
rect 1753 4238 1788 4246
rect 1020 4116 1055 4117
rect 719 4089 1055 4116
rect 1025 4088 1055 4089
rect 1135 4080 1720 4088
rect 1135 4060 1144 4080
rect 1164 4079 1720 4080
rect 1164 4060 1684 4079
rect 1135 4059 1684 4060
rect 1704 4059 1720 4079
rect 1135 4053 1720 4059
rect 959 4043 991 4044
rect 956 4038 991 4043
rect 956 4018 963 4038
rect 983 4018 991 4038
rect 1754 4032 1788 4238
rect 956 4010 991 4018
rect 338 3852 923 3860
rect 338 3832 347 3852
rect 367 3851 923 3852
rect 367 3832 887 3851
rect 338 3831 887 3832
rect 907 3831 923 3851
rect 338 3825 923 3831
rect 712 3801 751 3805
rect 957 3804 991 4010
rect 1520 4025 1555 4031
rect 1520 4006 1525 4025
rect 1546 4006 1555 4025
rect 1520 3997 1555 4006
rect 1732 4027 1788 4032
rect 1732 4007 1739 4027
rect 1759 4007 1788 4027
rect 1732 4000 1788 4007
rect 1732 3999 1767 4000
rect 1524 3929 1553 3997
rect 1524 3895 1870 3929
rect 712 3781 720 3801
rect 740 3781 751 3801
rect 712 3706 751 3781
rect 935 3799 991 3804
rect 935 3779 942 3799
rect 962 3779 991 3799
rect 935 3772 991 3779
rect 935 3771 970 3772
rect 1475 3711 1514 3724
rect 1475 3706 1480 3711
rect 712 3689 1480 3706
rect 1504 3706 1514 3711
rect 1504 3689 1515 3706
rect 712 3681 1515 3689
rect 714 3680 1000 3681
rect 1831 3658 1870 3895
rect 1831 3646 1842 3658
rect 1835 3638 1842 3646
rect 1862 3638 1870 3658
rect 1835 3630 1870 3638
rect 1217 3472 1802 3480
rect 1217 3452 1226 3472
rect 1246 3471 1802 3472
rect 1246 3452 1766 3471
rect 1217 3451 1766 3452
rect 1786 3451 1802 3471
rect 1217 3445 1802 3451
rect 941 3437 973 3438
rect 938 3432 973 3437
rect 938 3412 945 3432
rect 965 3412 973 3432
rect 1836 3424 1870 3630
rect 938 3404 973 3412
rect 320 3246 905 3254
rect 320 3226 329 3246
rect 349 3245 905 3246
rect 349 3226 869 3245
rect 320 3225 869 3226
rect 889 3225 905 3245
rect 320 3219 905 3225
rect 939 3198 973 3404
rect 1604 3418 1635 3424
rect 1604 3399 1609 3418
rect 1630 3399 1635 3418
rect 1604 3357 1635 3399
rect 1814 3419 1870 3424
rect 1814 3399 1821 3419
rect 1841 3399 1870 3419
rect 1814 3392 1870 3399
rect 1814 3391 1849 3392
rect 1604 3329 1943 3357
rect 703 3191 738 3198
rect 703 3171 711 3191
rect 731 3171 738 3191
rect 703 3098 738 3171
rect 917 3193 973 3198
rect 917 3173 924 3193
rect 944 3173 973 3193
rect 917 3166 973 3173
rect 1008 3300 1038 3302
rect 1737 3300 1770 3301
rect 1008 3274 1771 3300
rect 917 3165 952 3166
rect 1008 3099 1038 3274
rect 1737 3253 1771 3274
rect 1736 3248 1771 3253
rect 1736 3228 1743 3248
rect 1763 3228 1771 3248
rect 1736 3220 1771 3228
rect 1003 3098 1038 3099
rect 702 3071 1038 3098
rect 1008 3070 1038 3071
rect 1118 3062 1703 3070
rect 1118 3042 1127 3062
rect 1147 3061 1703 3062
rect 1147 3042 1667 3061
rect 1118 3041 1667 3042
rect 1687 3041 1703 3061
rect 1118 3035 1703 3041
rect 942 3025 974 3026
rect 939 3020 974 3025
rect 939 3000 946 3020
rect 966 3000 974 3020
rect 1737 3014 1771 3220
rect 939 2992 974 3000
rect 321 2834 906 2842
rect 321 2814 330 2834
rect 350 2833 906 2834
rect 350 2814 870 2833
rect 321 2813 870 2814
rect 890 2813 906 2833
rect 321 2807 906 2813
rect 695 2783 734 2787
rect 940 2786 974 2992
rect 1504 3004 1538 3012
rect 1504 2986 1511 3004
rect 1530 2986 1538 3004
rect 1504 2979 1538 2986
rect 1715 3009 1771 3014
rect 1715 2989 1722 3009
rect 1742 2989 1771 3009
rect 1715 2982 1771 2989
rect 1715 2981 1750 2982
rect 1508 2949 1537 2979
rect 1508 2941 1890 2949
rect 1508 2922 1861 2941
rect 1882 2922 1890 2941
rect 1508 2917 1890 2922
rect 695 2763 703 2783
rect 723 2763 734 2783
rect 695 2688 734 2763
rect 918 2781 974 2786
rect 918 2761 925 2781
rect 945 2761 974 2781
rect 918 2754 974 2761
rect 918 2753 953 2754
rect 1458 2693 1497 2706
rect 1458 2688 1463 2693
rect 695 2671 1463 2688
rect 1487 2688 1497 2693
rect 1487 2671 1498 2688
rect 695 2663 1498 2671
rect 697 2662 983 2663
rect 1914 2644 1943 3329
rect 2251 3083 2278 4783
rect 5095 4812 5103 4832
rect 5123 4812 5134 4832
rect 3314 4759 3600 4760
rect 2799 4751 3602 4759
rect 2799 4734 2810 4751
rect 2800 4729 2810 4734
rect 2834 4734 3602 4751
rect 2834 4729 2839 4734
rect 2800 4716 2839 4729
rect 3344 4668 3379 4669
rect 3323 4661 3379 4668
rect 3323 4641 3352 4661
rect 3372 4641 3379 4661
rect 3323 4636 3379 4641
rect 3563 4659 3602 4734
rect 5095 4737 5134 4812
rect 5318 4830 5374 4835
rect 5318 4810 5325 4830
rect 5345 4810 5374 4830
rect 5318 4803 5374 4810
rect 5318 4802 5353 4803
rect 5858 4742 5897 4755
rect 5858 4737 5863 4742
rect 5095 4720 5863 4737
rect 5887 4737 5897 4742
rect 5887 4720 5898 4737
rect 5095 4712 5898 4720
rect 5097 4711 5383 4712
rect 3563 4639 3574 4659
rect 3594 4639 3602 4659
rect 6419 4688 6446 6388
rect 6754 6142 6783 6827
rect 7714 6808 8000 6809
rect 7199 6800 8002 6808
rect 7199 6783 7210 6800
rect 7200 6778 7210 6783
rect 7234 6783 8002 6800
rect 7234 6778 7239 6783
rect 7200 6765 7239 6778
rect 7744 6717 7779 6718
rect 7723 6710 7779 6717
rect 7723 6690 7752 6710
rect 7772 6690 7779 6710
rect 7723 6685 7779 6690
rect 7963 6708 8002 6783
rect 9509 6785 9548 6860
rect 9732 6878 9788 6883
rect 9732 6858 9739 6878
rect 9759 6858 9788 6878
rect 9732 6851 9788 6858
rect 9732 6850 9767 6851
rect 10272 6790 10311 6803
rect 10272 6785 10277 6790
rect 9509 6768 10277 6785
rect 10301 6785 10311 6790
rect 10301 6768 10312 6785
rect 9509 6760 10312 6768
rect 9511 6759 9797 6760
rect 10728 6741 10757 7426
rect 11169 7359 11201 8168
rect 11477 8133 11503 8168
rect 11262 8127 11297 8128
rect 11241 8120 11297 8127
rect 11241 8100 11270 8120
rect 11290 8100 11297 8120
rect 11241 8095 11297 8100
rect 11473 8124 11509 8133
rect 11473 8107 11481 8124
rect 11500 8107 11509 8124
rect 11473 8098 11509 8107
rect 12138 8115 12172 8321
rect 13898 8319 13933 8326
rect 12206 8294 12791 8300
rect 12206 8274 12222 8294
rect 12242 8293 12791 8294
rect 12242 8274 12762 8293
rect 12206 8273 12762 8274
rect 12782 8273 12791 8293
rect 12206 8265 12791 8273
rect 13898 8299 13906 8319
rect 13926 8299 13933 8319
rect 13898 8226 13933 8299
rect 14112 8321 14168 8326
rect 14112 8301 14119 8321
rect 14139 8301 14168 8321
rect 14112 8294 14168 8301
rect 14203 8428 14233 8430
rect 14932 8428 14965 8429
rect 14203 8402 14966 8428
rect 14112 8293 14147 8294
rect 14203 8227 14233 8402
rect 14932 8381 14966 8402
rect 14931 8376 14966 8381
rect 14931 8356 14938 8376
rect 14958 8356 14966 8376
rect 14931 8348 14966 8356
rect 14198 8226 14233 8227
rect 13897 8199 14233 8226
rect 14203 8198 14233 8199
rect 14313 8190 14898 8198
rect 14313 8170 14322 8190
rect 14342 8189 14898 8190
rect 14342 8170 14862 8189
rect 14313 8169 14862 8170
rect 14882 8169 14898 8189
rect 14313 8163 14898 8169
rect 14137 8153 14169 8154
rect 14134 8148 14169 8153
rect 14134 8128 14141 8148
rect 14161 8128 14169 8148
rect 14932 8142 14966 8348
rect 15704 8312 15738 8518
rect 16501 8512 16509 8532
rect 16529 8512 16536 8532
rect 16501 8507 16536 8512
rect 16501 8506 16533 8507
rect 15772 8491 16357 8497
rect 15772 8471 15788 8491
rect 15808 8490 16357 8491
rect 15808 8471 16328 8490
rect 15772 8470 16328 8471
rect 16348 8470 16357 8490
rect 15772 8462 16357 8470
rect 16437 8461 16467 8462
rect 16437 8434 16773 8461
rect 16437 8433 16472 8434
rect 15704 8304 15739 8312
rect 15704 8284 15712 8304
rect 15732 8284 15739 8304
rect 15704 8279 15739 8284
rect 15704 8258 15738 8279
rect 16437 8258 16467 8433
rect 16523 8366 16558 8367
rect 15704 8232 16467 8258
rect 15705 8231 15738 8232
rect 16437 8230 16467 8232
rect 16502 8359 16558 8366
rect 16502 8339 16531 8359
rect 16551 8339 16558 8359
rect 16502 8334 16558 8339
rect 16737 8361 16772 8434
rect 16737 8341 16744 8361
rect 16764 8341 16772 8361
rect 16737 8334 16772 8341
rect 14134 8120 14169 8128
rect 12138 8107 12173 8115
rect 11241 7889 11275 8095
rect 12138 8087 12146 8107
rect 12166 8087 12173 8107
rect 12138 8082 12173 8087
rect 12138 8081 12170 8082
rect 11309 8068 11894 8074
rect 11309 8048 11325 8068
rect 11345 8067 11894 8068
rect 11345 8048 11865 8067
rect 11309 8047 11865 8048
rect 11885 8047 11894 8067
rect 11309 8039 11894 8047
rect 13516 7962 14101 7970
rect 13516 7942 13525 7962
rect 13545 7961 14101 7962
rect 13545 7942 14065 7961
rect 13516 7941 14065 7942
rect 14085 7941 14101 7961
rect 13516 7935 14101 7941
rect 13890 7911 13929 7915
rect 14135 7914 14169 8120
rect 14698 8135 14733 8141
rect 14698 8116 14703 8135
rect 14724 8116 14733 8135
rect 14698 8107 14733 8116
rect 14910 8137 14966 8142
rect 14910 8117 14917 8137
rect 14937 8117 14966 8137
rect 14910 8110 14966 8117
rect 15533 8181 15867 8209
rect 14910 8109 14945 8110
rect 14702 8039 14731 8107
rect 14702 8005 15048 8039
rect 13890 7891 13898 7911
rect 13918 7891 13929 7911
rect 11241 7881 11276 7889
rect 11241 7861 11249 7881
rect 11269 7873 11276 7881
rect 11269 7861 11280 7873
rect 11241 7624 11280 7861
rect 12111 7838 12397 7839
rect 11596 7830 12399 7838
rect 11596 7813 11607 7830
rect 11597 7808 11607 7813
rect 11631 7813 12399 7830
rect 11631 7808 11636 7813
rect 11597 7795 11636 7808
rect 12141 7747 12176 7748
rect 12120 7740 12176 7747
rect 12120 7720 12149 7740
rect 12169 7720 12176 7740
rect 12120 7715 12176 7720
rect 12360 7738 12399 7813
rect 13890 7816 13929 7891
rect 14113 7909 14169 7914
rect 14113 7889 14120 7909
rect 14140 7889 14169 7909
rect 14113 7882 14169 7889
rect 14113 7881 14148 7882
rect 14653 7821 14692 7834
rect 14653 7816 14658 7821
rect 13890 7799 14658 7816
rect 14682 7816 14692 7821
rect 14682 7799 14693 7816
rect 13890 7791 14693 7799
rect 13892 7790 14178 7791
rect 15009 7768 15048 8005
rect 15009 7756 15020 7768
rect 15013 7748 15020 7756
rect 15040 7748 15048 7768
rect 15013 7740 15048 7748
rect 12360 7718 12371 7738
rect 12391 7718 12399 7738
rect 11241 7590 11587 7624
rect 11558 7522 11587 7590
rect 11344 7519 11379 7520
rect 11169 7341 11172 7359
rect 11194 7341 11201 7359
rect 11169 7329 11201 7341
rect 11323 7512 11379 7519
rect 11323 7492 11352 7512
rect 11372 7492 11379 7512
rect 11323 7487 11379 7492
rect 11556 7513 11591 7522
rect 11556 7494 11565 7513
rect 11586 7494 11591 7513
rect 11556 7488 11591 7494
rect 12120 7509 12154 7715
rect 12360 7714 12399 7718
rect 12188 7688 12773 7694
rect 12188 7668 12204 7688
rect 12224 7687 12773 7688
rect 12224 7668 12744 7687
rect 12188 7667 12744 7668
rect 12764 7667 12773 7687
rect 12188 7659 12773 7667
rect 14395 7582 14980 7590
rect 14395 7562 14404 7582
rect 14424 7581 14980 7582
rect 14424 7562 14944 7581
rect 14395 7561 14944 7562
rect 14964 7561 14980 7581
rect 14395 7555 14980 7561
rect 14119 7547 14151 7548
rect 14116 7542 14151 7547
rect 14116 7522 14123 7542
rect 14143 7522 14151 7542
rect 15014 7534 15048 7740
rect 14116 7514 14151 7522
rect 12120 7501 12155 7509
rect 11323 7281 11357 7487
rect 12120 7481 12128 7501
rect 12148 7481 12155 7501
rect 12120 7476 12155 7481
rect 12120 7475 12152 7476
rect 11391 7460 11976 7466
rect 11391 7440 11407 7460
rect 11427 7459 11976 7460
rect 11427 7440 11947 7459
rect 11391 7439 11947 7440
rect 11967 7439 11976 7459
rect 11391 7431 11976 7439
rect 12056 7430 12086 7431
rect 12056 7403 12392 7430
rect 12056 7402 12091 7403
rect 11323 7273 11358 7281
rect 11323 7253 11331 7273
rect 11351 7253 11358 7273
rect 11323 7248 11358 7253
rect 11323 7227 11357 7248
rect 12056 7227 12086 7402
rect 12142 7335 12177 7336
rect 11323 7201 12086 7227
rect 11324 7200 11357 7201
rect 12056 7199 12086 7201
rect 12121 7328 12177 7335
rect 12121 7308 12150 7328
rect 12170 7308 12177 7328
rect 12121 7303 12177 7308
rect 12356 7330 12391 7403
rect 12356 7310 12363 7330
rect 12383 7310 12391 7330
rect 13498 7356 14083 7364
rect 13498 7336 13507 7356
rect 13527 7355 14083 7356
rect 13527 7336 14047 7355
rect 13498 7335 14047 7336
rect 14067 7335 14083 7355
rect 13498 7329 14083 7335
rect 12356 7303 12391 7310
rect 14117 7308 14151 7514
rect 14782 7528 14813 7534
rect 14782 7509 14787 7528
rect 14808 7509 14813 7528
rect 14782 7467 14813 7509
rect 14992 7529 15048 7534
rect 14992 7509 14999 7529
rect 15019 7509 15048 7529
rect 14992 7502 15048 7509
rect 14992 7501 15027 7502
rect 14782 7439 15121 7467
rect 10961 7167 11424 7175
rect 10961 7145 10973 7167
rect 10997 7145 11424 7167
rect 10961 7144 11424 7145
rect 10963 7132 11002 7144
rect 11397 7113 11424 7144
rect 11179 7111 11214 7112
rect 11158 7104 11214 7111
rect 11158 7084 11187 7104
rect 11207 7084 11214 7104
rect 11158 7079 11214 7084
rect 11393 7104 11426 7113
rect 11393 7082 11398 7104
rect 11421 7082 11426 7104
rect 11158 6873 11192 7079
rect 11393 7076 11426 7082
rect 12121 7097 12155 7303
rect 13881 7301 13916 7308
rect 12189 7276 12774 7282
rect 12189 7256 12205 7276
rect 12225 7275 12774 7276
rect 12225 7256 12745 7275
rect 12189 7255 12745 7256
rect 12765 7255 12774 7275
rect 12189 7247 12774 7255
rect 13881 7281 13889 7301
rect 13909 7281 13916 7301
rect 13881 7208 13916 7281
rect 14095 7303 14151 7308
rect 14095 7283 14102 7303
rect 14122 7283 14151 7303
rect 14095 7276 14151 7283
rect 14186 7410 14216 7412
rect 14915 7410 14948 7411
rect 14186 7384 14949 7410
rect 14095 7275 14130 7276
rect 14186 7209 14216 7384
rect 14915 7363 14949 7384
rect 14914 7358 14949 7363
rect 14914 7338 14921 7358
rect 14941 7338 14949 7358
rect 14914 7330 14949 7338
rect 14181 7208 14216 7209
rect 13880 7181 14216 7208
rect 14186 7180 14216 7181
rect 14296 7172 14881 7180
rect 14296 7152 14305 7172
rect 14325 7171 14881 7172
rect 14325 7152 14845 7171
rect 14296 7151 14845 7152
rect 14865 7151 14881 7171
rect 14296 7145 14881 7151
rect 14120 7135 14152 7136
rect 14117 7130 14152 7135
rect 14117 7110 14124 7130
rect 14144 7110 14152 7130
rect 14915 7124 14949 7330
rect 14117 7102 14152 7110
rect 12121 7089 12156 7097
rect 12121 7069 12129 7089
rect 12149 7069 12156 7089
rect 12121 7064 12156 7069
rect 12121 7063 12153 7064
rect 11226 7052 11811 7058
rect 11226 7032 11242 7052
rect 11262 7051 11811 7052
rect 11262 7032 11782 7051
rect 11226 7031 11782 7032
rect 11802 7031 11811 7051
rect 11226 7023 11811 7031
rect 13499 6944 14084 6952
rect 13499 6924 13508 6944
rect 13528 6943 14084 6944
rect 13528 6924 14048 6943
rect 13499 6923 14048 6924
rect 14068 6923 14084 6943
rect 13499 6917 14084 6923
rect 13873 6893 13912 6897
rect 14118 6896 14152 7102
rect 14682 7114 14716 7122
rect 14682 7096 14689 7114
rect 14708 7096 14716 7114
rect 14682 7089 14716 7096
rect 14893 7119 14949 7124
rect 14893 7099 14900 7119
rect 14920 7099 14949 7119
rect 14893 7092 14949 7099
rect 14893 7091 14928 7092
rect 14686 7059 14715 7089
rect 14686 7051 15068 7059
rect 14686 7032 15039 7051
rect 15060 7032 15068 7051
rect 14686 7027 15068 7032
rect 13873 6873 13881 6893
rect 13901 6873 13912 6893
rect 11158 6872 11193 6873
rect 11126 6865 11193 6872
rect 11126 6845 11166 6865
rect 11186 6845 11193 6865
rect 11126 6842 11193 6845
rect 11126 6839 11191 6842
rect 10697 6738 10762 6741
rect 7963 6688 7974 6708
rect 7994 6688 8002 6708
rect 10695 6735 10762 6738
rect 10695 6715 10702 6735
rect 10722 6715 10762 6735
rect 10695 6708 10762 6715
rect 10695 6707 10730 6708
rect 6807 6549 7189 6554
rect 6807 6530 6815 6549
rect 6836 6530 7189 6549
rect 6807 6522 7189 6530
rect 7160 6492 7189 6522
rect 6947 6489 6982 6490
rect 6926 6482 6982 6489
rect 6926 6462 6955 6482
rect 6975 6462 6982 6482
rect 6926 6457 6982 6462
rect 7159 6485 7193 6492
rect 7159 6467 7167 6485
rect 7186 6467 7193 6485
rect 7159 6459 7193 6467
rect 7723 6479 7757 6685
rect 7963 6684 8002 6688
rect 7791 6658 8376 6664
rect 7791 6638 7807 6658
rect 7827 6657 8376 6658
rect 7827 6638 8347 6657
rect 7791 6637 8347 6638
rect 8367 6637 8376 6657
rect 7791 6629 8376 6637
rect 10077 6549 10662 6557
rect 10077 6529 10086 6549
rect 10106 6548 10662 6549
rect 10106 6529 10626 6548
rect 10077 6528 10626 6529
rect 10646 6528 10662 6548
rect 10077 6522 10662 6528
rect 9735 6516 9767 6517
rect 9732 6511 9767 6516
rect 9732 6491 9739 6511
rect 9759 6491 9767 6511
rect 9732 6483 9767 6491
rect 7723 6471 7758 6479
rect 6926 6251 6960 6457
rect 7723 6451 7731 6471
rect 7751 6451 7758 6471
rect 7723 6446 7758 6451
rect 7723 6445 7755 6446
rect 6994 6430 7579 6436
rect 6994 6410 7010 6430
rect 7030 6429 7579 6430
rect 7030 6410 7550 6429
rect 6994 6409 7550 6410
rect 7570 6409 7579 6429
rect 6994 6401 7579 6409
rect 7659 6400 7689 6401
rect 7659 6373 7995 6400
rect 7659 6372 7694 6373
rect 6926 6243 6961 6251
rect 6926 6223 6934 6243
rect 6954 6223 6961 6243
rect 6926 6218 6961 6223
rect 6926 6197 6960 6218
rect 7659 6197 7689 6372
rect 7745 6305 7780 6306
rect 6926 6171 7689 6197
rect 6927 6170 6960 6171
rect 7659 6169 7689 6171
rect 7724 6298 7780 6305
rect 7724 6278 7753 6298
rect 7773 6278 7780 6298
rect 7724 6273 7780 6278
rect 7959 6300 7994 6373
rect 7959 6280 7966 6300
rect 7986 6280 7994 6300
rect 9114 6325 9699 6333
rect 9114 6305 9123 6325
rect 9143 6324 9699 6325
rect 9143 6305 9663 6324
rect 9114 6304 9663 6305
rect 9683 6304 9699 6324
rect 9114 6298 9699 6304
rect 7959 6273 7994 6280
rect 9733 6277 9767 6483
rect 10460 6493 10501 6504
rect 10696 6501 10730 6707
rect 10460 6475 10470 6493
rect 10488 6475 10501 6493
rect 10460 6467 10501 6475
rect 10674 6496 10730 6501
rect 10674 6476 10681 6496
rect 10701 6476 10730 6496
rect 10674 6469 10730 6476
rect 10674 6468 10709 6469
rect 10469 6437 10495 6467
rect 10469 6436 10807 6437
rect 10469 6400 10823 6436
rect 6754 6114 7093 6142
rect 6848 6079 6883 6080
rect 6827 6072 6883 6079
rect 6827 6052 6856 6072
rect 6876 6052 6883 6072
rect 6827 6047 6883 6052
rect 7062 6072 7093 6114
rect 7062 6053 7067 6072
rect 7088 6053 7093 6072
rect 7062 6047 7093 6053
rect 7724 6067 7758 6273
rect 9497 6270 9532 6277
rect 7792 6246 8377 6252
rect 7792 6226 7808 6246
rect 7828 6245 8377 6246
rect 7828 6226 8348 6245
rect 7792 6225 8348 6226
rect 8368 6225 8377 6245
rect 7792 6217 8377 6225
rect 9497 6250 9505 6270
rect 9525 6250 9532 6270
rect 9497 6177 9532 6250
rect 9711 6272 9767 6277
rect 9711 6252 9718 6272
rect 9738 6252 9767 6272
rect 9711 6245 9767 6252
rect 9802 6379 9832 6381
rect 10531 6379 10564 6380
rect 9802 6353 10565 6379
rect 9711 6244 9746 6245
rect 9802 6178 9832 6353
rect 10531 6332 10565 6353
rect 10530 6327 10565 6332
rect 10530 6307 10537 6327
rect 10557 6307 10565 6327
rect 10530 6299 10565 6307
rect 9797 6177 9832 6178
rect 9496 6150 9832 6177
rect 9802 6149 9832 6150
rect 9912 6141 10497 6149
rect 9912 6121 9921 6141
rect 9941 6140 10497 6141
rect 9941 6121 10461 6140
rect 9912 6120 10461 6121
rect 10481 6120 10497 6140
rect 9912 6114 10497 6120
rect 9736 6104 9768 6105
rect 9733 6099 9768 6104
rect 9733 6079 9740 6099
rect 9760 6079 9768 6099
rect 10531 6093 10565 6299
rect 9733 6071 9768 6079
rect 7724 6059 7759 6067
rect 6827 5841 6861 6047
rect 7724 6039 7732 6059
rect 7752 6039 7759 6059
rect 7724 6034 7759 6039
rect 7724 6033 7756 6034
rect 6895 6020 7480 6026
rect 6895 6000 6911 6020
rect 6931 6019 7480 6020
rect 6931 6000 7451 6019
rect 6895 5999 7451 6000
rect 7471 5999 7480 6019
rect 6895 5991 7480 5999
rect 9115 5913 9700 5921
rect 9115 5893 9124 5913
rect 9144 5912 9700 5913
rect 9144 5893 9664 5912
rect 9115 5892 9664 5893
rect 9684 5892 9700 5912
rect 9115 5886 9700 5892
rect 9489 5862 9528 5866
rect 9734 5865 9768 6071
rect 10297 6086 10332 6092
rect 10297 6067 10302 6086
rect 10323 6067 10332 6086
rect 10297 6058 10332 6067
rect 10509 6088 10565 6093
rect 10509 6068 10516 6088
rect 10536 6068 10565 6088
rect 10509 6061 10565 6068
rect 10509 6060 10544 6061
rect 10301 5990 10330 6058
rect 10301 5956 10647 5990
rect 9489 5842 9497 5862
rect 9517 5842 9528 5862
rect 6827 5833 6862 5841
rect 6827 5813 6835 5833
rect 6855 5825 6862 5833
rect 6855 5813 6866 5825
rect 6827 5576 6866 5813
rect 7697 5790 7983 5791
rect 7182 5782 7985 5790
rect 7182 5765 7193 5782
rect 7183 5760 7193 5765
rect 7217 5765 7985 5782
rect 7217 5760 7222 5765
rect 7183 5747 7222 5760
rect 7727 5699 7762 5700
rect 7706 5692 7762 5699
rect 7706 5672 7735 5692
rect 7755 5672 7762 5692
rect 7706 5667 7762 5672
rect 7946 5690 7985 5765
rect 9489 5767 9528 5842
rect 9712 5860 9768 5865
rect 9712 5840 9719 5860
rect 9739 5840 9768 5860
rect 9712 5833 9768 5840
rect 9712 5832 9747 5833
rect 10252 5772 10291 5785
rect 10252 5767 10257 5772
rect 9489 5750 10257 5767
rect 10281 5767 10291 5772
rect 10281 5750 10292 5767
rect 9489 5742 10292 5750
rect 9491 5741 9777 5742
rect 10608 5719 10647 5956
rect 10608 5707 10619 5719
rect 10612 5699 10619 5707
rect 10639 5699 10647 5719
rect 10612 5691 10647 5699
rect 7946 5670 7957 5690
rect 7977 5670 7985 5690
rect 6827 5542 7173 5576
rect 7144 5474 7173 5542
rect 6930 5471 6965 5472
rect 6909 5464 6965 5471
rect 6909 5444 6938 5464
rect 6958 5444 6965 5464
rect 6909 5439 6965 5444
rect 7142 5465 7177 5474
rect 7142 5446 7151 5465
rect 7172 5446 7177 5465
rect 7142 5440 7177 5446
rect 7706 5461 7740 5667
rect 7946 5666 7985 5670
rect 7774 5640 8359 5646
rect 7774 5620 7790 5640
rect 7810 5639 8359 5640
rect 7810 5620 8330 5639
rect 7774 5619 8330 5620
rect 8350 5619 8359 5639
rect 7774 5611 8359 5619
rect 9994 5533 10579 5541
rect 9994 5513 10003 5533
rect 10023 5532 10579 5533
rect 10023 5513 10543 5532
rect 9994 5512 10543 5513
rect 10563 5512 10579 5532
rect 9994 5506 10579 5512
rect 9718 5498 9750 5499
rect 9715 5493 9750 5498
rect 9715 5473 9722 5493
rect 9742 5473 9750 5493
rect 10613 5485 10647 5691
rect 9715 5465 9750 5473
rect 7706 5453 7741 5461
rect 6909 5233 6943 5439
rect 7706 5433 7714 5453
rect 7734 5433 7741 5453
rect 7706 5428 7741 5433
rect 7706 5427 7738 5428
rect 6977 5412 7562 5418
rect 6977 5392 6993 5412
rect 7013 5411 7562 5412
rect 7013 5392 7533 5411
rect 6977 5391 7533 5392
rect 7553 5391 7562 5411
rect 6977 5383 7562 5391
rect 7642 5382 7672 5383
rect 7642 5355 7978 5382
rect 7642 5354 7677 5355
rect 6909 5225 6944 5233
rect 6909 5205 6917 5225
rect 6937 5205 6944 5225
rect 6909 5200 6944 5205
rect 6909 5179 6943 5200
rect 7642 5179 7672 5354
rect 7728 5287 7763 5288
rect 6909 5153 7672 5179
rect 6910 5152 6943 5153
rect 7642 5151 7672 5153
rect 7707 5280 7763 5287
rect 7707 5260 7736 5280
rect 7756 5260 7763 5280
rect 7707 5255 7763 5260
rect 7942 5282 7977 5355
rect 7942 5262 7949 5282
rect 7969 5262 7977 5282
rect 9097 5307 9682 5315
rect 9097 5287 9106 5307
rect 9126 5306 9682 5307
rect 9126 5287 9646 5306
rect 9097 5286 9646 5287
rect 9666 5286 9682 5306
rect 9097 5280 9682 5286
rect 7942 5255 7977 5262
rect 9716 5259 9750 5465
rect 10379 5473 10415 5482
rect 10379 5456 10388 5473
rect 10407 5456 10415 5473
rect 10379 5447 10415 5456
rect 10591 5480 10647 5485
rect 10591 5460 10598 5480
rect 10618 5460 10647 5480
rect 10591 5453 10647 5460
rect 10591 5452 10626 5453
rect 10385 5412 10411 5447
rect 10693 5412 10725 5413
rect 10385 5407 10725 5412
rect 10385 5389 10700 5407
rect 10722 5389 10725 5407
rect 10385 5384 10725 5389
rect 10693 5383 10725 5384
rect 6561 5132 6878 5135
rect 6561 5105 6564 5132
rect 6591 5105 6878 5132
rect 6561 5099 6878 5105
rect 6561 5096 6597 5099
rect 6842 5069 6878 5099
rect 6626 5065 6661 5066
rect 6605 5058 6661 5065
rect 6605 5038 6634 5058
rect 6654 5038 6661 5058
rect 6605 5033 6661 5038
rect 6840 5063 6878 5069
rect 6840 5037 6846 5063
rect 6872 5037 6878 5063
rect 6605 4834 6639 5033
rect 6840 5029 6878 5037
rect 7707 5049 7741 5255
rect 9480 5252 9515 5259
rect 7775 5228 8360 5234
rect 7775 5208 7791 5228
rect 7811 5227 8360 5228
rect 7811 5208 8331 5227
rect 7775 5207 8331 5208
rect 8351 5207 8360 5227
rect 7775 5199 8360 5207
rect 9480 5232 9488 5252
rect 9508 5232 9515 5252
rect 9480 5159 9515 5232
rect 9694 5254 9750 5259
rect 9694 5234 9701 5254
rect 9721 5234 9750 5254
rect 9694 5227 9750 5234
rect 9785 5361 9815 5363
rect 10514 5361 10547 5362
rect 9785 5335 10548 5361
rect 9694 5226 9729 5227
rect 9785 5160 9815 5335
rect 10514 5314 10548 5335
rect 10513 5309 10548 5314
rect 10513 5289 10520 5309
rect 10540 5289 10548 5309
rect 10513 5281 10548 5289
rect 9780 5159 9815 5160
rect 9479 5132 9815 5159
rect 9785 5131 9815 5132
rect 9895 5123 10480 5131
rect 9895 5103 9904 5123
rect 9924 5122 10480 5123
rect 9924 5103 10444 5122
rect 9895 5102 10444 5103
rect 10464 5102 10480 5122
rect 9895 5096 10480 5102
rect 9719 5086 9751 5087
rect 9716 5081 9751 5086
rect 9716 5061 9723 5081
rect 9743 5061 9751 5081
rect 10514 5075 10548 5281
rect 9716 5053 9751 5061
rect 7707 5041 7742 5049
rect 7707 5021 7715 5041
rect 7735 5021 7742 5041
rect 7707 5016 7742 5021
rect 7707 5015 7739 5016
rect 6673 5006 7258 5012
rect 6673 4986 6689 5006
rect 6709 5005 7258 5006
rect 6709 4986 7229 5005
rect 6673 4985 7229 4986
rect 7249 4985 7258 5005
rect 6673 4977 7258 4985
rect 9098 4895 9683 4903
rect 9098 4875 9107 4895
rect 9127 4894 9683 4895
rect 9127 4875 9647 4894
rect 9098 4874 9647 4875
rect 9667 4874 9683 4894
rect 9098 4868 9683 4874
rect 9472 4844 9511 4848
rect 9717 4847 9751 5053
rect 10281 5065 10315 5073
rect 10281 5047 10288 5065
rect 10307 5047 10315 5065
rect 10281 5040 10315 5047
rect 10492 5070 10548 5075
rect 10492 5050 10499 5070
rect 10519 5050 10548 5070
rect 10492 5043 10548 5050
rect 10492 5042 10527 5043
rect 10285 5010 10314 5040
rect 10285 5002 10667 5010
rect 10285 4983 10638 5002
rect 10659 4983 10667 5002
rect 10285 4978 10667 4983
rect 6605 4819 6642 4834
rect 6605 4799 6613 4819
rect 6633 4799 6642 4819
rect 6605 4796 6642 4799
rect 6419 4685 6456 4688
rect 6419 4665 6428 4685
rect 6448 4665 6456 4685
rect 6419 4650 6456 4665
rect 2407 4500 2789 4505
rect 2407 4481 2415 4500
rect 2436 4481 2789 4500
rect 2407 4473 2789 4481
rect 2760 4443 2789 4473
rect 2547 4440 2582 4441
rect 2526 4433 2582 4440
rect 2526 4413 2555 4433
rect 2575 4413 2582 4433
rect 2526 4408 2582 4413
rect 2759 4436 2793 4443
rect 2759 4418 2767 4436
rect 2786 4418 2793 4436
rect 2759 4410 2793 4418
rect 3323 4430 3357 4636
rect 3563 4635 3602 4639
rect 3391 4609 3976 4615
rect 3391 4589 3407 4609
rect 3427 4608 3976 4609
rect 3427 4589 3947 4608
rect 3391 4588 3947 4589
rect 3967 4588 3976 4608
rect 3391 4580 3976 4588
rect 5803 4499 6388 4507
rect 5803 4479 5812 4499
rect 5832 4498 6388 4499
rect 5832 4479 6352 4498
rect 5803 4478 6352 4479
rect 6372 4478 6388 4498
rect 5803 4472 6388 4478
rect 5322 4468 5354 4469
rect 5319 4463 5354 4468
rect 5319 4443 5326 4463
rect 5346 4443 5354 4463
rect 6422 4451 6456 4650
rect 6400 4446 6456 4451
rect 5319 4435 5354 4443
rect 3323 4422 3358 4430
rect 2526 4202 2560 4408
rect 3323 4402 3331 4422
rect 3351 4402 3358 4422
rect 3323 4397 3358 4402
rect 3323 4396 3355 4397
rect 2594 4381 3179 4387
rect 2594 4361 2610 4381
rect 2630 4380 3179 4381
rect 2630 4361 3150 4380
rect 2594 4360 3150 4361
rect 3170 4360 3179 4380
rect 2594 4352 3179 4360
rect 3259 4351 3289 4352
rect 3259 4324 3595 4351
rect 3259 4323 3294 4324
rect 2526 4194 2561 4202
rect 2526 4174 2534 4194
rect 2554 4174 2561 4194
rect 2526 4169 2561 4174
rect 2526 4148 2560 4169
rect 3259 4148 3289 4323
rect 3345 4256 3380 4257
rect 2526 4122 3289 4148
rect 2527 4121 2560 4122
rect 3259 4120 3289 4122
rect 3324 4249 3380 4256
rect 3324 4229 3353 4249
rect 3373 4229 3380 4249
rect 3324 4224 3380 4229
rect 3559 4251 3594 4324
rect 3559 4231 3566 4251
rect 3586 4231 3594 4251
rect 4701 4277 5286 4285
rect 4701 4257 4710 4277
rect 4730 4276 5286 4277
rect 4730 4257 5250 4276
rect 4701 4256 5250 4257
rect 5270 4256 5286 4276
rect 4701 4250 5286 4256
rect 3559 4224 3594 4231
rect 5320 4229 5354 4435
rect 6182 4444 6217 4446
rect 6182 4438 6220 4444
rect 6182 4415 6190 4438
rect 6213 4415 6220 4438
rect 6400 4426 6407 4446
rect 6427 4426 6456 4446
rect 6400 4419 6456 4426
rect 6400 4418 6435 4419
rect 6182 4409 6220 4415
rect 6182 4396 6217 4409
rect 6180 4338 6217 4396
rect 2349 4099 2381 4100
rect 2349 4094 2689 4099
rect 2349 4076 2352 4094
rect 2374 4076 2689 4094
rect 2349 4071 2689 4076
rect 2349 4070 2381 4071
rect 2663 4036 2689 4071
rect 2448 4030 2483 4031
rect 2427 4023 2483 4030
rect 2427 4003 2456 4023
rect 2476 4003 2483 4023
rect 2427 3998 2483 4003
rect 2659 4027 2695 4036
rect 2659 4010 2667 4027
rect 2686 4010 2695 4027
rect 2659 4001 2695 4010
rect 3324 4018 3358 4224
rect 5084 4222 5119 4229
rect 3392 4197 3977 4203
rect 3392 4177 3408 4197
rect 3428 4196 3977 4197
rect 3428 4177 3948 4196
rect 3392 4176 3948 4177
rect 3968 4176 3977 4196
rect 3392 4168 3977 4176
rect 5084 4202 5092 4222
rect 5112 4202 5119 4222
rect 5084 4129 5119 4202
rect 5298 4224 5354 4229
rect 5298 4204 5305 4224
rect 5325 4204 5354 4224
rect 5298 4197 5354 4204
rect 5389 4331 5419 4333
rect 6118 4331 6151 4332
rect 5389 4305 6152 4331
rect 5298 4196 5333 4197
rect 5389 4130 5419 4305
rect 6118 4284 6152 4305
rect 6180 4321 6215 4338
rect 6180 4320 6474 4321
rect 6180 4319 6517 4320
rect 6180 4312 6522 4319
rect 6180 4286 6482 4312
rect 6513 4286 6522 4312
rect 6117 4279 6152 4284
rect 6473 4283 6522 4286
rect 6117 4259 6124 4279
rect 6144 4259 6152 4279
rect 6479 4278 6522 4283
rect 6117 4251 6152 4259
rect 5384 4129 5419 4130
rect 5083 4102 5419 4129
rect 5389 4101 5419 4102
rect 5499 4093 6084 4101
rect 5499 4073 5508 4093
rect 5528 4092 6084 4093
rect 5528 4073 6048 4092
rect 5499 4072 6048 4073
rect 6068 4072 6084 4092
rect 5499 4066 6084 4072
rect 5323 4056 5355 4057
rect 5320 4051 5355 4056
rect 5320 4031 5327 4051
rect 5347 4031 5355 4051
rect 6118 4045 6152 4251
rect 5320 4023 5355 4031
rect 3324 4010 3359 4018
rect 2427 3792 2461 3998
rect 3324 3990 3332 4010
rect 3352 3990 3359 4010
rect 3324 3985 3359 3990
rect 3324 3984 3356 3985
rect 2495 3971 3080 3977
rect 2495 3951 2511 3971
rect 2531 3970 3080 3971
rect 2531 3951 3051 3970
rect 2495 3950 3051 3951
rect 3071 3950 3080 3970
rect 2495 3942 3080 3950
rect 4702 3865 5287 3873
rect 4702 3845 4711 3865
rect 4731 3864 5287 3865
rect 4731 3845 5251 3864
rect 4702 3844 5251 3845
rect 5271 3844 5287 3864
rect 4702 3838 5287 3844
rect 5076 3814 5115 3818
rect 5321 3817 5355 4023
rect 5884 4038 5919 4044
rect 5884 4019 5889 4038
rect 5910 4019 5919 4038
rect 5884 4010 5919 4019
rect 6096 4040 6152 4045
rect 6096 4020 6103 4040
rect 6123 4020 6152 4040
rect 6096 4013 6152 4020
rect 6096 4012 6131 4013
rect 5888 3942 5917 4010
rect 5888 3908 6234 3942
rect 5076 3794 5084 3814
rect 5104 3794 5115 3814
rect 2427 3784 2462 3792
rect 2427 3764 2435 3784
rect 2455 3776 2462 3784
rect 2455 3764 2466 3776
rect 2427 3527 2466 3764
rect 3297 3741 3583 3742
rect 2782 3733 3585 3741
rect 2782 3716 2793 3733
rect 2783 3711 2793 3716
rect 2817 3716 3585 3733
rect 2817 3711 2822 3716
rect 2783 3698 2822 3711
rect 3327 3650 3362 3651
rect 3306 3643 3362 3650
rect 3306 3623 3335 3643
rect 3355 3623 3362 3643
rect 3306 3618 3362 3623
rect 3546 3641 3585 3716
rect 5076 3719 5115 3794
rect 5299 3812 5355 3817
rect 5299 3792 5306 3812
rect 5326 3792 5355 3812
rect 5299 3785 5355 3792
rect 5299 3784 5334 3785
rect 5839 3724 5878 3737
rect 5839 3719 5844 3724
rect 5076 3702 5844 3719
rect 5868 3719 5878 3724
rect 5868 3702 5879 3719
rect 5076 3694 5879 3702
rect 5078 3693 5364 3694
rect 6195 3671 6234 3908
rect 6195 3659 6206 3671
rect 6199 3651 6206 3659
rect 6226 3651 6234 3671
rect 6199 3643 6234 3651
rect 3546 3621 3557 3641
rect 3577 3621 3585 3641
rect 2427 3493 2773 3527
rect 2744 3425 2773 3493
rect 2530 3422 2565 3423
rect 2509 3415 2565 3422
rect 2509 3395 2538 3415
rect 2558 3395 2565 3415
rect 2509 3390 2565 3395
rect 2742 3416 2777 3425
rect 2742 3397 2751 3416
rect 2772 3397 2777 3416
rect 2742 3391 2777 3397
rect 3306 3412 3340 3618
rect 3546 3617 3585 3621
rect 3374 3591 3959 3597
rect 3374 3571 3390 3591
rect 3410 3590 3959 3591
rect 3410 3571 3930 3590
rect 3374 3570 3930 3571
rect 3950 3570 3959 3590
rect 3374 3562 3959 3570
rect 5581 3485 6166 3493
rect 5581 3465 5590 3485
rect 5610 3484 6166 3485
rect 5610 3465 6130 3484
rect 5581 3464 6130 3465
rect 6150 3464 6166 3484
rect 5581 3458 6166 3464
rect 5305 3450 5337 3451
rect 5302 3445 5337 3450
rect 5302 3425 5309 3445
rect 5329 3425 5337 3445
rect 6200 3437 6234 3643
rect 5302 3417 5337 3425
rect 3306 3404 3341 3412
rect 2509 3184 2543 3390
rect 3306 3384 3314 3404
rect 3334 3384 3341 3404
rect 3306 3379 3341 3384
rect 3306 3378 3338 3379
rect 2577 3363 3162 3369
rect 2577 3343 2593 3363
rect 2613 3362 3162 3363
rect 2613 3343 3133 3362
rect 2577 3342 3133 3343
rect 3153 3342 3162 3362
rect 2577 3334 3162 3342
rect 3242 3333 3272 3334
rect 3242 3306 3578 3333
rect 3242 3305 3277 3306
rect 2509 3176 2544 3184
rect 2509 3156 2517 3176
rect 2537 3156 2544 3176
rect 2509 3151 2544 3156
rect 2509 3130 2543 3151
rect 3242 3130 3272 3305
rect 3328 3238 3363 3239
rect 2509 3104 3272 3130
rect 2510 3103 2543 3104
rect 3242 3102 3272 3104
rect 3307 3231 3363 3238
rect 3307 3211 3336 3231
rect 3356 3211 3363 3231
rect 3307 3206 3363 3211
rect 3542 3233 3577 3306
rect 3542 3213 3549 3233
rect 3569 3213 3577 3233
rect 4684 3259 5269 3267
rect 4684 3239 4693 3259
rect 4713 3258 5269 3259
rect 4713 3239 5233 3258
rect 4684 3238 5233 3239
rect 5253 3238 5269 3258
rect 4684 3232 5269 3238
rect 3542 3206 3577 3213
rect 5303 3211 5337 3417
rect 5968 3431 5999 3437
rect 5968 3412 5973 3431
rect 5994 3412 5999 3431
rect 5968 3370 5999 3412
rect 6178 3432 6234 3437
rect 6178 3412 6185 3432
rect 6205 3412 6234 3432
rect 6178 3405 6234 3412
rect 6178 3404 6213 3405
rect 5968 3342 6307 3370
rect 2251 3047 2605 3083
rect 2267 3046 2605 3047
rect 2579 3016 2605 3046
rect 2365 3014 2400 3015
rect 2344 3007 2400 3014
rect 2344 2987 2373 3007
rect 2393 2987 2400 3007
rect 2344 2982 2400 2987
rect 2573 3008 2614 3016
rect 2573 2990 2586 3008
rect 2604 2990 2614 3008
rect 2344 2776 2378 2982
rect 2573 2979 2614 2990
rect 3307 3000 3341 3206
rect 5067 3204 5102 3211
rect 3375 3179 3960 3185
rect 3375 3159 3391 3179
rect 3411 3178 3960 3179
rect 3411 3159 3931 3178
rect 3375 3158 3931 3159
rect 3951 3158 3960 3178
rect 3375 3150 3960 3158
rect 5067 3184 5075 3204
rect 5095 3184 5102 3204
rect 5067 3111 5102 3184
rect 5281 3206 5337 3211
rect 5281 3186 5288 3206
rect 5308 3186 5337 3206
rect 5281 3179 5337 3186
rect 5372 3313 5402 3315
rect 6101 3313 6134 3314
rect 5372 3287 6135 3313
rect 5281 3178 5316 3179
rect 5372 3112 5402 3287
rect 6101 3266 6135 3287
rect 6100 3261 6135 3266
rect 6100 3241 6107 3261
rect 6127 3241 6135 3261
rect 6100 3233 6135 3241
rect 5367 3111 5402 3112
rect 5066 3084 5402 3111
rect 5372 3083 5402 3084
rect 5482 3075 6067 3083
rect 5482 3055 5491 3075
rect 5511 3074 6067 3075
rect 5511 3055 6031 3074
rect 5482 3054 6031 3055
rect 6051 3054 6067 3074
rect 5482 3048 6067 3054
rect 5306 3038 5338 3039
rect 5303 3033 5338 3038
rect 5303 3013 5310 3033
rect 5330 3013 5338 3033
rect 6101 3027 6135 3233
rect 5303 3005 5338 3013
rect 3307 2992 3342 3000
rect 3307 2972 3315 2992
rect 3335 2972 3342 2992
rect 3307 2967 3342 2972
rect 3307 2966 3339 2967
rect 2412 2955 2997 2961
rect 2412 2935 2428 2955
rect 2448 2954 2997 2955
rect 2448 2935 2968 2954
rect 2412 2934 2968 2935
rect 2988 2934 2997 2954
rect 2412 2926 2997 2934
rect 4685 2847 5270 2855
rect 4685 2827 4694 2847
rect 4714 2846 5270 2847
rect 4714 2827 5234 2846
rect 4685 2826 5234 2827
rect 5254 2826 5270 2846
rect 4685 2820 5270 2826
rect 5059 2796 5098 2800
rect 5304 2799 5338 3005
rect 5868 3017 5902 3025
rect 5868 2999 5875 3017
rect 5894 2999 5902 3017
rect 5868 2992 5902 2999
rect 6079 3022 6135 3027
rect 6079 3002 6086 3022
rect 6106 3002 6135 3022
rect 6079 2995 6135 3002
rect 6079 2994 6114 2995
rect 5872 2962 5901 2992
rect 5872 2954 6254 2962
rect 5872 2935 6225 2954
rect 6246 2935 6254 2954
rect 5872 2930 6254 2935
rect 5059 2776 5067 2796
rect 5087 2776 5098 2796
rect 2344 2775 2379 2776
rect 2312 2768 2379 2775
rect 2312 2748 2352 2768
rect 2372 2748 2379 2768
rect 2312 2745 2379 2748
rect 2312 2742 2377 2745
rect 1883 2641 1948 2644
rect 1881 2638 1948 2641
rect 1881 2618 1888 2638
rect 1908 2618 1948 2638
rect 1881 2611 1948 2618
rect 1881 2610 1916 2611
rect 1263 2452 1848 2460
rect 1263 2432 1272 2452
rect 1292 2451 1848 2452
rect 1292 2432 1812 2451
rect 1263 2431 1812 2432
rect 1832 2431 1848 2451
rect 1263 2425 1848 2431
rect 921 2419 953 2420
rect 918 2414 953 2419
rect 918 2394 925 2414
rect 945 2394 953 2414
rect 918 2386 953 2394
rect 300 2228 885 2236
rect 300 2208 309 2228
rect 329 2227 885 2228
rect 329 2208 849 2227
rect 300 2207 849 2208
rect 869 2207 885 2227
rect 300 2201 885 2207
rect 919 2180 953 2386
rect 1648 2401 1681 2407
rect 1882 2404 1916 2610
rect 1648 2379 1653 2401
rect 1676 2379 1681 2401
rect 1648 2370 1681 2379
rect 1860 2399 1916 2404
rect 1860 2379 1867 2399
rect 1887 2379 1916 2399
rect 1860 2372 1916 2379
rect 1860 2371 1895 2372
rect 1650 2339 1677 2370
rect 2072 2339 2111 2351
rect 1650 2338 2113 2339
rect 1650 2316 2077 2338
rect 2101 2316 2113 2338
rect 1650 2308 2113 2316
rect 683 2173 718 2180
rect 683 2153 691 2173
rect 711 2153 718 2173
rect 683 2080 718 2153
rect 897 2175 953 2180
rect 897 2155 904 2175
rect 924 2155 953 2175
rect 897 2148 953 2155
rect 988 2282 1018 2284
rect 1717 2282 1750 2283
rect 988 2256 1751 2282
rect 897 2147 932 2148
rect 988 2081 1018 2256
rect 1717 2235 1751 2256
rect 1716 2230 1751 2235
rect 1716 2210 1723 2230
rect 1743 2210 1751 2230
rect 1716 2202 1751 2210
rect 983 2080 1018 2081
rect 682 2053 1018 2080
rect 988 2052 1018 2053
rect 1098 2044 1683 2052
rect 1098 2024 1107 2044
rect 1127 2043 1683 2044
rect 1127 2024 1647 2043
rect 1098 2023 1647 2024
rect 1667 2023 1683 2043
rect 1098 2017 1683 2023
rect 922 2007 954 2008
rect 919 2002 954 2007
rect 919 1982 926 2002
rect 946 1982 954 2002
rect 1717 1996 1751 2202
rect 919 1974 954 1982
rect 301 1816 886 1824
rect 301 1796 310 1816
rect 330 1815 886 1816
rect 330 1796 850 1815
rect 301 1795 850 1796
rect 870 1795 886 1815
rect 301 1789 886 1795
rect 675 1765 714 1769
rect 920 1768 954 1974
rect 1483 1989 1518 1995
rect 1483 1970 1488 1989
rect 1509 1970 1518 1989
rect 1483 1961 1518 1970
rect 1695 1991 1751 1996
rect 1695 1971 1702 1991
rect 1722 1971 1751 1991
rect 1695 1964 1751 1971
rect 1873 2142 1905 2154
rect 1873 2124 1880 2142
rect 1902 2124 1905 2142
rect 1695 1963 1730 1964
rect 1487 1893 1516 1961
rect 1487 1859 1833 1893
rect 675 1745 683 1765
rect 703 1745 714 1765
rect 675 1670 714 1745
rect 898 1763 954 1768
rect 898 1743 905 1763
rect 925 1743 954 1763
rect 898 1736 954 1743
rect 898 1735 933 1736
rect 1438 1675 1477 1688
rect 1438 1670 1443 1675
rect 675 1653 1443 1670
rect 1467 1670 1477 1675
rect 1467 1653 1478 1670
rect 675 1645 1478 1653
rect 677 1644 963 1645
rect 1794 1622 1833 1859
rect 1794 1610 1805 1622
rect 1798 1602 1805 1610
rect 1825 1602 1833 1622
rect 1798 1594 1833 1602
rect 1180 1436 1765 1444
rect 1180 1416 1189 1436
rect 1209 1435 1765 1436
rect 1209 1416 1729 1435
rect 1180 1415 1729 1416
rect 1749 1415 1765 1435
rect 1180 1409 1765 1415
rect 904 1401 936 1402
rect 901 1396 936 1401
rect 901 1376 908 1396
rect 928 1376 936 1396
rect 1799 1388 1833 1594
rect 901 1368 936 1376
rect 283 1210 868 1218
rect 283 1190 292 1210
rect 312 1209 868 1210
rect 312 1190 832 1209
rect 283 1189 832 1190
rect 852 1189 868 1209
rect 283 1183 868 1189
rect 902 1162 936 1368
rect 1565 1376 1601 1385
rect 1565 1359 1574 1376
rect 1593 1359 1601 1376
rect 1565 1350 1601 1359
rect 1777 1383 1833 1388
rect 1777 1363 1784 1383
rect 1804 1363 1833 1383
rect 1777 1356 1833 1363
rect 1777 1355 1812 1356
rect 1571 1315 1597 1350
rect 1873 1315 1905 2124
rect 2317 2057 2346 2742
rect 3277 2723 3563 2724
rect 2762 2715 3565 2723
rect 2762 2698 2773 2715
rect 2763 2693 2773 2698
rect 2797 2698 3565 2715
rect 2797 2693 2802 2698
rect 2763 2680 2802 2693
rect 3307 2632 3342 2633
rect 3286 2625 3342 2632
rect 3286 2605 3315 2625
rect 3335 2605 3342 2625
rect 3286 2600 3342 2605
rect 3526 2623 3565 2698
rect 5059 2701 5098 2776
rect 5282 2794 5338 2799
rect 5282 2774 5289 2794
rect 5309 2774 5338 2794
rect 5282 2767 5338 2774
rect 5282 2766 5317 2767
rect 5822 2706 5861 2719
rect 5822 2701 5827 2706
rect 5059 2684 5827 2701
rect 5851 2701 5861 2706
rect 5851 2684 5862 2701
rect 5059 2676 5862 2684
rect 5061 2675 5347 2676
rect 6278 2657 6307 3342
rect 6615 3096 6642 4796
rect 9472 4824 9480 4844
rect 9500 4824 9511 4844
rect 7678 4772 7964 4773
rect 7163 4764 7966 4772
rect 7163 4747 7174 4764
rect 7164 4742 7174 4747
rect 7198 4747 7966 4764
rect 7198 4742 7203 4747
rect 7164 4729 7203 4742
rect 7708 4681 7743 4682
rect 7687 4674 7743 4681
rect 7687 4654 7716 4674
rect 7736 4654 7743 4674
rect 7687 4649 7743 4654
rect 7927 4672 7966 4747
rect 9472 4749 9511 4824
rect 9695 4842 9751 4847
rect 9695 4822 9702 4842
rect 9722 4822 9751 4842
rect 9695 4815 9751 4822
rect 9695 4814 9730 4815
rect 10235 4754 10274 4767
rect 10235 4749 10240 4754
rect 9472 4732 10240 4749
rect 10264 4749 10274 4754
rect 10264 4732 10275 4749
rect 9472 4724 10275 4732
rect 9474 4723 9760 4724
rect 7927 4652 7938 4672
rect 7958 4652 7966 4672
rect 10796 4700 10823 6400
rect 11131 6154 11160 6839
rect 12091 6820 12377 6821
rect 11576 6812 12379 6820
rect 11576 6795 11587 6812
rect 11577 6790 11587 6795
rect 11611 6795 12379 6812
rect 11611 6790 11616 6795
rect 11577 6777 11616 6790
rect 12121 6729 12156 6730
rect 12100 6722 12156 6729
rect 12100 6702 12129 6722
rect 12149 6702 12156 6722
rect 12100 6697 12156 6702
rect 12340 6720 12379 6795
rect 13873 6798 13912 6873
rect 14096 6891 14152 6896
rect 14096 6871 14103 6891
rect 14123 6871 14152 6891
rect 14096 6864 14152 6871
rect 14096 6863 14131 6864
rect 14636 6803 14675 6816
rect 14636 6798 14641 6803
rect 13873 6781 14641 6798
rect 14665 6798 14675 6803
rect 14665 6781 14676 6798
rect 13873 6773 14676 6781
rect 13875 6772 14161 6773
rect 15092 6754 15121 7439
rect 15533 7372 15565 8181
rect 15841 8146 15867 8181
rect 15626 8140 15661 8141
rect 15605 8133 15661 8140
rect 15605 8113 15634 8133
rect 15654 8113 15661 8133
rect 15605 8108 15661 8113
rect 15837 8137 15873 8146
rect 15837 8120 15845 8137
rect 15864 8120 15873 8137
rect 15837 8111 15873 8120
rect 16502 8128 16536 8334
rect 16570 8307 17155 8313
rect 16570 8287 16586 8307
rect 16606 8306 17155 8307
rect 16606 8287 17126 8306
rect 16570 8286 17126 8287
rect 17146 8286 17155 8306
rect 16570 8278 17155 8286
rect 16502 8120 16537 8128
rect 15605 7902 15639 8108
rect 16502 8100 16510 8120
rect 16530 8100 16537 8120
rect 16502 8095 16537 8100
rect 16502 8094 16534 8095
rect 15673 8081 16258 8087
rect 15673 8061 15689 8081
rect 15709 8080 16258 8081
rect 15709 8061 16229 8080
rect 15673 8060 16229 8061
rect 16249 8060 16258 8080
rect 15673 8052 16258 8060
rect 15605 7894 15640 7902
rect 15605 7874 15613 7894
rect 15633 7886 15640 7894
rect 15633 7874 15644 7886
rect 15605 7637 15644 7874
rect 16475 7851 16761 7852
rect 15960 7843 16763 7851
rect 15960 7826 15971 7843
rect 15961 7821 15971 7826
rect 15995 7826 16763 7843
rect 15995 7821 16000 7826
rect 15961 7808 16000 7821
rect 16505 7760 16540 7761
rect 16484 7753 16540 7760
rect 16484 7733 16513 7753
rect 16533 7733 16540 7753
rect 16484 7728 16540 7733
rect 16724 7751 16763 7826
rect 16724 7731 16735 7751
rect 16755 7731 16763 7751
rect 15605 7603 15951 7637
rect 15922 7535 15951 7603
rect 15708 7532 15743 7533
rect 15533 7354 15536 7372
rect 15558 7354 15565 7372
rect 15533 7342 15565 7354
rect 15687 7525 15743 7532
rect 15687 7505 15716 7525
rect 15736 7505 15743 7525
rect 15687 7500 15743 7505
rect 15920 7526 15955 7535
rect 15920 7507 15929 7526
rect 15950 7507 15955 7526
rect 15920 7501 15955 7507
rect 16484 7522 16518 7728
rect 16724 7727 16763 7731
rect 16552 7701 17137 7707
rect 16552 7681 16568 7701
rect 16588 7700 17137 7701
rect 16588 7681 17108 7700
rect 16552 7680 17108 7681
rect 17128 7680 17137 7700
rect 16552 7672 17137 7680
rect 16484 7514 16519 7522
rect 15687 7294 15721 7500
rect 16484 7494 16492 7514
rect 16512 7494 16519 7514
rect 16484 7489 16519 7494
rect 16484 7488 16516 7489
rect 15755 7473 16340 7479
rect 15755 7453 15771 7473
rect 15791 7472 16340 7473
rect 15791 7453 16311 7472
rect 15755 7452 16311 7453
rect 16331 7452 16340 7472
rect 15755 7444 16340 7452
rect 16420 7443 16450 7444
rect 16420 7416 16756 7443
rect 16420 7415 16455 7416
rect 15687 7286 15722 7294
rect 15687 7266 15695 7286
rect 15715 7266 15722 7286
rect 15687 7261 15722 7266
rect 15687 7240 15721 7261
rect 16420 7240 16450 7415
rect 16506 7348 16541 7349
rect 15687 7214 16450 7240
rect 15688 7213 15721 7214
rect 16420 7212 16450 7214
rect 16485 7341 16541 7348
rect 16485 7321 16514 7341
rect 16534 7321 16541 7341
rect 16485 7316 16541 7321
rect 16720 7343 16755 7416
rect 16720 7323 16727 7343
rect 16747 7323 16755 7343
rect 16720 7316 16755 7323
rect 15325 7180 15788 7188
rect 15325 7158 15337 7180
rect 15361 7158 15788 7180
rect 15325 7157 15788 7158
rect 15327 7145 15366 7157
rect 15761 7126 15788 7157
rect 15543 7124 15578 7125
rect 15522 7117 15578 7124
rect 15522 7097 15551 7117
rect 15571 7097 15578 7117
rect 15522 7092 15578 7097
rect 15757 7117 15790 7126
rect 15757 7095 15762 7117
rect 15785 7095 15790 7117
rect 15522 6886 15556 7092
rect 15757 7089 15790 7095
rect 16485 7110 16519 7316
rect 16553 7289 17138 7295
rect 16553 7269 16569 7289
rect 16589 7288 17138 7289
rect 16589 7269 17109 7288
rect 16553 7268 17109 7269
rect 17129 7268 17138 7288
rect 16553 7260 17138 7268
rect 16485 7102 16520 7110
rect 16485 7082 16493 7102
rect 16513 7082 16520 7102
rect 16485 7077 16520 7082
rect 16485 7076 16517 7077
rect 15590 7065 16175 7071
rect 15590 7045 15606 7065
rect 15626 7064 16175 7065
rect 15626 7045 16146 7064
rect 15590 7044 16146 7045
rect 16166 7044 16175 7064
rect 15590 7036 16175 7044
rect 15522 6885 15557 6886
rect 15490 6878 15557 6885
rect 15490 6858 15530 6878
rect 15550 6858 15557 6878
rect 15490 6855 15557 6858
rect 15490 6852 15555 6855
rect 15061 6751 15126 6754
rect 15059 6748 15126 6751
rect 15059 6728 15066 6748
rect 15086 6728 15126 6748
rect 15059 6721 15126 6728
rect 15059 6720 15094 6721
rect 12340 6700 12351 6720
rect 12371 6700 12379 6720
rect 11184 6561 11566 6566
rect 11184 6542 11192 6561
rect 11213 6542 11566 6561
rect 11184 6534 11566 6542
rect 11537 6504 11566 6534
rect 11324 6501 11359 6502
rect 11303 6494 11359 6501
rect 11303 6474 11332 6494
rect 11352 6474 11359 6494
rect 11303 6469 11359 6474
rect 11536 6497 11570 6504
rect 11536 6479 11544 6497
rect 11563 6479 11570 6497
rect 11536 6471 11570 6479
rect 12100 6491 12134 6697
rect 12340 6696 12379 6700
rect 12168 6670 12753 6676
rect 12168 6650 12184 6670
rect 12204 6669 12753 6670
rect 12204 6650 12724 6669
rect 12168 6649 12724 6650
rect 12744 6649 12753 6669
rect 12168 6641 12753 6649
rect 14441 6562 15026 6570
rect 14441 6542 14450 6562
rect 14470 6561 15026 6562
rect 14470 6542 14990 6561
rect 14441 6541 14990 6542
rect 15010 6541 15026 6561
rect 14441 6535 15026 6541
rect 14099 6529 14131 6530
rect 14096 6524 14131 6529
rect 14096 6504 14103 6524
rect 14123 6504 14131 6524
rect 14096 6496 14131 6504
rect 12100 6483 12135 6491
rect 11303 6263 11337 6469
rect 12100 6463 12108 6483
rect 12128 6463 12135 6483
rect 12100 6458 12135 6463
rect 12100 6457 12132 6458
rect 11371 6442 11956 6448
rect 11371 6422 11387 6442
rect 11407 6441 11956 6442
rect 11407 6422 11927 6441
rect 11371 6421 11927 6422
rect 11947 6421 11956 6441
rect 11371 6413 11956 6421
rect 12036 6412 12066 6413
rect 12036 6385 12372 6412
rect 12036 6384 12071 6385
rect 11303 6255 11338 6263
rect 11303 6235 11311 6255
rect 11331 6235 11338 6255
rect 11303 6230 11338 6235
rect 11303 6209 11337 6230
rect 12036 6209 12066 6384
rect 12122 6317 12157 6318
rect 11303 6183 12066 6209
rect 11304 6182 11337 6183
rect 12036 6181 12066 6183
rect 12101 6310 12157 6317
rect 12101 6290 12130 6310
rect 12150 6290 12157 6310
rect 12101 6285 12157 6290
rect 12336 6312 12371 6385
rect 12336 6292 12343 6312
rect 12363 6292 12371 6312
rect 13478 6338 14063 6346
rect 13478 6318 13487 6338
rect 13507 6337 14063 6338
rect 13507 6318 14027 6337
rect 13478 6317 14027 6318
rect 14047 6317 14063 6337
rect 13478 6311 14063 6317
rect 12336 6285 12371 6292
rect 14097 6290 14131 6496
rect 14824 6506 14865 6517
rect 15060 6514 15094 6720
rect 14824 6488 14834 6506
rect 14852 6488 14865 6506
rect 14824 6480 14865 6488
rect 15038 6509 15094 6514
rect 15038 6489 15045 6509
rect 15065 6489 15094 6509
rect 15038 6482 15094 6489
rect 15038 6481 15073 6482
rect 14833 6450 14859 6480
rect 14833 6449 15171 6450
rect 14833 6413 15187 6449
rect 11131 6126 11470 6154
rect 11225 6091 11260 6092
rect 11204 6084 11260 6091
rect 11204 6064 11233 6084
rect 11253 6064 11260 6084
rect 11204 6059 11260 6064
rect 11439 6084 11470 6126
rect 11439 6065 11444 6084
rect 11465 6065 11470 6084
rect 11439 6059 11470 6065
rect 12101 6079 12135 6285
rect 13861 6283 13896 6290
rect 12169 6258 12754 6264
rect 12169 6238 12185 6258
rect 12205 6257 12754 6258
rect 12205 6238 12725 6257
rect 12169 6237 12725 6238
rect 12745 6237 12754 6257
rect 12169 6229 12754 6237
rect 13861 6263 13869 6283
rect 13889 6263 13896 6283
rect 13861 6190 13896 6263
rect 14075 6285 14131 6290
rect 14075 6265 14082 6285
rect 14102 6265 14131 6285
rect 14075 6258 14131 6265
rect 14166 6392 14196 6394
rect 14895 6392 14928 6393
rect 14166 6366 14929 6392
rect 14075 6257 14110 6258
rect 14166 6191 14196 6366
rect 14895 6345 14929 6366
rect 14894 6340 14929 6345
rect 14894 6320 14901 6340
rect 14921 6320 14929 6340
rect 14894 6312 14929 6320
rect 14161 6190 14196 6191
rect 13860 6163 14196 6190
rect 14166 6162 14196 6163
rect 14276 6154 14861 6162
rect 14276 6134 14285 6154
rect 14305 6153 14861 6154
rect 14305 6134 14825 6153
rect 14276 6133 14825 6134
rect 14845 6133 14861 6153
rect 14276 6127 14861 6133
rect 14100 6117 14132 6118
rect 14097 6112 14132 6117
rect 14097 6092 14104 6112
rect 14124 6092 14132 6112
rect 14895 6106 14929 6312
rect 14097 6084 14132 6092
rect 12101 6071 12136 6079
rect 11204 5853 11238 6059
rect 12101 6051 12109 6071
rect 12129 6051 12136 6071
rect 12101 6046 12136 6051
rect 12101 6045 12133 6046
rect 11272 6032 11857 6038
rect 11272 6012 11288 6032
rect 11308 6031 11857 6032
rect 11308 6012 11828 6031
rect 11272 6011 11828 6012
rect 11848 6011 11857 6031
rect 11272 6003 11857 6011
rect 13479 5926 14064 5934
rect 13479 5906 13488 5926
rect 13508 5925 14064 5926
rect 13508 5906 14028 5925
rect 13479 5905 14028 5906
rect 14048 5905 14064 5925
rect 13479 5899 14064 5905
rect 13853 5875 13892 5879
rect 14098 5878 14132 6084
rect 14661 6099 14696 6105
rect 14661 6080 14666 6099
rect 14687 6080 14696 6099
rect 14661 6071 14696 6080
rect 14873 6101 14929 6106
rect 14873 6081 14880 6101
rect 14900 6081 14929 6101
rect 14873 6074 14929 6081
rect 14873 6073 14908 6074
rect 14665 6003 14694 6071
rect 14665 5969 15011 6003
rect 13853 5855 13861 5875
rect 13881 5855 13892 5875
rect 11204 5845 11239 5853
rect 11204 5825 11212 5845
rect 11232 5837 11239 5845
rect 11232 5825 11243 5837
rect 11204 5588 11243 5825
rect 12074 5802 12360 5803
rect 11559 5794 12362 5802
rect 11559 5777 11570 5794
rect 11560 5772 11570 5777
rect 11594 5777 12362 5794
rect 11594 5772 11599 5777
rect 11560 5759 11599 5772
rect 12104 5711 12139 5712
rect 12083 5704 12139 5711
rect 12083 5684 12112 5704
rect 12132 5684 12139 5704
rect 12083 5679 12139 5684
rect 12323 5702 12362 5777
rect 13853 5780 13892 5855
rect 14076 5873 14132 5878
rect 14076 5853 14083 5873
rect 14103 5853 14132 5873
rect 14076 5846 14132 5853
rect 14076 5845 14111 5846
rect 14616 5785 14655 5798
rect 14616 5780 14621 5785
rect 13853 5763 14621 5780
rect 14645 5780 14655 5785
rect 14645 5763 14656 5780
rect 13853 5755 14656 5763
rect 13855 5754 14141 5755
rect 14972 5732 15011 5969
rect 14972 5720 14983 5732
rect 14976 5712 14983 5720
rect 15003 5712 15011 5732
rect 14976 5704 15011 5712
rect 12323 5682 12334 5702
rect 12354 5682 12362 5702
rect 11204 5554 11550 5588
rect 11521 5486 11550 5554
rect 11307 5483 11342 5484
rect 11286 5476 11342 5483
rect 11286 5456 11315 5476
rect 11335 5456 11342 5476
rect 11286 5451 11342 5456
rect 11519 5477 11554 5486
rect 11519 5458 11528 5477
rect 11549 5458 11554 5477
rect 11519 5452 11554 5458
rect 12083 5473 12117 5679
rect 12323 5678 12362 5682
rect 12151 5652 12736 5658
rect 12151 5632 12167 5652
rect 12187 5651 12736 5652
rect 12187 5632 12707 5651
rect 12151 5631 12707 5632
rect 12727 5631 12736 5651
rect 12151 5623 12736 5631
rect 14358 5546 14943 5554
rect 14358 5526 14367 5546
rect 14387 5545 14943 5546
rect 14387 5526 14907 5545
rect 14358 5525 14907 5526
rect 14927 5525 14943 5545
rect 14358 5519 14943 5525
rect 14082 5511 14114 5512
rect 14079 5506 14114 5511
rect 14079 5486 14086 5506
rect 14106 5486 14114 5506
rect 14977 5498 15011 5704
rect 14079 5478 14114 5486
rect 12083 5465 12118 5473
rect 11286 5245 11320 5451
rect 12083 5445 12091 5465
rect 12111 5445 12118 5465
rect 12083 5440 12118 5445
rect 12083 5439 12115 5440
rect 11354 5424 11939 5430
rect 11354 5404 11370 5424
rect 11390 5423 11939 5424
rect 11390 5404 11910 5423
rect 11354 5403 11910 5404
rect 11930 5403 11939 5423
rect 11354 5395 11939 5403
rect 12019 5394 12049 5395
rect 12019 5367 12355 5394
rect 12019 5366 12054 5367
rect 11286 5237 11321 5245
rect 11286 5217 11294 5237
rect 11314 5217 11321 5237
rect 11286 5212 11321 5217
rect 11286 5191 11320 5212
rect 12019 5191 12049 5366
rect 12105 5299 12140 5300
rect 11286 5165 12049 5191
rect 11287 5164 11320 5165
rect 12019 5163 12049 5165
rect 12084 5292 12140 5299
rect 12084 5272 12113 5292
rect 12133 5272 12140 5292
rect 12084 5267 12140 5272
rect 12319 5294 12354 5367
rect 12319 5274 12326 5294
rect 12346 5274 12354 5294
rect 13461 5320 14046 5328
rect 13461 5300 13470 5320
rect 13490 5319 14046 5320
rect 13490 5300 14010 5319
rect 13461 5299 14010 5300
rect 14030 5299 14046 5319
rect 13461 5293 14046 5299
rect 12319 5267 12354 5274
rect 14080 5272 14114 5478
rect 14743 5486 14779 5495
rect 14743 5469 14752 5486
rect 14771 5469 14779 5486
rect 14743 5460 14779 5469
rect 14955 5493 15011 5498
rect 14955 5473 14962 5493
rect 14982 5473 15011 5493
rect 14955 5466 15011 5473
rect 14955 5465 14990 5466
rect 14749 5425 14775 5460
rect 15057 5425 15089 5426
rect 14749 5420 15089 5425
rect 14749 5402 15064 5420
rect 15086 5402 15089 5420
rect 14749 5397 15089 5402
rect 15057 5396 15089 5397
rect 10938 5144 11255 5147
rect 10938 5117 10941 5144
rect 10968 5117 11255 5144
rect 10938 5111 11255 5117
rect 10938 5108 10974 5111
rect 11219 5081 11255 5111
rect 11003 5077 11038 5078
rect 10982 5070 11038 5077
rect 10982 5050 11011 5070
rect 11031 5050 11038 5070
rect 10982 5045 11038 5050
rect 11217 5075 11255 5081
rect 11217 5049 11223 5075
rect 11249 5049 11255 5075
rect 10982 4846 11016 5045
rect 11217 5041 11255 5049
rect 12084 5061 12118 5267
rect 13844 5265 13879 5272
rect 12152 5240 12737 5246
rect 12152 5220 12168 5240
rect 12188 5239 12737 5240
rect 12188 5220 12708 5239
rect 12152 5219 12708 5220
rect 12728 5219 12737 5239
rect 12152 5211 12737 5219
rect 13844 5245 13852 5265
rect 13872 5245 13879 5265
rect 13844 5172 13879 5245
rect 14058 5267 14114 5272
rect 14058 5247 14065 5267
rect 14085 5247 14114 5267
rect 14058 5240 14114 5247
rect 14149 5374 14179 5376
rect 14878 5374 14911 5375
rect 14149 5348 14912 5374
rect 14058 5239 14093 5240
rect 14149 5173 14179 5348
rect 14878 5327 14912 5348
rect 14877 5322 14912 5327
rect 14877 5302 14884 5322
rect 14904 5302 14912 5322
rect 14877 5294 14912 5302
rect 14144 5172 14179 5173
rect 13843 5145 14179 5172
rect 14149 5144 14179 5145
rect 14259 5136 14844 5144
rect 14259 5116 14268 5136
rect 14288 5135 14844 5136
rect 14288 5116 14808 5135
rect 14259 5115 14808 5116
rect 14828 5115 14844 5135
rect 14259 5109 14844 5115
rect 14083 5099 14115 5100
rect 14080 5094 14115 5099
rect 14080 5074 14087 5094
rect 14107 5074 14115 5094
rect 14878 5088 14912 5294
rect 14080 5066 14115 5074
rect 12084 5053 12119 5061
rect 12084 5033 12092 5053
rect 12112 5033 12119 5053
rect 12084 5028 12119 5033
rect 12084 5027 12116 5028
rect 11050 5018 11635 5024
rect 11050 4998 11066 5018
rect 11086 5017 11635 5018
rect 11086 4998 11606 5017
rect 11050 4997 11606 4998
rect 11626 4997 11635 5017
rect 11050 4989 11635 4997
rect 13462 4908 14047 4916
rect 13462 4888 13471 4908
rect 13491 4907 14047 4908
rect 13491 4888 14011 4907
rect 13462 4887 14011 4888
rect 14031 4887 14047 4907
rect 13462 4881 14047 4887
rect 13836 4857 13875 4861
rect 14081 4860 14115 5066
rect 14645 5078 14679 5086
rect 14645 5060 14652 5078
rect 14671 5060 14679 5078
rect 14645 5053 14679 5060
rect 14856 5083 14912 5088
rect 14856 5063 14863 5083
rect 14883 5063 14912 5083
rect 14856 5056 14912 5063
rect 14856 5055 14891 5056
rect 14649 5023 14678 5053
rect 14649 5015 15031 5023
rect 14649 4996 15002 5015
rect 15023 4996 15031 5015
rect 14649 4991 15031 4996
rect 10982 4831 11019 4846
rect 10982 4811 10990 4831
rect 11010 4811 11019 4831
rect 10982 4808 11019 4811
rect 10796 4697 10833 4700
rect 10796 4677 10805 4697
rect 10825 4677 10833 4697
rect 10796 4662 10833 4677
rect 6771 4513 7153 4518
rect 6771 4494 6779 4513
rect 6800 4494 7153 4513
rect 6771 4486 7153 4494
rect 7124 4456 7153 4486
rect 6911 4453 6946 4454
rect 6890 4446 6946 4453
rect 6890 4426 6919 4446
rect 6939 4426 6946 4446
rect 6890 4421 6946 4426
rect 7123 4449 7157 4456
rect 7123 4431 7131 4449
rect 7150 4431 7157 4449
rect 7123 4423 7157 4431
rect 7687 4443 7721 4649
rect 7927 4648 7966 4652
rect 7755 4622 8340 4628
rect 7755 4602 7771 4622
rect 7791 4621 8340 4622
rect 7791 4602 8311 4621
rect 7755 4601 8311 4602
rect 8331 4601 8340 4621
rect 7755 4593 8340 4601
rect 10180 4511 10765 4519
rect 10180 4491 10189 4511
rect 10209 4510 10765 4511
rect 10209 4491 10729 4510
rect 10180 4490 10729 4491
rect 10749 4490 10765 4510
rect 10180 4484 10765 4490
rect 9699 4480 9731 4481
rect 9696 4475 9731 4480
rect 9696 4455 9703 4475
rect 9723 4455 9731 4475
rect 10799 4463 10833 4662
rect 10777 4458 10833 4463
rect 9696 4447 9731 4455
rect 7687 4435 7722 4443
rect 6890 4215 6924 4421
rect 7687 4415 7695 4435
rect 7715 4415 7722 4435
rect 7687 4410 7722 4415
rect 7687 4409 7719 4410
rect 6958 4394 7543 4400
rect 6958 4374 6974 4394
rect 6994 4393 7543 4394
rect 6994 4374 7514 4393
rect 6958 4373 7514 4374
rect 7534 4373 7543 4393
rect 6958 4365 7543 4373
rect 7623 4364 7653 4365
rect 7623 4337 7959 4364
rect 7623 4336 7658 4337
rect 6890 4207 6925 4215
rect 6890 4187 6898 4207
rect 6918 4187 6925 4207
rect 6890 4182 6925 4187
rect 6890 4161 6924 4182
rect 7623 4161 7653 4336
rect 7709 4269 7744 4270
rect 6890 4135 7653 4161
rect 6891 4134 6924 4135
rect 7623 4133 7653 4135
rect 7688 4262 7744 4269
rect 7688 4242 7717 4262
rect 7737 4242 7744 4262
rect 7688 4237 7744 4242
rect 7923 4264 7958 4337
rect 7923 4244 7930 4264
rect 7950 4244 7958 4264
rect 9078 4289 9663 4297
rect 9078 4269 9087 4289
rect 9107 4288 9663 4289
rect 9107 4269 9627 4288
rect 9078 4268 9627 4269
rect 9647 4268 9663 4288
rect 9078 4262 9663 4268
rect 7923 4237 7958 4244
rect 9697 4241 9731 4447
rect 10559 4456 10594 4458
rect 10559 4450 10597 4456
rect 10559 4427 10567 4450
rect 10590 4427 10597 4450
rect 10777 4438 10784 4458
rect 10804 4438 10833 4458
rect 10777 4431 10833 4438
rect 10777 4430 10812 4431
rect 10559 4421 10597 4427
rect 10559 4408 10594 4421
rect 10557 4350 10594 4408
rect 6713 4112 6745 4113
rect 6713 4107 7053 4112
rect 6713 4089 6716 4107
rect 6738 4089 7053 4107
rect 6713 4084 7053 4089
rect 6713 4083 6745 4084
rect 7027 4049 7053 4084
rect 6812 4043 6847 4044
rect 6791 4036 6847 4043
rect 6791 4016 6820 4036
rect 6840 4016 6847 4036
rect 6791 4011 6847 4016
rect 7023 4040 7059 4049
rect 7023 4023 7031 4040
rect 7050 4023 7059 4040
rect 7023 4014 7059 4023
rect 7688 4031 7722 4237
rect 9461 4234 9496 4241
rect 7756 4210 8341 4216
rect 7756 4190 7772 4210
rect 7792 4209 8341 4210
rect 7792 4190 8312 4209
rect 7756 4189 8312 4190
rect 8332 4189 8341 4209
rect 7756 4181 8341 4189
rect 9461 4214 9469 4234
rect 9489 4214 9496 4234
rect 9461 4141 9496 4214
rect 9675 4236 9731 4241
rect 9675 4216 9682 4236
rect 9702 4216 9731 4236
rect 9675 4209 9731 4216
rect 9766 4343 9796 4345
rect 10495 4343 10528 4344
rect 9766 4317 10529 4343
rect 9675 4208 9710 4209
rect 9766 4142 9796 4317
rect 10495 4296 10529 4317
rect 10557 4333 10592 4350
rect 10557 4332 10851 4333
rect 10557 4331 10894 4332
rect 10557 4324 10899 4331
rect 10557 4298 10859 4324
rect 10890 4298 10899 4324
rect 10494 4291 10529 4296
rect 10850 4295 10899 4298
rect 10494 4271 10501 4291
rect 10521 4271 10529 4291
rect 10856 4290 10899 4295
rect 10494 4263 10529 4271
rect 9761 4141 9796 4142
rect 9460 4114 9796 4141
rect 9766 4113 9796 4114
rect 9876 4105 10461 4113
rect 9876 4085 9885 4105
rect 9905 4104 10461 4105
rect 9905 4085 10425 4104
rect 9876 4084 10425 4085
rect 10445 4084 10461 4104
rect 9876 4078 10461 4084
rect 9700 4068 9732 4069
rect 9697 4063 9732 4068
rect 9697 4043 9704 4063
rect 9724 4043 9732 4063
rect 10495 4057 10529 4263
rect 9697 4035 9732 4043
rect 7688 4023 7723 4031
rect 6791 3805 6825 4011
rect 7688 4003 7696 4023
rect 7716 4003 7723 4023
rect 7688 3998 7723 4003
rect 7688 3997 7720 3998
rect 6859 3984 7444 3990
rect 6859 3964 6875 3984
rect 6895 3983 7444 3984
rect 6895 3964 7415 3983
rect 6859 3963 7415 3964
rect 7435 3963 7444 3983
rect 6859 3955 7444 3963
rect 9079 3877 9664 3885
rect 9079 3857 9088 3877
rect 9108 3876 9664 3877
rect 9108 3857 9628 3876
rect 9079 3856 9628 3857
rect 9648 3856 9664 3876
rect 9079 3850 9664 3856
rect 9453 3826 9492 3830
rect 9698 3829 9732 4035
rect 10261 4050 10296 4056
rect 10261 4031 10266 4050
rect 10287 4031 10296 4050
rect 10261 4022 10296 4031
rect 10473 4052 10529 4057
rect 10473 4032 10480 4052
rect 10500 4032 10529 4052
rect 10473 4025 10529 4032
rect 10473 4024 10508 4025
rect 10265 3954 10294 4022
rect 10265 3920 10611 3954
rect 9453 3806 9461 3826
rect 9481 3806 9492 3826
rect 6791 3797 6826 3805
rect 6791 3777 6799 3797
rect 6819 3789 6826 3797
rect 6819 3777 6830 3789
rect 6791 3540 6830 3777
rect 7661 3754 7947 3755
rect 7146 3746 7949 3754
rect 7146 3729 7157 3746
rect 7147 3724 7157 3729
rect 7181 3729 7949 3746
rect 7181 3724 7186 3729
rect 7147 3711 7186 3724
rect 7691 3663 7726 3664
rect 7670 3656 7726 3663
rect 7670 3636 7699 3656
rect 7719 3636 7726 3656
rect 7670 3631 7726 3636
rect 7910 3654 7949 3729
rect 9453 3731 9492 3806
rect 9676 3824 9732 3829
rect 9676 3804 9683 3824
rect 9703 3804 9732 3824
rect 9676 3797 9732 3804
rect 9676 3796 9711 3797
rect 10216 3736 10255 3749
rect 10216 3731 10221 3736
rect 9453 3714 10221 3731
rect 10245 3731 10255 3736
rect 10245 3714 10256 3731
rect 9453 3706 10256 3714
rect 9455 3705 9741 3706
rect 10572 3683 10611 3920
rect 10572 3671 10583 3683
rect 10576 3663 10583 3671
rect 10603 3663 10611 3683
rect 10576 3655 10611 3663
rect 7910 3634 7921 3654
rect 7941 3634 7949 3654
rect 6791 3506 7137 3540
rect 7108 3438 7137 3506
rect 6894 3435 6929 3436
rect 6873 3428 6929 3435
rect 6873 3408 6902 3428
rect 6922 3408 6929 3428
rect 6873 3403 6929 3408
rect 7106 3429 7141 3438
rect 7106 3410 7115 3429
rect 7136 3410 7141 3429
rect 7106 3404 7141 3410
rect 7670 3425 7704 3631
rect 7910 3630 7949 3634
rect 7738 3604 8323 3610
rect 7738 3584 7754 3604
rect 7774 3603 8323 3604
rect 7774 3584 8294 3603
rect 7738 3583 8294 3584
rect 8314 3583 8323 3603
rect 7738 3575 8323 3583
rect 9958 3497 10543 3505
rect 9958 3477 9967 3497
rect 9987 3496 10543 3497
rect 9987 3477 10507 3496
rect 9958 3476 10507 3477
rect 10527 3476 10543 3496
rect 9958 3470 10543 3476
rect 9682 3462 9714 3463
rect 9679 3457 9714 3462
rect 9679 3437 9686 3457
rect 9706 3437 9714 3457
rect 10577 3449 10611 3655
rect 9679 3429 9714 3437
rect 7670 3417 7705 3425
rect 6873 3197 6907 3403
rect 7670 3397 7678 3417
rect 7698 3397 7705 3417
rect 7670 3392 7705 3397
rect 7670 3391 7702 3392
rect 6941 3376 7526 3382
rect 6941 3356 6957 3376
rect 6977 3375 7526 3376
rect 6977 3356 7497 3375
rect 6941 3355 7497 3356
rect 7517 3355 7526 3375
rect 6941 3347 7526 3355
rect 7606 3346 7636 3347
rect 7606 3319 7942 3346
rect 7606 3318 7641 3319
rect 6873 3189 6908 3197
rect 6873 3169 6881 3189
rect 6901 3169 6908 3189
rect 6873 3164 6908 3169
rect 6873 3143 6907 3164
rect 7606 3143 7636 3318
rect 7692 3251 7727 3252
rect 6873 3117 7636 3143
rect 6874 3116 6907 3117
rect 7606 3115 7636 3117
rect 7671 3244 7727 3251
rect 7671 3224 7700 3244
rect 7720 3224 7727 3244
rect 7671 3219 7727 3224
rect 7906 3246 7941 3319
rect 7906 3226 7913 3246
rect 7933 3226 7941 3246
rect 9061 3271 9646 3279
rect 9061 3251 9070 3271
rect 9090 3270 9646 3271
rect 9090 3251 9610 3270
rect 9061 3250 9610 3251
rect 9630 3250 9646 3270
rect 9061 3244 9646 3250
rect 7906 3219 7941 3226
rect 9680 3223 9714 3429
rect 10345 3443 10376 3449
rect 10345 3424 10350 3443
rect 10371 3424 10376 3443
rect 10345 3382 10376 3424
rect 10555 3444 10611 3449
rect 10555 3424 10562 3444
rect 10582 3424 10611 3444
rect 10555 3417 10611 3424
rect 10555 3416 10590 3417
rect 10345 3354 10684 3382
rect 6615 3060 6969 3096
rect 6631 3059 6969 3060
rect 6943 3029 6969 3059
rect 6729 3027 6764 3028
rect 6708 3020 6764 3027
rect 6708 3000 6737 3020
rect 6757 3000 6764 3020
rect 6708 2995 6764 3000
rect 6937 3021 6978 3029
rect 6937 3003 6950 3021
rect 6968 3003 6978 3021
rect 6708 2789 6742 2995
rect 6937 2992 6978 3003
rect 7671 3013 7705 3219
rect 9444 3216 9479 3223
rect 7739 3192 8324 3198
rect 7739 3172 7755 3192
rect 7775 3191 8324 3192
rect 7775 3172 8295 3191
rect 7739 3171 8295 3172
rect 8315 3171 8324 3191
rect 7739 3163 8324 3171
rect 9444 3196 9452 3216
rect 9472 3196 9479 3216
rect 9444 3123 9479 3196
rect 9658 3218 9714 3223
rect 9658 3198 9665 3218
rect 9685 3198 9714 3218
rect 9658 3191 9714 3198
rect 9749 3325 9779 3327
rect 10478 3325 10511 3326
rect 9749 3299 10512 3325
rect 9658 3190 9693 3191
rect 9749 3124 9779 3299
rect 10478 3278 10512 3299
rect 10477 3273 10512 3278
rect 10477 3253 10484 3273
rect 10504 3253 10512 3273
rect 10477 3245 10512 3253
rect 9744 3123 9779 3124
rect 9443 3096 9779 3123
rect 9749 3095 9779 3096
rect 9859 3087 10444 3095
rect 9859 3067 9868 3087
rect 9888 3086 10444 3087
rect 9888 3067 10408 3086
rect 9859 3066 10408 3067
rect 10428 3066 10444 3086
rect 9859 3060 10444 3066
rect 9683 3050 9715 3051
rect 9680 3045 9715 3050
rect 9680 3025 9687 3045
rect 9707 3025 9715 3045
rect 10478 3039 10512 3245
rect 9680 3017 9715 3025
rect 7671 3005 7706 3013
rect 7671 2985 7679 3005
rect 7699 2985 7706 3005
rect 7671 2980 7706 2985
rect 7671 2979 7703 2980
rect 6776 2968 7361 2974
rect 6776 2948 6792 2968
rect 6812 2967 7361 2968
rect 6812 2948 7332 2967
rect 6776 2947 7332 2948
rect 7352 2947 7361 2967
rect 6776 2939 7361 2947
rect 9062 2859 9647 2867
rect 9062 2839 9071 2859
rect 9091 2858 9647 2859
rect 9091 2839 9611 2858
rect 9062 2838 9611 2839
rect 9631 2838 9647 2858
rect 9062 2832 9647 2838
rect 9436 2808 9475 2812
rect 9681 2811 9715 3017
rect 10245 3029 10279 3037
rect 10245 3011 10252 3029
rect 10271 3011 10279 3029
rect 10245 3004 10279 3011
rect 10456 3034 10512 3039
rect 10456 3014 10463 3034
rect 10483 3014 10512 3034
rect 10456 3007 10512 3014
rect 10456 3006 10491 3007
rect 10249 2974 10278 3004
rect 10249 2966 10631 2974
rect 10249 2947 10602 2966
rect 10623 2947 10631 2966
rect 10249 2942 10631 2947
rect 6708 2788 6743 2789
rect 6676 2781 6743 2788
rect 6676 2761 6716 2781
rect 6736 2761 6743 2781
rect 6676 2758 6743 2761
rect 9436 2788 9444 2808
rect 9464 2788 9475 2808
rect 6676 2755 6741 2758
rect 6247 2654 6312 2657
rect 6245 2651 6312 2654
rect 6245 2631 6252 2651
rect 6272 2631 6312 2651
rect 6245 2624 6312 2631
rect 6245 2623 6280 2624
rect 3526 2603 3537 2623
rect 3557 2603 3565 2623
rect 2370 2464 2752 2469
rect 2370 2445 2378 2464
rect 2399 2445 2752 2464
rect 2370 2437 2752 2445
rect 2723 2407 2752 2437
rect 2510 2404 2545 2405
rect 2489 2397 2545 2404
rect 2489 2377 2518 2397
rect 2538 2377 2545 2397
rect 2489 2372 2545 2377
rect 2722 2400 2756 2407
rect 2722 2382 2730 2400
rect 2749 2382 2756 2400
rect 2722 2374 2756 2382
rect 3286 2394 3320 2600
rect 3526 2599 3565 2603
rect 3354 2573 3939 2579
rect 3354 2553 3370 2573
rect 3390 2572 3939 2573
rect 3390 2553 3910 2572
rect 3354 2552 3910 2553
rect 3930 2552 3939 2572
rect 3354 2544 3939 2552
rect 5627 2465 6212 2473
rect 5627 2445 5636 2465
rect 5656 2464 6212 2465
rect 5656 2445 6176 2464
rect 5627 2444 6176 2445
rect 6196 2444 6212 2464
rect 5627 2438 6212 2444
rect 5285 2432 5317 2433
rect 5282 2427 5317 2432
rect 5282 2407 5289 2427
rect 5309 2407 5317 2427
rect 5282 2399 5317 2407
rect 3286 2386 3321 2394
rect 2489 2166 2523 2372
rect 3286 2366 3294 2386
rect 3314 2366 3321 2386
rect 3286 2361 3321 2366
rect 3286 2360 3318 2361
rect 2557 2345 3142 2351
rect 2557 2325 2573 2345
rect 2593 2344 3142 2345
rect 2593 2325 3113 2344
rect 2557 2324 3113 2325
rect 3133 2324 3142 2344
rect 2557 2316 3142 2324
rect 3222 2315 3252 2316
rect 3222 2288 3558 2315
rect 3222 2287 3257 2288
rect 2489 2158 2524 2166
rect 2489 2138 2497 2158
rect 2517 2138 2524 2158
rect 2489 2133 2524 2138
rect 2489 2112 2523 2133
rect 3222 2112 3252 2287
rect 3308 2220 3343 2221
rect 2489 2086 3252 2112
rect 2490 2085 2523 2086
rect 3222 2084 3252 2086
rect 3287 2213 3343 2220
rect 3287 2193 3316 2213
rect 3336 2193 3343 2213
rect 3287 2188 3343 2193
rect 3522 2215 3557 2288
rect 3522 2195 3529 2215
rect 3549 2195 3557 2215
rect 4664 2241 5249 2249
rect 4664 2221 4673 2241
rect 4693 2240 5249 2241
rect 4693 2221 5213 2240
rect 4664 2220 5213 2221
rect 5233 2220 5249 2240
rect 4664 2214 5249 2220
rect 3522 2188 3557 2195
rect 5283 2193 5317 2399
rect 6012 2414 6045 2420
rect 6246 2417 6280 2623
rect 6012 2392 6017 2414
rect 6040 2392 6045 2414
rect 6012 2383 6045 2392
rect 6224 2412 6280 2417
rect 6224 2392 6231 2412
rect 6251 2392 6280 2412
rect 6224 2385 6280 2392
rect 6224 2384 6259 2385
rect 6014 2352 6041 2383
rect 6436 2352 6475 2364
rect 6014 2351 6477 2352
rect 6014 2329 6441 2351
rect 6465 2329 6477 2351
rect 6014 2321 6477 2329
rect 2317 2029 2656 2057
rect 2411 1994 2446 1995
rect 2390 1987 2446 1994
rect 2390 1967 2419 1987
rect 2439 1967 2446 1987
rect 2390 1962 2446 1967
rect 2625 1987 2656 2029
rect 2625 1968 2630 1987
rect 2651 1968 2656 1987
rect 2625 1962 2656 1968
rect 3287 1982 3321 2188
rect 5047 2186 5082 2193
rect 3355 2161 3940 2167
rect 3355 2141 3371 2161
rect 3391 2160 3940 2161
rect 3391 2141 3911 2160
rect 3355 2140 3911 2141
rect 3931 2140 3940 2160
rect 3355 2132 3940 2140
rect 5047 2166 5055 2186
rect 5075 2166 5082 2186
rect 5047 2093 5082 2166
rect 5261 2188 5317 2193
rect 5261 2168 5268 2188
rect 5288 2168 5317 2188
rect 5261 2161 5317 2168
rect 5352 2295 5382 2297
rect 6081 2295 6114 2296
rect 5352 2269 6115 2295
rect 5261 2160 5296 2161
rect 5352 2094 5382 2269
rect 6081 2248 6115 2269
rect 6080 2243 6115 2248
rect 6080 2223 6087 2243
rect 6107 2223 6115 2243
rect 6080 2215 6115 2223
rect 5347 2093 5382 2094
rect 5046 2066 5382 2093
rect 5352 2065 5382 2066
rect 5462 2057 6047 2065
rect 5462 2037 5471 2057
rect 5491 2056 6047 2057
rect 5491 2037 6011 2056
rect 5462 2036 6011 2037
rect 6031 2036 6047 2056
rect 5462 2030 6047 2036
rect 5286 2020 5318 2021
rect 5283 2015 5318 2020
rect 5283 1995 5290 2015
rect 5310 1995 5318 2015
rect 6081 2009 6115 2215
rect 5283 1987 5318 1995
rect 3287 1974 3322 1982
rect 2390 1756 2424 1962
rect 3287 1954 3295 1974
rect 3315 1954 3322 1974
rect 3287 1949 3322 1954
rect 3287 1948 3319 1949
rect 2458 1935 3043 1941
rect 2458 1915 2474 1935
rect 2494 1934 3043 1935
rect 2494 1915 3014 1934
rect 2458 1914 3014 1915
rect 3034 1914 3043 1934
rect 2458 1906 3043 1914
rect 4665 1829 5250 1837
rect 4665 1809 4674 1829
rect 4694 1828 5250 1829
rect 4694 1809 5214 1828
rect 4665 1808 5214 1809
rect 5234 1808 5250 1828
rect 4665 1802 5250 1808
rect 5039 1778 5078 1782
rect 5284 1781 5318 1987
rect 5847 2002 5882 2008
rect 5847 1983 5852 2002
rect 5873 1983 5882 2002
rect 5847 1974 5882 1983
rect 6059 2004 6115 2009
rect 6059 1984 6066 2004
rect 6086 1984 6115 2004
rect 6059 1977 6115 1984
rect 6237 2155 6269 2167
rect 6237 2137 6244 2155
rect 6266 2137 6269 2155
rect 6059 1976 6094 1977
rect 5851 1906 5880 1974
rect 5851 1872 6197 1906
rect 5039 1758 5047 1778
rect 5067 1758 5078 1778
rect 2390 1748 2425 1756
rect 2390 1728 2398 1748
rect 2418 1740 2425 1748
rect 2418 1728 2429 1740
rect 2390 1491 2429 1728
rect 3260 1705 3546 1706
rect 2745 1697 3548 1705
rect 2745 1680 2756 1697
rect 2746 1675 2756 1680
rect 2780 1680 3548 1697
rect 2780 1675 2785 1680
rect 2746 1662 2785 1675
rect 3290 1614 3325 1615
rect 3269 1607 3325 1614
rect 3269 1587 3298 1607
rect 3318 1587 3325 1607
rect 3269 1582 3325 1587
rect 3509 1605 3548 1680
rect 5039 1683 5078 1758
rect 5262 1776 5318 1781
rect 5262 1756 5269 1776
rect 5289 1756 5318 1776
rect 5262 1749 5318 1756
rect 5262 1748 5297 1749
rect 5802 1688 5841 1701
rect 5802 1683 5807 1688
rect 5039 1666 5807 1683
rect 5831 1683 5841 1688
rect 5831 1666 5842 1683
rect 5039 1658 5842 1666
rect 5041 1657 5327 1658
rect 6158 1635 6197 1872
rect 6158 1623 6169 1635
rect 6162 1615 6169 1623
rect 6189 1615 6197 1635
rect 6162 1607 6197 1615
rect 3509 1585 3520 1605
rect 3540 1585 3548 1605
rect 2390 1457 2736 1491
rect 2707 1389 2736 1457
rect 2493 1386 2528 1387
rect 1571 1287 1905 1315
rect 2472 1379 2528 1386
rect 2472 1359 2501 1379
rect 2521 1359 2528 1379
rect 2472 1354 2528 1359
rect 2705 1380 2740 1389
rect 2705 1361 2714 1380
rect 2735 1361 2740 1380
rect 2705 1355 2740 1361
rect 3269 1376 3303 1582
rect 3509 1581 3548 1585
rect 3337 1555 3922 1561
rect 3337 1535 3353 1555
rect 3373 1554 3922 1555
rect 3373 1535 3893 1554
rect 3337 1534 3893 1535
rect 3913 1534 3922 1554
rect 3337 1526 3922 1534
rect 5544 1449 6129 1457
rect 5544 1429 5553 1449
rect 5573 1448 6129 1449
rect 5573 1429 6093 1448
rect 5544 1428 6093 1429
rect 6113 1428 6129 1448
rect 5544 1422 6129 1428
rect 5268 1414 5300 1415
rect 5265 1409 5300 1414
rect 5265 1389 5272 1409
rect 5292 1389 5300 1409
rect 6163 1401 6197 1607
rect 5265 1381 5300 1389
rect 3269 1368 3304 1376
rect 666 1155 701 1162
rect 666 1135 674 1155
rect 694 1135 701 1155
rect 666 1062 701 1135
rect 880 1157 936 1162
rect 880 1137 887 1157
rect 907 1137 936 1157
rect 880 1130 936 1137
rect 971 1264 1001 1266
rect 1700 1264 1733 1265
rect 971 1238 1734 1264
rect 880 1129 915 1130
rect 971 1063 1001 1238
rect 1700 1217 1734 1238
rect 1699 1212 1734 1217
rect 1699 1192 1706 1212
rect 1726 1192 1734 1212
rect 1699 1184 1734 1192
rect 966 1062 1001 1063
rect 665 1035 1001 1062
rect 971 1034 1001 1035
rect 1081 1026 1666 1034
rect 1081 1006 1090 1026
rect 1110 1025 1666 1026
rect 1110 1006 1630 1025
rect 1081 1005 1630 1006
rect 1650 1005 1666 1025
rect 1081 999 1666 1005
rect 905 989 937 990
rect 902 984 937 989
rect 902 964 909 984
rect 929 964 937 984
rect 1700 978 1734 1184
rect 2472 1148 2506 1354
rect 3269 1348 3277 1368
rect 3297 1348 3304 1368
rect 3269 1343 3304 1348
rect 3269 1342 3301 1343
rect 2540 1327 3125 1333
rect 2540 1307 2556 1327
rect 2576 1326 3125 1327
rect 2576 1307 3096 1326
rect 2540 1306 3096 1307
rect 3116 1306 3125 1326
rect 2540 1298 3125 1306
rect 3205 1297 3235 1298
rect 3205 1270 3541 1297
rect 3205 1269 3240 1270
rect 2472 1140 2507 1148
rect 2472 1120 2480 1140
rect 2500 1120 2507 1140
rect 2472 1115 2507 1120
rect 2472 1094 2506 1115
rect 3205 1094 3235 1269
rect 3291 1202 3326 1203
rect 2472 1068 3235 1094
rect 2473 1067 2506 1068
rect 3205 1066 3235 1068
rect 3270 1195 3326 1202
rect 3270 1175 3299 1195
rect 3319 1175 3326 1195
rect 3270 1170 3326 1175
rect 3505 1197 3540 1270
rect 3505 1177 3512 1197
rect 3532 1177 3540 1197
rect 4647 1223 5232 1231
rect 4647 1203 4656 1223
rect 4676 1222 5232 1223
rect 4676 1203 5196 1222
rect 4647 1202 5196 1203
rect 5216 1202 5232 1222
rect 4647 1196 5232 1202
rect 3505 1170 3540 1177
rect 5266 1175 5300 1381
rect 5929 1389 5965 1398
rect 5929 1372 5938 1389
rect 5957 1372 5965 1389
rect 5929 1363 5965 1372
rect 6141 1396 6197 1401
rect 6141 1376 6148 1396
rect 6168 1376 6197 1396
rect 6141 1369 6197 1376
rect 6141 1368 6176 1369
rect 5935 1328 5961 1363
rect 6237 1328 6269 2137
rect 6681 2070 6710 2755
rect 7641 2736 7927 2737
rect 7126 2728 7929 2736
rect 7126 2711 7137 2728
rect 7127 2706 7137 2711
rect 7161 2711 7929 2728
rect 7161 2706 7166 2711
rect 7127 2693 7166 2706
rect 7671 2645 7706 2646
rect 7650 2638 7706 2645
rect 7650 2618 7679 2638
rect 7699 2618 7706 2638
rect 7650 2613 7706 2618
rect 7890 2636 7929 2711
rect 9436 2713 9475 2788
rect 9659 2806 9715 2811
rect 9659 2786 9666 2806
rect 9686 2786 9715 2806
rect 9659 2779 9715 2786
rect 9659 2778 9694 2779
rect 10199 2718 10238 2731
rect 10199 2713 10204 2718
rect 9436 2696 10204 2713
rect 10228 2713 10238 2718
rect 10228 2696 10239 2713
rect 9436 2688 10239 2696
rect 9438 2687 9724 2688
rect 10655 2669 10684 3354
rect 10992 3108 11019 4808
rect 13836 4837 13844 4857
rect 13864 4837 13875 4857
rect 12055 4784 12341 4785
rect 11540 4776 12343 4784
rect 11540 4759 11551 4776
rect 11541 4754 11551 4759
rect 11575 4759 12343 4776
rect 11575 4754 11580 4759
rect 11541 4741 11580 4754
rect 12085 4693 12120 4694
rect 12064 4686 12120 4693
rect 12064 4666 12093 4686
rect 12113 4666 12120 4686
rect 12064 4661 12120 4666
rect 12304 4684 12343 4759
rect 13836 4762 13875 4837
rect 14059 4855 14115 4860
rect 14059 4835 14066 4855
rect 14086 4835 14115 4855
rect 14059 4828 14115 4835
rect 14059 4827 14094 4828
rect 14599 4767 14638 4780
rect 14599 4762 14604 4767
rect 13836 4745 14604 4762
rect 14628 4762 14638 4767
rect 14628 4745 14639 4762
rect 13836 4737 14639 4745
rect 13838 4736 14124 4737
rect 12304 4664 12315 4684
rect 12335 4664 12343 4684
rect 15160 4713 15187 6413
rect 15495 6167 15524 6852
rect 16455 6833 16741 6834
rect 15940 6825 16743 6833
rect 15940 6808 15951 6825
rect 15941 6803 15951 6808
rect 15975 6808 16743 6825
rect 15975 6803 15980 6808
rect 15941 6790 15980 6803
rect 16485 6742 16520 6743
rect 16464 6735 16520 6742
rect 16464 6715 16493 6735
rect 16513 6715 16520 6735
rect 16464 6710 16520 6715
rect 16704 6733 16743 6808
rect 16704 6713 16715 6733
rect 16735 6713 16743 6733
rect 15548 6574 15930 6579
rect 15548 6555 15556 6574
rect 15577 6555 15930 6574
rect 15548 6547 15930 6555
rect 15901 6517 15930 6547
rect 15688 6514 15723 6515
rect 15667 6507 15723 6514
rect 15667 6487 15696 6507
rect 15716 6487 15723 6507
rect 15667 6482 15723 6487
rect 15900 6510 15934 6517
rect 15900 6492 15908 6510
rect 15927 6492 15934 6510
rect 15900 6484 15934 6492
rect 16464 6504 16498 6710
rect 16704 6709 16743 6713
rect 16532 6683 17117 6689
rect 16532 6663 16548 6683
rect 16568 6682 17117 6683
rect 16568 6663 17088 6682
rect 16532 6662 17088 6663
rect 17108 6662 17117 6682
rect 16532 6654 17117 6662
rect 16464 6496 16499 6504
rect 15667 6276 15701 6482
rect 16464 6476 16472 6496
rect 16492 6476 16499 6496
rect 16464 6471 16499 6476
rect 16464 6470 16496 6471
rect 15735 6455 16320 6461
rect 15735 6435 15751 6455
rect 15771 6454 16320 6455
rect 15771 6435 16291 6454
rect 15735 6434 16291 6435
rect 16311 6434 16320 6454
rect 15735 6426 16320 6434
rect 16400 6425 16430 6426
rect 16400 6398 16736 6425
rect 16400 6397 16435 6398
rect 15667 6268 15702 6276
rect 15667 6248 15675 6268
rect 15695 6248 15702 6268
rect 15667 6243 15702 6248
rect 15667 6222 15701 6243
rect 16400 6222 16430 6397
rect 16486 6330 16521 6331
rect 15667 6196 16430 6222
rect 15668 6195 15701 6196
rect 16400 6194 16430 6196
rect 16465 6323 16521 6330
rect 16465 6303 16494 6323
rect 16514 6303 16521 6323
rect 16465 6298 16521 6303
rect 16700 6325 16735 6398
rect 16700 6305 16707 6325
rect 16727 6305 16735 6325
rect 16700 6298 16735 6305
rect 15495 6139 15834 6167
rect 15589 6104 15624 6105
rect 15568 6097 15624 6104
rect 15568 6077 15597 6097
rect 15617 6077 15624 6097
rect 15568 6072 15624 6077
rect 15803 6097 15834 6139
rect 15803 6078 15808 6097
rect 15829 6078 15834 6097
rect 15803 6072 15834 6078
rect 16465 6092 16499 6298
rect 16533 6271 17118 6277
rect 16533 6251 16549 6271
rect 16569 6270 17118 6271
rect 16569 6251 17089 6270
rect 16533 6250 17089 6251
rect 17109 6250 17118 6270
rect 16533 6242 17118 6250
rect 16465 6084 16500 6092
rect 15568 5866 15602 6072
rect 16465 6064 16473 6084
rect 16493 6064 16500 6084
rect 16465 6059 16500 6064
rect 16465 6058 16497 6059
rect 15636 6045 16221 6051
rect 15636 6025 15652 6045
rect 15672 6044 16221 6045
rect 15672 6025 16192 6044
rect 15636 6024 16192 6025
rect 16212 6024 16221 6044
rect 15636 6016 16221 6024
rect 15568 5858 15603 5866
rect 15568 5838 15576 5858
rect 15596 5850 15603 5858
rect 15596 5838 15607 5850
rect 15568 5601 15607 5838
rect 16438 5815 16724 5816
rect 15923 5807 16726 5815
rect 15923 5790 15934 5807
rect 15924 5785 15934 5790
rect 15958 5790 16726 5807
rect 15958 5785 15963 5790
rect 15924 5772 15963 5785
rect 16468 5724 16503 5725
rect 16447 5717 16503 5724
rect 16447 5697 16476 5717
rect 16496 5697 16503 5717
rect 16447 5692 16503 5697
rect 16687 5715 16726 5790
rect 16687 5695 16698 5715
rect 16718 5695 16726 5715
rect 15568 5567 15914 5601
rect 15885 5499 15914 5567
rect 15671 5496 15706 5497
rect 15650 5489 15706 5496
rect 15650 5469 15679 5489
rect 15699 5469 15706 5489
rect 15650 5464 15706 5469
rect 15883 5490 15918 5499
rect 15883 5471 15892 5490
rect 15913 5471 15918 5490
rect 15883 5465 15918 5471
rect 16447 5486 16481 5692
rect 16687 5691 16726 5695
rect 16515 5665 17100 5671
rect 16515 5645 16531 5665
rect 16551 5664 17100 5665
rect 16551 5645 17071 5664
rect 16515 5644 17071 5645
rect 17091 5644 17100 5664
rect 16515 5636 17100 5644
rect 16447 5478 16482 5486
rect 15650 5258 15684 5464
rect 16447 5458 16455 5478
rect 16475 5458 16482 5478
rect 16447 5453 16482 5458
rect 16447 5452 16479 5453
rect 15718 5437 16303 5443
rect 15718 5417 15734 5437
rect 15754 5436 16303 5437
rect 15754 5417 16274 5436
rect 15718 5416 16274 5417
rect 16294 5416 16303 5436
rect 15718 5408 16303 5416
rect 16383 5407 16413 5408
rect 16383 5380 16719 5407
rect 16383 5379 16418 5380
rect 15650 5250 15685 5258
rect 15650 5230 15658 5250
rect 15678 5230 15685 5250
rect 15650 5225 15685 5230
rect 15650 5204 15684 5225
rect 16383 5204 16413 5379
rect 16469 5312 16504 5313
rect 15650 5178 16413 5204
rect 15651 5177 15684 5178
rect 16383 5176 16413 5178
rect 16448 5305 16504 5312
rect 16448 5285 16477 5305
rect 16497 5285 16504 5305
rect 16448 5280 16504 5285
rect 16683 5307 16718 5380
rect 16683 5287 16690 5307
rect 16710 5287 16718 5307
rect 16683 5280 16718 5287
rect 15302 5157 15619 5160
rect 15302 5130 15305 5157
rect 15332 5130 15619 5157
rect 15302 5124 15619 5130
rect 15302 5121 15338 5124
rect 15583 5094 15619 5124
rect 15367 5090 15402 5091
rect 15346 5083 15402 5090
rect 15346 5063 15375 5083
rect 15395 5063 15402 5083
rect 15346 5058 15402 5063
rect 15581 5088 15619 5094
rect 15581 5062 15587 5088
rect 15613 5062 15619 5088
rect 15346 4859 15380 5058
rect 15581 5054 15619 5062
rect 16448 5074 16482 5280
rect 16516 5253 17101 5259
rect 16516 5233 16532 5253
rect 16552 5252 17101 5253
rect 16552 5233 17072 5252
rect 16516 5232 17072 5233
rect 17092 5232 17101 5252
rect 16516 5224 17101 5232
rect 16448 5066 16483 5074
rect 16448 5046 16456 5066
rect 16476 5046 16483 5066
rect 16448 5041 16483 5046
rect 16448 5040 16480 5041
rect 15414 5031 15999 5037
rect 15414 5011 15430 5031
rect 15450 5030 15999 5031
rect 15450 5011 15970 5030
rect 15414 5010 15970 5011
rect 15990 5010 15999 5030
rect 15414 5002 15999 5010
rect 15346 4844 15383 4859
rect 15346 4824 15354 4844
rect 15374 4824 15383 4844
rect 15346 4821 15383 4824
rect 15160 4710 15197 4713
rect 15160 4690 15169 4710
rect 15189 4690 15197 4710
rect 15160 4675 15197 4690
rect 11148 4525 11530 4530
rect 11148 4506 11156 4525
rect 11177 4506 11530 4525
rect 11148 4498 11530 4506
rect 11501 4468 11530 4498
rect 11288 4465 11323 4466
rect 11267 4458 11323 4465
rect 11267 4438 11296 4458
rect 11316 4438 11323 4458
rect 11267 4433 11323 4438
rect 11500 4461 11534 4468
rect 11500 4443 11508 4461
rect 11527 4443 11534 4461
rect 11500 4435 11534 4443
rect 12064 4455 12098 4661
rect 12304 4660 12343 4664
rect 12132 4634 12717 4640
rect 12132 4614 12148 4634
rect 12168 4633 12717 4634
rect 12168 4614 12688 4633
rect 12132 4613 12688 4614
rect 12708 4613 12717 4633
rect 12132 4605 12717 4613
rect 14544 4524 15129 4532
rect 14544 4504 14553 4524
rect 14573 4523 15129 4524
rect 14573 4504 15093 4523
rect 14544 4503 15093 4504
rect 15113 4503 15129 4523
rect 14544 4497 15129 4503
rect 14063 4493 14095 4494
rect 14060 4488 14095 4493
rect 14060 4468 14067 4488
rect 14087 4468 14095 4488
rect 15163 4476 15197 4675
rect 15141 4471 15197 4476
rect 14060 4460 14095 4468
rect 12064 4447 12099 4455
rect 11267 4227 11301 4433
rect 12064 4427 12072 4447
rect 12092 4427 12099 4447
rect 12064 4422 12099 4427
rect 12064 4421 12096 4422
rect 11335 4406 11920 4412
rect 11335 4386 11351 4406
rect 11371 4405 11920 4406
rect 11371 4386 11891 4405
rect 11335 4385 11891 4386
rect 11911 4385 11920 4405
rect 11335 4377 11920 4385
rect 12000 4376 12030 4377
rect 12000 4349 12336 4376
rect 12000 4348 12035 4349
rect 11267 4219 11302 4227
rect 11267 4199 11275 4219
rect 11295 4199 11302 4219
rect 11267 4194 11302 4199
rect 11267 4173 11301 4194
rect 12000 4173 12030 4348
rect 12086 4281 12121 4282
rect 11267 4147 12030 4173
rect 11268 4146 11301 4147
rect 12000 4145 12030 4147
rect 12065 4274 12121 4281
rect 12065 4254 12094 4274
rect 12114 4254 12121 4274
rect 12065 4249 12121 4254
rect 12300 4276 12335 4349
rect 12300 4256 12307 4276
rect 12327 4256 12335 4276
rect 13442 4302 14027 4310
rect 13442 4282 13451 4302
rect 13471 4301 14027 4302
rect 13471 4282 13991 4301
rect 13442 4281 13991 4282
rect 14011 4281 14027 4301
rect 13442 4275 14027 4281
rect 12300 4249 12335 4256
rect 14061 4254 14095 4460
rect 14923 4469 14958 4471
rect 14923 4463 14961 4469
rect 14923 4440 14931 4463
rect 14954 4440 14961 4463
rect 15141 4451 15148 4471
rect 15168 4451 15197 4471
rect 15141 4444 15197 4451
rect 15141 4443 15176 4444
rect 14923 4434 14961 4440
rect 14923 4421 14958 4434
rect 14921 4363 14958 4421
rect 11090 4124 11122 4125
rect 11090 4119 11430 4124
rect 11090 4101 11093 4119
rect 11115 4101 11430 4119
rect 11090 4096 11430 4101
rect 11090 4095 11122 4096
rect 11404 4061 11430 4096
rect 11189 4055 11224 4056
rect 11168 4048 11224 4055
rect 11168 4028 11197 4048
rect 11217 4028 11224 4048
rect 11168 4023 11224 4028
rect 11400 4052 11436 4061
rect 11400 4035 11408 4052
rect 11427 4035 11436 4052
rect 11400 4026 11436 4035
rect 12065 4043 12099 4249
rect 13825 4247 13860 4254
rect 12133 4222 12718 4228
rect 12133 4202 12149 4222
rect 12169 4221 12718 4222
rect 12169 4202 12689 4221
rect 12133 4201 12689 4202
rect 12709 4201 12718 4221
rect 12133 4193 12718 4201
rect 13825 4227 13833 4247
rect 13853 4227 13860 4247
rect 13825 4154 13860 4227
rect 14039 4249 14095 4254
rect 14039 4229 14046 4249
rect 14066 4229 14095 4249
rect 14039 4222 14095 4229
rect 14130 4356 14160 4358
rect 14859 4356 14892 4357
rect 14130 4330 14893 4356
rect 14039 4221 14074 4222
rect 14130 4155 14160 4330
rect 14859 4309 14893 4330
rect 14921 4346 14956 4363
rect 14921 4345 15215 4346
rect 14921 4344 15258 4345
rect 14921 4337 15263 4344
rect 14921 4311 15223 4337
rect 15254 4311 15263 4337
rect 14858 4304 14893 4309
rect 15214 4308 15263 4311
rect 14858 4284 14865 4304
rect 14885 4284 14893 4304
rect 15220 4303 15263 4308
rect 14858 4276 14893 4284
rect 14125 4154 14160 4155
rect 13824 4127 14160 4154
rect 14130 4126 14160 4127
rect 14240 4118 14825 4126
rect 14240 4098 14249 4118
rect 14269 4117 14825 4118
rect 14269 4098 14789 4117
rect 14240 4097 14789 4098
rect 14809 4097 14825 4117
rect 14240 4091 14825 4097
rect 14064 4081 14096 4082
rect 14061 4076 14096 4081
rect 14061 4056 14068 4076
rect 14088 4056 14096 4076
rect 14859 4070 14893 4276
rect 14061 4048 14096 4056
rect 12065 4035 12100 4043
rect 11168 3817 11202 4023
rect 12065 4015 12073 4035
rect 12093 4015 12100 4035
rect 12065 4010 12100 4015
rect 12065 4009 12097 4010
rect 11236 3996 11821 4002
rect 11236 3976 11252 3996
rect 11272 3995 11821 3996
rect 11272 3976 11792 3995
rect 11236 3975 11792 3976
rect 11812 3975 11821 3995
rect 11236 3967 11821 3975
rect 13443 3890 14028 3898
rect 13443 3870 13452 3890
rect 13472 3889 14028 3890
rect 13472 3870 13992 3889
rect 13443 3869 13992 3870
rect 14012 3869 14028 3889
rect 13443 3863 14028 3869
rect 13817 3839 13856 3843
rect 14062 3842 14096 4048
rect 14625 4063 14660 4069
rect 14625 4044 14630 4063
rect 14651 4044 14660 4063
rect 14625 4035 14660 4044
rect 14837 4065 14893 4070
rect 14837 4045 14844 4065
rect 14864 4045 14893 4065
rect 14837 4038 14893 4045
rect 14837 4037 14872 4038
rect 14629 3967 14658 4035
rect 14629 3933 14975 3967
rect 13817 3819 13825 3839
rect 13845 3819 13856 3839
rect 11168 3809 11203 3817
rect 11168 3789 11176 3809
rect 11196 3801 11203 3809
rect 11196 3789 11207 3801
rect 11168 3552 11207 3789
rect 12038 3766 12324 3767
rect 11523 3758 12326 3766
rect 11523 3741 11534 3758
rect 11524 3736 11534 3741
rect 11558 3741 12326 3758
rect 11558 3736 11563 3741
rect 11524 3723 11563 3736
rect 12068 3675 12103 3676
rect 12047 3668 12103 3675
rect 12047 3648 12076 3668
rect 12096 3648 12103 3668
rect 12047 3643 12103 3648
rect 12287 3666 12326 3741
rect 13817 3744 13856 3819
rect 14040 3837 14096 3842
rect 14040 3817 14047 3837
rect 14067 3817 14096 3837
rect 14040 3810 14096 3817
rect 14040 3809 14075 3810
rect 14580 3749 14619 3762
rect 14580 3744 14585 3749
rect 13817 3727 14585 3744
rect 14609 3744 14619 3749
rect 14609 3727 14620 3744
rect 13817 3719 14620 3727
rect 13819 3718 14105 3719
rect 14936 3696 14975 3933
rect 14936 3684 14947 3696
rect 14940 3676 14947 3684
rect 14967 3676 14975 3696
rect 14940 3668 14975 3676
rect 12287 3646 12298 3666
rect 12318 3646 12326 3666
rect 11168 3518 11514 3552
rect 11485 3450 11514 3518
rect 11271 3447 11306 3448
rect 11250 3440 11306 3447
rect 11250 3420 11279 3440
rect 11299 3420 11306 3440
rect 11250 3415 11306 3420
rect 11483 3441 11518 3450
rect 11483 3422 11492 3441
rect 11513 3422 11518 3441
rect 11483 3416 11518 3422
rect 12047 3437 12081 3643
rect 12287 3642 12326 3646
rect 12115 3616 12700 3622
rect 12115 3596 12131 3616
rect 12151 3615 12700 3616
rect 12151 3596 12671 3615
rect 12115 3595 12671 3596
rect 12691 3595 12700 3615
rect 12115 3587 12700 3595
rect 14322 3510 14907 3518
rect 14322 3490 14331 3510
rect 14351 3509 14907 3510
rect 14351 3490 14871 3509
rect 14322 3489 14871 3490
rect 14891 3489 14907 3509
rect 14322 3483 14907 3489
rect 14046 3475 14078 3476
rect 14043 3470 14078 3475
rect 14043 3450 14050 3470
rect 14070 3450 14078 3470
rect 14941 3462 14975 3668
rect 14043 3442 14078 3450
rect 12047 3429 12082 3437
rect 11250 3209 11284 3415
rect 12047 3409 12055 3429
rect 12075 3409 12082 3429
rect 12047 3404 12082 3409
rect 12047 3403 12079 3404
rect 11318 3388 11903 3394
rect 11318 3368 11334 3388
rect 11354 3387 11903 3388
rect 11354 3368 11874 3387
rect 11318 3367 11874 3368
rect 11894 3367 11903 3387
rect 11318 3359 11903 3367
rect 11983 3358 12013 3359
rect 11983 3331 12319 3358
rect 11983 3330 12018 3331
rect 11250 3201 11285 3209
rect 11250 3181 11258 3201
rect 11278 3181 11285 3201
rect 11250 3176 11285 3181
rect 11250 3155 11284 3176
rect 11983 3155 12013 3330
rect 12069 3263 12104 3264
rect 11250 3129 12013 3155
rect 11251 3128 11284 3129
rect 11983 3127 12013 3129
rect 12048 3256 12104 3263
rect 12048 3236 12077 3256
rect 12097 3236 12104 3256
rect 12048 3231 12104 3236
rect 12283 3258 12318 3331
rect 12283 3238 12290 3258
rect 12310 3238 12318 3258
rect 13425 3284 14010 3292
rect 13425 3264 13434 3284
rect 13454 3283 14010 3284
rect 13454 3264 13974 3283
rect 13425 3263 13974 3264
rect 13994 3263 14010 3283
rect 13425 3257 14010 3263
rect 12283 3231 12318 3238
rect 14044 3236 14078 3442
rect 14709 3456 14740 3462
rect 14709 3437 14714 3456
rect 14735 3437 14740 3456
rect 14709 3395 14740 3437
rect 14919 3457 14975 3462
rect 14919 3437 14926 3457
rect 14946 3437 14975 3457
rect 14919 3430 14975 3437
rect 14919 3429 14954 3430
rect 14709 3367 15048 3395
rect 10992 3072 11346 3108
rect 11008 3071 11346 3072
rect 11320 3041 11346 3071
rect 11106 3039 11141 3040
rect 11085 3032 11141 3039
rect 11085 3012 11114 3032
rect 11134 3012 11141 3032
rect 11085 3007 11141 3012
rect 11314 3033 11355 3041
rect 11314 3015 11327 3033
rect 11345 3015 11355 3033
rect 11085 2801 11119 3007
rect 11314 3004 11355 3015
rect 12048 3025 12082 3231
rect 13808 3229 13843 3236
rect 12116 3204 12701 3210
rect 12116 3184 12132 3204
rect 12152 3203 12701 3204
rect 12152 3184 12672 3203
rect 12116 3183 12672 3184
rect 12692 3183 12701 3203
rect 12116 3175 12701 3183
rect 13808 3209 13816 3229
rect 13836 3209 13843 3229
rect 13808 3136 13843 3209
rect 14022 3231 14078 3236
rect 14022 3211 14029 3231
rect 14049 3211 14078 3231
rect 14022 3204 14078 3211
rect 14113 3338 14143 3340
rect 14842 3338 14875 3339
rect 14113 3312 14876 3338
rect 14022 3203 14057 3204
rect 14113 3137 14143 3312
rect 14842 3291 14876 3312
rect 14841 3286 14876 3291
rect 14841 3266 14848 3286
rect 14868 3266 14876 3286
rect 14841 3258 14876 3266
rect 14108 3136 14143 3137
rect 13807 3109 14143 3136
rect 14113 3108 14143 3109
rect 14223 3100 14808 3108
rect 14223 3080 14232 3100
rect 14252 3099 14808 3100
rect 14252 3080 14772 3099
rect 14223 3079 14772 3080
rect 14792 3079 14808 3099
rect 14223 3073 14808 3079
rect 14047 3063 14079 3064
rect 14044 3058 14079 3063
rect 14044 3038 14051 3058
rect 14071 3038 14079 3058
rect 14842 3052 14876 3258
rect 14044 3030 14079 3038
rect 12048 3017 12083 3025
rect 12048 2997 12056 3017
rect 12076 2997 12083 3017
rect 12048 2992 12083 2997
rect 12048 2991 12080 2992
rect 11153 2980 11738 2986
rect 11153 2960 11169 2980
rect 11189 2979 11738 2980
rect 11189 2960 11709 2979
rect 11153 2959 11709 2960
rect 11729 2959 11738 2979
rect 11153 2951 11738 2959
rect 13426 2872 14011 2880
rect 13426 2852 13435 2872
rect 13455 2871 14011 2872
rect 13455 2852 13975 2871
rect 13426 2851 13975 2852
rect 13995 2851 14011 2871
rect 13426 2845 14011 2851
rect 13800 2821 13839 2825
rect 14045 2824 14079 3030
rect 14609 3042 14643 3050
rect 14609 3024 14616 3042
rect 14635 3024 14643 3042
rect 14609 3017 14643 3024
rect 14820 3047 14876 3052
rect 14820 3027 14827 3047
rect 14847 3027 14876 3047
rect 14820 3020 14876 3027
rect 14820 3019 14855 3020
rect 14613 2987 14642 3017
rect 14613 2979 14995 2987
rect 14613 2960 14966 2979
rect 14987 2960 14995 2979
rect 14613 2955 14995 2960
rect 13800 2801 13808 2821
rect 13828 2801 13839 2821
rect 11085 2800 11120 2801
rect 11053 2793 11120 2800
rect 11053 2773 11093 2793
rect 11113 2773 11120 2793
rect 11053 2770 11120 2773
rect 11053 2767 11118 2770
rect 10624 2666 10689 2669
rect 7890 2616 7901 2636
rect 7921 2616 7929 2636
rect 10622 2663 10689 2666
rect 10622 2643 10629 2663
rect 10649 2643 10689 2663
rect 10622 2636 10689 2643
rect 10622 2635 10657 2636
rect 6734 2477 7116 2482
rect 6734 2458 6742 2477
rect 6763 2458 7116 2477
rect 6734 2450 7116 2458
rect 7087 2420 7116 2450
rect 6874 2417 6909 2418
rect 6853 2410 6909 2417
rect 6853 2390 6882 2410
rect 6902 2390 6909 2410
rect 6853 2385 6909 2390
rect 7086 2413 7120 2420
rect 7086 2395 7094 2413
rect 7113 2395 7120 2413
rect 7086 2387 7120 2395
rect 7650 2407 7684 2613
rect 7890 2612 7929 2616
rect 7718 2586 8303 2592
rect 7718 2566 7734 2586
rect 7754 2585 8303 2586
rect 7754 2566 8274 2585
rect 7718 2565 8274 2566
rect 8294 2565 8303 2585
rect 7718 2557 8303 2565
rect 10004 2477 10589 2485
rect 10004 2457 10013 2477
rect 10033 2476 10589 2477
rect 10033 2457 10553 2476
rect 10004 2456 10553 2457
rect 10573 2456 10589 2476
rect 10004 2450 10589 2456
rect 9662 2444 9694 2445
rect 9659 2439 9694 2444
rect 9659 2419 9666 2439
rect 9686 2419 9694 2439
rect 9659 2411 9694 2419
rect 7650 2399 7685 2407
rect 6853 2179 6887 2385
rect 7650 2379 7658 2399
rect 7678 2379 7685 2399
rect 7650 2374 7685 2379
rect 7650 2373 7682 2374
rect 6921 2358 7506 2364
rect 6921 2338 6937 2358
rect 6957 2357 7506 2358
rect 6957 2338 7477 2357
rect 6921 2337 7477 2338
rect 7497 2337 7506 2357
rect 6921 2329 7506 2337
rect 7586 2328 7616 2329
rect 7586 2301 7922 2328
rect 7586 2300 7621 2301
rect 6853 2171 6888 2179
rect 6853 2151 6861 2171
rect 6881 2151 6888 2171
rect 6853 2146 6888 2151
rect 6853 2125 6887 2146
rect 7586 2125 7616 2300
rect 7672 2233 7707 2234
rect 6853 2099 7616 2125
rect 6854 2098 6887 2099
rect 7586 2097 7616 2099
rect 7651 2226 7707 2233
rect 7651 2206 7680 2226
rect 7700 2206 7707 2226
rect 7651 2201 7707 2206
rect 7886 2228 7921 2301
rect 7886 2208 7893 2228
rect 7913 2208 7921 2228
rect 9041 2253 9626 2261
rect 9041 2233 9050 2253
rect 9070 2252 9626 2253
rect 9070 2233 9590 2252
rect 9041 2232 9590 2233
rect 9610 2232 9626 2252
rect 9041 2226 9626 2232
rect 7886 2201 7921 2208
rect 9660 2205 9694 2411
rect 10389 2426 10422 2432
rect 10623 2429 10657 2635
rect 10389 2404 10394 2426
rect 10417 2404 10422 2426
rect 10389 2395 10422 2404
rect 10601 2424 10657 2429
rect 10601 2404 10608 2424
rect 10628 2404 10657 2424
rect 10601 2397 10657 2404
rect 10601 2396 10636 2397
rect 10391 2364 10418 2395
rect 10813 2364 10852 2376
rect 10391 2363 10854 2364
rect 10391 2341 10818 2363
rect 10842 2341 10854 2363
rect 10391 2333 10854 2341
rect 6681 2042 7020 2070
rect 6775 2007 6810 2008
rect 6754 2000 6810 2007
rect 6754 1980 6783 2000
rect 6803 1980 6810 2000
rect 6754 1975 6810 1980
rect 6989 2000 7020 2042
rect 6989 1981 6994 2000
rect 7015 1981 7020 2000
rect 6989 1975 7020 1981
rect 7651 1995 7685 2201
rect 9424 2198 9459 2205
rect 7719 2174 8304 2180
rect 7719 2154 7735 2174
rect 7755 2173 8304 2174
rect 7755 2154 8275 2173
rect 7719 2153 8275 2154
rect 8295 2153 8304 2173
rect 7719 2145 8304 2153
rect 9424 2178 9432 2198
rect 9452 2178 9459 2198
rect 9424 2105 9459 2178
rect 9638 2200 9694 2205
rect 9638 2180 9645 2200
rect 9665 2180 9694 2200
rect 9638 2173 9694 2180
rect 9729 2307 9759 2309
rect 10458 2307 10491 2308
rect 9729 2281 10492 2307
rect 9638 2172 9673 2173
rect 9729 2106 9759 2281
rect 10458 2260 10492 2281
rect 10457 2255 10492 2260
rect 10457 2235 10464 2255
rect 10484 2235 10492 2255
rect 10457 2227 10492 2235
rect 9724 2105 9759 2106
rect 9423 2078 9759 2105
rect 9729 2077 9759 2078
rect 9839 2069 10424 2077
rect 9839 2049 9848 2069
rect 9868 2068 10424 2069
rect 9868 2049 10388 2068
rect 9839 2048 10388 2049
rect 10408 2048 10424 2068
rect 9839 2042 10424 2048
rect 9663 2032 9695 2033
rect 9660 2027 9695 2032
rect 9660 2007 9667 2027
rect 9687 2007 9695 2027
rect 10458 2021 10492 2227
rect 9660 1999 9695 2007
rect 7651 1987 7686 1995
rect 6754 1769 6788 1975
rect 7651 1967 7659 1987
rect 7679 1967 7686 1987
rect 7651 1962 7686 1967
rect 7651 1961 7683 1962
rect 6822 1948 7407 1954
rect 6822 1928 6838 1948
rect 6858 1947 7407 1948
rect 6858 1928 7378 1947
rect 6822 1927 7378 1928
rect 7398 1927 7407 1947
rect 6822 1919 7407 1927
rect 9042 1841 9627 1849
rect 9042 1821 9051 1841
rect 9071 1840 9627 1841
rect 9071 1821 9591 1840
rect 9042 1820 9591 1821
rect 9611 1820 9627 1840
rect 9042 1814 9627 1820
rect 9416 1790 9455 1794
rect 9661 1793 9695 1999
rect 10224 2014 10259 2020
rect 10224 1995 10229 2014
rect 10250 1995 10259 2014
rect 10224 1986 10259 1995
rect 10436 2016 10492 2021
rect 10436 1996 10443 2016
rect 10463 1996 10492 2016
rect 10436 1989 10492 1996
rect 10614 2167 10646 2179
rect 10614 2149 10621 2167
rect 10643 2149 10646 2167
rect 10436 1988 10471 1989
rect 10228 1918 10257 1986
rect 10228 1884 10574 1918
rect 9416 1770 9424 1790
rect 9444 1770 9455 1790
rect 6754 1761 6789 1769
rect 6754 1741 6762 1761
rect 6782 1753 6789 1761
rect 6782 1741 6793 1753
rect 6754 1504 6793 1741
rect 7624 1718 7910 1719
rect 7109 1710 7912 1718
rect 7109 1693 7120 1710
rect 7110 1688 7120 1693
rect 7144 1693 7912 1710
rect 7144 1688 7149 1693
rect 7110 1675 7149 1688
rect 7654 1627 7689 1628
rect 7633 1620 7689 1627
rect 7633 1600 7662 1620
rect 7682 1600 7689 1620
rect 7633 1595 7689 1600
rect 7873 1618 7912 1693
rect 9416 1695 9455 1770
rect 9639 1788 9695 1793
rect 9639 1768 9646 1788
rect 9666 1768 9695 1788
rect 9639 1761 9695 1768
rect 9639 1760 9674 1761
rect 10179 1700 10218 1713
rect 10179 1695 10184 1700
rect 9416 1678 10184 1695
rect 10208 1695 10218 1700
rect 10208 1678 10219 1695
rect 9416 1670 10219 1678
rect 9418 1669 9704 1670
rect 10535 1647 10574 1884
rect 10535 1635 10546 1647
rect 10539 1627 10546 1635
rect 10566 1627 10574 1647
rect 10539 1619 10574 1627
rect 7873 1598 7884 1618
rect 7904 1598 7912 1618
rect 6754 1470 7100 1504
rect 7071 1402 7100 1470
rect 6857 1399 6892 1400
rect 5935 1300 6269 1328
rect 6836 1392 6892 1399
rect 6836 1372 6865 1392
rect 6885 1372 6892 1392
rect 6836 1367 6892 1372
rect 7069 1393 7104 1402
rect 7069 1374 7078 1393
rect 7099 1374 7104 1393
rect 7069 1368 7104 1374
rect 7633 1389 7667 1595
rect 7873 1594 7912 1598
rect 7701 1568 8286 1574
rect 7701 1548 7717 1568
rect 7737 1567 8286 1568
rect 7737 1548 8257 1567
rect 7701 1547 8257 1548
rect 8277 1547 8286 1567
rect 7701 1539 8286 1547
rect 9921 1461 10506 1469
rect 9921 1441 9930 1461
rect 9950 1460 10506 1461
rect 9950 1441 10470 1460
rect 9921 1440 10470 1441
rect 10490 1440 10506 1460
rect 9921 1434 10506 1440
rect 9645 1426 9677 1427
rect 9642 1421 9677 1426
rect 9642 1401 9649 1421
rect 9669 1401 9677 1421
rect 10540 1413 10574 1619
rect 9642 1393 9677 1401
rect 7633 1381 7668 1389
rect 902 956 937 964
rect 284 798 869 806
rect 284 778 293 798
rect 313 797 869 798
rect 313 778 833 797
rect 284 777 833 778
rect 853 777 869 797
rect 284 771 869 777
rect 658 747 697 751
rect 903 750 937 956
rect 1467 968 1501 976
rect 1467 950 1474 968
rect 1493 950 1501 968
rect 1467 943 1501 950
rect 1678 973 1734 978
rect 1678 953 1685 973
rect 1705 953 1734 973
rect 1678 946 1734 953
rect 3270 964 3304 1170
rect 5030 1168 5065 1175
rect 3338 1143 3923 1149
rect 3338 1123 3354 1143
rect 3374 1142 3923 1143
rect 3374 1123 3894 1142
rect 3338 1122 3894 1123
rect 3914 1122 3923 1142
rect 3338 1114 3923 1122
rect 5030 1148 5038 1168
rect 5058 1148 5065 1168
rect 5030 1075 5065 1148
rect 5244 1170 5300 1175
rect 5244 1150 5251 1170
rect 5271 1150 5300 1170
rect 5244 1143 5300 1150
rect 5335 1277 5365 1279
rect 6064 1277 6097 1278
rect 5335 1251 6098 1277
rect 5244 1142 5279 1143
rect 5335 1076 5365 1251
rect 6064 1230 6098 1251
rect 6063 1225 6098 1230
rect 6063 1205 6070 1225
rect 6090 1205 6098 1225
rect 6063 1197 6098 1205
rect 5330 1075 5365 1076
rect 5029 1048 5365 1075
rect 5335 1047 5365 1048
rect 5445 1039 6030 1047
rect 5445 1019 5454 1039
rect 5474 1038 6030 1039
rect 5474 1019 5994 1038
rect 5445 1018 5994 1019
rect 6014 1018 6030 1038
rect 5445 1012 6030 1018
rect 5269 1002 5301 1003
rect 5266 997 5301 1002
rect 5266 977 5273 997
rect 5293 977 5301 997
rect 6064 991 6098 1197
rect 6836 1161 6870 1367
rect 7633 1361 7641 1381
rect 7661 1361 7668 1381
rect 7633 1356 7668 1361
rect 7633 1355 7665 1356
rect 6904 1340 7489 1346
rect 6904 1320 6920 1340
rect 6940 1339 7489 1340
rect 6940 1320 7460 1339
rect 6904 1319 7460 1320
rect 7480 1319 7489 1339
rect 6904 1311 7489 1319
rect 7569 1310 7599 1311
rect 7569 1283 7905 1310
rect 7569 1282 7604 1283
rect 6836 1153 6871 1161
rect 6836 1133 6844 1153
rect 6864 1133 6871 1153
rect 6836 1128 6871 1133
rect 6836 1107 6870 1128
rect 7569 1107 7599 1282
rect 7655 1215 7690 1216
rect 6836 1081 7599 1107
rect 6837 1080 6870 1081
rect 7569 1079 7599 1081
rect 7634 1208 7690 1215
rect 7634 1188 7663 1208
rect 7683 1188 7690 1208
rect 7634 1183 7690 1188
rect 7869 1210 7904 1283
rect 7869 1190 7876 1210
rect 7896 1190 7904 1210
rect 9024 1235 9609 1243
rect 9024 1215 9033 1235
rect 9053 1234 9609 1235
rect 9053 1215 9573 1234
rect 9024 1214 9573 1215
rect 9593 1214 9609 1234
rect 9024 1208 9609 1214
rect 7869 1183 7904 1190
rect 9643 1187 9677 1393
rect 10306 1401 10342 1410
rect 10306 1384 10315 1401
rect 10334 1384 10342 1401
rect 10306 1375 10342 1384
rect 10518 1408 10574 1413
rect 10518 1388 10525 1408
rect 10545 1388 10574 1408
rect 10518 1381 10574 1388
rect 10518 1380 10553 1381
rect 10312 1340 10338 1375
rect 10614 1340 10646 2149
rect 11058 2082 11087 2767
rect 12018 2748 12304 2749
rect 11503 2740 12306 2748
rect 11503 2723 11514 2740
rect 11504 2718 11514 2723
rect 11538 2723 12306 2740
rect 11538 2718 11543 2723
rect 11504 2705 11543 2718
rect 12048 2657 12083 2658
rect 12027 2650 12083 2657
rect 12027 2630 12056 2650
rect 12076 2630 12083 2650
rect 12027 2625 12083 2630
rect 12267 2648 12306 2723
rect 13800 2726 13839 2801
rect 14023 2819 14079 2824
rect 14023 2799 14030 2819
rect 14050 2799 14079 2819
rect 14023 2792 14079 2799
rect 14023 2791 14058 2792
rect 14563 2731 14602 2744
rect 14563 2726 14568 2731
rect 13800 2709 14568 2726
rect 14592 2726 14602 2731
rect 14592 2709 14603 2726
rect 13800 2701 14603 2709
rect 13802 2700 14088 2701
rect 15019 2682 15048 3367
rect 15356 3121 15383 4821
rect 16419 4797 16705 4798
rect 15904 4789 16707 4797
rect 15904 4772 15915 4789
rect 15905 4767 15915 4772
rect 15939 4772 16707 4789
rect 15939 4767 15944 4772
rect 15905 4754 15944 4767
rect 16449 4706 16484 4707
rect 16428 4699 16484 4706
rect 16428 4679 16457 4699
rect 16477 4679 16484 4699
rect 16428 4674 16484 4679
rect 16668 4697 16707 4772
rect 16668 4677 16679 4697
rect 16699 4677 16707 4697
rect 15512 4538 15894 4543
rect 15512 4519 15520 4538
rect 15541 4519 15894 4538
rect 15512 4511 15894 4519
rect 15865 4481 15894 4511
rect 15652 4478 15687 4479
rect 15631 4471 15687 4478
rect 15631 4451 15660 4471
rect 15680 4451 15687 4471
rect 15631 4446 15687 4451
rect 15864 4474 15898 4481
rect 15864 4456 15872 4474
rect 15891 4456 15898 4474
rect 15864 4448 15898 4456
rect 16428 4468 16462 4674
rect 16668 4673 16707 4677
rect 16496 4647 17081 4653
rect 16496 4627 16512 4647
rect 16532 4646 17081 4647
rect 16532 4627 17052 4646
rect 16496 4626 17052 4627
rect 17072 4626 17081 4646
rect 16496 4618 17081 4626
rect 16428 4460 16463 4468
rect 15631 4240 15665 4446
rect 16428 4440 16436 4460
rect 16456 4440 16463 4460
rect 16428 4435 16463 4440
rect 16428 4434 16460 4435
rect 15699 4419 16284 4425
rect 15699 4399 15715 4419
rect 15735 4418 16284 4419
rect 15735 4399 16255 4418
rect 15699 4398 16255 4399
rect 16275 4398 16284 4418
rect 15699 4390 16284 4398
rect 16364 4389 16394 4390
rect 16364 4362 16700 4389
rect 16364 4361 16399 4362
rect 15631 4232 15666 4240
rect 15631 4212 15639 4232
rect 15659 4212 15666 4232
rect 15631 4207 15666 4212
rect 15631 4186 15665 4207
rect 16364 4186 16394 4361
rect 16450 4294 16485 4295
rect 15631 4160 16394 4186
rect 15632 4159 15665 4160
rect 16364 4158 16394 4160
rect 16429 4287 16485 4294
rect 16429 4267 16458 4287
rect 16478 4267 16485 4287
rect 16429 4262 16485 4267
rect 16664 4289 16699 4362
rect 16664 4269 16671 4289
rect 16691 4269 16699 4289
rect 16664 4262 16699 4269
rect 15454 4137 15486 4138
rect 15454 4132 15794 4137
rect 15454 4114 15457 4132
rect 15479 4114 15794 4132
rect 15454 4109 15794 4114
rect 15454 4108 15486 4109
rect 15768 4074 15794 4109
rect 15553 4068 15588 4069
rect 15532 4061 15588 4068
rect 15532 4041 15561 4061
rect 15581 4041 15588 4061
rect 15532 4036 15588 4041
rect 15764 4065 15800 4074
rect 15764 4048 15772 4065
rect 15791 4048 15800 4065
rect 15764 4039 15800 4048
rect 16429 4056 16463 4262
rect 16497 4235 17082 4241
rect 16497 4215 16513 4235
rect 16533 4234 17082 4235
rect 16533 4215 17053 4234
rect 16497 4214 17053 4215
rect 17073 4214 17082 4234
rect 16497 4206 17082 4214
rect 16429 4048 16464 4056
rect 15532 3830 15566 4036
rect 16429 4028 16437 4048
rect 16457 4028 16464 4048
rect 16429 4023 16464 4028
rect 16429 4022 16461 4023
rect 15600 4009 16185 4015
rect 15600 3989 15616 4009
rect 15636 4008 16185 4009
rect 15636 3989 16156 4008
rect 15600 3988 16156 3989
rect 16176 3988 16185 4008
rect 15600 3980 16185 3988
rect 15532 3822 15567 3830
rect 15532 3802 15540 3822
rect 15560 3814 15567 3822
rect 15560 3802 15571 3814
rect 15532 3565 15571 3802
rect 16402 3779 16688 3780
rect 15887 3771 16690 3779
rect 15887 3754 15898 3771
rect 15888 3749 15898 3754
rect 15922 3754 16690 3771
rect 15922 3749 15927 3754
rect 15888 3736 15927 3749
rect 16432 3688 16467 3689
rect 16411 3681 16467 3688
rect 16411 3661 16440 3681
rect 16460 3661 16467 3681
rect 16411 3656 16467 3661
rect 16651 3679 16690 3754
rect 16651 3659 16662 3679
rect 16682 3659 16690 3679
rect 15532 3531 15878 3565
rect 15849 3463 15878 3531
rect 15635 3460 15670 3461
rect 15614 3453 15670 3460
rect 15614 3433 15643 3453
rect 15663 3433 15670 3453
rect 15614 3428 15670 3433
rect 15847 3454 15882 3463
rect 15847 3435 15856 3454
rect 15877 3435 15882 3454
rect 15847 3429 15882 3435
rect 16411 3450 16445 3656
rect 16651 3655 16690 3659
rect 16479 3629 17064 3635
rect 16479 3609 16495 3629
rect 16515 3628 17064 3629
rect 16515 3609 17035 3628
rect 16479 3608 17035 3609
rect 17055 3608 17064 3628
rect 16479 3600 17064 3608
rect 16411 3442 16446 3450
rect 15614 3222 15648 3428
rect 16411 3422 16419 3442
rect 16439 3422 16446 3442
rect 16411 3417 16446 3422
rect 16411 3416 16443 3417
rect 15682 3401 16267 3407
rect 15682 3381 15698 3401
rect 15718 3400 16267 3401
rect 15718 3381 16238 3400
rect 15682 3380 16238 3381
rect 16258 3380 16267 3400
rect 15682 3372 16267 3380
rect 16347 3371 16377 3372
rect 16347 3344 16683 3371
rect 16347 3343 16382 3344
rect 15614 3214 15649 3222
rect 15614 3194 15622 3214
rect 15642 3194 15649 3214
rect 15614 3189 15649 3194
rect 15614 3168 15648 3189
rect 16347 3168 16377 3343
rect 16433 3276 16468 3277
rect 15614 3142 16377 3168
rect 15615 3141 15648 3142
rect 16347 3140 16377 3142
rect 16412 3269 16468 3276
rect 16412 3249 16441 3269
rect 16461 3249 16468 3269
rect 16412 3244 16468 3249
rect 16647 3271 16682 3344
rect 16647 3251 16654 3271
rect 16674 3251 16682 3271
rect 16647 3244 16682 3251
rect 15356 3085 15710 3121
rect 15372 3084 15710 3085
rect 15684 3054 15710 3084
rect 15470 3052 15505 3053
rect 15449 3045 15505 3052
rect 15449 3025 15478 3045
rect 15498 3025 15505 3045
rect 15449 3020 15505 3025
rect 15678 3046 15719 3054
rect 15678 3028 15691 3046
rect 15709 3028 15719 3046
rect 15449 2814 15483 3020
rect 15678 3017 15719 3028
rect 16412 3038 16446 3244
rect 16480 3217 17065 3223
rect 16480 3197 16496 3217
rect 16516 3216 17065 3217
rect 16516 3197 17036 3216
rect 16480 3196 17036 3197
rect 17056 3196 17065 3216
rect 16480 3188 17065 3196
rect 16412 3030 16447 3038
rect 16412 3010 16420 3030
rect 16440 3010 16447 3030
rect 16412 3005 16447 3010
rect 16412 3004 16444 3005
rect 15517 2993 16102 2999
rect 15517 2973 15533 2993
rect 15553 2992 16102 2993
rect 15553 2973 16073 2992
rect 15517 2972 16073 2973
rect 16093 2972 16102 2992
rect 15517 2964 16102 2972
rect 15449 2813 15484 2814
rect 15417 2806 15484 2813
rect 15417 2786 15457 2806
rect 15477 2786 15484 2806
rect 15417 2783 15484 2786
rect 15417 2780 15482 2783
rect 14988 2679 15053 2682
rect 14986 2676 15053 2679
rect 14986 2656 14993 2676
rect 15013 2656 15053 2676
rect 14986 2649 15053 2656
rect 14986 2648 15021 2649
rect 12267 2628 12278 2648
rect 12298 2628 12306 2648
rect 11111 2489 11493 2494
rect 11111 2470 11119 2489
rect 11140 2470 11493 2489
rect 11111 2462 11493 2470
rect 11464 2432 11493 2462
rect 11251 2429 11286 2430
rect 11230 2422 11286 2429
rect 11230 2402 11259 2422
rect 11279 2402 11286 2422
rect 11230 2397 11286 2402
rect 11463 2425 11497 2432
rect 11463 2407 11471 2425
rect 11490 2407 11497 2425
rect 11463 2399 11497 2407
rect 12027 2419 12061 2625
rect 12267 2624 12306 2628
rect 12095 2598 12680 2604
rect 12095 2578 12111 2598
rect 12131 2597 12680 2598
rect 12131 2578 12651 2597
rect 12095 2577 12651 2578
rect 12671 2577 12680 2597
rect 12095 2569 12680 2577
rect 14368 2490 14953 2498
rect 14368 2470 14377 2490
rect 14397 2489 14953 2490
rect 14397 2470 14917 2489
rect 14368 2469 14917 2470
rect 14937 2469 14953 2489
rect 14368 2463 14953 2469
rect 14026 2457 14058 2458
rect 14023 2452 14058 2457
rect 14023 2432 14030 2452
rect 14050 2432 14058 2452
rect 14023 2424 14058 2432
rect 12027 2411 12062 2419
rect 11230 2191 11264 2397
rect 12027 2391 12035 2411
rect 12055 2391 12062 2411
rect 12027 2386 12062 2391
rect 12027 2385 12059 2386
rect 11298 2370 11883 2376
rect 11298 2350 11314 2370
rect 11334 2369 11883 2370
rect 11334 2350 11854 2369
rect 11298 2349 11854 2350
rect 11874 2349 11883 2369
rect 11298 2341 11883 2349
rect 11963 2340 11993 2341
rect 11963 2313 12299 2340
rect 11963 2312 11998 2313
rect 11230 2183 11265 2191
rect 11230 2163 11238 2183
rect 11258 2163 11265 2183
rect 11230 2158 11265 2163
rect 11230 2137 11264 2158
rect 11963 2137 11993 2312
rect 12049 2245 12084 2246
rect 11230 2111 11993 2137
rect 11231 2110 11264 2111
rect 11963 2109 11993 2111
rect 12028 2238 12084 2245
rect 12028 2218 12057 2238
rect 12077 2218 12084 2238
rect 12028 2213 12084 2218
rect 12263 2240 12298 2313
rect 12263 2220 12270 2240
rect 12290 2220 12298 2240
rect 13405 2266 13990 2274
rect 13405 2246 13414 2266
rect 13434 2265 13990 2266
rect 13434 2246 13954 2265
rect 13405 2245 13954 2246
rect 13974 2245 13990 2265
rect 13405 2239 13990 2245
rect 12263 2213 12298 2220
rect 14024 2218 14058 2424
rect 14753 2439 14786 2445
rect 14987 2442 15021 2648
rect 14753 2417 14758 2439
rect 14781 2417 14786 2439
rect 14753 2408 14786 2417
rect 14965 2437 15021 2442
rect 14965 2417 14972 2437
rect 14992 2417 15021 2437
rect 14965 2410 15021 2417
rect 14965 2409 15000 2410
rect 14755 2377 14782 2408
rect 15177 2377 15216 2389
rect 14755 2376 15218 2377
rect 14755 2354 15182 2376
rect 15206 2354 15218 2376
rect 14755 2346 15218 2354
rect 11058 2054 11397 2082
rect 11152 2019 11187 2020
rect 11131 2012 11187 2019
rect 11131 1992 11160 2012
rect 11180 1992 11187 2012
rect 11131 1987 11187 1992
rect 11366 2012 11397 2054
rect 11366 1993 11371 2012
rect 11392 1993 11397 2012
rect 11366 1987 11397 1993
rect 12028 2007 12062 2213
rect 13788 2211 13823 2218
rect 12096 2186 12681 2192
rect 12096 2166 12112 2186
rect 12132 2185 12681 2186
rect 12132 2166 12652 2185
rect 12096 2165 12652 2166
rect 12672 2165 12681 2185
rect 12096 2157 12681 2165
rect 13788 2191 13796 2211
rect 13816 2191 13823 2211
rect 13788 2118 13823 2191
rect 14002 2213 14058 2218
rect 14002 2193 14009 2213
rect 14029 2193 14058 2213
rect 14002 2186 14058 2193
rect 14093 2320 14123 2322
rect 14822 2320 14855 2321
rect 14093 2294 14856 2320
rect 14002 2185 14037 2186
rect 14093 2119 14123 2294
rect 14822 2273 14856 2294
rect 14821 2268 14856 2273
rect 14821 2248 14828 2268
rect 14848 2248 14856 2268
rect 14821 2240 14856 2248
rect 14088 2118 14123 2119
rect 13787 2091 14123 2118
rect 14093 2090 14123 2091
rect 14203 2082 14788 2090
rect 14203 2062 14212 2082
rect 14232 2081 14788 2082
rect 14232 2062 14752 2081
rect 14203 2061 14752 2062
rect 14772 2061 14788 2081
rect 14203 2055 14788 2061
rect 14027 2045 14059 2046
rect 14024 2040 14059 2045
rect 14024 2020 14031 2040
rect 14051 2020 14059 2040
rect 14822 2034 14856 2240
rect 14024 2012 14059 2020
rect 12028 1999 12063 2007
rect 11131 1781 11165 1987
rect 12028 1979 12036 1999
rect 12056 1979 12063 1999
rect 12028 1974 12063 1979
rect 12028 1973 12060 1974
rect 11199 1960 11784 1966
rect 11199 1940 11215 1960
rect 11235 1959 11784 1960
rect 11235 1940 11755 1959
rect 11199 1939 11755 1940
rect 11775 1939 11784 1959
rect 11199 1931 11784 1939
rect 13406 1854 13991 1862
rect 13406 1834 13415 1854
rect 13435 1853 13991 1854
rect 13435 1834 13955 1853
rect 13406 1833 13955 1834
rect 13975 1833 13991 1853
rect 13406 1827 13991 1833
rect 13780 1803 13819 1807
rect 14025 1806 14059 2012
rect 14588 2027 14623 2033
rect 14588 2008 14593 2027
rect 14614 2008 14623 2027
rect 14588 1999 14623 2008
rect 14800 2029 14856 2034
rect 14800 2009 14807 2029
rect 14827 2009 14856 2029
rect 14800 2002 14856 2009
rect 14978 2180 15010 2192
rect 14978 2162 14985 2180
rect 15007 2162 15010 2180
rect 14800 2001 14835 2002
rect 14592 1931 14621 1999
rect 14592 1897 14938 1931
rect 13780 1783 13788 1803
rect 13808 1783 13819 1803
rect 11131 1773 11166 1781
rect 11131 1753 11139 1773
rect 11159 1765 11166 1773
rect 11159 1753 11170 1765
rect 11131 1516 11170 1753
rect 12001 1730 12287 1731
rect 11486 1722 12289 1730
rect 11486 1705 11497 1722
rect 11487 1700 11497 1705
rect 11521 1705 12289 1722
rect 11521 1700 11526 1705
rect 11487 1687 11526 1700
rect 12031 1639 12066 1640
rect 12010 1632 12066 1639
rect 12010 1612 12039 1632
rect 12059 1612 12066 1632
rect 12010 1607 12066 1612
rect 12250 1630 12289 1705
rect 13780 1708 13819 1783
rect 14003 1801 14059 1806
rect 14003 1781 14010 1801
rect 14030 1781 14059 1801
rect 14003 1774 14059 1781
rect 14003 1773 14038 1774
rect 14543 1713 14582 1726
rect 14543 1708 14548 1713
rect 13780 1691 14548 1708
rect 14572 1708 14582 1713
rect 14572 1691 14583 1708
rect 13780 1683 14583 1691
rect 13782 1682 14068 1683
rect 14899 1660 14938 1897
rect 14899 1648 14910 1660
rect 14903 1640 14910 1648
rect 14930 1640 14938 1660
rect 14903 1632 14938 1640
rect 12250 1610 12261 1630
rect 12281 1610 12289 1630
rect 11131 1482 11477 1516
rect 11448 1414 11477 1482
rect 11234 1411 11269 1412
rect 10312 1312 10646 1340
rect 11213 1404 11269 1411
rect 11213 1384 11242 1404
rect 11262 1384 11269 1404
rect 11213 1379 11269 1384
rect 11446 1405 11481 1414
rect 11446 1386 11455 1405
rect 11476 1386 11481 1405
rect 11446 1380 11481 1386
rect 12010 1401 12044 1607
rect 12250 1606 12289 1610
rect 12078 1580 12663 1586
rect 12078 1560 12094 1580
rect 12114 1579 12663 1580
rect 12114 1560 12634 1579
rect 12078 1559 12634 1560
rect 12654 1559 12663 1579
rect 12078 1551 12663 1559
rect 14285 1474 14870 1482
rect 14285 1454 14294 1474
rect 14314 1473 14870 1474
rect 14314 1454 14834 1473
rect 14285 1453 14834 1454
rect 14854 1453 14870 1473
rect 14285 1447 14870 1453
rect 14009 1439 14041 1440
rect 14006 1434 14041 1439
rect 14006 1414 14013 1434
rect 14033 1414 14041 1434
rect 14904 1426 14938 1632
rect 14006 1406 14041 1414
rect 12010 1393 12045 1401
rect 5266 969 5301 977
rect 3270 956 3305 964
rect 1678 945 1713 946
rect 1471 913 1500 943
rect 3270 936 3278 956
rect 3298 936 3305 956
rect 3270 931 3305 936
rect 3270 930 3302 931
rect 1471 905 1853 913
rect 1471 886 1824 905
rect 1845 886 1853 905
rect 1471 881 1853 886
rect 4648 811 5233 819
rect 4648 791 4657 811
rect 4677 810 5233 811
rect 4677 791 5197 810
rect 4648 790 5197 791
rect 5217 790 5233 810
rect 4648 784 5233 790
rect 658 727 666 747
rect 686 727 697 747
rect 658 652 697 727
rect 881 745 937 750
rect 881 725 888 745
rect 908 725 937 745
rect 881 718 937 725
rect 5022 760 5061 764
rect 5267 763 5301 969
rect 5831 981 5865 989
rect 5831 963 5838 981
rect 5857 963 5865 981
rect 5831 956 5865 963
rect 6042 986 6098 991
rect 6042 966 6049 986
rect 6069 966 6098 986
rect 6042 959 6098 966
rect 7634 977 7668 1183
rect 9407 1180 9442 1187
rect 7702 1156 8287 1162
rect 7702 1136 7718 1156
rect 7738 1155 8287 1156
rect 7738 1136 8258 1155
rect 7702 1135 8258 1136
rect 8278 1135 8287 1155
rect 7702 1127 8287 1135
rect 9407 1160 9415 1180
rect 9435 1160 9442 1180
rect 9407 1087 9442 1160
rect 9621 1182 9677 1187
rect 9621 1162 9628 1182
rect 9648 1162 9677 1182
rect 9621 1155 9677 1162
rect 9712 1289 9742 1291
rect 10441 1289 10474 1290
rect 9712 1263 10475 1289
rect 9621 1154 9656 1155
rect 9712 1088 9742 1263
rect 10441 1242 10475 1263
rect 10440 1237 10475 1242
rect 10440 1217 10447 1237
rect 10467 1217 10475 1237
rect 10440 1209 10475 1217
rect 9707 1087 9742 1088
rect 9406 1060 9742 1087
rect 9712 1059 9742 1060
rect 9822 1051 10407 1059
rect 9822 1031 9831 1051
rect 9851 1050 10407 1051
rect 9851 1031 10371 1050
rect 9822 1030 10371 1031
rect 10391 1030 10407 1050
rect 9822 1024 10407 1030
rect 9646 1014 9678 1015
rect 9643 1009 9678 1014
rect 9643 989 9650 1009
rect 9670 989 9678 1009
rect 10441 1003 10475 1209
rect 11213 1173 11247 1379
rect 12010 1373 12018 1393
rect 12038 1373 12045 1393
rect 12010 1368 12045 1373
rect 12010 1367 12042 1368
rect 11281 1352 11866 1358
rect 11281 1332 11297 1352
rect 11317 1351 11866 1352
rect 11317 1332 11837 1351
rect 11281 1331 11837 1332
rect 11857 1331 11866 1351
rect 11281 1323 11866 1331
rect 11946 1322 11976 1323
rect 11946 1295 12282 1322
rect 11946 1294 11981 1295
rect 11213 1165 11248 1173
rect 11213 1145 11221 1165
rect 11241 1145 11248 1165
rect 11213 1140 11248 1145
rect 11213 1119 11247 1140
rect 11946 1119 11976 1294
rect 12032 1227 12067 1228
rect 11213 1093 11976 1119
rect 11214 1092 11247 1093
rect 11946 1091 11976 1093
rect 12011 1220 12067 1227
rect 12011 1200 12040 1220
rect 12060 1200 12067 1220
rect 12011 1195 12067 1200
rect 12246 1222 12281 1295
rect 12246 1202 12253 1222
rect 12273 1202 12281 1222
rect 13388 1248 13973 1256
rect 13388 1228 13397 1248
rect 13417 1247 13973 1248
rect 13417 1228 13937 1247
rect 13388 1227 13937 1228
rect 13957 1227 13973 1247
rect 13388 1221 13973 1227
rect 12246 1195 12281 1202
rect 14007 1200 14041 1406
rect 14670 1414 14706 1423
rect 14670 1397 14679 1414
rect 14698 1397 14706 1414
rect 14670 1388 14706 1397
rect 14882 1421 14938 1426
rect 14882 1401 14889 1421
rect 14909 1401 14938 1421
rect 14882 1394 14938 1401
rect 14882 1393 14917 1394
rect 14676 1353 14702 1388
rect 14978 1353 15010 2162
rect 15422 2095 15451 2780
rect 16382 2761 16668 2762
rect 15867 2753 16670 2761
rect 15867 2736 15878 2753
rect 15868 2731 15878 2736
rect 15902 2736 16670 2753
rect 15902 2731 15907 2736
rect 15868 2718 15907 2731
rect 16412 2670 16447 2671
rect 16391 2663 16447 2670
rect 16391 2643 16420 2663
rect 16440 2643 16447 2663
rect 16391 2638 16447 2643
rect 16631 2661 16670 2736
rect 16631 2641 16642 2661
rect 16662 2641 16670 2661
rect 15475 2502 15857 2507
rect 15475 2483 15483 2502
rect 15504 2483 15857 2502
rect 15475 2475 15857 2483
rect 15828 2445 15857 2475
rect 15615 2442 15650 2443
rect 15594 2435 15650 2442
rect 15594 2415 15623 2435
rect 15643 2415 15650 2435
rect 15594 2410 15650 2415
rect 15827 2438 15861 2445
rect 15827 2420 15835 2438
rect 15854 2420 15861 2438
rect 15827 2412 15861 2420
rect 16391 2432 16425 2638
rect 16631 2637 16670 2641
rect 16459 2611 17044 2617
rect 16459 2591 16475 2611
rect 16495 2610 17044 2611
rect 16495 2591 17015 2610
rect 16459 2590 17015 2591
rect 17035 2590 17044 2610
rect 16459 2582 17044 2590
rect 16391 2424 16426 2432
rect 15594 2204 15628 2410
rect 16391 2404 16399 2424
rect 16419 2404 16426 2424
rect 16391 2399 16426 2404
rect 16391 2398 16423 2399
rect 15662 2383 16247 2389
rect 15662 2363 15678 2383
rect 15698 2382 16247 2383
rect 15698 2363 16218 2382
rect 15662 2362 16218 2363
rect 16238 2362 16247 2382
rect 15662 2354 16247 2362
rect 16327 2353 16357 2354
rect 16327 2326 16663 2353
rect 16327 2325 16362 2326
rect 15594 2196 15629 2204
rect 15594 2176 15602 2196
rect 15622 2176 15629 2196
rect 15594 2171 15629 2176
rect 15594 2150 15628 2171
rect 16327 2150 16357 2325
rect 16413 2258 16448 2259
rect 15594 2124 16357 2150
rect 15595 2123 15628 2124
rect 16327 2122 16357 2124
rect 16392 2251 16448 2258
rect 16392 2231 16421 2251
rect 16441 2231 16448 2251
rect 16392 2226 16448 2231
rect 16627 2253 16662 2326
rect 16627 2233 16634 2253
rect 16654 2233 16662 2253
rect 16627 2226 16662 2233
rect 15422 2067 15761 2095
rect 15516 2032 15551 2033
rect 15495 2025 15551 2032
rect 15495 2005 15524 2025
rect 15544 2005 15551 2025
rect 15495 2000 15551 2005
rect 15730 2025 15761 2067
rect 15730 2006 15735 2025
rect 15756 2006 15761 2025
rect 15730 2000 15761 2006
rect 16392 2020 16426 2226
rect 16460 2199 17045 2205
rect 16460 2179 16476 2199
rect 16496 2198 17045 2199
rect 16496 2179 17016 2198
rect 16460 2178 17016 2179
rect 17036 2178 17045 2198
rect 16460 2170 17045 2178
rect 16392 2012 16427 2020
rect 15495 1794 15529 2000
rect 16392 1992 16400 2012
rect 16420 1992 16427 2012
rect 16392 1987 16427 1992
rect 16392 1986 16424 1987
rect 15563 1973 16148 1979
rect 15563 1953 15579 1973
rect 15599 1972 16148 1973
rect 15599 1953 16119 1972
rect 15563 1952 16119 1953
rect 16139 1952 16148 1972
rect 15563 1944 16148 1952
rect 15495 1786 15530 1794
rect 15495 1766 15503 1786
rect 15523 1778 15530 1786
rect 15523 1766 15534 1778
rect 15495 1529 15534 1766
rect 16365 1743 16651 1744
rect 15850 1735 16653 1743
rect 15850 1718 15861 1735
rect 15851 1713 15861 1718
rect 15885 1718 16653 1735
rect 15885 1713 15890 1718
rect 15851 1700 15890 1713
rect 16395 1652 16430 1653
rect 16374 1645 16430 1652
rect 16374 1625 16403 1645
rect 16423 1625 16430 1645
rect 16374 1620 16430 1625
rect 16614 1643 16653 1718
rect 16614 1623 16625 1643
rect 16645 1623 16653 1643
rect 15495 1495 15841 1529
rect 15812 1427 15841 1495
rect 15598 1424 15633 1425
rect 14676 1325 15010 1353
rect 15577 1417 15633 1424
rect 15577 1397 15606 1417
rect 15626 1397 15633 1417
rect 15577 1392 15633 1397
rect 15810 1418 15845 1427
rect 15810 1399 15819 1418
rect 15840 1399 15845 1418
rect 15810 1393 15845 1399
rect 16374 1414 16408 1620
rect 16614 1619 16653 1623
rect 16442 1593 17027 1599
rect 16442 1573 16458 1593
rect 16478 1592 17027 1593
rect 16478 1573 16998 1592
rect 16442 1572 16998 1573
rect 17018 1572 17027 1592
rect 16442 1564 17027 1572
rect 16374 1406 16409 1414
rect 9643 981 9678 989
rect 7634 969 7669 977
rect 6042 958 6077 959
rect 5835 926 5864 956
rect 7634 949 7642 969
rect 7662 949 7669 969
rect 7634 944 7669 949
rect 7634 943 7666 944
rect 5835 918 6217 926
rect 5835 899 6188 918
rect 6209 899 6217 918
rect 5835 894 6217 899
rect 9025 823 9610 831
rect 9025 803 9034 823
rect 9054 822 9610 823
rect 9054 803 9574 822
rect 9025 802 9574 803
rect 9594 802 9610 822
rect 9025 796 9610 802
rect 5022 740 5030 760
rect 5050 740 5061 760
rect 881 717 916 718
rect 2116 670 2167 701
rect 1421 657 1460 670
rect 1421 652 1426 657
rect 658 635 1426 652
rect 1450 652 1460 657
rect 1450 635 1461 652
rect 658 627 1461 635
rect 2116 644 2133 670
rect 2161 644 2167 670
rect 660 626 946 627
rect 2116 621 2167 644
rect 2196 676 2242 707
rect 4040 705 4083 713
rect 2196 645 2210 676
rect 2238 645 2242 676
rect 2196 638 2242 645
rect 4034 698 4089 705
rect 4034 673 4047 698
rect 4079 673 4089 698
rect 498 610 559 619
rect 498 583 506 610
rect 542 604 559 610
rect 600 604 675 608
rect 542 602 675 604
rect 542 583 606 602
rect 498 566 606 583
rect 651 566 675 602
rect 498 564 675 566
rect 600 534 675 564
rect 2129 429 2160 621
rect 2115 408 2161 429
rect 2115 387 2122 408
rect 2143 387 2161 408
rect 2115 383 2161 387
rect 2115 380 2150 383
rect 1497 222 2082 230
rect 1497 202 1506 222
rect 1526 221 2082 222
rect 1526 202 2046 221
rect 1497 201 2046 202
rect 2066 201 2082 221
rect 1497 195 2082 201
rect 2116 174 2150 380
rect 2198 314 2232 638
rect 4034 581 4089 673
rect 5022 665 5061 740
rect 5245 758 5301 763
rect 5245 738 5252 758
rect 5272 738 5301 758
rect 5245 731 5301 738
rect 9399 772 9438 776
rect 9644 775 9678 981
rect 10208 993 10242 1001
rect 10208 975 10215 993
rect 10234 975 10242 993
rect 10208 968 10242 975
rect 10419 998 10475 1003
rect 10419 978 10426 998
rect 10446 978 10475 998
rect 10419 971 10475 978
rect 12011 989 12045 1195
rect 13771 1193 13806 1200
rect 12079 1168 12664 1174
rect 12079 1148 12095 1168
rect 12115 1167 12664 1168
rect 12115 1148 12635 1167
rect 12079 1147 12635 1148
rect 12655 1147 12664 1167
rect 12079 1139 12664 1147
rect 13771 1173 13779 1193
rect 13799 1173 13806 1193
rect 13771 1100 13806 1173
rect 13985 1195 14041 1200
rect 13985 1175 13992 1195
rect 14012 1175 14041 1195
rect 13985 1168 14041 1175
rect 14076 1302 14106 1304
rect 14805 1302 14838 1303
rect 14076 1276 14839 1302
rect 13985 1167 14020 1168
rect 14076 1101 14106 1276
rect 14805 1255 14839 1276
rect 14804 1250 14839 1255
rect 14804 1230 14811 1250
rect 14831 1230 14839 1250
rect 14804 1222 14839 1230
rect 14071 1100 14106 1101
rect 13770 1073 14106 1100
rect 14076 1072 14106 1073
rect 14186 1064 14771 1072
rect 14186 1044 14195 1064
rect 14215 1063 14771 1064
rect 14215 1044 14735 1063
rect 14186 1043 14735 1044
rect 14755 1043 14771 1063
rect 14186 1037 14771 1043
rect 14010 1027 14042 1028
rect 14007 1022 14042 1027
rect 14007 1002 14014 1022
rect 14034 1002 14042 1022
rect 14805 1016 14839 1222
rect 15577 1186 15611 1392
rect 16374 1386 16382 1406
rect 16402 1386 16409 1406
rect 16374 1381 16409 1386
rect 16374 1380 16406 1381
rect 15645 1365 16230 1371
rect 15645 1345 15661 1365
rect 15681 1364 16230 1365
rect 15681 1345 16201 1364
rect 15645 1344 16201 1345
rect 16221 1344 16230 1364
rect 15645 1336 16230 1344
rect 16310 1335 16340 1336
rect 16310 1308 16646 1335
rect 16310 1307 16345 1308
rect 15577 1178 15612 1186
rect 15577 1158 15585 1178
rect 15605 1158 15612 1178
rect 15577 1153 15612 1158
rect 15577 1132 15611 1153
rect 16310 1132 16340 1307
rect 16396 1240 16431 1241
rect 15577 1106 16340 1132
rect 15578 1105 15611 1106
rect 16310 1104 16340 1106
rect 16375 1233 16431 1240
rect 16375 1213 16404 1233
rect 16424 1213 16431 1233
rect 16375 1208 16431 1213
rect 16610 1235 16645 1308
rect 16610 1215 16617 1235
rect 16637 1215 16645 1235
rect 16610 1208 16645 1215
rect 14007 994 14042 1002
rect 12011 981 12046 989
rect 10419 970 10454 971
rect 10212 938 10241 968
rect 12011 961 12019 981
rect 12039 961 12046 981
rect 12011 956 12046 961
rect 12011 955 12043 956
rect 10212 930 10594 938
rect 10212 911 10565 930
rect 10586 911 10594 930
rect 10212 906 10594 911
rect 13389 836 13974 844
rect 13389 816 13398 836
rect 13418 835 13974 836
rect 13418 816 13938 835
rect 13389 815 13938 816
rect 13958 815 13974 835
rect 13389 809 13974 815
rect 9399 752 9407 772
rect 9427 752 9438 772
rect 5245 730 5280 731
rect 6480 683 6531 714
rect 5785 670 5824 683
rect 5785 665 5790 670
rect 5022 648 5790 665
rect 5814 665 5824 670
rect 5814 648 5825 665
rect 5022 640 5825 648
rect 6480 657 6497 683
rect 6525 657 6531 683
rect 5024 639 5310 640
rect 6480 634 6531 657
rect 6560 689 6606 720
rect 8404 718 8447 726
rect 6560 658 6574 689
rect 6602 658 6606 689
rect 6560 651 6606 658
rect 8398 711 8453 718
rect 8398 686 8411 711
rect 8443 686 8453 711
rect 4034 549 4045 581
rect 4085 549 4089 581
rect 4862 623 4923 632
rect 4862 596 4870 623
rect 4906 617 4923 623
rect 4964 617 5039 621
rect 4906 615 5039 617
rect 4906 596 4970 615
rect 4862 579 4970 596
rect 5015 579 5039 615
rect 4862 577 5039 579
rect 4034 536 4089 549
rect 4964 547 5039 577
rect 6493 442 6524 634
rect 6479 421 6525 442
rect 6479 400 6486 421
rect 6507 400 6525 421
rect 6479 396 6525 400
rect 6479 393 6514 396
rect 4618 356 4649 361
rect 2198 294 2204 314
rect 2224 294 2232 314
rect 2198 288 2232 294
rect 3820 336 4654 356
rect 1877 168 1920 172
rect 1877 144 1888 168
rect 1911 144 1920 168
rect 1877 140 1920 144
rect 2094 169 2150 174
rect 2094 149 2101 169
rect 2121 149 2150 169
rect 2094 142 2150 149
rect 2094 141 2129 142
rect 1884 76 1915 140
rect 3820 76 3846 336
rect 4604 334 4650 336
rect 4604 313 4611 334
rect 4632 313 4650 334
rect 4684 326 5777 359
rect 4604 309 4650 313
rect 4604 306 4639 309
rect 3986 148 4571 156
rect 3986 128 3995 148
rect 4015 147 4571 148
rect 4015 128 4535 147
rect 3986 127 4535 128
rect 4555 127 4571 147
rect 3986 121 4571 127
rect 4605 100 4639 306
rect 4686 240 4729 326
rect 4686 220 4693 240
rect 4713 220 4729 240
rect 4686 209 4729 220
rect 4583 95 4639 100
rect 4373 90 4405 95
rect 1884 53 3847 76
rect 1892 51 3847 53
rect 4373 69 4380 90
rect 4397 69 4405 90
rect 4373 62 4405 69
rect 4583 75 4590 95
rect 4610 75 4639 95
rect 4583 68 4639 75
rect 5746 83 5775 326
rect 5861 235 6446 243
rect 5861 215 5870 235
rect 5890 234 6446 235
rect 5890 215 6410 234
rect 5861 214 6410 215
rect 6430 214 6446 234
rect 5861 208 6446 214
rect 6243 188 6286 190
rect 6239 182 6290 188
rect 6480 187 6514 393
rect 6562 327 6596 651
rect 8398 594 8453 686
rect 9399 677 9438 752
rect 9622 770 9678 775
rect 9622 750 9629 770
rect 9649 750 9678 770
rect 9622 743 9678 750
rect 13763 785 13802 789
rect 14008 788 14042 994
rect 14572 1006 14606 1014
rect 14572 988 14579 1006
rect 14598 988 14606 1006
rect 14572 981 14606 988
rect 14783 1011 14839 1016
rect 14783 991 14790 1011
rect 14810 991 14839 1011
rect 14783 984 14839 991
rect 16375 1002 16409 1208
rect 16443 1181 17028 1187
rect 16443 1161 16459 1181
rect 16479 1180 17028 1181
rect 16479 1161 16999 1180
rect 16443 1160 16999 1161
rect 17019 1160 17028 1180
rect 16443 1152 17028 1160
rect 16375 994 16410 1002
rect 14783 983 14818 984
rect 14576 951 14605 981
rect 16375 974 16383 994
rect 16403 974 16410 994
rect 16375 969 16410 974
rect 16375 968 16407 969
rect 14576 943 14958 951
rect 14576 924 14929 943
rect 14950 924 14958 943
rect 14576 919 14958 924
rect 13763 765 13771 785
rect 13791 765 13802 785
rect 9622 742 9657 743
rect 10857 695 10908 726
rect 10162 682 10201 695
rect 10162 677 10167 682
rect 9399 660 10167 677
rect 10191 677 10201 682
rect 10191 660 10202 677
rect 9399 652 10202 660
rect 10857 669 10874 695
rect 10902 669 10908 695
rect 9401 651 9687 652
rect 10857 646 10908 669
rect 10937 701 10983 732
rect 12781 730 12824 738
rect 10937 670 10951 701
rect 10979 670 10983 701
rect 10937 663 10983 670
rect 12775 723 12830 730
rect 12775 698 12788 723
rect 12820 698 12830 723
rect 8398 562 8409 594
rect 8449 562 8453 594
rect 9239 635 9300 644
rect 9239 608 9247 635
rect 9283 629 9300 635
rect 9341 629 9416 633
rect 9283 627 9416 629
rect 9283 608 9347 627
rect 9239 591 9347 608
rect 9392 591 9416 627
rect 9239 589 9416 591
rect 8398 549 8453 562
rect 9341 559 9416 589
rect 10870 454 10901 646
rect 10856 433 10902 454
rect 10856 412 10863 433
rect 10884 412 10902 433
rect 10856 408 10902 412
rect 10856 405 10891 408
rect 9066 380 9097 385
rect 6562 307 6568 327
rect 6588 307 6596 327
rect 6562 301 6596 307
rect 8268 360 9102 380
rect 6239 158 6255 182
rect 6278 158 6290 182
rect 6239 149 6290 158
rect 6458 182 6514 187
rect 6458 162 6465 182
rect 6485 162 6514 182
rect 6458 155 6514 162
rect 6458 154 6493 155
rect 6243 83 6286 149
rect 4583 67 4618 68
rect 4373 2 4401 62
rect 5746 55 6286 83
rect 5749 53 6286 55
rect 6243 51 6286 53
rect 8268 2 8294 360
rect 9052 358 9098 360
rect 9052 337 9059 358
rect 9080 337 9098 358
rect 9132 350 10061 383
rect 9052 333 9098 337
rect 9052 330 9087 333
rect 8434 172 9019 180
rect 8434 152 8443 172
rect 8463 171 9019 172
rect 8463 152 8983 171
rect 8434 151 8983 152
rect 9003 151 9019 171
rect 8434 145 9019 151
rect 9053 124 9087 330
rect 9134 264 9177 350
rect 9261 344 10061 350
rect 9134 244 9141 264
rect 9161 244 9177 264
rect 9134 233 9177 244
rect 9031 119 9087 124
rect 9031 99 9038 119
rect 9058 99 9087 119
rect 9031 92 9087 99
rect 9031 91 9066 92
rect 4373 -32 8299 2
rect 10022 -69 10061 344
rect 10238 247 10823 255
rect 10238 227 10247 247
rect 10267 246 10823 247
rect 10267 227 10787 246
rect 10238 226 10787 227
rect 10807 226 10823 246
rect 10238 220 10823 226
rect 10857 199 10891 405
rect 10939 339 10973 663
rect 12775 606 12830 698
rect 13763 690 13802 765
rect 13986 783 14042 788
rect 13986 763 13993 783
rect 14013 763 14042 783
rect 13986 756 14042 763
rect 13986 755 14021 756
rect 15221 708 15272 739
rect 14526 695 14565 708
rect 14526 690 14531 695
rect 13763 673 14531 690
rect 14555 690 14565 695
rect 14555 673 14566 690
rect 13763 665 14566 673
rect 15221 682 15238 708
rect 15266 682 15272 708
rect 13765 664 14051 665
rect 15221 659 15272 682
rect 15301 714 15347 745
rect 17145 743 17188 751
rect 15301 683 15315 714
rect 15343 683 15347 714
rect 15301 676 15347 683
rect 17139 736 17194 743
rect 17139 711 17152 736
rect 17184 711 17194 736
rect 12775 574 12786 606
rect 12826 574 12830 606
rect 13603 648 13664 657
rect 13603 621 13611 648
rect 13647 642 13664 648
rect 13705 642 13780 646
rect 13647 640 13780 642
rect 13647 621 13711 640
rect 13603 604 13711 621
rect 13756 604 13780 640
rect 13603 602 13780 604
rect 12775 561 12830 574
rect 13705 572 13780 602
rect 15234 467 15265 659
rect 15220 446 15266 467
rect 15220 425 15227 446
rect 15248 425 15266 446
rect 15220 421 15266 425
rect 15220 418 15255 421
rect 13359 381 13390 386
rect 10939 319 10945 339
rect 10965 319 10973 339
rect 10939 313 10973 319
rect 12561 361 13395 381
rect 10618 193 10661 197
rect 10618 169 10629 193
rect 10652 169 10661 193
rect 10618 165 10661 169
rect 10835 194 10891 199
rect 10835 174 10842 194
rect 10862 174 10891 194
rect 10835 167 10891 174
rect 10835 166 10870 167
rect 10625 101 10656 165
rect 12561 101 12587 361
rect 13345 359 13391 361
rect 13345 338 13352 359
rect 13373 338 13391 359
rect 13425 351 14518 384
rect 13345 334 13391 338
rect 13345 331 13380 334
rect 12727 173 13312 181
rect 12727 153 12736 173
rect 12756 172 13312 173
rect 12756 153 13276 172
rect 12727 152 13276 153
rect 13296 152 13312 172
rect 12727 146 13312 152
rect 13346 125 13380 331
rect 13427 265 13470 351
rect 13427 245 13434 265
rect 13454 245 13470 265
rect 13427 234 13470 245
rect 13105 118 13157 124
rect 10625 78 12588 101
rect 10633 76 12588 78
rect 13105 96 13117 118
rect 13138 96 13157 118
rect 13105 -69 13157 96
rect 13324 120 13380 125
rect 13324 100 13331 120
rect 13351 100 13380 120
rect 13324 93 13380 100
rect 14487 108 14516 351
rect 14602 260 15187 268
rect 14602 240 14611 260
rect 14631 259 15187 260
rect 14631 240 15151 259
rect 14602 239 15151 240
rect 15171 239 15187 259
rect 14602 233 15187 239
rect 14984 213 15027 215
rect 14980 207 15031 213
rect 15221 212 15255 418
rect 15303 352 15337 676
rect 17139 619 17194 711
rect 17139 587 17150 619
rect 17190 587 17194 619
rect 17139 574 17194 587
rect 15303 332 15309 352
rect 15329 332 15337 352
rect 15303 326 15337 332
rect 14980 183 14996 207
rect 15019 183 15031 207
rect 14980 174 15031 183
rect 15199 207 15255 212
rect 15199 187 15206 207
rect 15226 187 15255 207
rect 15199 180 15255 187
rect 15199 179 15234 180
rect 14984 108 15027 174
rect 13324 92 13359 93
rect 14487 80 15027 108
rect 14490 78 15027 80
rect 14984 76 15027 78
rect 10022 -113 13157 -69
rect 10022 -115 13102 -113
<< via1 >>
rect 2200 5092 2227 5119
rect 2118 4273 2149 4299
rect 6564 5105 6591 5132
rect 6482 4286 6513 4312
rect 10941 5117 10968 5144
rect 10859 4298 10890 4324
rect 15305 5130 15332 5157
rect 15223 4311 15254 4337
rect 2133 644 2161 670
rect 2210 645 2238 676
rect 606 566 651 602
rect 6497 657 6525 683
rect 6574 658 6602 689
rect 4045 549 4085 581
rect 4970 579 5015 615
rect 10874 669 10902 695
rect 10951 670 10979 701
rect 8409 562 8449 594
rect 9347 591 9392 627
rect 15238 682 15266 708
rect 15315 683 15343 714
rect 12786 574 12826 606
rect 13711 604 13756 640
rect 17150 587 17190 619
<< metal2 >>
rect 15300 5157 15337 5161
rect 10936 5144 10973 5148
rect 6559 5132 6596 5136
rect 2195 5119 2232 5123
rect 2195 5092 2200 5119
rect 2227 5092 2232 5119
rect 6559 5105 6564 5132
rect 6591 5105 6596 5132
rect 10936 5117 10941 5144
rect 10968 5117 10973 5144
rect 15300 5130 15305 5157
rect 15332 5130 15337 5157
rect 15300 5120 15337 5130
rect 10936 5107 10973 5117
rect 6559 5095 6596 5105
rect 2195 5082 2232 5092
rect 2110 4299 2158 4317
rect 2110 4273 2118 4299
rect 2149 4273 2158 4299
rect 2110 4241 2158 4273
rect 2118 695 2158 4241
rect 2199 2345 2225 5082
rect 6474 4312 6522 4330
rect 6474 4286 6482 4312
rect 6513 4286 6522 4312
rect 6474 4254 6522 4286
rect 2197 707 2225 2345
rect 6482 708 6522 4254
rect 6563 2358 6589 5095
rect 10851 4324 10899 4342
rect 10851 4298 10859 4324
rect 10890 4298 10899 4324
rect 10851 4266 10899 4298
rect 6561 720 6589 2358
rect 10859 720 10899 4266
rect 10940 2370 10966 5107
rect 15215 4337 15263 4355
rect 15215 4311 15223 4337
rect 15254 4311 15263 4337
rect 15215 4279 15263 4311
rect 10938 732 10966 2370
rect 15223 733 15263 4279
rect 15304 2383 15330 5120
rect 15302 745 15330 2383
rect 2118 670 2164 695
rect 2118 644 2133 670
rect 2161 644 2164 670
rect 2118 625 2164 644
rect 2196 676 2242 707
rect 2196 645 2210 676
rect 2238 645 2242 676
rect 2196 638 2242 645
rect 6482 683 6528 708
rect 6482 657 6497 683
rect 6525 657 6528 683
rect 6482 638 6528 657
rect 6560 689 6606 720
rect 6560 658 6574 689
rect 6602 658 6606 689
rect 6560 651 6606 658
rect 10859 695 10905 720
rect 10859 669 10874 695
rect 10902 669 10905 695
rect 10859 650 10905 669
rect 10937 701 10983 732
rect 10937 670 10951 701
rect 10979 670 10983 701
rect 10937 663 10983 670
rect 15223 708 15269 733
rect 15223 682 15238 708
rect 15266 682 15269 708
rect 15223 663 15269 682
rect 15301 714 15347 745
rect 15301 683 15315 714
rect 15343 683 15347 714
rect 15301 676 15347 683
rect 15227 659 15269 663
rect 10863 646 10905 650
rect 13697 640 13772 652
rect 6486 634 6528 638
rect 9333 627 9408 639
rect 2122 621 2164 625
rect 4956 615 5031 627
rect 592 602 667 614
rect 592 566 606 602
rect 651 589 667 602
rect 2109 589 2203 594
rect 651 581 4089 589
rect 651 566 4045 581
rect 592 549 4045 566
rect 4085 549 4089 581
rect 4956 579 4970 615
rect 5015 602 5031 615
rect 6473 602 6567 607
rect 5015 594 8453 602
rect 5015 579 8409 594
rect 4956 562 8409 579
rect 8449 562 8453 594
rect 9333 591 9347 627
rect 9392 614 9408 627
rect 10850 614 10944 619
rect 9392 606 12830 614
rect 9392 591 12786 606
rect 9333 574 12786 591
rect 12826 574 12830 606
rect 13697 604 13711 640
rect 13756 627 13772 640
rect 15214 627 15308 632
rect 13756 619 17194 627
rect 13756 604 17150 619
rect 13697 587 17150 604
rect 17190 587 17194 619
rect 13697 578 17194 587
rect 15214 575 15308 578
rect 9333 565 12830 574
rect 10850 562 10944 565
rect 4956 553 8453 562
rect 6473 550 6567 553
rect 592 540 4089 549
rect 2109 537 2203 540
<< labels >>
rlabel locali 3939 128 3962 144 1 d6
rlabel locali 4003 318 4032 324 1 vdd
rlabel locali 4000 19 4029 25 1 gnd
rlabel space 4106 37 4135 46 1 gnd
rlabel nwell 4138 295 4161 298 1 vdd
rlabel locali 5820 218 5835 231 1 d5
rlabel locali 5878 405 5907 411 1 vdd
rlabel locali 5875 106 5904 112 1 gnd
rlabel space 5981 124 6010 133 1 gnd
rlabel nwell 6013 382 6036 385 1 vdd
rlabel locali 8302 1138 8324 1153 5 d0
rlabel locali 8241 959 8270 965 5 vdd
rlabel locali 8244 1258 8273 1264 5 gnd
rlabel space 8138 1237 8167 1246 5 gnd
rlabel nwell 8112 985 8135 988 5 vdd
rlabel locali 8301 1550 8323 1565 5 d0
rlabel locali 8240 1371 8269 1377 5 vdd
rlabel locali 8243 1670 8272 1676 5 gnd
rlabel space 8137 1649 8166 1658 5 gnd
rlabel nwell 8111 1397 8134 1400 5 vdd
rlabel locali 8319 2156 8341 2171 5 d0
rlabel locali 8258 1977 8287 1983 5 vdd
rlabel locali 8261 2276 8290 2282 5 gnd
rlabel space 8155 2255 8184 2264 5 gnd
rlabel nwell 8129 2003 8152 2006 5 vdd
rlabel locali 8318 2568 8340 2583 5 d0
rlabel locali 8257 2389 8286 2395 5 vdd
rlabel locali 8260 2688 8289 2694 5 gnd
rlabel space 8154 2667 8183 2676 5 gnd
rlabel nwell 8128 2415 8151 2418 5 vdd
rlabel locali 7443 1143 7472 1149 5 vdd
rlabel locali 7446 1442 7475 1448 5 gnd
rlabel space 7340 1421 7369 1430 5 gnd
rlabel nwell 7314 1169 7337 1172 5 vdd
rlabel locali 7510 1324 7532 1341 5 d1
rlabel locali 7460 2161 7489 2167 5 vdd
rlabel locali 7463 2460 7492 2466 5 gnd
rlabel space 7357 2439 7386 2448 5 gnd
rlabel nwell 7331 2187 7354 2190 5 vdd
rlabel locali 7527 2342 7549 2359 5 d1
rlabel locali 7361 1751 7390 1757 5 vdd
rlabel locali 7364 2050 7393 2056 5 gnd
rlabel space 7258 2029 7287 2038 5 gnd
rlabel nwell 7232 1777 7255 1780 5 vdd
rlabel locali 7428 1925 7448 1949 5 d2
rlabel locali 8339 3174 8361 3189 5 d0
rlabel locali 8278 2995 8307 3001 5 vdd
rlabel locali 8281 3294 8310 3300 5 gnd
rlabel space 8175 3273 8204 3282 5 gnd
rlabel nwell 8149 3021 8172 3024 5 vdd
rlabel locali 8338 3586 8360 3601 5 d0
rlabel locali 8277 3407 8306 3413 5 vdd
rlabel locali 8280 3706 8309 3712 5 gnd
rlabel space 8174 3685 8203 3694 5 gnd
rlabel nwell 8148 3433 8171 3436 5 vdd
rlabel locali 8356 4192 8378 4207 5 d0
rlabel locali 8295 4013 8324 4019 5 vdd
rlabel locali 8298 4312 8327 4318 5 gnd
rlabel space 8192 4291 8221 4300 5 gnd
rlabel nwell 8166 4039 8189 4042 5 vdd
rlabel locali 8355 4604 8377 4619 5 d0
rlabel locali 8294 4425 8323 4431 5 vdd
rlabel locali 8297 4724 8326 4730 5 gnd
rlabel space 8191 4703 8220 4712 5 gnd
rlabel nwell 8165 4451 8188 4454 5 vdd
rlabel locali 7480 3179 7509 3185 5 vdd
rlabel locali 7483 3478 7512 3484 5 gnd
rlabel space 7377 3457 7406 3466 5 gnd
rlabel nwell 7351 3205 7374 3208 5 vdd
rlabel locali 7547 3360 7569 3377 5 d1
rlabel locali 7497 4197 7526 4203 5 vdd
rlabel locali 7500 4496 7529 4502 5 gnd
rlabel space 7394 4475 7423 4484 5 gnd
rlabel nwell 7368 4223 7391 4226 5 vdd
rlabel locali 7564 4378 7586 4395 5 d1
rlabel locali 7398 3787 7427 3793 5 vdd
rlabel locali 7401 4086 7430 4092 5 gnd
rlabel space 7295 4065 7324 4074 5 gnd
rlabel nwell 7269 3813 7292 3816 5 vdd
rlabel locali 7465 3961 7485 3985 5 d2
rlabel locali 7315 2771 7344 2777 5 vdd
rlabel locali 7318 3070 7347 3076 5 gnd
rlabel space 7212 3049 7241 3058 5 gnd
rlabel nwell 7186 2797 7209 2800 5 vdd
rlabel locali 7380 2950 7400 2963 5 d3
rlabel locali 8375 5210 8397 5225 5 d0
rlabel locali 8314 5031 8343 5037 5 vdd
rlabel locali 8317 5330 8346 5336 5 gnd
rlabel space 8211 5309 8240 5318 5 gnd
rlabel nwell 8185 5057 8208 5060 5 vdd
rlabel locali 8374 5622 8396 5637 5 d0
rlabel locali 8313 5443 8342 5449 5 vdd
rlabel locali 8316 5742 8345 5748 5 gnd
rlabel space 8210 5721 8239 5730 5 gnd
rlabel nwell 8184 5469 8207 5472 5 vdd
rlabel locali 8392 6228 8414 6243 5 d0
rlabel locali 8331 6049 8360 6055 5 vdd
rlabel locali 8334 6348 8363 6354 5 gnd
rlabel space 8228 6327 8257 6336 5 gnd
rlabel nwell 8202 6075 8225 6078 5 vdd
rlabel locali 8391 6640 8413 6655 5 d0
rlabel locali 8330 6461 8359 6467 5 vdd
rlabel locali 8333 6760 8362 6766 5 gnd
rlabel space 8227 6739 8256 6748 5 gnd
rlabel nwell 8201 6487 8224 6490 5 vdd
rlabel locali 7516 5215 7545 5221 5 vdd
rlabel locali 7519 5514 7548 5520 5 gnd
rlabel space 7413 5493 7442 5502 5 gnd
rlabel nwell 7387 5241 7410 5244 5 vdd
rlabel locali 7583 5396 7605 5413 5 d1
rlabel locali 7533 6233 7562 6239 5 vdd
rlabel locali 7536 6532 7565 6538 5 gnd
rlabel space 7430 6511 7459 6520 5 gnd
rlabel nwell 7404 6259 7427 6262 5 vdd
rlabel locali 7600 6414 7622 6431 5 d1
rlabel locali 7434 5823 7463 5829 5 vdd
rlabel locali 7437 6122 7466 6128 5 gnd
rlabel space 7331 6101 7360 6110 5 gnd
rlabel nwell 7305 5849 7328 5852 5 vdd
rlabel locali 7501 5997 7521 6021 5 d2
rlabel locali 8412 7246 8434 7261 5 d0
rlabel locali 8351 7067 8380 7073 5 vdd
rlabel locali 8354 7366 8383 7372 5 gnd
rlabel space 8248 7345 8277 7354 5 gnd
rlabel nwell 8222 7093 8245 7096 5 vdd
rlabel locali 8411 7658 8433 7673 5 d0
rlabel locali 8350 7479 8379 7485 5 vdd
rlabel locali 8353 7778 8382 7784 5 gnd
rlabel space 8247 7757 8276 7766 5 gnd
rlabel nwell 8221 7505 8244 7508 5 vdd
rlabel locali 8429 8264 8451 8279 5 d0
rlabel locali 8368 8085 8397 8091 5 vdd
rlabel locali 8371 8384 8400 8390 5 gnd
rlabel space 8265 8363 8294 8372 5 gnd
rlabel nwell 8239 8111 8262 8114 5 vdd
rlabel locali 8428 8676 8450 8691 5 d0
rlabel locali 8367 8497 8396 8503 5 vdd
rlabel locali 8370 8796 8399 8802 5 gnd
rlabel space 8264 8775 8293 8784 5 gnd
rlabel nwell 8238 8523 8261 8526 5 vdd
rlabel locali 7553 7251 7582 7257 5 vdd
rlabel locali 7556 7550 7585 7556 5 gnd
rlabel space 7450 7529 7479 7538 5 gnd
rlabel nwell 7424 7277 7447 7280 5 vdd
rlabel locali 7620 7432 7642 7449 5 d1
rlabel locali 7570 8269 7599 8275 5 vdd
rlabel locali 7573 8568 7602 8574 5 gnd
rlabel space 7467 8547 7496 8556 5 gnd
rlabel nwell 7441 8295 7464 8298 5 vdd
rlabel locali 7637 8450 7659 8467 5 d1
rlabel locali 7471 7859 7500 7865 5 vdd
rlabel locali 7474 8158 7503 8164 5 gnd
rlabel space 7368 8137 7397 8146 5 gnd
rlabel nwell 7342 7885 7365 7888 5 vdd
rlabel locali 7538 8033 7558 8057 5 d2
rlabel locali 7388 6843 7417 6849 5 vdd
rlabel locali 7391 7142 7420 7148 5 gnd
rlabel space 7285 7121 7314 7130 5 gnd
rlabel nwell 7259 6869 7282 6872 5 vdd
rlabel locali 7453 7022 7473 7035 5 d3
rlabel locali 7212 4809 7241 4815 5 vdd
rlabel locali 7215 5108 7244 5114 5 gnd
rlabel space 7109 5087 7138 5096 5 gnd
rlabel nwell 7083 4835 7106 4838 5 vdd
rlabel locali 7276 4988 7295 5005 5 d4
rlabel locali 5766 4479 5785 4496 1 d4
rlabel nwell 5955 4646 5978 4649 1 vdd
rlabel space 5923 4388 5952 4397 1 gnd
rlabel locali 5817 4370 5846 4376 1 gnd
rlabel locali 5820 4669 5849 4675 1 vdd
rlabel locali 5588 2449 5608 2462 1 d3
rlabel nwell 5779 2612 5802 2615 1 vdd
rlabel space 5747 2354 5776 2363 1 gnd
rlabel locali 5641 2336 5670 2342 1 gnd
rlabel locali 5644 2635 5673 2641 1 vdd
rlabel locali 5503 1427 5523 1451 1 d2
rlabel nwell 5696 1596 5719 1599 1 vdd
rlabel space 5664 1338 5693 1347 1 gnd
rlabel locali 5558 1320 5587 1326 1 gnd
rlabel locali 5561 1619 5590 1625 1 vdd
rlabel locali 5402 1017 5424 1034 1 d1
rlabel nwell 5597 1186 5620 1189 1 vdd
rlabel space 5565 928 5594 937 1 gnd
rlabel locali 5459 910 5488 916 1 gnd
rlabel locali 5462 1209 5491 1215 1 vdd
rlabel locali 5419 2035 5441 2052 1 d1
rlabel nwell 5614 2204 5637 2207 1 vdd
rlabel space 5582 1946 5611 1955 1 gnd
rlabel locali 5476 1928 5505 1934 1 gnd
rlabel locali 5479 2227 5508 2233 1 vdd
rlabel nwell 4800 958 4823 961 1 vdd
rlabel space 4768 700 4797 709 1 gnd
rlabel locali 4662 682 4691 688 1 gnd
rlabel locali 4665 981 4694 987 1 vdd
rlabel locali 4611 793 4633 808 1 d0
rlabel nwell 4799 1370 4822 1373 1 vdd
rlabel space 4767 1112 4796 1121 1 gnd
rlabel locali 4661 1094 4690 1100 1 gnd
rlabel locali 4664 1393 4693 1399 1 vdd
rlabel locali 4610 1205 4632 1220 1 d0
rlabel nwell 4817 1976 4840 1979 1 vdd
rlabel space 4785 1718 4814 1727 1 gnd
rlabel locali 4679 1700 4708 1706 1 gnd
rlabel locali 4682 1999 4711 2005 1 vdd
rlabel locali 4628 1811 4650 1826 1 d0
rlabel nwell 4816 2388 4839 2391 1 vdd
rlabel space 4784 2130 4813 2139 1 gnd
rlabel locali 4678 2112 4707 2118 1 gnd
rlabel locali 4681 2411 4710 2417 1 vdd
rlabel locali 4627 2223 4649 2238 1 d0
rlabel locali 5540 3463 5560 3487 1 d2
rlabel nwell 5733 3632 5756 3635 1 vdd
rlabel space 5701 3374 5730 3383 1 gnd
rlabel locali 5595 3356 5624 3362 1 gnd
rlabel locali 5598 3655 5627 3661 1 vdd
rlabel locali 5439 3053 5461 3070 1 d1
rlabel nwell 5634 3222 5657 3225 1 vdd
rlabel space 5602 2964 5631 2973 1 gnd
rlabel locali 5496 2946 5525 2952 1 gnd
rlabel locali 5499 3245 5528 3251 1 vdd
rlabel locali 5456 4071 5478 4088 1 d1
rlabel nwell 5651 4240 5674 4243 1 vdd
rlabel space 5619 3982 5648 3991 1 gnd
rlabel locali 5513 3964 5542 3970 1 gnd
rlabel locali 5516 4263 5545 4269 1 vdd
rlabel nwell 4837 2994 4860 2997 1 vdd
rlabel space 4805 2736 4834 2745 1 gnd
rlabel locali 4699 2718 4728 2724 1 gnd
rlabel locali 4702 3017 4731 3023 1 vdd
rlabel locali 4648 2829 4670 2844 1 d0
rlabel nwell 4836 3406 4859 3409 1 vdd
rlabel space 4804 3148 4833 3157 1 gnd
rlabel locali 4698 3130 4727 3136 1 gnd
rlabel locali 4701 3429 4730 3435 1 vdd
rlabel locali 4647 3241 4669 3256 1 d0
rlabel nwell 4854 4012 4877 4015 1 vdd
rlabel space 4822 3754 4851 3763 1 gnd
rlabel locali 4716 3736 4745 3742 1 gnd
rlabel locali 4719 4035 4748 4041 1 vdd
rlabel locali 4665 3847 4687 3862 1 d0
rlabel nwell 4853 4424 4876 4427 1 vdd
rlabel space 4821 4166 4850 4175 1 gnd
rlabel locali 4715 4148 4744 4154 1 gnd
rlabel locali 4718 4447 4747 4453 1 vdd
rlabel locali 4664 4259 4686 4274 1 d0
rlabel locali 5661 6521 5681 6534 1 d3
rlabel nwell 5852 6684 5875 6687 1 vdd
rlabel space 5820 6426 5849 6435 1 gnd
rlabel locali 5714 6408 5743 6414 1 gnd
rlabel locali 5717 6707 5746 6713 1 vdd
rlabel locali 5576 5499 5596 5523 1 d2
rlabel nwell 5769 5668 5792 5671 1 vdd
rlabel space 5737 5410 5766 5419 1 gnd
rlabel locali 5631 5392 5660 5398 1 gnd
rlabel locali 5634 5691 5663 5697 1 vdd
rlabel locali 5475 5089 5497 5106 1 d1
rlabel nwell 5670 5258 5693 5261 1 vdd
rlabel space 5638 5000 5667 5009 1 gnd
rlabel locali 5532 4982 5561 4988 1 gnd
rlabel locali 5535 5281 5564 5287 1 vdd
rlabel locali 5492 6107 5514 6124 1 d1
rlabel nwell 5687 6276 5710 6279 1 vdd
rlabel space 5655 6018 5684 6027 1 gnd
rlabel locali 5549 6000 5578 6006 1 gnd
rlabel locali 5552 6299 5581 6305 1 vdd
rlabel nwell 4873 5030 4896 5033 1 vdd
rlabel space 4841 4772 4870 4781 1 gnd
rlabel locali 4735 4754 4764 4760 1 gnd
rlabel locali 4738 5053 4767 5059 1 vdd
rlabel locali 4684 4865 4706 4880 1 d0
rlabel nwell 4872 5442 4895 5445 1 vdd
rlabel space 4840 5184 4869 5193 1 gnd
rlabel locali 4734 5166 4763 5172 1 gnd
rlabel locali 4737 5465 4766 5471 1 vdd
rlabel locali 4683 5277 4705 5292 1 d0
rlabel nwell 4890 6048 4913 6051 1 vdd
rlabel space 4858 5790 4887 5799 1 gnd
rlabel locali 4752 5772 4781 5778 1 gnd
rlabel locali 4755 6071 4784 6077 1 vdd
rlabel locali 4701 5883 4723 5898 1 d0
rlabel nwell 4889 6460 4912 6463 1 vdd
rlabel space 4857 6202 4886 6211 1 gnd
rlabel locali 4751 6184 4780 6190 1 gnd
rlabel locali 4754 6483 4783 6489 1 vdd
rlabel locali 4700 6295 4722 6310 1 d0
rlabel locali 5613 7535 5633 7559 1 d2
rlabel nwell 5806 7704 5829 7707 1 vdd
rlabel space 5774 7446 5803 7455 1 gnd
rlabel locali 5668 7428 5697 7434 1 gnd
rlabel locali 5671 7727 5700 7733 1 vdd
rlabel locali 5512 7125 5534 7142 1 d1
rlabel nwell 5707 7294 5730 7297 1 vdd
rlabel space 5675 7036 5704 7045 1 gnd
rlabel locali 5569 7018 5598 7024 1 gnd
rlabel locali 5572 7317 5601 7323 1 vdd
rlabel locali 5529 8143 5551 8160 1 d1
rlabel nwell 5724 8312 5747 8315 1 vdd
rlabel space 5692 8054 5721 8063 1 gnd
rlabel locali 5586 8036 5615 8042 1 gnd
rlabel locali 5589 8335 5618 8341 1 vdd
rlabel nwell 4910 7066 4933 7069 1 vdd
rlabel space 4878 6808 4907 6817 1 gnd
rlabel locali 4772 6790 4801 6796 1 gnd
rlabel locali 4775 7089 4804 7095 1 vdd
rlabel locali 4721 6901 4743 6916 1 d0
rlabel nwell 4909 7478 4932 7481 1 vdd
rlabel space 4877 7220 4906 7229 1 gnd
rlabel locali 4771 7202 4800 7208 1 gnd
rlabel locali 4774 7501 4803 7507 1 vdd
rlabel locali 4720 7313 4742 7328 1 d0
rlabel nwell 4927 8084 4950 8087 1 vdd
rlabel space 4895 7826 4924 7835 1 gnd
rlabel locali 4789 7808 4818 7814 1 gnd
rlabel locali 4792 8107 4821 8113 1 vdd
rlabel locali 4738 7919 4760 7934 1 d0
rlabel nwell 4926 8496 4949 8499 1 vdd
rlabel space 4894 8238 4923 8247 1 gnd
rlabel locali 4788 8220 4817 8226 1 gnd
rlabel locali 4791 8519 4820 8525 1 vdd
rlabel locali 4737 8331 4759 8346 1 d0
rlabel locali 1456 205 1471 218 1 d5
rlabel locali 1514 392 1543 398 1 vdd
rlabel locali 1511 93 1540 99 1 gnd
rlabel space 1617 111 1646 120 1 gnd
rlabel nwell 1649 369 1672 372 1 vdd
rlabel locali 3938 1125 3960 1140 5 d0
rlabel locali 3877 946 3906 952 5 vdd
rlabel locali 3880 1245 3909 1251 5 gnd
rlabel space 3774 1224 3803 1233 5 gnd
rlabel nwell 3748 972 3771 975 5 vdd
rlabel locali 3937 1537 3959 1552 5 d0
rlabel locali 3876 1358 3905 1364 5 vdd
rlabel locali 3879 1657 3908 1663 5 gnd
rlabel space 3773 1636 3802 1645 5 gnd
rlabel nwell 3747 1384 3770 1387 5 vdd
rlabel locali 3955 2143 3977 2158 5 d0
rlabel locali 3894 1964 3923 1970 5 vdd
rlabel locali 3897 2263 3926 2269 5 gnd
rlabel space 3791 2242 3820 2251 5 gnd
rlabel nwell 3765 1990 3788 1993 5 vdd
rlabel locali 3954 2555 3976 2570 5 d0
rlabel locali 3893 2376 3922 2382 5 vdd
rlabel locali 3896 2675 3925 2681 5 gnd
rlabel space 3790 2654 3819 2663 5 gnd
rlabel nwell 3764 2402 3787 2405 5 vdd
rlabel locali 3079 1130 3108 1136 5 vdd
rlabel locali 3082 1429 3111 1435 5 gnd
rlabel space 2976 1408 3005 1417 5 gnd
rlabel nwell 2950 1156 2973 1159 5 vdd
rlabel locali 3146 1311 3168 1328 5 d1
rlabel locali 3096 2148 3125 2154 5 vdd
rlabel locali 3099 2447 3128 2453 5 gnd
rlabel space 2993 2426 3022 2435 5 gnd
rlabel nwell 2967 2174 2990 2177 5 vdd
rlabel locali 3163 2329 3185 2346 5 d1
rlabel locali 2997 1738 3026 1744 5 vdd
rlabel locali 3000 2037 3029 2043 5 gnd
rlabel space 2894 2016 2923 2025 5 gnd
rlabel nwell 2868 1764 2891 1767 5 vdd
rlabel locali 3064 1912 3084 1936 5 d2
rlabel locali 3975 3161 3997 3176 5 d0
rlabel locali 3914 2982 3943 2988 5 vdd
rlabel locali 3917 3281 3946 3287 5 gnd
rlabel space 3811 3260 3840 3269 5 gnd
rlabel nwell 3785 3008 3808 3011 5 vdd
rlabel locali 3974 3573 3996 3588 5 d0
rlabel locali 3913 3394 3942 3400 5 vdd
rlabel locali 3916 3693 3945 3699 5 gnd
rlabel space 3810 3672 3839 3681 5 gnd
rlabel nwell 3784 3420 3807 3423 5 vdd
rlabel locali 3992 4179 4014 4194 5 d0
rlabel locali 3931 4000 3960 4006 5 vdd
rlabel locali 3934 4299 3963 4305 5 gnd
rlabel space 3828 4278 3857 4287 5 gnd
rlabel nwell 3802 4026 3825 4029 5 vdd
rlabel locali 3991 4591 4013 4606 5 d0
rlabel locali 3930 4412 3959 4418 5 vdd
rlabel locali 3933 4711 3962 4717 5 gnd
rlabel space 3827 4690 3856 4699 5 gnd
rlabel nwell 3801 4438 3824 4441 5 vdd
rlabel locali 3116 3166 3145 3172 5 vdd
rlabel locali 3119 3465 3148 3471 5 gnd
rlabel space 3013 3444 3042 3453 5 gnd
rlabel nwell 2987 3192 3010 3195 5 vdd
rlabel locali 3183 3347 3205 3364 5 d1
rlabel locali 3133 4184 3162 4190 5 vdd
rlabel locali 3136 4483 3165 4489 5 gnd
rlabel space 3030 4462 3059 4471 5 gnd
rlabel nwell 3004 4210 3027 4213 5 vdd
rlabel locali 3200 4365 3222 4382 5 d1
rlabel locali 3034 3774 3063 3780 5 vdd
rlabel locali 3037 4073 3066 4079 5 gnd
rlabel space 2931 4052 2960 4061 5 gnd
rlabel nwell 2905 3800 2928 3803 5 vdd
rlabel locali 3101 3948 3121 3972 5 d2
rlabel locali 2951 2758 2980 2764 5 vdd
rlabel locali 2954 3057 2983 3063 5 gnd
rlabel space 2848 3036 2877 3045 5 gnd
rlabel nwell 2822 2784 2845 2787 5 vdd
rlabel locali 3016 2937 3036 2950 5 d3
rlabel locali 4011 5197 4033 5212 5 d0
rlabel locali 3950 5018 3979 5024 5 vdd
rlabel locali 3953 5317 3982 5323 5 gnd
rlabel space 3847 5296 3876 5305 5 gnd
rlabel nwell 3821 5044 3844 5047 5 vdd
rlabel locali 4010 5609 4032 5624 5 d0
rlabel locali 3949 5430 3978 5436 5 vdd
rlabel locali 3952 5729 3981 5735 5 gnd
rlabel space 3846 5708 3875 5717 5 gnd
rlabel nwell 3820 5456 3843 5459 5 vdd
rlabel locali 4028 6215 4050 6230 5 d0
rlabel locali 3967 6036 3996 6042 5 vdd
rlabel locali 3970 6335 3999 6341 5 gnd
rlabel space 3864 6314 3893 6323 5 gnd
rlabel nwell 3838 6062 3861 6065 5 vdd
rlabel locali 4027 6627 4049 6642 5 d0
rlabel locali 3966 6448 3995 6454 5 vdd
rlabel locali 3969 6747 3998 6753 5 gnd
rlabel space 3863 6726 3892 6735 5 gnd
rlabel nwell 3837 6474 3860 6477 5 vdd
rlabel locali 3152 5202 3181 5208 5 vdd
rlabel locali 3155 5501 3184 5507 5 gnd
rlabel space 3049 5480 3078 5489 5 gnd
rlabel nwell 3023 5228 3046 5231 5 vdd
rlabel locali 3219 5383 3241 5400 5 d1
rlabel locali 3169 6220 3198 6226 5 vdd
rlabel locali 3172 6519 3201 6525 5 gnd
rlabel space 3066 6498 3095 6507 5 gnd
rlabel nwell 3040 6246 3063 6249 5 vdd
rlabel locali 3236 6401 3258 6418 5 d1
rlabel locali 3070 5810 3099 5816 5 vdd
rlabel locali 3073 6109 3102 6115 5 gnd
rlabel space 2967 6088 2996 6097 5 gnd
rlabel nwell 2941 5836 2964 5839 5 vdd
rlabel locali 3137 5984 3157 6008 5 d2
rlabel locali 4048 7233 4070 7248 5 d0
rlabel locali 3987 7054 4016 7060 5 vdd
rlabel locali 3990 7353 4019 7359 5 gnd
rlabel space 3884 7332 3913 7341 5 gnd
rlabel nwell 3858 7080 3881 7083 5 vdd
rlabel locali 4047 7645 4069 7660 5 d0
rlabel locali 3986 7466 4015 7472 5 vdd
rlabel locali 3989 7765 4018 7771 5 gnd
rlabel space 3883 7744 3912 7753 5 gnd
rlabel nwell 3857 7492 3880 7495 5 vdd
rlabel locali 4065 8251 4087 8266 5 d0
rlabel locali 4004 8072 4033 8078 5 vdd
rlabel locali 4007 8371 4036 8377 5 gnd
rlabel space 3901 8350 3930 8359 5 gnd
rlabel nwell 3875 8098 3898 8101 5 vdd
rlabel locali 4064 8663 4086 8678 5 d0
rlabel locali 4003 8484 4032 8490 5 vdd
rlabel locali 4006 8783 4035 8789 5 gnd
rlabel space 3900 8762 3929 8771 5 gnd
rlabel nwell 3874 8510 3897 8513 5 vdd
rlabel locali 3189 7238 3218 7244 5 vdd
rlabel locali 3192 7537 3221 7543 5 gnd
rlabel space 3086 7516 3115 7525 5 gnd
rlabel nwell 3060 7264 3083 7267 5 vdd
rlabel locali 3256 7419 3278 7436 5 d1
rlabel locali 3206 8256 3235 8262 5 vdd
rlabel locali 3209 8555 3238 8561 5 gnd
rlabel space 3103 8534 3132 8543 5 gnd
rlabel nwell 3077 8282 3100 8285 5 vdd
rlabel locali 3273 8437 3295 8454 5 d1
rlabel locali 3107 7846 3136 7852 5 vdd
rlabel locali 3110 8145 3139 8151 5 gnd
rlabel space 3004 8124 3033 8133 5 gnd
rlabel nwell 2978 7872 3001 7875 5 vdd
rlabel locali 3174 8020 3194 8044 5 d2
rlabel locali 3024 6830 3053 6836 5 vdd
rlabel locali 3027 7129 3056 7135 5 gnd
rlabel space 2921 7108 2950 7117 5 gnd
rlabel nwell 2895 6856 2918 6859 5 vdd
rlabel locali 3089 7009 3109 7022 5 d3
rlabel locali 2848 4796 2877 4802 5 vdd
rlabel locali 2851 5095 2880 5101 5 gnd
rlabel space 2745 5074 2774 5083 5 gnd
rlabel nwell 2719 4822 2742 4825 5 vdd
rlabel locali 2912 4975 2931 4992 5 d4
rlabel locali 1402 4466 1421 4483 1 d4
rlabel nwell 1591 4633 1614 4636 1 vdd
rlabel space 1559 4375 1588 4384 1 gnd
rlabel locali 1453 4357 1482 4363 1 gnd
rlabel locali 1456 4656 1485 4662 1 vdd
rlabel locali 1224 2436 1244 2449 1 d3
rlabel nwell 1415 2599 1438 2602 1 vdd
rlabel space 1383 2341 1412 2350 1 gnd
rlabel locali 1277 2323 1306 2329 1 gnd
rlabel locali 1280 2622 1309 2628 1 vdd
rlabel locali 1139 1414 1159 1438 1 d2
rlabel nwell 1332 1583 1355 1586 1 vdd
rlabel space 1300 1325 1329 1334 1 gnd
rlabel locali 1194 1307 1223 1313 1 gnd
rlabel locali 1197 1606 1226 1612 1 vdd
rlabel locali 1038 1004 1060 1021 1 d1
rlabel nwell 1233 1173 1256 1176 1 vdd
rlabel space 1201 915 1230 924 1 gnd
rlabel locali 1095 897 1124 903 1 gnd
rlabel locali 1098 1196 1127 1202 1 vdd
rlabel locali 1055 2022 1077 2039 1 d1
rlabel nwell 1250 2191 1273 2194 1 vdd
rlabel space 1218 1933 1247 1942 1 gnd
rlabel locali 1112 1915 1141 1921 1 gnd
rlabel locali 1115 2214 1144 2220 1 vdd
rlabel nwell 436 945 459 948 1 vdd
rlabel space 404 687 433 696 1 gnd
rlabel locali 298 669 327 675 1 gnd
rlabel locali 301 968 330 974 1 vdd
rlabel locali 247 780 269 795 1 d0
rlabel nwell 435 1357 458 1360 1 vdd
rlabel space 403 1099 432 1108 1 gnd
rlabel locali 297 1081 326 1087 1 gnd
rlabel locali 300 1380 329 1386 1 vdd
rlabel locali 246 1192 268 1207 1 d0
rlabel nwell 453 1963 476 1966 1 vdd
rlabel space 421 1705 450 1714 1 gnd
rlabel locali 315 1687 344 1693 1 gnd
rlabel locali 318 1986 347 1992 1 vdd
rlabel locali 264 1798 286 1813 1 d0
rlabel nwell 452 2375 475 2378 1 vdd
rlabel space 420 2117 449 2126 1 gnd
rlabel locali 314 2099 343 2105 1 gnd
rlabel locali 317 2398 346 2404 1 vdd
rlabel locali 263 2210 285 2225 1 d0
rlabel locali 1176 3450 1196 3474 1 d2
rlabel nwell 1369 3619 1392 3622 1 vdd
rlabel space 1337 3361 1366 3370 1 gnd
rlabel locali 1231 3343 1260 3349 1 gnd
rlabel locali 1234 3642 1263 3648 1 vdd
rlabel locali 1075 3040 1097 3057 1 d1
rlabel nwell 1270 3209 1293 3212 1 vdd
rlabel space 1238 2951 1267 2960 1 gnd
rlabel locali 1132 2933 1161 2939 1 gnd
rlabel locali 1135 3232 1164 3238 1 vdd
rlabel locali 1092 4058 1114 4075 1 d1
rlabel nwell 1287 4227 1310 4230 1 vdd
rlabel space 1255 3969 1284 3978 1 gnd
rlabel locali 1149 3951 1178 3957 1 gnd
rlabel locali 1152 4250 1181 4256 1 vdd
rlabel nwell 473 2981 496 2984 1 vdd
rlabel space 441 2723 470 2732 1 gnd
rlabel locali 335 2705 364 2711 1 gnd
rlabel locali 338 3004 367 3010 1 vdd
rlabel locali 284 2816 306 2831 1 d0
rlabel nwell 472 3393 495 3396 1 vdd
rlabel space 440 3135 469 3144 1 gnd
rlabel locali 334 3117 363 3123 1 gnd
rlabel locali 337 3416 366 3422 1 vdd
rlabel locali 283 3228 305 3243 1 d0
rlabel nwell 490 3999 513 4002 1 vdd
rlabel space 458 3741 487 3750 1 gnd
rlabel locali 352 3723 381 3729 1 gnd
rlabel locali 355 4022 384 4028 1 vdd
rlabel locali 301 3834 323 3849 1 d0
rlabel nwell 489 4411 512 4414 1 vdd
rlabel space 457 4153 486 4162 1 gnd
rlabel locali 351 4135 380 4141 1 gnd
rlabel locali 354 4434 383 4440 1 vdd
rlabel locali 300 4246 322 4261 1 d0
rlabel locali 1297 6508 1317 6521 1 d3
rlabel nwell 1488 6671 1511 6674 1 vdd
rlabel space 1456 6413 1485 6422 1 gnd
rlabel locali 1350 6395 1379 6401 1 gnd
rlabel locali 1353 6694 1382 6700 1 vdd
rlabel locali 1212 5486 1232 5510 1 d2
rlabel nwell 1405 5655 1428 5658 1 vdd
rlabel space 1373 5397 1402 5406 1 gnd
rlabel locali 1267 5379 1296 5385 1 gnd
rlabel locali 1270 5678 1299 5684 1 vdd
rlabel locali 1111 5076 1133 5093 1 d1
rlabel nwell 1306 5245 1329 5248 1 vdd
rlabel space 1274 4987 1303 4996 1 gnd
rlabel locali 1168 4969 1197 4975 1 gnd
rlabel locali 1171 5268 1200 5274 1 vdd
rlabel locali 1128 6094 1150 6111 1 d1
rlabel nwell 1323 6263 1346 6266 1 vdd
rlabel space 1291 6005 1320 6014 1 gnd
rlabel locali 1185 5987 1214 5993 1 gnd
rlabel locali 1188 6286 1217 6292 1 vdd
rlabel nwell 509 5017 532 5020 1 vdd
rlabel space 477 4759 506 4768 1 gnd
rlabel locali 371 4741 400 4747 1 gnd
rlabel locali 374 5040 403 5046 1 vdd
rlabel locali 320 4852 342 4867 1 d0
rlabel nwell 508 5429 531 5432 1 vdd
rlabel space 476 5171 505 5180 1 gnd
rlabel locali 370 5153 399 5159 1 gnd
rlabel locali 373 5452 402 5458 1 vdd
rlabel locali 319 5264 341 5279 1 d0
rlabel nwell 526 6035 549 6038 1 vdd
rlabel space 494 5777 523 5786 1 gnd
rlabel locali 388 5759 417 5765 1 gnd
rlabel locali 391 6058 420 6064 1 vdd
rlabel locali 337 5870 359 5885 1 d0
rlabel nwell 525 6447 548 6450 1 vdd
rlabel space 493 6189 522 6198 1 gnd
rlabel locali 387 6171 416 6177 1 gnd
rlabel locali 390 6470 419 6476 1 vdd
rlabel locali 336 6282 358 6297 1 d0
rlabel locali 1249 7522 1269 7546 1 d2
rlabel nwell 1442 7691 1465 7694 1 vdd
rlabel space 1410 7433 1439 7442 1 gnd
rlabel locali 1304 7415 1333 7421 1 gnd
rlabel locali 1307 7714 1336 7720 1 vdd
rlabel locali 1148 7112 1170 7129 1 d1
rlabel nwell 1343 7281 1366 7284 1 vdd
rlabel space 1311 7023 1340 7032 1 gnd
rlabel locali 1205 7005 1234 7011 1 gnd
rlabel locali 1208 7304 1237 7310 1 vdd
rlabel locali 1165 8130 1187 8147 1 d1
rlabel nwell 1360 8299 1383 8302 1 vdd
rlabel space 1328 8041 1357 8050 1 gnd
rlabel locali 1222 8023 1251 8029 1 gnd
rlabel locali 1225 8322 1254 8328 1 vdd
rlabel nwell 546 7053 569 7056 1 vdd
rlabel space 514 6795 543 6804 1 gnd
rlabel locali 408 6777 437 6783 1 gnd
rlabel locali 411 7076 440 7082 1 vdd
rlabel locali 357 6888 379 6903 1 d0
rlabel nwell 545 7465 568 7468 1 vdd
rlabel space 513 7207 542 7216 1 gnd
rlabel locali 407 7189 436 7195 1 gnd
rlabel locali 410 7488 439 7494 1 vdd
rlabel locali 356 7300 378 7315 1 d0
rlabel locali 264 8751 288 8781 1 vref
rlabel nwell 563 8071 586 8074 1 vdd
rlabel space 531 7813 560 7822 1 gnd
rlabel locali 425 7795 454 7801 1 gnd
rlabel locali 428 8094 457 8100 1 vdd
rlabel locali 374 7906 396 7921 1 d0
rlabel nwell 562 8483 585 8486 1 vdd
rlabel space 530 8225 559 8234 1 gnd
rlabel locali 424 8207 453 8213 1 gnd
rlabel locali 427 8506 456 8512 1 vdd
rlabel locali 373 8318 395 8333 1 d0
rlabel locali 12680 153 12703 169 1 d6
rlabel locali 12744 343 12773 349 1 vdd
rlabel locali 12741 44 12770 50 1 gnd
rlabel space 12847 62 12876 71 1 gnd
rlabel nwell 12879 320 12902 323 1 vdd
rlabel locali 14561 243 14576 256 1 d5
rlabel locali 14619 430 14648 436 1 vdd
rlabel locali 14616 131 14645 137 1 gnd
rlabel space 14722 149 14751 158 1 gnd
rlabel nwell 14754 407 14777 410 1 vdd
rlabel locali 17043 1163 17065 1178 5 d0
rlabel locali 16982 984 17011 990 5 vdd
rlabel locali 16985 1283 17014 1289 5 gnd
rlabel space 16879 1262 16908 1271 5 gnd
rlabel nwell 16853 1010 16876 1013 5 vdd
rlabel locali 17042 1575 17064 1590 5 d0
rlabel locali 16981 1396 17010 1402 5 vdd
rlabel locali 16984 1695 17013 1701 5 gnd
rlabel space 16878 1674 16907 1683 5 gnd
rlabel nwell 16852 1422 16875 1425 5 vdd
rlabel locali 17060 2181 17082 2196 5 d0
rlabel locali 16999 2002 17028 2008 5 vdd
rlabel locali 17002 2301 17031 2307 5 gnd
rlabel space 16896 2280 16925 2289 5 gnd
rlabel nwell 16870 2028 16893 2031 5 vdd
rlabel locali 17059 2593 17081 2608 5 d0
rlabel locali 16998 2414 17027 2420 5 vdd
rlabel locali 17001 2713 17030 2719 5 gnd
rlabel space 16895 2692 16924 2701 5 gnd
rlabel nwell 16869 2440 16892 2443 5 vdd
rlabel locali 16184 1168 16213 1174 5 vdd
rlabel locali 16187 1467 16216 1473 5 gnd
rlabel space 16081 1446 16110 1455 5 gnd
rlabel nwell 16055 1194 16078 1197 5 vdd
rlabel locali 16251 1349 16273 1366 5 d1
rlabel locali 16201 2186 16230 2192 5 vdd
rlabel locali 16204 2485 16233 2491 5 gnd
rlabel space 16098 2464 16127 2473 5 gnd
rlabel nwell 16072 2212 16095 2215 5 vdd
rlabel locali 16268 2367 16290 2384 5 d1
rlabel locali 16102 1776 16131 1782 5 vdd
rlabel locali 16105 2075 16134 2081 5 gnd
rlabel space 15999 2054 16028 2063 5 gnd
rlabel nwell 15973 1802 15996 1805 5 vdd
rlabel locali 16169 1950 16189 1974 5 d2
rlabel locali 17080 3199 17102 3214 5 d0
rlabel locali 17019 3020 17048 3026 5 vdd
rlabel locali 17022 3319 17051 3325 5 gnd
rlabel space 16916 3298 16945 3307 5 gnd
rlabel nwell 16890 3046 16913 3049 5 vdd
rlabel locali 17079 3611 17101 3626 5 d0
rlabel locali 17018 3432 17047 3438 5 vdd
rlabel locali 17021 3731 17050 3737 5 gnd
rlabel space 16915 3710 16944 3719 5 gnd
rlabel nwell 16889 3458 16912 3461 5 vdd
rlabel locali 17097 4217 17119 4232 5 d0
rlabel locali 17036 4038 17065 4044 5 vdd
rlabel locali 17039 4337 17068 4343 5 gnd
rlabel space 16933 4316 16962 4325 5 gnd
rlabel nwell 16907 4064 16930 4067 5 vdd
rlabel locali 17096 4629 17118 4644 5 d0
rlabel locali 17035 4450 17064 4456 5 vdd
rlabel locali 17038 4749 17067 4755 5 gnd
rlabel space 16932 4728 16961 4737 5 gnd
rlabel nwell 16906 4476 16929 4479 5 vdd
rlabel locali 16221 3204 16250 3210 5 vdd
rlabel locali 16224 3503 16253 3509 5 gnd
rlabel space 16118 3482 16147 3491 5 gnd
rlabel nwell 16092 3230 16115 3233 5 vdd
rlabel locali 16288 3385 16310 3402 5 d1
rlabel locali 16238 4222 16267 4228 5 vdd
rlabel locali 16241 4521 16270 4527 5 gnd
rlabel space 16135 4500 16164 4509 5 gnd
rlabel nwell 16109 4248 16132 4251 5 vdd
rlabel locali 16305 4403 16327 4420 5 d1
rlabel locali 16139 3812 16168 3818 5 vdd
rlabel locali 16142 4111 16171 4117 5 gnd
rlabel space 16036 4090 16065 4099 5 gnd
rlabel nwell 16010 3838 16033 3841 5 vdd
rlabel locali 16206 3986 16226 4010 5 d2
rlabel locali 16056 2796 16085 2802 5 vdd
rlabel locali 16059 3095 16088 3101 5 gnd
rlabel space 15953 3074 15982 3083 5 gnd
rlabel nwell 15927 2822 15950 2825 5 vdd
rlabel locali 16121 2975 16141 2988 5 d3
rlabel locali 17116 5235 17138 5250 5 d0
rlabel locali 17055 5056 17084 5062 5 vdd
rlabel locali 17058 5355 17087 5361 5 gnd
rlabel space 16952 5334 16981 5343 5 gnd
rlabel nwell 16926 5082 16949 5085 5 vdd
rlabel locali 17115 5647 17137 5662 5 d0
rlabel locali 17054 5468 17083 5474 5 vdd
rlabel locali 17057 5767 17086 5773 5 gnd
rlabel space 16951 5746 16980 5755 5 gnd
rlabel nwell 16925 5494 16948 5497 5 vdd
rlabel locali 17133 6253 17155 6268 5 d0
rlabel locali 17072 6074 17101 6080 5 vdd
rlabel locali 17075 6373 17104 6379 5 gnd
rlabel space 16969 6352 16998 6361 5 gnd
rlabel nwell 16943 6100 16966 6103 5 vdd
rlabel locali 17132 6665 17154 6680 5 d0
rlabel locali 17071 6486 17100 6492 5 vdd
rlabel locali 17074 6785 17103 6791 5 gnd
rlabel space 16968 6764 16997 6773 5 gnd
rlabel nwell 16942 6512 16965 6515 5 vdd
rlabel locali 16257 5240 16286 5246 5 vdd
rlabel locali 16260 5539 16289 5545 5 gnd
rlabel space 16154 5518 16183 5527 5 gnd
rlabel nwell 16128 5266 16151 5269 5 vdd
rlabel locali 16324 5421 16346 5438 5 d1
rlabel locali 16274 6258 16303 6264 5 vdd
rlabel locali 16277 6557 16306 6563 5 gnd
rlabel space 16171 6536 16200 6545 5 gnd
rlabel nwell 16145 6284 16168 6287 5 vdd
rlabel locali 16341 6439 16363 6456 5 d1
rlabel locali 16175 5848 16204 5854 5 vdd
rlabel locali 16178 6147 16207 6153 5 gnd
rlabel space 16072 6126 16101 6135 5 gnd
rlabel nwell 16046 5874 16069 5877 5 vdd
rlabel locali 16242 6022 16262 6046 5 d2
rlabel locali 17153 7271 17175 7286 5 d0
rlabel locali 17092 7092 17121 7098 5 vdd
rlabel locali 17095 7391 17124 7397 5 gnd
rlabel space 16989 7370 17018 7379 5 gnd
rlabel nwell 16963 7118 16986 7121 5 vdd
rlabel locali 17152 7683 17174 7698 5 d0
rlabel locali 17091 7504 17120 7510 5 vdd
rlabel locali 17094 7803 17123 7809 5 gnd
rlabel space 16988 7782 17017 7791 5 gnd
rlabel nwell 16962 7530 16985 7533 5 vdd
rlabel locali 17170 8289 17192 8304 5 d0
rlabel locali 17109 8110 17138 8116 5 vdd
rlabel locali 17112 8409 17141 8415 5 gnd
rlabel space 17006 8388 17035 8397 5 gnd
rlabel nwell 16980 8136 17003 8139 5 vdd
rlabel locali 17169 8701 17191 8716 5 d0
rlabel locali 17108 8522 17137 8528 5 vdd
rlabel locali 17111 8821 17140 8827 5 gnd
rlabel space 17005 8800 17034 8809 5 gnd
rlabel nwell 16979 8548 17002 8551 5 vdd
rlabel locali 17297 8810 17325 8828 5 gnd
rlabel locali 16294 7276 16323 7282 5 vdd
rlabel locali 16297 7575 16326 7581 5 gnd
rlabel space 16191 7554 16220 7563 5 gnd
rlabel nwell 16165 7302 16188 7305 5 vdd
rlabel locali 16361 7457 16383 7474 5 d1
rlabel locali 16311 8294 16340 8300 5 vdd
rlabel locali 16314 8593 16343 8599 5 gnd
rlabel space 16208 8572 16237 8581 5 gnd
rlabel nwell 16182 8320 16205 8323 5 vdd
rlabel locali 16378 8475 16400 8492 5 d1
rlabel locali 16212 7884 16241 7890 5 vdd
rlabel locali 16215 8183 16244 8189 5 gnd
rlabel space 16109 8162 16138 8171 5 gnd
rlabel nwell 16083 7910 16106 7913 5 vdd
rlabel locali 16279 8058 16299 8082 5 d2
rlabel locali 16129 6868 16158 6874 5 vdd
rlabel locali 16132 7167 16161 7173 5 gnd
rlabel space 16026 7146 16055 7155 5 gnd
rlabel nwell 16000 6894 16023 6897 5 vdd
rlabel locali 16194 7047 16214 7060 5 d3
rlabel locali 15953 4834 15982 4840 5 vdd
rlabel locali 15956 5133 15985 5139 5 gnd
rlabel space 15850 5112 15879 5121 5 gnd
rlabel nwell 15824 4860 15847 4863 5 vdd
rlabel locali 16017 5013 16036 5030 5 d4
rlabel locali 14507 4504 14526 4521 1 d4
rlabel nwell 14696 4671 14719 4674 1 vdd
rlabel space 14664 4413 14693 4422 1 gnd
rlabel locali 14558 4395 14587 4401 1 gnd
rlabel locali 14561 4694 14590 4700 1 vdd
rlabel locali 14329 2474 14349 2487 1 d3
rlabel nwell 14520 2637 14543 2640 1 vdd
rlabel space 14488 2379 14517 2388 1 gnd
rlabel locali 14382 2361 14411 2367 1 gnd
rlabel locali 14385 2660 14414 2666 1 vdd
rlabel locali 14244 1452 14264 1476 1 d2
rlabel nwell 14437 1621 14460 1624 1 vdd
rlabel space 14405 1363 14434 1372 1 gnd
rlabel locali 14299 1345 14328 1351 1 gnd
rlabel locali 14302 1644 14331 1650 1 vdd
rlabel locali 14143 1042 14165 1059 1 d1
rlabel nwell 14338 1211 14361 1214 1 vdd
rlabel space 14306 953 14335 962 1 gnd
rlabel locali 14200 935 14229 941 1 gnd
rlabel locali 14203 1234 14232 1240 1 vdd
rlabel locali 14160 2060 14182 2077 1 d1
rlabel nwell 14355 2229 14378 2232 1 vdd
rlabel space 14323 1971 14352 1980 1 gnd
rlabel locali 14217 1953 14246 1959 1 gnd
rlabel locali 14220 2252 14249 2258 1 vdd
rlabel nwell 13541 983 13564 986 1 vdd
rlabel space 13509 725 13538 734 1 gnd
rlabel locali 13403 707 13432 713 1 gnd
rlabel locali 13406 1006 13435 1012 1 vdd
rlabel locali 13352 818 13374 833 1 d0
rlabel nwell 13540 1395 13563 1398 1 vdd
rlabel space 13508 1137 13537 1146 1 gnd
rlabel locali 13402 1119 13431 1125 1 gnd
rlabel locali 13405 1418 13434 1424 1 vdd
rlabel locali 13351 1230 13373 1245 1 d0
rlabel nwell 13558 2001 13581 2004 1 vdd
rlabel space 13526 1743 13555 1752 1 gnd
rlabel locali 13420 1725 13449 1731 1 gnd
rlabel locali 13423 2024 13452 2030 1 vdd
rlabel locali 13369 1836 13391 1851 1 d0
rlabel nwell 13557 2413 13580 2416 1 vdd
rlabel space 13525 2155 13554 2164 1 gnd
rlabel locali 13419 2137 13448 2143 1 gnd
rlabel locali 13422 2436 13451 2442 1 vdd
rlabel locali 13368 2248 13390 2263 1 d0
rlabel locali 14281 3488 14301 3512 1 d2
rlabel nwell 14474 3657 14497 3660 1 vdd
rlabel space 14442 3399 14471 3408 1 gnd
rlabel locali 14336 3381 14365 3387 1 gnd
rlabel locali 14339 3680 14368 3686 1 vdd
rlabel locali 14180 3078 14202 3095 1 d1
rlabel nwell 14375 3247 14398 3250 1 vdd
rlabel space 14343 2989 14372 2998 1 gnd
rlabel locali 14237 2971 14266 2977 1 gnd
rlabel locali 14240 3270 14269 3276 1 vdd
rlabel locali 14197 4096 14219 4113 1 d1
rlabel nwell 14392 4265 14415 4268 1 vdd
rlabel space 14360 4007 14389 4016 1 gnd
rlabel locali 14254 3989 14283 3995 1 gnd
rlabel locali 14257 4288 14286 4294 1 vdd
rlabel nwell 13578 3019 13601 3022 1 vdd
rlabel space 13546 2761 13575 2770 1 gnd
rlabel locali 13440 2743 13469 2749 1 gnd
rlabel locali 13443 3042 13472 3048 1 vdd
rlabel locali 13389 2854 13411 2869 1 d0
rlabel nwell 13577 3431 13600 3434 1 vdd
rlabel space 13545 3173 13574 3182 1 gnd
rlabel locali 13439 3155 13468 3161 1 gnd
rlabel locali 13442 3454 13471 3460 1 vdd
rlabel locali 13388 3266 13410 3281 1 d0
rlabel nwell 13595 4037 13618 4040 1 vdd
rlabel space 13563 3779 13592 3788 1 gnd
rlabel locali 13457 3761 13486 3767 1 gnd
rlabel locali 13460 4060 13489 4066 1 vdd
rlabel locali 13406 3872 13428 3887 1 d0
rlabel nwell 13594 4449 13617 4452 1 vdd
rlabel space 13562 4191 13591 4200 1 gnd
rlabel locali 13456 4173 13485 4179 1 gnd
rlabel locali 13459 4472 13488 4478 1 vdd
rlabel locali 13405 4284 13427 4299 1 d0
rlabel locali 14402 6546 14422 6559 1 d3
rlabel nwell 14593 6709 14616 6712 1 vdd
rlabel space 14561 6451 14590 6460 1 gnd
rlabel locali 14455 6433 14484 6439 1 gnd
rlabel locali 14458 6732 14487 6738 1 vdd
rlabel locali 14317 5524 14337 5548 1 d2
rlabel nwell 14510 5693 14533 5696 1 vdd
rlabel space 14478 5435 14507 5444 1 gnd
rlabel locali 14372 5417 14401 5423 1 gnd
rlabel locali 14375 5716 14404 5722 1 vdd
rlabel locali 14216 5114 14238 5131 1 d1
rlabel nwell 14411 5283 14434 5286 1 vdd
rlabel space 14379 5025 14408 5034 1 gnd
rlabel locali 14273 5007 14302 5013 1 gnd
rlabel locali 14276 5306 14305 5312 1 vdd
rlabel locali 14233 6132 14255 6149 1 d1
rlabel nwell 14428 6301 14451 6304 1 vdd
rlabel space 14396 6043 14425 6052 1 gnd
rlabel locali 14290 6025 14319 6031 1 gnd
rlabel locali 14293 6324 14322 6330 1 vdd
rlabel nwell 13614 5055 13637 5058 1 vdd
rlabel space 13582 4797 13611 4806 1 gnd
rlabel locali 13476 4779 13505 4785 1 gnd
rlabel locali 13479 5078 13508 5084 1 vdd
rlabel locali 13425 4890 13447 4905 1 d0
rlabel nwell 13613 5467 13636 5470 1 vdd
rlabel space 13581 5209 13610 5218 1 gnd
rlabel locali 13475 5191 13504 5197 1 gnd
rlabel locali 13478 5490 13507 5496 1 vdd
rlabel locali 13424 5302 13446 5317 1 d0
rlabel nwell 13631 6073 13654 6076 1 vdd
rlabel space 13599 5815 13628 5824 1 gnd
rlabel locali 13493 5797 13522 5803 1 gnd
rlabel locali 13496 6096 13525 6102 1 vdd
rlabel locali 13442 5908 13464 5923 1 d0
rlabel nwell 13630 6485 13653 6488 1 vdd
rlabel space 13598 6227 13627 6236 1 gnd
rlabel locali 13492 6209 13521 6215 1 gnd
rlabel locali 13495 6508 13524 6514 1 vdd
rlabel locali 13441 6320 13463 6335 1 d0
rlabel locali 14354 7560 14374 7584 1 d2
rlabel nwell 14547 7729 14570 7732 1 vdd
rlabel space 14515 7471 14544 7480 1 gnd
rlabel locali 14409 7453 14438 7459 1 gnd
rlabel locali 14412 7752 14441 7758 1 vdd
rlabel locali 14253 7150 14275 7167 1 d1
rlabel nwell 14448 7319 14471 7322 1 vdd
rlabel space 14416 7061 14445 7070 1 gnd
rlabel locali 14310 7043 14339 7049 1 gnd
rlabel locali 14313 7342 14342 7348 1 vdd
rlabel locali 14270 8168 14292 8185 1 d1
rlabel nwell 14465 8337 14488 8340 1 vdd
rlabel space 14433 8079 14462 8088 1 gnd
rlabel locali 14327 8061 14356 8067 1 gnd
rlabel locali 14330 8360 14359 8366 1 vdd
rlabel nwell 13651 7091 13674 7094 1 vdd
rlabel space 13619 6833 13648 6842 1 gnd
rlabel locali 13513 6815 13542 6821 1 gnd
rlabel locali 13516 7114 13545 7120 1 vdd
rlabel locali 13462 6926 13484 6941 1 d0
rlabel nwell 13650 7503 13673 7506 1 vdd
rlabel space 13618 7245 13647 7254 1 gnd
rlabel locali 13512 7227 13541 7233 1 gnd
rlabel locali 13515 7526 13544 7532 1 vdd
rlabel locali 13461 7338 13483 7353 1 d0
rlabel nwell 13668 8109 13691 8112 1 vdd
rlabel space 13636 7851 13665 7860 1 gnd
rlabel locali 13530 7833 13559 7839 1 gnd
rlabel locali 13533 8132 13562 8138 1 vdd
rlabel locali 13479 7944 13501 7959 1 d0
rlabel nwell 13667 8521 13690 8524 1 vdd
rlabel space 13635 8263 13664 8272 1 gnd
rlabel locali 13529 8245 13558 8251 1 gnd
rlabel locali 13532 8544 13561 8550 1 vdd
rlabel locali 13478 8356 13500 8371 1 d0
rlabel locali 10197 230 10212 243 1 d5
rlabel locali 10255 417 10284 423 1 vdd
rlabel locali 10252 118 10281 124 1 gnd
rlabel space 10358 136 10387 145 1 gnd
rlabel nwell 10390 394 10413 397 1 vdd
rlabel locali 12679 1150 12701 1165 5 d0
rlabel locali 12618 971 12647 977 5 vdd
rlabel locali 12621 1270 12650 1276 5 gnd
rlabel space 12515 1249 12544 1258 5 gnd
rlabel nwell 12489 997 12512 1000 5 vdd
rlabel locali 12678 1562 12700 1577 5 d0
rlabel locali 12617 1383 12646 1389 5 vdd
rlabel locali 12620 1682 12649 1688 5 gnd
rlabel space 12514 1661 12543 1670 5 gnd
rlabel nwell 12488 1409 12511 1412 5 vdd
rlabel locali 12696 2168 12718 2183 5 d0
rlabel locali 12635 1989 12664 1995 5 vdd
rlabel locali 12638 2288 12667 2294 5 gnd
rlabel space 12532 2267 12561 2276 5 gnd
rlabel nwell 12506 2015 12529 2018 5 vdd
rlabel locali 12695 2580 12717 2595 5 d0
rlabel locali 12634 2401 12663 2407 5 vdd
rlabel locali 12637 2700 12666 2706 5 gnd
rlabel space 12531 2679 12560 2688 5 gnd
rlabel nwell 12505 2427 12528 2430 5 vdd
rlabel locali 11820 1155 11849 1161 5 vdd
rlabel locali 11823 1454 11852 1460 5 gnd
rlabel space 11717 1433 11746 1442 5 gnd
rlabel nwell 11691 1181 11714 1184 5 vdd
rlabel locali 11887 1336 11909 1353 5 d1
rlabel locali 11837 2173 11866 2179 5 vdd
rlabel locali 11840 2472 11869 2478 5 gnd
rlabel space 11734 2451 11763 2460 5 gnd
rlabel nwell 11708 2199 11731 2202 5 vdd
rlabel locali 11904 2354 11926 2371 5 d1
rlabel locali 11738 1763 11767 1769 5 vdd
rlabel locali 11741 2062 11770 2068 5 gnd
rlabel space 11635 2041 11664 2050 5 gnd
rlabel nwell 11609 1789 11632 1792 5 vdd
rlabel locali 11805 1937 11825 1961 5 d2
rlabel locali 12716 3186 12738 3201 5 d0
rlabel locali 12655 3007 12684 3013 5 vdd
rlabel locali 12658 3306 12687 3312 5 gnd
rlabel space 12552 3285 12581 3294 5 gnd
rlabel nwell 12526 3033 12549 3036 5 vdd
rlabel locali 12715 3598 12737 3613 5 d0
rlabel locali 12654 3419 12683 3425 5 vdd
rlabel locali 12657 3718 12686 3724 5 gnd
rlabel space 12551 3697 12580 3706 5 gnd
rlabel nwell 12525 3445 12548 3448 5 vdd
rlabel locali 12733 4204 12755 4219 5 d0
rlabel locali 12672 4025 12701 4031 5 vdd
rlabel locali 12675 4324 12704 4330 5 gnd
rlabel space 12569 4303 12598 4312 5 gnd
rlabel nwell 12543 4051 12566 4054 5 vdd
rlabel locali 12732 4616 12754 4631 5 d0
rlabel locali 12671 4437 12700 4443 5 vdd
rlabel locali 12674 4736 12703 4742 5 gnd
rlabel space 12568 4715 12597 4724 5 gnd
rlabel nwell 12542 4463 12565 4466 5 vdd
rlabel locali 11857 3191 11886 3197 5 vdd
rlabel locali 11860 3490 11889 3496 5 gnd
rlabel space 11754 3469 11783 3478 5 gnd
rlabel nwell 11728 3217 11751 3220 5 vdd
rlabel locali 11924 3372 11946 3389 5 d1
rlabel locali 11874 4209 11903 4215 5 vdd
rlabel locali 11877 4508 11906 4514 5 gnd
rlabel space 11771 4487 11800 4496 5 gnd
rlabel nwell 11745 4235 11768 4238 5 vdd
rlabel locali 11941 4390 11963 4407 5 d1
rlabel locali 11775 3799 11804 3805 5 vdd
rlabel locali 11778 4098 11807 4104 5 gnd
rlabel space 11672 4077 11701 4086 5 gnd
rlabel nwell 11646 3825 11669 3828 5 vdd
rlabel locali 11842 3973 11862 3997 5 d2
rlabel locali 11692 2783 11721 2789 5 vdd
rlabel locali 11695 3082 11724 3088 5 gnd
rlabel space 11589 3061 11618 3070 5 gnd
rlabel nwell 11563 2809 11586 2812 5 vdd
rlabel locali 11757 2962 11777 2975 5 d3
rlabel locali 12752 5222 12774 5237 5 d0
rlabel locali 12691 5043 12720 5049 5 vdd
rlabel locali 12694 5342 12723 5348 5 gnd
rlabel space 12588 5321 12617 5330 5 gnd
rlabel nwell 12562 5069 12585 5072 5 vdd
rlabel locali 12751 5634 12773 5649 5 d0
rlabel locali 12690 5455 12719 5461 5 vdd
rlabel locali 12693 5754 12722 5760 5 gnd
rlabel space 12587 5733 12616 5742 5 gnd
rlabel nwell 12561 5481 12584 5484 5 vdd
rlabel locali 12769 6240 12791 6255 5 d0
rlabel locali 12708 6061 12737 6067 5 vdd
rlabel locali 12711 6360 12740 6366 5 gnd
rlabel space 12605 6339 12634 6348 5 gnd
rlabel nwell 12579 6087 12602 6090 5 vdd
rlabel locali 12768 6652 12790 6667 5 d0
rlabel locali 12707 6473 12736 6479 5 vdd
rlabel locali 12710 6772 12739 6778 5 gnd
rlabel space 12604 6751 12633 6760 5 gnd
rlabel nwell 12578 6499 12601 6502 5 vdd
rlabel locali 11893 5227 11922 5233 5 vdd
rlabel locali 11896 5526 11925 5532 5 gnd
rlabel space 11790 5505 11819 5514 5 gnd
rlabel nwell 11764 5253 11787 5256 5 vdd
rlabel locali 11960 5408 11982 5425 5 d1
rlabel locali 11910 6245 11939 6251 5 vdd
rlabel locali 11913 6544 11942 6550 5 gnd
rlabel space 11807 6523 11836 6532 5 gnd
rlabel nwell 11781 6271 11804 6274 5 vdd
rlabel locali 11977 6426 11999 6443 5 d1
rlabel locali 11811 5835 11840 5841 5 vdd
rlabel locali 11814 6134 11843 6140 5 gnd
rlabel space 11708 6113 11737 6122 5 gnd
rlabel nwell 11682 5861 11705 5864 5 vdd
rlabel locali 11878 6009 11898 6033 5 d2
rlabel locali 12789 7258 12811 7273 5 d0
rlabel locali 12728 7079 12757 7085 5 vdd
rlabel locali 12731 7378 12760 7384 5 gnd
rlabel space 12625 7357 12654 7366 5 gnd
rlabel nwell 12599 7105 12622 7108 5 vdd
rlabel locali 12788 7670 12810 7685 5 d0
rlabel locali 12727 7491 12756 7497 5 vdd
rlabel locali 12730 7790 12759 7796 5 gnd
rlabel space 12624 7769 12653 7778 5 gnd
rlabel nwell 12598 7517 12621 7520 5 vdd
rlabel locali 12806 8276 12828 8291 5 d0
rlabel locali 12745 8097 12774 8103 5 vdd
rlabel locali 12748 8396 12777 8402 5 gnd
rlabel space 12642 8375 12671 8384 5 gnd
rlabel nwell 12616 8123 12639 8126 5 vdd
rlabel locali 12805 8688 12827 8703 5 d0
rlabel locali 12744 8509 12773 8515 5 vdd
rlabel locali 12747 8808 12776 8814 5 gnd
rlabel space 12641 8787 12670 8796 5 gnd
rlabel nwell 12615 8535 12638 8538 5 vdd
rlabel locali 11930 7263 11959 7269 5 vdd
rlabel locali 11933 7562 11962 7568 5 gnd
rlabel space 11827 7541 11856 7550 5 gnd
rlabel nwell 11801 7289 11824 7292 5 vdd
rlabel locali 11997 7444 12019 7461 5 d1
rlabel locali 11947 8281 11976 8287 5 vdd
rlabel locali 11950 8580 11979 8586 5 gnd
rlabel space 11844 8559 11873 8568 5 gnd
rlabel nwell 11818 8307 11841 8310 5 vdd
rlabel locali 12014 8462 12036 8479 5 d1
rlabel locali 11848 7871 11877 7877 5 vdd
rlabel locali 11851 8170 11880 8176 5 gnd
rlabel space 11745 8149 11774 8158 5 gnd
rlabel nwell 11719 7897 11742 7900 5 vdd
rlabel locali 11915 8045 11935 8069 5 d2
rlabel locali 11765 6855 11794 6861 5 vdd
rlabel locali 11768 7154 11797 7160 5 gnd
rlabel space 11662 7133 11691 7142 5 gnd
rlabel nwell 11636 6881 11659 6884 5 vdd
rlabel locali 11830 7034 11850 7047 5 d3
rlabel locali 11589 4821 11618 4827 5 vdd
rlabel locali 11592 5120 11621 5126 5 gnd
rlabel space 11486 5099 11515 5108 5 gnd
rlabel nwell 11460 4847 11483 4850 5 vdd
rlabel locali 11653 5000 11672 5017 5 d4
rlabel locali 10143 4491 10162 4508 1 d4
rlabel nwell 10332 4658 10355 4661 1 vdd
rlabel space 10300 4400 10329 4409 1 gnd
rlabel locali 10194 4382 10223 4388 1 gnd
rlabel locali 10197 4681 10226 4687 1 vdd
rlabel locali 9965 2461 9985 2474 1 d3
rlabel nwell 10156 2624 10179 2627 1 vdd
rlabel space 10124 2366 10153 2375 1 gnd
rlabel locali 10018 2348 10047 2354 1 gnd
rlabel locali 10021 2647 10050 2653 1 vdd
rlabel locali 9880 1439 9900 1463 1 d2
rlabel nwell 10073 1608 10096 1611 1 vdd
rlabel space 10041 1350 10070 1359 1 gnd
rlabel locali 9935 1332 9964 1338 1 gnd
rlabel locali 9938 1631 9967 1637 1 vdd
rlabel locali 9779 1029 9801 1046 1 d1
rlabel nwell 9974 1198 9997 1201 1 vdd
rlabel space 9942 940 9971 949 1 gnd
rlabel locali 9836 922 9865 928 1 gnd
rlabel locali 9839 1221 9868 1227 1 vdd
rlabel locali 9796 2047 9818 2064 1 d1
rlabel nwell 9991 2216 10014 2219 1 vdd
rlabel space 9959 1958 9988 1967 1 gnd
rlabel locali 9853 1940 9882 1946 1 gnd
rlabel locali 9856 2239 9885 2245 1 vdd
rlabel nwell 9177 970 9200 973 1 vdd
rlabel space 9145 712 9174 721 1 gnd
rlabel locali 9039 694 9068 700 1 gnd
rlabel locali 9042 993 9071 999 1 vdd
rlabel locali 8988 805 9010 820 1 d0
rlabel nwell 9176 1382 9199 1385 1 vdd
rlabel space 9144 1124 9173 1133 1 gnd
rlabel locali 9038 1106 9067 1112 1 gnd
rlabel locali 9041 1405 9070 1411 1 vdd
rlabel locali 8987 1217 9009 1232 1 d0
rlabel nwell 9194 1988 9217 1991 1 vdd
rlabel space 9162 1730 9191 1739 1 gnd
rlabel locali 9056 1712 9085 1718 1 gnd
rlabel locali 9059 2011 9088 2017 1 vdd
rlabel locali 9005 1823 9027 1838 1 d0
rlabel nwell 9193 2400 9216 2403 1 vdd
rlabel space 9161 2142 9190 2151 1 gnd
rlabel locali 9055 2124 9084 2130 1 gnd
rlabel locali 9058 2423 9087 2429 1 vdd
rlabel locali 9004 2235 9026 2250 1 d0
rlabel locali 9917 3475 9937 3499 1 d2
rlabel nwell 10110 3644 10133 3647 1 vdd
rlabel space 10078 3386 10107 3395 1 gnd
rlabel locali 9972 3368 10001 3374 1 gnd
rlabel locali 9975 3667 10004 3673 1 vdd
rlabel locali 9816 3065 9838 3082 1 d1
rlabel nwell 10011 3234 10034 3237 1 vdd
rlabel space 9979 2976 10008 2985 1 gnd
rlabel locali 9873 2958 9902 2964 1 gnd
rlabel locali 9876 3257 9905 3263 1 vdd
rlabel locali 9833 4083 9855 4100 1 d1
rlabel nwell 10028 4252 10051 4255 1 vdd
rlabel space 9996 3994 10025 4003 1 gnd
rlabel locali 9890 3976 9919 3982 1 gnd
rlabel locali 9893 4275 9922 4281 1 vdd
rlabel nwell 9214 3006 9237 3009 1 vdd
rlabel space 9182 2748 9211 2757 1 gnd
rlabel locali 9076 2730 9105 2736 1 gnd
rlabel locali 9079 3029 9108 3035 1 vdd
rlabel locali 9025 2841 9047 2856 1 d0
rlabel nwell 9213 3418 9236 3421 1 vdd
rlabel space 9181 3160 9210 3169 1 gnd
rlabel locali 9075 3142 9104 3148 1 gnd
rlabel locali 9078 3441 9107 3447 1 vdd
rlabel locali 9024 3253 9046 3268 1 d0
rlabel nwell 9231 4024 9254 4027 1 vdd
rlabel space 9199 3766 9228 3775 1 gnd
rlabel locali 9093 3748 9122 3754 1 gnd
rlabel locali 9096 4047 9125 4053 1 vdd
rlabel locali 9042 3859 9064 3874 1 d0
rlabel nwell 9230 4436 9253 4439 1 vdd
rlabel space 9198 4178 9227 4187 1 gnd
rlabel locali 9092 4160 9121 4166 1 gnd
rlabel locali 9095 4459 9124 4465 1 vdd
rlabel locali 9041 4271 9063 4286 1 d0
rlabel locali 10038 6533 10058 6546 1 d3
rlabel nwell 10229 6696 10252 6699 1 vdd
rlabel space 10197 6438 10226 6447 1 gnd
rlabel locali 10091 6420 10120 6426 1 gnd
rlabel locali 10094 6719 10123 6725 1 vdd
rlabel locali 9953 5511 9973 5535 1 d2
rlabel nwell 10146 5680 10169 5683 1 vdd
rlabel space 10114 5422 10143 5431 1 gnd
rlabel locali 10008 5404 10037 5410 1 gnd
rlabel locali 10011 5703 10040 5709 1 vdd
rlabel locali 9852 5101 9874 5118 1 d1
rlabel nwell 10047 5270 10070 5273 1 vdd
rlabel space 10015 5012 10044 5021 1 gnd
rlabel locali 9909 4994 9938 5000 1 gnd
rlabel locali 9912 5293 9941 5299 1 vdd
rlabel locali 9869 6119 9891 6136 1 d1
rlabel nwell 10064 6288 10087 6291 1 vdd
rlabel space 10032 6030 10061 6039 1 gnd
rlabel locali 9926 6012 9955 6018 1 gnd
rlabel locali 9929 6311 9958 6317 1 vdd
rlabel nwell 9250 5042 9273 5045 1 vdd
rlabel space 9218 4784 9247 4793 1 gnd
rlabel locali 9112 4766 9141 4772 1 gnd
rlabel locali 9115 5065 9144 5071 1 vdd
rlabel locali 9061 4877 9083 4892 1 d0
rlabel nwell 9249 5454 9272 5457 1 vdd
rlabel space 9217 5196 9246 5205 1 gnd
rlabel locali 9111 5178 9140 5184 1 gnd
rlabel locali 9114 5477 9143 5483 1 vdd
rlabel locali 9060 5289 9082 5304 1 d0
rlabel nwell 9267 6060 9290 6063 1 vdd
rlabel space 9235 5802 9264 5811 1 gnd
rlabel locali 9129 5784 9158 5790 1 gnd
rlabel locali 9132 6083 9161 6089 1 vdd
rlabel locali 9078 5895 9100 5910 1 d0
rlabel nwell 9266 6472 9289 6475 1 vdd
rlabel space 9234 6214 9263 6223 1 gnd
rlabel locali 9128 6196 9157 6202 1 gnd
rlabel locali 9131 6495 9160 6501 1 vdd
rlabel locali 9077 6307 9099 6322 1 d0
rlabel locali 9990 7547 10010 7571 1 d2
rlabel nwell 10183 7716 10206 7719 1 vdd
rlabel space 10151 7458 10180 7467 1 gnd
rlabel locali 10045 7440 10074 7446 1 gnd
rlabel locali 10048 7739 10077 7745 1 vdd
rlabel locali 9889 7137 9911 7154 1 d1
rlabel nwell 10084 7306 10107 7309 1 vdd
rlabel space 10052 7048 10081 7057 1 gnd
rlabel locali 9946 7030 9975 7036 1 gnd
rlabel locali 9949 7329 9978 7335 1 vdd
rlabel locali 9906 8155 9928 8172 1 d1
rlabel nwell 10101 8324 10124 8327 1 vdd
rlabel space 10069 8066 10098 8075 1 gnd
rlabel locali 9963 8048 9992 8054 1 gnd
rlabel locali 9966 8347 9995 8353 1 vdd
rlabel nwell 9287 7078 9310 7081 1 vdd
rlabel space 9255 6820 9284 6829 1 gnd
rlabel locali 9149 6802 9178 6808 1 gnd
rlabel locali 9152 7101 9181 7107 1 vdd
rlabel locali 9098 6913 9120 6928 1 d0
rlabel nwell 9286 7490 9309 7493 1 vdd
rlabel space 9254 7232 9283 7241 1 gnd
rlabel locali 9148 7214 9177 7220 1 gnd
rlabel locali 9151 7513 9180 7519 1 vdd
rlabel locali 9097 7325 9119 7340 1 d0
rlabel nwell 9304 8096 9327 8099 1 vdd
rlabel space 9272 7838 9301 7847 1 gnd
rlabel locali 9166 7820 9195 7826 1 gnd
rlabel locali 9169 8119 9198 8125 1 vdd
rlabel locali 9115 7931 9137 7946 1 d0
rlabel nwell 9303 8508 9326 8511 1 vdd
rlabel space 9271 8250 9300 8259 1 gnd
rlabel locali 9165 8232 9194 8238 1 gnd
rlabel locali 9168 8531 9197 8537 1 vdd
rlabel locali 9114 8343 9136 8358 1 d0
rlabel locali 8451 342 8480 348 1 vdd
rlabel locali 8448 43 8477 49 1 gnd
rlabel space 8554 61 8583 70 1 gnd
rlabel nwell 8586 319 8609 322 1 vdd
rlabel locali 8824 189 8846 204 1 vout
rlabel locali 8390 155 8412 170 1 d7
<< end >>

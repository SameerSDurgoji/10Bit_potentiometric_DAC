magic
tech sky130A
timestamp 1616089871
<< nwell >>
rect 328 3648 936 3798
rect 1126 3464 1734 3614
rect 329 3236 937 3386
rect 1208 2856 1816 3006
rect 311 2630 919 2780
rect 1109 2446 1717 2596
rect 312 2218 920 2368
rect 1254 1836 1862 1986
rect 291 1612 899 1762
rect 1089 1428 1697 1578
rect 292 1200 900 1350
rect 1171 820 1779 970
rect 274 594 882 744
rect 1072 410 1680 560
rect 275 182 883 332
rect 1357 -202 1965 -52
rect 255 -424 863 -274
rect 1053 -608 1661 -458
rect 256 -836 864 -686
rect 1135 -1216 1743 -1066
rect 238 -1442 846 -1292
rect 1036 -1626 1644 -1476
rect 239 -1854 847 -1704
rect 1181 -2236 1789 -2086
rect 218 -2460 826 -2310
rect 1016 -2644 1624 -2494
rect 219 -2872 827 -2722
rect 1098 -3252 1706 -3102
rect 201 -3478 809 -3328
rect 999 -3662 1607 -3512
rect 202 -3890 810 -3740
<< nmos >>
rect 392 3547 442 3589
rect 610 3547 660 3589
rect 818 3547 868 3589
rect 1190 3363 1240 3405
rect 1408 3363 1458 3405
rect 1616 3363 1666 3405
rect 393 3135 443 3177
rect 611 3135 661 3177
rect 819 3135 869 3177
rect 1272 2755 1322 2797
rect 1490 2755 1540 2797
rect 1698 2755 1748 2797
rect 375 2529 425 2571
rect 593 2529 643 2571
rect 801 2529 851 2571
rect 1173 2345 1223 2387
rect 1391 2345 1441 2387
rect 1599 2345 1649 2387
rect 376 2117 426 2159
rect 594 2117 644 2159
rect 802 2117 852 2159
rect 1318 1735 1368 1777
rect 1536 1735 1586 1777
rect 1744 1735 1794 1777
rect 355 1511 405 1553
rect 573 1511 623 1553
rect 781 1511 831 1553
rect 1153 1327 1203 1369
rect 1371 1327 1421 1369
rect 1579 1327 1629 1369
rect 356 1099 406 1141
rect 574 1099 624 1141
rect 782 1099 832 1141
rect 1235 719 1285 761
rect 1453 719 1503 761
rect 1661 719 1711 761
rect 338 493 388 535
rect 556 493 606 535
rect 764 493 814 535
rect 1136 309 1186 351
rect 1354 309 1404 351
rect 1562 309 1612 351
rect 339 81 389 123
rect 557 81 607 123
rect 765 81 815 123
rect 1421 -303 1471 -261
rect 1639 -303 1689 -261
rect 1847 -303 1897 -261
rect 319 -525 369 -483
rect 537 -525 587 -483
rect 745 -525 795 -483
rect 1117 -709 1167 -667
rect 1335 -709 1385 -667
rect 1543 -709 1593 -667
rect 320 -937 370 -895
rect 538 -937 588 -895
rect 746 -937 796 -895
rect 1199 -1317 1249 -1275
rect 1417 -1317 1467 -1275
rect 1625 -1317 1675 -1275
rect 302 -1543 352 -1501
rect 520 -1543 570 -1501
rect 728 -1543 778 -1501
rect 1100 -1727 1150 -1685
rect 1318 -1727 1368 -1685
rect 1526 -1727 1576 -1685
rect 303 -1955 353 -1913
rect 521 -1955 571 -1913
rect 729 -1955 779 -1913
rect 1245 -2337 1295 -2295
rect 1463 -2337 1513 -2295
rect 1671 -2337 1721 -2295
rect 282 -2561 332 -2519
rect 500 -2561 550 -2519
rect 708 -2561 758 -2519
rect 1080 -2745 1130 -2703
rect 1298 -2745 1348 -2703
rect 1506 -2745 1556 -2703
rect 283 -2973 333 -2931
rect 501 -2973 551 -2931
rect 709 -2973 759 -2931
rect 1162 -3353 1212 -3311
rect 1380 -3353 1430 -3311
rect 1588 -3353 1638 -3311
rect 265 -3579 315 -3537
rect 483 -3579 533 -3537
rect 691 -3579 741 -3537
rect 1063 -3763 1113 -3721
rect 1281 -3763 1331 -3721
rect 1489 -3763 1539 -3721
rect 266 -3991 316 -3949
rect 484 -3991 534 -3949
rect 692 -3991 742 -3949
<< pmos >>
rect 392 3666 442 3766
rect 610 3666 660 3766
rect 818 3666 868 3766
rect 1190 3482 1240 3582
rect 1408 3482 1458 3582
rect 1616 3482 1666 3582
rect 393 3254 443 3354
rect 611 3254 661 3354
rect 819 3254 869 3354
rect 1272 2874 1322 2974
rect 1490 2874 1540 2974
rect 1698 2874 1748 2974
rect 375 2648 425 2748
rect 593 2648 643 2748
rect 801 2648 851 2748
rect 1173 2464 1223 2564
rect 1391 2464 1441 2564
rect 1599 2464 1649 2564
rect 376 2236 426 2336
rect 594 2236 644 2336
rect 802 2236 852 2336
rect 1318 1854 1368 1954
rect 1536 1854 1586 1954
rect 1744 1854 1794 1954
rect 355 1630 405 1730
rect 573 1630 623 1730
rect 781 1630 831 1730
rect 1153 1446 1203 1546
rect 1371 1446 1421 1546
rect 1579 1446 1629 1546
rect 356 1218 406 1318
rect 574 1218 624 1318
rect 782 1218 832 1318
rect 1235 838 1285 938
rect 1453 838 1503 938
rect 1661 838 1711 938
rect 338 612 388 712
rect 556 612 606 712
rect 764 612 814 712
rect 1136 428 1186 528
rect 1354 428 1404 528
rect 1562 428 1612 528
rect 339 200 389 300
rect 557 200 607 300
rect 765 200 815 300
rect 1421 -184 1471 -84
rect 1639 -184 1689 -84
rect 1847 -184 1897 -84
rect 319 -406 369 -306
rect 537 -406 587 -306
rect 745 -406 795 -306
rect 1117 -590 1167 -490
rect 1335 -590 1385 -490
rect 1543 -590 1593 -490
rect 320 -818 370 -718
rect 538 -818 588 -718
rect 746 -818 796 -718
rect 1199 -1198 1249 -1098
rect 1417 -1198 1467 -1098
rect 1625 -1198 1675 -1098
rect 302 -1424 352 -1324
rect 520 -1424 570 -1324
rect 728 -1424 778 -1324
rect 1100 -1608 1150 -1508
rect 1318 -1608 1368 -1508
rect 1526 -1608 1576 -1508
rect 303 -1836 353 -1736
rect 521 -1836 571 -1736
rect 729 -1836 779 -1736
rect 1245 -2218 1295 -2118
rect 1463 -2218 1513 -2118
rect 1671 -2218 1721 -2118
rect 282 -2442 332 -2342
rect 500 -2442 550 -2342
rect 708 -2442 758 -2342
rect 1080 -2626 1130 -2526
rect 1298 -2626 1348 -2526
rect 1506 -2626 1556 -2526
rect 283 -2854 333 -2754
rect 501 -2854 551 -2754
rect 709 -2854 759 -2754
rect 1162 -3234 1212 -3134
rect 1380 -3234 1430 -3134
rect 1588 -3234 1638 -3134
rect 265 -3460 315 -3360
rect 483 -3460 533 -3360
rect 691 -3460 741 -3360
rect 1063 -3644 1113 -3544
rect 1281 -3644 1331 -3544
rect 1489 -3644 1539 -3544
rect 266 -3872 316 -3772
rect 484 -3872 534 -3772
rect 692 -3872 742 -3772
<< ndiff >>
rect 343 3579 392 3589
rect 343 3559 354 3579
rect 374 3559 392 3579
rect 343 3547 392 3559
rect 442 3583 486 3589
rect 442 3563 457 3583
rect 477 3563 486 3583
rect 442 3547 486 3563
rect 561 3579 610 3589
rect 561 3559 572 3579
rect 592 3559 610 3579
rect 561 3547 610 3559
rect 660 3583 704 3589
rect 660 3563 675 3583
rect 695 3563 704 3583
rect 660 3547 704 3563
rect 774 3583 818 3589
rect 774 3563 783 3583
rect 803 3563 818 3583
rect 774 3547 818 3563
rect 868 3579 917 3589
rect 868 3559 886 3579
rect 906 3559 917 3579
rect 868 3547 917 3559
rect 1141 3395 1190 3405
rect 1141 3375 1152 3395
rect 1172 3375 1190 3395
rect 1141 3363 1190 3375
rect 1240 3399 1284 3405
rect 1240 3379 1255 3399
rect 1275 3379 1284 3399
rect 1240 3363 1284 3379
rect 1359 3395 1408 3405
rect 1359 3375 1370 3395
rect 1390 3375 1408 3395
rect 1359 3363 1408 3375
rect 1458 3399 1502 3405
rect 1458 3379 1473 3399
rect 1493 3379 1502 3399
rect 1458 3363 1502 3379
rect 1572 3399 1616 3405
rect 1572 3379 1581 3399
rect 1601 3379 1616 3399
rect 1572 3363 1616 3379
rect 1666 3395 1715 3405
rect 1666 3375 1684 3395
rect 1704 3375 1715 3395
rect 1666 3363 1715 3375
rect 344 3167 393 3177
rect 344 3147 355 3167
rect 375 3147 393 3167
rect 344 3135 393 3147
rect 443 3171 487 3177
rect 443 3151 458 3171
rect 478 3151 487 3171
rect 443 3135 487 3151
rect 562 3167 611 3177
rect 562 3147 573 3167
rect 593 3147 611 3167
rect 562 3135 611 3147
rect 661 3171 705 3177
rect 661 3151 676 3171
rect 696 3151 705 3171
rect 661 3135 705 3151
rect 775 3171 819 3177
rect 775 3151 784 3171
rect 804 3151 819 3171
rect 775 3135 819 3151
rect 869 3167 918 3177
rect 869 3147 887 3167
rect 907 3147 918 3167
rect 869 3135 918 3147
rect 1223 2787 1272 2797
rect 1223 2767 1234 2787
rect 1254 2767 1272 2787
rect 1223 2755 1272 2767
rect 1322 2791 1366 2797
rect 1322 2771 1337 2791
rect 1357 2771 1366 2791
rect 1322 2755 1366 2771
rect 1441 2787 1490 2797
rect 1441 2767 1452 2787
rect 1472 2767 1490 2787
rect 1441 2755 1490 2767
rect 1540 2791 1584 2797
rect 1540 2771 1555 2791
rect 1575 2771 1584 2791
rect 1540 2755 1584 2771
rect 1654 2791 1698 2797
rect 1654 2771 1663 2791
rect 1683 2771 1698 2791
rect 1654 2755 1698 2771
rect 1748 2787 1797 2797
rect 1748 2767 1766 2787
rect 1786 2767 1797 2787
rect 1748 2755 1797 2767
rect 326 2561 375 2571
rect 326 2541 337 2561
rect 357 2541 375 2561
rect 326 2529 375 2541
rect 425 2565 469 2571
rect 425 2545 440 2565
rect 460 2545 469 2565
rect 425 2529 469 2545
rect 544 2561 593 2571
rect 544 2541 555 2561
rect 575 2541 593 2561
rect 544 2529 593 2541
rect 643 2565 687 2571
rect 643 2545 658 2565
rect 678 2545 687 2565
rect 643 2529 687 2545
rect 757 2565 801 2571
rect 757 2545 766 2565
rect 786 2545 801 2565
rect 757 2529 801 2545
rect 851 2561 900 2571
rect 851 2541 869 2561
rect 889 2541 900 2561
rect 851 2529 900 2541
rect 1124 2377 1173 2387
rect 1124 2357 1135 2377
rect 1155 2357 1173 2377
rect 1124 2345 1173 2357
rect 1223 2381 1267 2387
rect 1223 2361 1238 2381
rect 1258 2361 1267 2381
rect 1223 2345 1267 2361
rect 1342 2377 1391 2387
rect 1342 2357 1353 2377
rect 1373 2357 1391 2377
rect 1342 2345 1391 2357
rect 1441 2381 1485 2387
rect 1441 2361 1456 2381
rect 1476 2361 1485 2381
rect 1441 2345 1485 2361
rect 1555 2381 1599 2387
rect 1555 2361 1564 2381
rect 1584 2361 1599 2381
rect 1555 2345 1599 2361
rect 1649 2377 1698 2387
rect 1649 2357 1667 2377
rect 1687 2357 1698 2377
rect 1649 2345 1698 2357
rect 327 2149 376 2159
rect 327 2129 338 2149
rect 358 2129 376 2149
rect 327 2117 376 2129
rect 426 2153 470 2159
rect 426 2133 441 2153
rect 461 2133 470 2153
rect 426 2117 470 2133
rect 545 2149 594 2159
rect 545 2129 556 2149
rect 576 2129 594 2149
rect 545 2117 594 2129
rect 644 2153 688 2159
rect 644 2133 659 2153
rect 679 2133 688 2153
rect 644 2117 688 2133
rect 758 2153 802 2159
rect 758 2133 767 2153
rect 787 2133 802 2153
rect 758 2117 802 2133
rect 852 2149 901 2159
rect 852 2129 870 2149
rect 890 2129 901 2149
rect 852 2117 901 2129
rect 1269 1767 1318 1777
rect 1269 1747 1280 1767
rect 1300 1747 1318 1767
rect 1269 1735 1318 1747
rect 1368 1771 1412 1777
rect 1368 1751 1383 1771
rect 1403 1751 1412 1771
rect 1368 1735 1412 1751
rect 1487 1767 1536 1777
rect 1487 1747 1498 1767
rect 1518 1747 1536 1767
rect 1487 1735 1536 1747
rect 1586 1771 1630 1777
rect 1586 1751 1601 1771
rect 1621 1751 1630 1771
rect 1586 1735 1630 1751
rect 1700 1771 1744 1777
rect 1700 1751 1709 1771
rect 1729 1751 1744 1771
rect 1700 1735 1744 1751
rect 1794 1767 1843 1777
rect 1794 1747 1812 1767
rect 1832 1747 1843 1767
rect 1794 1735 1843 1747
rect 306 1543 355 1553
rect 306 1523 317 1543
rect 337 1523 355 1543
rect 306 1511 355 1523
rect 405 1547 449 1553
rect 405 1527 420 1547
rect 440 1527 449 1547
rect 405 1511 449 1527
rect 524 1543 573 1553
rect 524 1523 535 1543
rect 555 1523 573 1543
rect 524 1511 573 1523
rect 623 1547 667 1553
rect 623 1527 638 1547
rect 658 1527 667 1547
rect 623 1511 667 1527
rect 737 1547 781 1553
rect 737 1527 746 1547
rect 766 1527 781 1547
rect 737 1511 781 1527
rect 831 1543 880 1553
rect 831 1523 849 1543
rect 869 1523 880 1543
rect 831 1511 880 1523
rect 1104 1359 1153 1369
rect 1104 1339 1115 1359
rect 1135 1339 1153 1359
rect 1104 1327 1153 1339
rect 1203 1363 1247 1369
rect 1203 1343 1218 1363
rect 1238 1343 1247 1363
rect 1203 1327 1247 1343
rect 1322 1359 1371 1369
rect 1322 1339 1333 1359
rect 1353 1339 1371 1359
rect 1322 1327 1371 1339
rect 1421 1363 1465 1369
rect 1421 1343 1436 1363
rect 1456 1343 1465 1363
rect 1421 1327 1465 1343
rect 1535 1363 1579 1369
rect 1535 1343 1544 1363
rect 1564 1343 1579 1363
rect 1535 1327 1579 1343
rect 1629 1359 1678 1369
rect 1629 1339 1647 1359
rect 1667 1339 1678 1359
rect 1629 1327 1678 1339
rect 307 1131 356 1141
rect 307 1111 318 1131
rect 338 1111 356 1131
rect 307 1099 356 1111
rect 406 1135 450 1141
rect 406 1115 421 1135
rect 441 1115 450 1135
rect 406 1099 450 1115
rect 525 1131 574 1141
rect 525 1111 536 1131
rect 556 1111 574 1131
rect 525 1099 574 1111
rect 624 1135 668 1141
rect 624 1115 639 1135
rect 659 1115 668 1135
rect 624 1099 668 1115
rect 738 1135 782 1141
rect 738 1115 747 1135
rect 767 1115 782 1135
rect 738 1099 782 1115
rect 832 1131 881 1141
rect 832 1111 850 1131
rect 870 1111 881 1131
rect 832 1099 881 1111
rect 1186 751 1235 761
rect 1186 731 1197 751
rect 1217 731 1235 751
rect 1186 719 1235 731
rect 1285 755 1329 761
rect 1285 735 1300 755
rect 1320 735 1329 755
rect 1285 719 1329 735
rect 1404 751 1453 761
rect 1404 731 1415 751
rect 1435 731 1453 751
rect 1404 719 1453 731
rect 1503 755 1547 761
rect 1503 735 1518 755
rect 1538 735 1547 755
rect 1503 719 1547 735
rect 1617 755 1661 761
rect 1617 735 1626 755
rect 1646 735 1661 755
rect 1617 719 1661 735
rect 1711 751 1760 761
rect 1711 731 1729 751
rect 1749 731 1760 751
rect 1711 719 1760 731
rect 289 525 338 535
rect 289 505 300 525
rect 320 505 338 525
rect 289 493 338 505
rect 388 529 432 535
rect 388 509 403 529
rect 423 509 432 529
rect 388 493 432 509
rect 507 525 556 535
rect 507 505 518 525
rect 538 505 556 525
rect 507 493 556 505
rect 606 529 650 535
rect 606 509 621 529
rect 641 509 650 529
rect 606 493 650 509
rect 720 529 764 535
rect 720 509 729 529
rect 749 509 764 529
rect 720 493 764 509
rect 814 525 863 535
rect 814 505 832 525
rect 852 505 863 525
rect 814 493 863 505
rect 1087 341 1136 351
rect 1087 321 1098 341
rect 1118 321 1136 341
rect 1087 309 1136 321
rect 1186 345 1230 351
rect 1186 325 1201 345
rect 1221 325 1230 345
rect 1186 309 1230 325
rect 1305 341 1354 351
rect 1305 321 1316 341
rect 1336 321 1354 341
rect 1305 309 1354 321
rect 1404 345 1448 351
rect 1404 325 1419 345
rect 1439 325 1448 345
rect 1404 309 1448 325
rect 1518 345 1562 351
rect 1518 325 1527 345
rect 1547 325 1562 345
rect 1518 309 1562 325
rect 1612 341 1661 351
rect 1612 321 1630 341
rect 1650 321 1661 341
rect 1612 309 1661 321
rect 290 113 339 123
rect 290 93 301 113
rect 321 93 339 113
rect 290 81 339 93
rect 389 117 433 123
rect 389 97 404 117
rect 424 97 433 117
rect 389 81 433 97
rect 508 113 557 123
rect 508 93 519 113
rect 539 93 557 113
rect 508 81 557 93
rect 607 117 651 123
rect 607 97 622 117
rect 642 97 651 117
rect 607 81 651 97
rect 721 117 765 123
rect 721 97 730 117
rect 750 97 765 117
rect 721 81 765 97
rect 815 113 864 123
rect 815 93 833 113
rect 853 93 864 113
rect 815 81 864 93
rect 1372 -271 1421 -261
rect 1372 -291 1383 -271
rect 1403 -291 1421 -271
rect 1372 -303 1421 -291
rect 1471 -267 1515 -261
rect 1471 -287 1486 -267
rect 1506 -287 1515 -267
rect 1471 -303 1515 -287
rect 1590 -271 1639 -261
rect 1590 -291 1601 -271
rect 1621 -291 1639 -271
rect 1590 -303 1639 -291
rect 1689 -267 1733 -261
rect 1689 -287 1704 -267
rect 1724 -287 1733 -267
rect 1689 -303 1733 -287
rect 1803 -267 1847 -261
rect 1803 -287 1812 -267
rect 1832 -287 1847 -267
rect 1803 -303 1847 -287
rect 1897 -271 1946 -261
rect 1897 -291 1915 -271
rect 1935 -291 1946 -271
rect 1897 -303 1946 -291
rect 270 -493 319 -483
rect 270 -513 281 -493
rect 301 -513 319 -493
rect 270 -525 319 -513
rect 369 -489 413 -483
rect 369 -509 384 -489
rect 404 -509 413 -489
rect 369 -525 413 -509
rect 488 -493 537 -483
rect 488 -513 499 -493
rect 519 -513 537 -493
rect 488 -525 537 -513
rect 587 -489 631 -483
rect 587 -509 602 -489
rect 622 -509 631 -489
rect 587 -525 631 -509
rect 701 -489 745 -483
rect 701 -509 710 -489
rect 730 -509 745 -489
rect 701 -525 745 -509
rect 795 -493 844 -483
rect 795 -513 813 -493
rect 833 -513 844 -493
rect 795 -525 844 -513
rect 1068 -677 1117 -667
rect 1068 -697 1079 -677
rect 1099 -697 1117 -677
rect 1068 -709 1117 -697
rect 1167 -673 1211 -667
rect 1167 -693 1182 -673
rect 1202 -693 1211 -673
rect 1167 -709 1211 -693
rect 1286 -677 1335 -667
rect 1286 -697 1297 -677
rect 1317 -697 1335 -677
rect 1286 -709 1335 -697
rect 1385 -673 1429 -667
rect 1385 -693 1400 -673
rect 1420 -693 1429 -673
rect 1385 -709 1429 -693
rect 1499 -673 1543 -667
rect 1499 -693 1508 -673
rect 1528 -693 1543 -673
rect 1499 -709 1543 -693
rect 1593 -677 1642 -667
rect 1593 -697 1611 -677
rect 1631 -697 1642 -677
rect 1593 -709 1642 -697
rect 271 -905 320 -895
rect 271 -925 282 -905
rect 302 -925 320 -905
rect 271 -937 320 -925
rect 370 -901 414 -895
rect 370 -921 385 -901
rect 405 -921 414 -901
rect 370 -937 414 -921
rect 489 -905 538 -895
rect 489 -925 500 -905
rect 520 -925 538 -905
rect 489 -937 538 -925
rect 588 -901 632 -895
rect 588 -921 603 -901
rect 623 -921 632 -901
rect 588 -937 632 -921
rect 702 -901 746 -895
rect 702 -921 711 -901
rect 731 -921 746 -901
rect 702 -937 746 -921
rect 796 -905 845 -895
rect 796 -925 814 -905
rect 834 -925 845 -905
rect 796 -937 845 -925
rect 1150 -1285 1199 -1275
rect 1150 -1305 1161 -1285
rect 1181 -1305 1199 -1285
rect 1150 -1317 1199 -1305
rect 1249 -1281 1293 -1275
rect 1249 -1301 1264 -1281
rect 1284 -1301 1293 -1281
rect 1249 -1317 1293 -1301
rect 1368 -1285 1417 -1275
rect 1368 -1305 1379 -1285
rect 1399 -1305 1417 -1285
rect 1368 -1317 1417 -1305
rect 1467 -1281 1511 -1275
rect 1467 -1301 1482 -1281
rect 1502 -1301 1511 -1281
rect 1467 -1317 1511 -1301
rect 1581 -1281 1625 -1275
rect 1581 -1301 1590 -1281
rect 1610 -1301 1625 -1281
rect 1581 -1317 1625 -1301
rect 1675 -1285 1724 -1275
rect 1675 -1305 1693 -1285
rect 1713 -1305 1724 -1285
rect 1675 -1317 1724 -1305
rect 253 -1511 302 -1501
rect 253 -1531 264 -1511
rect 284 -1531 302 -1511
rect 253 -1543 302 -1531
rect 352 -1507 396 -1501
rect 352 -1527 367 -1507
rect 387 -1527 396 -1507
rect 352 -1543 396 -1527
rect 471 -1511 520 -1501
rect 471 -1531 482 -1511
rect 502 -1531 520 -1511
rect 471 -1543 520 -1531
rect 570 -1507 614 -1501
rect 570 -1527 585 -1507
rect 605 -1527 614 -1507
rect 570 -1543 614 -1527
rect 684 -1507 728 -1501
rect 684 -1527 693 -1507
rect 713 -1527 728 -1507
rect 684 -1543 728 -1527
rect 778 -1511 827 -1501
rect 778 -1531 796 -1511
rect 816 -1531 827 -1511
rect 778 -1543 827 -1531
rect 1051 -1695 1100 -1685
rect 1051 -1715 1062 -1695
rect 1082 -1715 1100 -1695
rect 1051 -1727 1100 -1715
rect 1150 -1691 1194 -1685
rect 1150 -1711 1165 -1691
rect 1185 -1711 1194 -1691
rect 1150 -1727 1194 -1711
rect 1269 -1695 1318 -1685
rect 1269 -1715 1280 -1695
rect 1300 -1715 1318 -1695
rect 1269 -1727 1318 -1715
rect 1368 -1691 1412 -1685
rect 1368 -1711 1383 -1691
rect 1403 -1711 1412 -1691
rect 1368 -1727 1412 -1711
rect 1482 -1691 1526 -1685
rect 1482 -1711 1491 -1691
rect 1511 -1711 1526 -1691
rect 1482 -1727 1526 -1711
rect 1576 -1695 1625 -1685
rect 1576 -1715 1594 -1695
rect 1614 -1715 1625 -1695
rect 1576 -1727 1625 -1715
rect 254 -1923 303 -1913
rect 254 -1943 265 -1923
rect 285 -1943 303 -1923
rect 254 -1955 303 -1943
rect 353 -1919 397 -1913
rect 353 -1939 368 -1919
rect 388 -1939 397 -1919
rect 353 -1955 397 -1939
rect 472 -1923 521 -1913
rect 472 -1943 483 -1923
rect 503 -1943 521 -1923
rect 472 -1955 521 -1943
rect 571 -1919 615 -1913
rect 571 -1939 586 -1919
rect 606 -1939 615 -1919
rect 571 -1955 615 -1939
rect 685 -1919 729 -1913
rect 685 -1939 694 -1919
rect 714 -1939 729 -1919
rect 685 -1955 729 -1939
rect 779 -1923 828 -1913
rect 779 -1943 797 -1923
rect 817 -1943 828 -1923
rect 779 -1955 828 -1943
rect 1196 -2305 1245 -2295
rect 1196 -2325 1207 -2305
rect 1227 -2325 1245 -2305
rect 1196 -2337 1245 -2325
rect 1295 -2301 1339 -2295
rect 1295 -2321 1310 -2301
rect 1330 -2321 1339 -2301
rect 1295 -2337 1339 -2321
rect 1414 -2305 1463 -2295
rect 1414 -2325 1425 -2305
rect 1445 -2325 1463 -2305
rect 1414 -2337 1463 -2325
rect 1513 -2301 1557 -2295
rect 1513 -2321 1528 -2301
rect 1548 -2321 1557 -2301
rect 1513 -2337 1557 -2321
rect 1627 -2301 1671 -2295
rect 1627 -2321 1636 -2301
rect 1656 -2321 1671 -2301
rect 1627 -2337 1671 -2321
rect 1721 -2305 1770 -2295
rect 1721 -2325 1739 -2305
rect 1759 -2325 1770 -2305
rect 1721 -2337 1770 -2325
rect 233 -2529 282 -2519
rect 233 -2549 244 -2529
rect 264 -2549 282 -2529
rect 233 -2561 282 -2549
rect 332 -2525 376 -2519
rect 332 -2545 347 -2525
rect 367 -2545 376 -2525
rect 332 -2561 376 -2545
rect 451 -2529 500 -2519
rect 451 -2549 462 -2529
rect 482 -2549 500 -2529
rect 451 -2561 500 -2549
rect 550 -2525 594 -2519
rect 550 -2545 565 -2525
rect 585 -2545 594 -2525
rect 550 -2561 594 -2545
rect 664 -2525 708 -2519
rect 664 -2545 673 -2525
rect 693 -2545 708 -2525
rect 664 -2561 708 -2545
rect 758 -2529 807 -2519
rect 758 -2549 776 -2529
rect 796 -2549 807 -2529
rect 758 -2561 807 -2549
rect 1031 -2713 1080 -2703
rect 1031 -2733 1042 -2713
rect 1062 -2733 1080 -2713
rect 1031 -2745 1080 -2733
rect 1130 -2709 1174 -2703
rect 1130 -2729 1145 -2709
rect 1165 -2729 1174 -2709
rect 1130 -2745 1174 -2729
rect 1249 -2713 1298 -2703
rect 1249 -2733 1260 -2713
rect 1280 -2733 1298 -2713
rect 1249 -2745 1298 -2733
rect 1348 -2709 1392 -2703
rect 1348 -2729 1363 -2709
rect 1383 -2729 1392 -2709
rect 1348 -2745 1392 -2729
rect 1462 -2709 1506 -2703
rect 1462 -2729 1471 -2709
rect 1491 -2729 1506 -2709
rect 1462 -2745 1506 -2729
rect 1556 -2713 1605 -2703
rect 1556 -2733 1574 -2713
rect 1594 -2733 1605 -2713
rect 1556 -2745 1605 -2733
rect 234 -2941 283 -2931
rect 234 -2961 245 -2941
rect 265 -2961 283 -2941
rect 234 -2973 283 -2961
rect 333 -2937 377 -2931
rect 333 -2957 348 -2937
rect 368 -2957 377 -2937
rect 333 -2973 377 -2957
rect 452 -2941 501 -2931
rect 452 -2961 463 -2941
rect 483 -2961 501 -2941
rect 452 -2973 501 -2961
rect 551 -2937 595 -2931
rect 551 -2957 566 -2937
rect 586 -2957 595 -2937
rect 551 -2973 595 -2957
rect 665 -2937 709 -2931
rect 665 -2957 674 -2937
rect 694 -2957 709 -2937
rect 665 -2973 709 -2957
rect 759 -2941 808 -2931
rect 759 -2961 777 -2941
rect 797 -2961 808 -2941
rect 759 -2973 808 -2961
rect 1113 -3321 1162 -3311
rect 1113 -3341 1124 -3321
rect 1144 -3341 1162 -3321
rect 1113 -3353 1162 -3341
rect 1212 -3317 1256 -3311
rect 1212 -3337 1227 -3317
rect 1247 -3337 1256 -3317
rect 1212 -3353 1256 -3337
rect 1331 -3321 1380 -3311
rect 1331 -3341 1342 -3321
rect 1362 -3341 1380 -3321
rect 1331 -3353 1380 -3341
rect 1430 -3317 1474 -3311
rect 1430 -3337 1445 -3317
rect 1465 -3337 1474 -3317
rect 1430 -3353 1474 -3337
rect 1544 -3317 1588 -3311
rect 1544 -3337 1553 -3317
rect 1573 -3337 1588 -3317
rect 1544 -3353 1588 -3337
rect 1638 -3321 1687 -3311
rect 1638 -3341 1656 -3321
rect 1676 -3341 1687 -3321
rect 1638 -3353 1687 -3341
rect 216 -3547 265 -3537
rect 216 -3567 227 -3547
rect 247 -3567 265 -3547
rect 216 -3579 265 -3567
rect 315 -3543 359 -3537
rect 315 -3563 330 -3543
rect 350 -3563 359 -3543
rect 315 -3579 359 -3563
rect 434 -3547 483 -3537
rect 434 -3567 445 -3547
rect 465 -3567 483 -3547
rect 434 -3579 483 -3567
rect 533 -3543 577 -3537
rect 533 -3563 548 -3543
rect 568 -3563 577 -3543
rect 533 -3579 577 -3563
rect 647 -3543 691 -3537
rect 647 -3563 656 -3543
rect 676 -3563 691 -3543
rect 647 -3579 691 -3563
rect 741 -3547 790 -3537
rect 741 -3567 759 -3547
rect 779 -3567 790 -3547
rect 741 -3579 790 -3567
rect 1014 -3731 1063 -3721
rect 1014 -3751 1025 -3731
rect 1045 -3751 1063 -3731
rect 1014 -3763 1063 -3751
rect 1113 -3727 1157 -3721
rect 1113 -3747 1128 -3727
rect 1148 -3747 1157 -3727
rect 1113 -3763 1157 -3747
rect 1232 -3731 1281 -3721
rect 1232 -3751 1243 -3731
rect 1263 -3751 1281 -3731
rect 1232 -3763 1281 -3751
rect 1331 -3727 1375 -3721
rect 1331 -3747 1346 -3727
rect 1366 -3747 1375 -3727
rect 1331 -3763 1375 -3747
rect 1445 -3727 1489 -3721
rect 1445 -3747 1454 -3727
rect 1474 -3747 1489 -3727
rect 1445 -3763 1489 -3747
rect 1539 -3731 1588 -3721
rect 1539 -3751 1557 -3731
rect 1577 -3751 1588 -3731
rect 1539 -3763 1588 -3751
rect 217 -3959 266 -3949
rect 217 -3979 228 -3959
rect 248 -3979 266 -3959
rect 217 -3991 266 -3979
rect 316 -3955 360 -3949
rect 316 -3975 331 -3955
rect 351 -3975 360 -3955
rect 316 -3991 360 -3975
rect 435 -3959 484 -3949
rect 435 -3979 446 -3959
rect 466 -3979 484 -3959
rect 435 -3991 484 -3979
rect 534 -3955 578 -3949
rect 534 -3975 549 -3955
rect 569 -3975 578 -3955
rect 534 -3991 578 -3975
rect 648 -3955 692 -3949
rect 648 -3975 657 -3955
rect 677 -3975 692 -3955
rect 648 -3991 692 -3975
rect 742 -3959 791 -3949
rect 742 -3979 760 -3959
rect 780 -3979 791 -3959
rect 742 -3991 791 -3979
<< pdiff >>
rect 348 3728 392 3766
rect 348 3708 360 3728
rect 380 3708 392 3728
rect 348 3666 392 3708
rect 442 3728 484 3766
rect 442 3708 456 3728
rect 476 3708 484 3728
rect 442 3666 484 3708
rect 566 3728 610 3766
rect 566 3708 578 3728
rect 598 3708 610 3728
rect 566 3666 610 3708
rect 660 3728 702 3766
rect 660 3708 674 3728
rect 694 3708 702 3728
rect 660 3666 702 3708
rect 776 3728 818 3766
rect 776 3708 784 3728
rect 804 3708 818 3728
rect 776 3666 818 3708
rect 868 3735 913 3766
rect 868 3728 912 3735
rect 868 3708 880 3728
rect 900 3708 912 3728
rect 868 3666 912 3708
rect 1146 3544 1190 3582
rect 1146 3524 1158 3544
rect 1178 3524 1190 3544
rect 1146 3482 1190 3524
rect 1240 3544 1282 3582
rect 1240 3524 1254 3544
rect 1274 3524 1282 3544
rect 1240 3482 1282 3524
rect 1364 3544 1408 3582
rect 1364 3524 1376 3544
rect 1396 3524 1408 3544
rect 1364 3482 1408 3524
rect 1458 3544 1500 3582
rect 1458 3524 1472 3544
rect 1492 3524 1500 3544
rect 1458 3482 1500 3524
rect 1574 3544 1616 3582
rect 1574 3524 1582 3544
rect 1602 3524 1616 3544
rect 1574 3482 1616 3524
rect 1666 3551 1711 3582
rect 1666 3544 1710 3551
rect 1666 3524 1678 3544
rect 1698 3524 1710 3544
rect 1666 3482 1710 3524
rect 349 3316 393 3354
rect 349 3296 361 3316
rect 381 3296 393 3316
rect 349 3254 393 3296
rect 443 3316 485 3354
rect 443 3296 457 3316
rect 477 3296 485 3316
rect 443 3254 485 3296
rect 567 3316 611 3354
rect 567 3296 579 3316
rect 599 3296 611 3316
rect 567 3254 611 3296
rect 661 3316 703 3354
rect 661 3296 675 3316
rect 695 3296 703 3316
rect 661 3254 703 3296
rect 777 3316 819 3354
rect 777 3296 785 3316
rect 805 3296 819 3316
rect 777 3254 819 3296
rect 869 3323 914 3354
rect 869 3316 913 3323
rect 869 3296 881 3316
rect 901 3296 913 3316
rect 869 3254 913 3296
rect 1228 2936 1272 2974
rect 1228 2916 1240 2936
rect 1260 2916 1272 2936
rect 1228 2874 1272 2916
rect 1322 2936 1364 2974
rect 1322 2916 1336 2936
rect 1356 2916 1364 2936
rect 1322 2874 1364 2916
rect 1446 2936 1490 2974
rect 1446 2916 1458 2936
rect 1478 2916 1490 2936
rect 1446 2874 1490 2916
rect 1540 2936 1582 2974
rect 1540 2916 1554 2936
rect 1574 2916 1582 2936
rect 1540 2874 1582 2916
rect 1656 2936 1698 2974
rect 1656 2916 1664 2936
rect 1684 2916 1698 2936
rect 1656 2874 1698 2916
rect 1748 2943 1793 2974
rect 1748 2936 1792 2943
rect 1748 2916 1760 2936
rect 1780 2916 1792 2936
rect 1748 2874 1792 2916
rect 331 2710 375 2748
rect 331 2690 343 2710
rect 363 2690 375 2710
rect 331 2648 375 2690
rect 425 2710 467 2748
rect 425 2690 439 2710
rect 459 2690 467 2710
rect 425 2648 467 2690
rect 549 2710 593 2748
rect 549 2690 561 2710
rect 581 2690 593 2710
rect 549 2648 593 2690
rect 643 2710 685 2748
rect 643 2690 657 2710
rect 677 2690 685 2710
rect 643 2648 685 2690
rect 759 2710 801 2748
rect 759 2690 767 2710
rect 787 2690 801 2710
rect 759 2648 801 2690
rect 851 2717 896 2748
rect 851 2710 895 2717
rect 851 2690 863 2710
rect 883 2690 895 2710
rect 851 2648 895 2690
rect 1129 2526 1173 2564
rect 1129 2506 1141 2526
rect 1161 2506 1173 2526
rect 1129 2464 1173 2506
rect 1223 2526 1265 2564
rect 1223 2506 1237 2526
rect 1257 2506 1265 2526
rect 1223 2464 1265 2506
rect 1347 2526 1391 2564
rect 1347 2506 1359 2526
rect 1379 2506 1391 2526
rect 1347 2464 1391 2506
rect 1441 2526 1483 2564
rect 1441 2506 1455 2526
rect 1475 2506 1483 2526
rect 1441 2464 1483 2506
rect 1557 2526 1599 2564
rect 1557 2506 1565 2526
rect 1585 2506 1599 2526
rect 1557 2464 1599 2506
rect 1649 2533 1694 2564
rect 1649 2526 1693 2533
rect 1649 2506 1661 2526
rect 1681 2506 1693 2526
rect 1649 2464 1693 2506
rect 332 2298 376 2336
rect 332 2278 344 2298
rect 364 2278 376 2298
rect 332 2236 376 2278
rect 426 2298 468 2336
rect 426 2278 440 2298
rect 460 2278 468 2298
rect 426 2236 468 2278
rect 550 2298 594 2336
rect 550 2278 562 2298
rect 582 2278 594 2298
rect 550 2236 594 2278
rect 644 2298 686 2336
rect 644 2278 658 2298
rect 678 2278 686 2298
rect 644 2236 686 2278
rect 760 2298 802 2336
rect 760 2278 768 2298
rect 788 2278 802 2298
rect 760 2236 802 2278
rect 852 2305 897 2336
rect 852 2298 896 2305
rect 852 2278 864 2298
rect 884 2278 896 2298
rect 852 2236 896 2278
rect 1274 1916 1318 1954
rect 1274 1896 1286 1916
rect 1306 1896 1318 1916
rect 1274 1854 1318 1896
rect 1368 1916 1410 1954
rect 1368 1896 1382 1916
rect 1402 1896 1410 1916
rect 1368 1854 1410 1896
rect 1492 1916 1536 1954
rect 1492 1896 1504 1916
rect 1524 1896 1536 1916
rect 1492 1854 1536 1896
rect 1586 1916 1628 1954
rect 1586 1896 1600 1916
rect 1620 1896 1628 1916
rect 1586 1854 1628 1896
rect 1702 1916 1744 1954
rect 1702 1896 1710 1916
rect 1730 1896 1744 1916
rect 1702 1854 1744 1896
rect 1794 1923 1839 1954
rect 1794 1916 1838 1923
rect 1794 1896 1806 1916
rect 1826 1896 1838 1916
rect 1794 1854 1838 1896
rect 311 1692 355 1730
rect 311 1672 323 1692
rect 343 1672 355 1692
rect 311 1630 355 1672
rect 405 1692 447 1730
rect 405 1672 419 1692
rect 439 1672 447 1692
rect 405 1630 447 1672
rect 529 1692 573 1730
rect 529 1672 541 1692
rect 561 1672 573 1692
rect 529 1630 573 1672
rect 623 1692 665 1730
rect 623 1672 637 1692
rect 657 1672 665 1692
rect 623 1630 665 1672
rect 739 1692 781 1730
rect 739 1672 747 1692
rect 767 1672 781 1692
rect 739 1630 781 1672
rect 831 1699 876 1730
rect 831 1692 875 1699
rect 831 1672 843 1692
rect 863 1672 875 1692
rect 831 1630 875 1672
rect 1109 1508 1153 1546
rect 1109 1488 1121 1508
rect 1141 1488 1153 1508
rect 1109 1446 1153 1488
rect 1203 1508 1245 1546
rect 1203 1488 1217 1508
rect 1237 1488 1245 1508
rect 1203 1446 1245 1488
rect 1327 1508 1371 1546
rect 1327 1488 1339 1508
rect 1359 1488 1371 1508
rect 1327 1446 1371 1488
rect 1421 1508 1463 1546
rect 1421 1488 1435 1508
rect 1455 1488 1463 1508
rect 1421 1446 1463 1488
rect 1537 1508 1579 1546
rect 1537 1488 1545 1508
rect 1565 1488 1579 1508
rect 1537 1446 1579 1488
rect 1629 1515 1674 1546
rect 1629 1508 1673 1515
rect 1629 1488 1641 1508
rect 1661 1488 1673 1508
rect 1629 1446 1673 1488
rect 312 1280 356 1318
rect 312 1260 324 1280
rect 344 1260 356 1280
rect 312 1218 356 1260
rect 406 1280 448 1318
rect 406 1260 420 1280
rect 440 1260 448 1280
rect 406 1218 448 1260
rect 530 1280 574 1318
rect 530 1260 542 1280
rect 562 1260 574 1280
rect 530 1218 574 1260
rect 624 1280 666 1318
rect 624 1260 638 1280
rect 658 1260 666 1280
rect 624 1218 666 1260
rect 740 1280 782 1318
rect 740 1260 748 1280
rect 768 1260 782 1280
rect 740 1218 782 1260
rect 832 1287 877 1318
rect 832 1280 876 1287
rect 832 1260 844 1280
rect 864 1260 876 1280
rect 832 1218 876 1260
rect 1191 900 1235 938
rect 1191 880 1203 900
rect 1223 880 1235 900
rect 1191 838 1235 880
rect 1285 900 1327 938
rect 1285 880 1299 900
rect 1319 880 1327 900
rect 1285 838 1327 880
rect 1409 900 1453 938
rect 1409 880 1421 900
rect 1441 880 1453 900
rect 1409 838 1453 880
rect 1503 900 1545 938
rect 1503 880 1517 900
rect 1537 880 1545 900
rect 1503 838 1545 880
rect 1619 900 1661 938
rect 1619 880 1627 900
rect 1647 880 1661 900
rect 1619 838 1661 880
rect 1711 907 1756 938
rect 1711 900 1755 907
rect 1711 880 1723 900
rect 1743 880 1755 900
rect 1711 838 1755 880
rect 294 674 338 712
rect 294 654 306 674
rect 326 654 338 674
rect 294 612 338 654
rect 388 674 430 712
rect 388 654 402 674
rect 422 654 430 674
rect 388 612 430 654
rect 512 674 556 712
rect 512 654 524 674
rect 544 654 556 674
rect 512 612 556 654
rect 606 674 648 712
rect 606 654 620 674
rect 640 654 648 674
rect 606 612 648 654
rect 722 674 764 712
rect 722 654 730 674
rect 750 654 764 674
rect 722 612 764 654
rect 814 681 859 712
rect 814 674 858 681
rect 814 654 826 674
rect 846 654 858 674
rect 814 612 858 654
rect 1092 490 1136 528
rect 1092 470 1104 490
rect 1124 470 1136 490
rect 1092 428 1136 470
rect 1186 490 1228 528
rect 1186 470 1200 490
rect 1220 470 1228 490
rect 1186 428 1228 470
rect 1310 490 1354 528
rect 1310 470 1322 490
rect 1342 470 1354 490
rect 1310 428 1354 470
rect 1404 490 1446 528
rect 1404 470 1418 490
rect 1438 470 1446 490
rect 1404 428 1446 470
rect 1520 490 1562 528
rect 1520 470 1528 490
rect 1548 470 1562 490
rect 1520 428 1562 470
rect 1612 497 1657 528
rect 1612 490 1656 497
rect 1612 470 1624 490
rect 1644 470 1656 490
rect 1612 428 1656 470
rect 295 262 339 300
rect 295 242 307 262
rect 327 242 339 262
rect 295 200 339 242
rect 389 262 431 300
rect 389 242 403 262
rect 423 242 431 262
rect 389 200 431 242
rect 513 262 557 300
rect 513 242 525 262
rect 545 242 557 262
rect 513 200 557 242
rect 607 262 649 300
rect 607 242 621 262
rect 641 242 649 262
rect 607 200 649 242
rect 723 262 765 300
rect 723 242 731 262
rect 751 242 765 262
rect 723 200 765 242
rect 815 269 860 300
rect 815 262 859 269
rect 815 242 827 262
rect 847 242 859 262
rect 815 200 859 242
rect 1377 -122 1421 -84
rect 1377 -142 1389 -122
rect 1409 -142 1421 -122
rect 1377 -184 1421 -142
rect 1471 -122 1513 -84
rect 1471 -142 1485 -122
rect 1505 -142 1513 -122
rect 1471 -184 1513 -142
rect 1595 -122 1639 -84
rect 1595 -142 1607 -122
rect 1627 -142 1639 -122
rect 1595 -184 1639 -142
rect 1689 -122 1731 -84
rect 1689 -142 1703 -122
rect 1723 -142 1731 -122
rect 1689 -184 1731 -142
rect 1805 -122 1847 -84
rect 1805 -142 1813 -122
rect 1833 -142 1847 -122
rect 1805 -184 1847 -142
rect 1897 -115 1942 -84
rect 1897 -122 1941 -115
rect 1897 -142 1909 -122
rect 1929 -142 1941 -122
rect 1897 -184 1941 -142
rect 275 -344 319 -306
rect 275 -364 287 -344
rect 307 -364 319 -344
rect 275 -406 319 -364
rect 369 -344 411 -306
rect 369 -364 383 -344
rect 403 -364 411 -344
rect 369 -406 411 -364
rect 493 -344 537 -306
rect 493 -364 505 -344
rect 525 -364 537 -344
rect 493 -406 537 -364
rect 587 -344 629 -306
rect 587 -364 601 -344
rect 621 -364 629 -344
rect 587 -406 629 -364
rect 703 -344 745 -306
rect 703 -364 711 -344
rect 731 -364 745 -344
rect 703 -406 745 -364
rect 795 -337 840 -306
rect 795 -344 839 -337
rect 795 -364 807 -344
rect 827 -364 839 -344
rect 795 -406 839 -364
rect 1073 -528 1117 -490
rect 1073 -548 1085 -528
rect 1105 -548 1117 -528
rect 1073 -590 1117 -548
rect 1167 -528 1209 -490
rect 1167 -548 1181 -528
rect 1201 -548 1209 -528
rect 1167 -590 1209 -548
rect 1291 -528 1335 -490
rect 1291 -548 1303 -528
rect 1323 -548 1335 -528
rect 1291 -590 1335 -548
rect 1385 -528 1427 -490
rect 1385 -548 1399 -528
rect 1419 -548 1427 -528
rect 1385 -590 1427 -548
rect 1501 -528 1543 -490
rect 1501 -548 1509 -528
rect 1529 -548 1543 -528
rect 1501 -590 1543 -548
rect 1593 -521 1638 -490
rect 1593 -528 1637 -521
rect 1593 -548 1605 -528
rect 1625 -548 1637 -528
rect 1593 -590 1637 -548
rect 276 -756 320 -718
rect 276 -776 288 -756
rect 308 -776 320 -756
rect 276 -818 320 -776
rect 370 -756 412 -718
rect 370 -776 384 -756
rect 404 -776 412 -756
rect 370 -818 412 -776
rect 494 -756 538 -718
rect 494 -776 506 -756
rect 526 -776 538 -756
rect 494 -818 538 -776
rect 588 -756 630 -718
rect 588 -776 602 -756
rect 622 -776 630 -756
rect 588 -818 630 -776
rect 704 -756 746 -718
rect 704 -776 712 -756
rect 732 -776 746 -756
rect 704 -818 746 -776
rect 796 -749 841 -718
rect 796 -756 840 -749
rect 796 -776 808 -756
rect 828 -776 840 -756
rect 796 -818 840 -776
rect 1155 -1136 1199 -1098
rect 1155 -1156 1167 -1136
rect 1187 -1156 1199 -1136
rect 1155 -1198 1199 -1156
rect 1249 -1136 1291 -1098
rect 1249 -1156 1263 -1136
rect 1283 -1156 1291 -1136
rect 1249 -1198 1291 -1156
rect 1373 -1136 1417 -1098
rect 1373 -1156 1385 -1136
rect 1405 -1156 1417 -1136
rect 1373 -1198 1417 -1156
rect 1467 -1136 1509 -1098
rect 1467 -1156 1481 -1136
rect 1501 -1156 1509 -1136
rect 1467 -1198 1509 -1156
rect 1583 -1136 1625 -1098
rect 1583 -1156 1591 -1136
rect 1611 -1156 1625 -1136
rect 1583 -1198 1625 -1156
rect 1675 -1129 1720 -1098
rect 1675 -1136 1719 -1129
rect 1675 -1156 1687 -1136
rect 1707 -1156 1719 -1136
rect 1675 -1198 1719 -1156
rect 258 -1362 302 -1324
rect 258 -1382 270 -1362
rect 290 -1382 302 -1362
rect 258 -1424 302 -1382
rect 352 -1362 394 -1324
rect 352 -1382 366 -1362
rect 386 -1382 394 -1362
rect 352 -1424 394 -1382
rect 476 -1362 520 -1324
rect 476 -1382 488 -1362
rect 508 -1382 520 -1362
rect 476 -1424 520 -1382
rect 570 -1362 612 -1324
rect 570 -1382 584 -1362
rect 604 -1382 612 -1362
rect 570 -1424 612 -1382
rect 686 -1362 728 -1324
rect 686 -1382 694 -1362
rect 714 -1382 728 -1362
rect 686 -1424 728 -1382
rect 778 -1355 823 -1324
rect 778 -1362 822 -1355
rect 778 -1382 790 -1362
rect 810 -1382 822 -1362
rect 778 -1424 822 -1382
rect 1056 -1546 1100 -1508
rect 1056 -1566 1068 -1546
rect 1088 -1566 1100 -1546
rect 1056 -1608 1100 -1566
rect 1150 -1546 1192 -1508
rect 1150 -1566 1164 -1546
rect 1184 -1566 1192 -1546
rect 1150 -1608 1192 -1566
rect 1274 -1546 1318 -1508
rect 1274 -1566 1286 -1546
rect 1306 -1566 1318 -1546
rect 1274 -1608 1318 -1566
rect 1368 -1546 1410 -1508
rect 1368 -1566 1382 -1546
rect 1402 -1566 1410 -1546
rect 1368 -1608 1410 -1566
rect 1484 -1546 1526 -1508
rect 1484 -1566 1492 -1546
rect 1512 -1566 1526 -1546
rect 1484 -1608 1526 -1566
rect 1576 -1539 1621 -1508
rect 1576 -1546 1620 -1539
rect 1576 -1566 1588 -1546
rect 1608 -1566 1620 -1546
rect 1576 -1608 1620 -1566
rect 259 -1774 303 -1736
rect 259 -1794 271 -1774
rect 291 -1794 303 -1774
rect 259 -1836 303 -1794
rect 353 -1774 395 -1736
rect 353 -1794 367 -1774
rect 387 -1794 395 -1774
rect 353 -1836 395 -1794
rect 477 -1774 521 -1736
rect 477 -1794 489 -1774
rect 509 -1794 521 -1774
rect 477 -1836 521 -1794
rect 571 -1774 613 -1736
rect 571 -1794 585 -1774
rect 605 -1794 613 -1774
rect 571 -1836 613 -1794
rect 687 -1774 729 -1736
rect 687 -1794 695 -1774
rect 715 -1794 729 -1774
rect 687 -1836 729 -1794
rect 779 -1767 824 -1736
rect 779 -1774 823 -1767
rect 779 -1794 791 -1774
rect 811 -1794 823 -1774
rect 779 -1836 823 -1794
rect 1201 -2156 1245 -2118
rect 1201 -2176 1213 -2156
rect 1233 -2176 1245 -2156
rect 1201 -2218 1245 -2176
rect 1295 -2156 1337 -2118
rect 1295 -2176 1309 -2156
rect 1329 -2176 1337 -2156
rect 1295 -2218 1337 -2176
rect 1419 -2156 1463 -2118
rect 1419 -2176 1431 -2156
rect 1451 -2176 1463 -2156
rect 1419 -2218 1463 -2176
rect 1513 -2156 1555 -2118
rect 1513 -2176 1527 -2156
rect 1547 -2176 1555 -2156
rect 1513 -2218 1555 -2176
rect 1629 -2156 1671 -2118
rect 1629 -2176 1637 -2156
rect 1657 -2176 1671 -2156
rect 1629 -2218 1671 -2176
rect 1721 -2149 1766 -2118
rect 1721 -2156 1765 -2149
rect 1721 -2176 1733 -2156
rect 1753 -2176 1765 -2156
rect 1721 -2218 1765 -2176
rect 238 -2380 282 -2342
rect 238 -2400 250 -2380
rect 270 -2400 282 -2380
rect 238 -2442 282 -2400
rect 332 -2380 374 -2342
rect 332 -2400 346 -2380
rect 366 -2400 374 -2380
rect 332 -2442 374 -2400
rect 456 -2380 500 -2342
rect 456 -2400 468 -2380
rect 488 -2400 500 -2380
rect 456 -2442 500 -2400
rect 550 -2380 592 -2342
rect 550 -2400 564 -2380
rect 584 -2400 592 -2380
rect 550 -2442 592 -2400
rect 666 -2380 708 -2342
rect 666 -2400 674 -2380
rect 694 -2400 708 -2380
rect 666 -2442 708 -2400
rect 758 -2373 803 -2342
rect 758 -2380 802 -2373
rect 758 -2400 770 -2380
rect 790 -2400 802 -2380
rect 758 -2442 802 -2400
rect 1036 -2564 1080 -2526
rect 1036 -2584 1048 -2564
rect 1068 -2584 1080 -2564
rect 1036 -2626 1080 -2584
rect 1130 -2564 1172 -2526
rect 1130 -2584 1144 -2564
rect 1164 -2584 1172 -2564
rect 1130 -2626 1172 -2584
rect 1254 -2564 1298 -2526
rect 1254 -2584 1266 -2564
rect 1286 -2584 1298 -2564
rect 1254 -2626 1298 -2584
rect 1348 -2564 1390 -2526
rect 1348 -2584 1362 -2564
rect 1382 -2584 1390 -2564
rect 1348 -2626 1390 -2584
rect 1464 -2564 1506 -2526
rect 1464 -2584 1472 -2564
rect 1492 -2584 1506 -2564
rect 1464 -2626 1506 -2584
rect 1556 -2557 1601 -2526
rect 1556 -2564 1600 -2557
rect 1556 -2584 1568 -2564
rect 1588 -2584 1600 -2564
rect 1556 -2626 1600 -2584
rect 239 -2792 283 -2754
rect 239 -2812 251 -2792
rect 271 -2812 283 -2792
rect 239 -2854 283 -2812
rect 333 -2792 375 -2754
rect 333 -2812 347 -2792
rect 367 -2812 375 -2792
rect 333 -2854 375 -2812
rect 457 -2792 501 -2754
rect 457 -2812 469 -2792
rect 489 -2812 501 -2792
rect 457 -2854 501 -2812
rect 551 -2792 593 -2754
rect 551 -2812 565 -2792
rect 585 -2812 593 -2792
rect 551 -2854 593 -2812
rect 667 -2792 709 -2754
rect 667 -2812 675 -2792
rect 695 -2812 709 -2792
rect 667 -2854 709 -2812
rect 759 -2785 804 -2754
rect 759 -2792 803 -2785
rect 759 -2812 771 -2792
rect 791 -2812 803 -2792
rect 759 -2854 803 -2812
rect 1118 -3172 1162 -3134
rect 1118 -3192 1130 -3172
rect 1150 -3192 1162 -3172
rect 1118 -3234 1162 -3192
rect 1212 -3172 1254 -3134
rect 1212 -3192 1226 -3172
rect 1246 -3192 1254 -3172
rect 1212 -3234 1254 -3192
rect 1336 -3172 1380 -3134
rect 1336 -3192 1348 -3172
rect 1368 -3192 1380 -3172
rect 1336 -3234 1380 -3192
rect 1430 -3172 1472 -3134
rect 1430 -3192 1444 -3172
rect 1464 -3192 1472 -3172
rect 1430 -3234 1472 -3192
rect 1546 -3172 1588 -3134
rect 1546 -3192 1554 -3172
rect 1574 -3192 1588 -3172
rect 1546 -3234 1588 -3192
rect 1638 -3165 1683 -3134
rect 1638 -3172 1682 -3165
rect 1638 -3192 1650 -3172
rect 1670 -3192 1682 -3172
rect 1638 -3234 1682 -3192
rect 221 -3398 265 -3360
rect 221 -3418 233 -3398
rect 253 -3418 265 -3398
rect 221 -3460 265 -3418
rect 315 -3398 357 -3360
rect 315 -3418 329 -3398
rect 349 -3418 357 -3398
rect 315 -3460 357 -3418
rect 439 -3398 483 -3360
rect 439 -3418 451 -3398
rect 471 -3418 483 -3398
rect 439 -3460 483 -3418
rect 533 -3398 575 -3360
rect 533 -3418 547 -3398
rect 567 -3418 575 -3398
rect 533 -3460 575 -3418
rect 649 -3398 691 -3360
rect 649 -3418 657 -3398
rect 677 -3418 691 -3398
rect 649 -3460 691 -3418
rect 741 -3391 786 -3360
rect 741 -3398 785 -3391
rect 741 -3418 753 -3398
rect 773 -3418 785 -3398
rect 741 -3460 785 -3418
rect 1019 -3582 1063 -3544
rect 1019 -3602 1031 -3582
rect 1051 -3602 1063 -3582
rect 1019 -3644 1063 -3602
rect 1113 -3582 1155 -3544
rect 1113 -3602 1127 -3582
rect 1147 -3602 1155 -3582
rect 1113 -3644 1155 -3602
rect 1237 -3582 1281 -3544
rect 1237 -3602 1249 -3582
rect 1269 -3602 1281 -3582
rect 1237 -3644 1281 -3602
rect 1331 -3582 1373 -3544
rect 1331 -3602 1345 -3582
rect 1365 -3602 1373 -3582
rect 1331 -3644 1373 -3602
rect 1447 -3582 1489 -3544
rect 1447 -3602 1455 -3582
rect 1475 -3602 1489 -3582
rect 1447 -3644 1489 -3602
rect 1539 -3575 1584 -3544
rect 1539 -3582 1583 -3575
rect 1539 -3602 1551 -3582
rect 1571 -3602 1583 -3582
rect 1539 -3644 1583 -3602
rect 222 -3810 266 -3772
rect 222 -3830 234 -3810
rect 254 -3830 266 -3810
rect 222 -3872 266 -3830
rect 316 -3810 358 -3772
rect 316 -3830 330 -3810
rect 350 -3830 358 -3810
rect 316 -3872 358 -3830
rect 440 -3810 484 -3772
rect 440 -3830 452 -3810
rect 472 -3830 484 -3810
rect 440 -3872 484 -3830
rect 534 -3810 576 -3772
rect 534 -3830 548 -3810
rect 568 -3830 576 -3810
rect 534 -3872 576 -3830
rect 650 -3810 692 -3772
rect 650 -3830 658 -3810
rect 678 -3830 692 -3810
rect 650 -3872 692 -3830
rect 742 -3803 787 -3772
rect 742 -3810 786 -3803
rect 742 -3830 754 -3810
rect 774 -3830 786 -3810
rect 742 -3872 786 -3830
<< ndiffc >>
rect 190 3966 208 3984
rect 188 3867 206 3885
rect 185 3642 203 3660
rect 183 3543 201 3561
rect 354 3559 374 3579
rect 457 3563 477 3583
rect 572 3559 592 3579
rect 675 3563 695 3583
rect 783 3563 803 3583
rect 886 3559 906 3579
rect 179 3459 197 3477
rect 177 3360 195 3378
rect 1152 3375 1172 3395
rect 1255 3379 1275 3399
rect 1370 3375 1390 3395
rect 1473 3379 1493 3399
rect 1581 3379 1601 3399
rect 1684 3375 1704 3395
rect 172 3241 190 3259
rect 170 3142 188 3160
rect 355 3147 375 3167
rect 458 3151 478 3171
rect 573 3147 593 3167
rect 676 3151 696 3171
rect 784 3151 804 3171
rect 887 3147 907 3167
rect 173 2948 191 2966
rect 171 2849 189 2867
rect 1234 2767 1254 2787
rect 1337 2771 1357 2791
rect 1452 2767 1472 2787
rect 1555 2771 1575 2791
rect 1663 2771 1683 2791
rect 1766 2767 1786 2787
rect 168 2624 186 2642
rect 166 2525 184 2543
rect 337 2541 357 2561
rect 440 2545 460 2565
rect 555 2541 575 2561
rect 658 2545 678 2565
rect 766 2545 786 2565
rect 869 2541 889 2561
rect 162 2441 180 2459
rect 160 2342 178 2360
rect 1135 2357 1155 2377
rect 1238 2361 1258 2381
rect 1353 2357 1373 2377
rect 1456 2361 1476 2381
rect 1564 2361 1584 2381
rect 1667 2357 1687 2377
rect 155 2223 173 2241
rect 153 2124 171 2142
rect 338 2129 358 2149
rect 441 2133 461 2153
rect 556 2129 576 2149
rect 659 2133 679 2153
rect 767 2133 787 2153
rect 870 2129 890 2149
rect 153 1930 171 1948
rect 151 1831 169 1849
rect 1280 1747 1300 1767
rect 1383 1751 1403 1771
rect 1498 1747 1518 1767
rect 1601 1751 1621 1771
rect 1709 1751 1729 1771
rect 1812 1747 1832 1767
rect 148 1606 166 1624
rect 146 1507 164 1525
rect 317 1523 337 1543
rect 420 1527 440 1547
rect 535 1523 555 1543
rect 638 1527 658 1547
rect 746 1527 766 1547
rect 849 1523 869 1543
rect 142 1423 160 1441
rect 140 1324 158 1342
rect 1115 1339 1135 1359
rect 1218 1343 1238 1363
rect 1333 1339 1353 1359
rect 1436 1343 1456 1363
rect 1544 1343 1564 1363
rect 1647 1339 1667 1359
rect 135 1205 153 1223
rect 133 1106 151 1124
rect 318 1111 338 1131
rect 421 1115 441 1135
rect 536 1111 556 1131
rect 639 1115 659 1135
rect 747 1115 767 1135
rect 850 1111 870 1131
rect 136 912 154 930
rect 134 813 152 831
rect 1197 731 1217 751
rect 1300 735 1320 755
rect 1415 731 1435 751
rect 1518 735 1538 755
rect 1626 735 1646 755
rect 1729 731 1749 751
rect 131 588 149 606
rect 129 489 147 507
rect 300 505 320 525
rect 403 509 423 529
rect 518 505 538 525
rect 621 509 641 529
rect 729 509 749 529
rect 832 505 852 525
rect 125 405 143 423
rect 123 306 141 324
rect 1098 321 1118 341
rect 1201 325 1221 345
rect 1316 321 1336 341
rect 1419 325 1439 345
rect 1527 325 1547 345
rect 1630 321 1650 341
rect 118 187 136 205
rect 116 88 134 106
rect 301 93 321 113
rect 404 97 424 117
rect 519 93 539 113
rect 622 97 642 117
rect 730 97 750 117
rect 833 93 853 113
rect 117 -106 135 -88
rect 115 -205 133 -187
rect 1383 -291 1403 -271
rect 1486 -287 1506 -267
rect 1601 -291 1621 -271
rect 1704 -287 1724 -267
rect 1812 -287 1832 -267
rect 1915 -291 1935 -271
rect 112 -430 130 -412
rect 110 -529 128 -511
rect 281 -513 301 -493
rect 384 -509 404 -489
rect 499 -513 519 -493
rect 602 -509 622 -489
rect 710 -509 730 -489
rect 813 -513 833 -493
rect 106 -613 124 -595
rect 104 -712 122 -694
rect 1079 -697 1099 -677
rect 1182 -693 1202 -673
rect 1297 -697 1317 -677
rect 1400 -693 1420 -673
rect 1508 -693 1528 -673
rect 1611 -697 1631 -677
rect 99 -831 117 -813
rect 97 -930 115 -912
rect 282 -925 302 -905
rect 385 -921 405 -901
rect 500 -925 520 -905
rect 603 -921 623 -901
rect 711 -921 731 -901
rect 814 -925 834 -905
rect 100 -1124 118 -1106
rect 98 -1223 116 -1205
rect 1161 -1305 1181 -1285
rect 1264 -1301 1284 -1281
rect 1379 -1305 1399 -1285
rect 1482 -1301 1502 -1281
rect 1590 -1301 1610 -1281
rect 1693 -1305 1713 -1285
rect 95 -1448 113 -1430
rect 93 -1547 111 -1529
rect 264 -1531 284 -1511
rect 367 -1527 387 -1507
rect 482 -1531 502 -1511
rect 585 -1527 605 -1507
rect 693 -1527 713 -1507
rect 796 -1531 816 -1511
rect 89 -1631 107 -1613
rect 87 -1730 105 -1712
rect 1062 -1715 1082 -1695
rect 1165 -1711 1185 -1691
rect 1280 -1715 1300 -1695
rect 1383 -1711 1403 -1691
rect 1491 -1711 1511 -1691
rect 1594 -1715 1614 -1695
rect 82 -1849 100 -1831
rect 80 -1948 98 -1930
rect 265 -1943 285 -1923
rect 368 -1939 388 -1919
rect 483 -1943 503 -1923
rect 586 -1939 606 -1919
rect 694 -1939 714 -1919
rect 797 -1943 817 -1923
rect 80 -2142 98 -2124
rect 78 -2241 96 -2223
rect 1207 -2325 1227 -2305
rect 1310 -2321 1330 -2301
rect 1425 -2325 1445 -2305
rect 1528 -2321 1548 -2301
rect 1636 -2321 1656 -2301
rect 1739 -2325 1759 -2305
rect 75 -2466 93 -2448
rect 73 -2565 91 -2547
rect 244 -2549 264 -2529
rect 347 -2545 367 -2525
rect 462 -2549 482 -2529
rect 565 -2545 585 -2525
rect 673 -2545 693 -2525
rect 776 -2549 796 -2529
rect 69 -2649 87 -2631
rect 67 -2748 85 -2730
rect 1042 -2733 1062 -2713
rect 1145 -2729 1165 -2709
rect 1260 -2733 1280 -2713
rect 1363 -2729 1383 -2709
rect 1471 -2729 1491 -2709
rect 1574 -2733 1594 -2713
rect 62 -2867 80 -2849
rect 60 -2966 78 -2948
rect 245 -2961 265 -2941
rect 348 -2957 368 -2937
rect 463 -2961 483 -2941
rect 566 -2957 586 -2937
rect 674 -2957 694 -2937
rect 777 -2961 797 -2941
rect 63 -3160 81 -3142
rect 61 -3259 79 -3241
rect 1124 -3341 1144 -3321
rect 1227 -3337 1247 -3317
rect 1342 -3341 1362 -3321
rect 1445 -3337 1465 -3317
rect 1553 -3337 1573 -3317
rect 1656 -3341 1676 -3321
rect 58 -3484 76 -3466
rect 56 -3583 74 -3565
rect 227 -3567 247 -3547
rect 330 -3563 350 -3543
rect 445 -3567 465 -3547
rect 548 -3563 568 -3543
rect 656 -3563 676 -3543
rect 759 -3567 779 -3547
rect 52 -3667 70 -3649
rect 50 -3766 68 -3748
rect 1025 -3751 1045 -3731
rect 1128 -3747 1148 -3727
rect 1243 -3751 1263 -3731
rect 1346 -3747 1366 -3727
rect 1454 -3747 1474 -3727
rect 1557 -3751 1577 -3731
rect 45 -3885 63 -3867
rect 43 -3984 61 -3966
rect 228 -3979 248 -3959
rect 331 -3975 351 -3955
rect 446 -3979 466 -3959
rect 549 -3975 569 -3955
rect 657 -3975 677 -3955
rect 760 -3979 780 -3959
<< pdiffc >>
rect 360 3708 380 3728
rect 456 3708 476 3728
rect 578 3708 598 3728
rect 674 3708 694 3728
rect 784 3708 804 3728
rect 880 3708 900 3728
rect 1158 3524 1178 3544
rect 1254 3524 1274 3544
rect 1376 3524 1396 3544
rect 1472 3524 1492 3544
rect 1582 3524 1602 3544
rect 1678 3524 1698 3544
rect 361 3296 381 3316
rect 457 3296 477 3316
rect 579 3296 599 3316
rect 675 3296 695 3316
rect 785 3296 805 3316
rect 881 3296 901 3316
rect 1240 2916 1260 2936
rect 1336 2916 1356 2936
rect 1458 2916 1478 2936
rect 1554 2916 1574 2936
rect 1664 2916 1684 2936
rect 1760 2916 1780 2936
rect 343 2690 363 2710
rect 439 2690 459 2710
rect 561 2690 581 2710
rect 657 2690 677 2710
rect 767 2690 787 2710
rect 863 2690 883 2710
rect 1141 2506 1161 2526
rect 1237 2506 1257 2526
rect 1359 2506 1379 2526
rect 1455 2506 1475 2526
rect 1565 2506 1585 2526
rect 1661 2506 1681 2526
rect 344 2278 364 2298
rect 440 2278 460 2298
rect 562 2278 582 2298
rect 658 2278 678 2298
rect 768 2278 788 2298
rect 864 2278 884 2298
rect 1286 1896 1306 1916
rect 1382 1896 1402 1916
rect 1504 1896 1524 1916
rect 1600 1896 1620 1916
rect 1710 1896 1730 1916
rect 1806 1896 1826 1916
rect 323 1672 343 1692
rect 419 1672 439 1692
rect 541 1672 561 1692
rect 637 1672 657 1692
rect 747 1672 767 1692
rect 843 1672 863 1692
rect 1121 1488 1141 1508
rect 1217 1488 1237 1508
rect 1339 1488 1359 1508
rect 1435 1488 1455 1508
rect 1545 1488 1565 1508
rect 1641 1488 1661 1508
rect 324 1260 344 1280
rect 420 1260 440 1280
rect 542 1260 562 1280
rect 638 1260 658 1280
rect 748 1260 768 1280
rect 844 1260 864 1280
rect 1203 880 1223 900
rect 1299 880 1319 900
rect 1421 880 1441 900
rect 1517 880 1537 900
rect 1627 880 1647 900
rect 1723 880 1743 900
rect 306 654 326 674
rect 402 654 422 674
rect 524 654 544 674
rect 620 654 640 674
rect 730 654 750 674
rect 826 654 846 674
rect 1104 470 1124 490
rect 1200 470 1220 490
rect 1322 470 1342 490
rect 1418 470 1438 490
rect 1528 470 1548 490
rect 1624 470 1644 490
rect 307 242 327 262
rect 403 242 423 262
rect 525 242 545 262
rect 621 242 641 262
rect 731 242 751 262
rect 827 242 847 262
rect 1389 -142 1409 -122
rect 1485 -142 1505 -122
rect 1607 -142 1627 -122
rect 1703 -142 1723 -122
rect 1813 -142 1833 -122
rect 1909 -142 1929 -122
rect 287 -364 307 -344
rect 383 -364 403 -344
rect 505 -364 525 -344
rect 601 -364 621 -344
rect 711 -364 731 -344
rect 807 -364 827 -344
rect 1085 -548 1105 -528
rect 1181 -548 1201 -528
rect 1303 -548 1323 -528
rect 1399 -548 1419 -528
rect 1509 -548 1529 -528
rect 1605 -548 1625 -528
rect 288 -776 308 -756
rect 384 -776 404 -756
rect 506 -776 526 -756
rect 602 -776 622 -756
rect 712 -776 732 -756
rect 808 -776 828 -756
rect 1167 -1156 1187 -1136
rect 1263 -1156 1283 -1136
rect 1385 -1156 1405 -1136
rect 1481 -1156 1501 -1136
rect 1591 -1156 1611 -1136
rect 1687 -1156 1707 -1136
rect 270 -1382 290 -1362
rect 366 -1382 386 -1362
rect 488 -1382 508 -1362
rect 584 -1382 604 -1362
rect 694 -1382 714 -1362
rect 790 -1382 810 -1362
rect 1068 -1566 1088 -1546
rect 1164 -1566 1184 -1546
rect 1286 -1566 1306 -1546
rect 1382 -1566 1402 -1546
rect 1492 -1566 1512 -1546
rect 1588 -1566 1608 -1546
rect 271 -1794 291 -1774
rect 367 -1794 387 -1774
rect 489 -1794 509 -1774
rect 585 -1794 605 -1774
rect 695 -1794 715 -1774
rect 791 -1794 811 -1774
rect 1213 -2176 1233 -2156
rect 1309 -2176 1329 -2156
rect 1431 -2176 1451 -2156
rect 1527 -2176 1547 -2156
rect 1637 -2176 1657 -2156
rect 1733 -2176 1753 -2156
rect 250 -2400 270 -2380
rect 346 -2400 366 -2380
rect 468 -2400 488 -2380
rect 564 -2400 584 -2380
rect 674 -2400 694 -2380
rect 770 -2400 790 -2380
rect 1048 -2584 1068 -2564
rect 1144 -2584 1164 -2564
rect 1266 -2584 1286 -2564
rect 1362 -2584 1382 -2564
rect 1472 -2584 1492 -2564
rect 1568 -2584 1588 -2564
rect 251 -2812 271 -2792
rect 347 -2812 367 -2792
rect 469 -2812 489 -2792
rect 565 -2812 585 -2792
rect 675 -2812 695 -2792
rect 771 -2812 791 -2792
rect 1130 -3192 1150 -3172
rect 1226 -3192 1246 -3172
rect 1348 -3192 1368 -3172
rect 1444 -3192 1464 -3172
rect 1554 -3192 1574 -3172
rect 1650 -3192 1670 -3172
rect 233 -3418 253 -3398
rect 329 -3418 349 -3398
rect 451 -3418 471 -3398
rect 547 -3418 567 -3398
rect 657 -3418 677 -3398
rect 753 -3418 773 -3398
rect 1031 -3602 1051 -3582
rect 1127 -3602 1147 -3582
rect 1249 -3602 1269 -3582
rect 1345 -3602 1365 -3582
rect 1455 -3602 1475 -3582
rect 1551 -3602 1571 -3582
rect 234 -3830 254 -3810
rect 330 -3830 350 -3810
rect 452 -3830 472 -3810
rect 548 -3830 568 -3810
rect 658 -3830 678 -3810
rect 754 -3830 774 -3810
<< poly >>
rect 392 3766 442 3779
rect 610 3766 660 3779
rect 818 3766 868 3779
rect 392 3638 442 3666
rect 392 3618 405 3638
rect 425 3618 442 3638
rect 392 3589 442 3618
rect 610 3641 660 3666
rect 610 3621 623 3641
rect 643 3621 660 3641
rect 610 3589 660 3621
rect 818 3639 868 3666
rect 818 3619 841 3639
rect 861 3619 868 3639
rect 818 3589 868 3619
rect 1190 3582 1240 3595
rect 1408 3582 1458 3595
rect 1616 3582 1666 3595
rect 392 3531 442 3547
rect 610 3531 660 3547
rect 818 3531 868 3547
rect 1190 3454 1240 3482
rect 1190 3434 1203 3454
rect 1223 3434 1240 3454
rect 1190 3405 1240 3434
rect 1408 3457 1458 3482
rect 1408 3437 1421 3457
rect 1441 3437 1458 3457
rect 1408 3405 1458 3437
rect 1616 3455 1666 3482
rect 1616 3435 1639 3455
rect 1659 3435 1666 3455
rect 1616 3405 1666 3435
rect 393 3354 443 3367
rect 611 3354 661 3367
rect 819 3354 869 3367
rect 1190 3347 1240 3363
rect 1408 3347 1458 3363
rect 1616 3347 1666 3363
rect 393 3226 443 3254
rect 393 3206 406 3226
rect 426 3206 443 3226
rect 393 3177 443 3206
rect 611 3229 661 3254
rect 611 3209 624 3229
rect 644 3209 661 3229
rect 611 3177 661 3209
rect 819 3227 869 3254
rect 819 3207 842 3227
rect 862 3207 869 3227
rect 819 3177 869 3207
rect 393 3119 443 3135
rect 611 3119 661 3135
rect 819 3119 869 3135
rect 1272 2974 1322 2987
rect 1490 2974 1540 2987
rect 1698 2974 1748 2987
rect 1272 2846 1322 2874
rect 1272 2826 1285 2846
rect 1305 2826 1322 2846
rect 1272 2797 1322 2826
rect 1490 2849 1540 2874
rect 1490 2829 1503 2849
rect 1523 2829 1540 2849
rect 1490 2797 1540 2829
rect 1698 2847 1748 2874
rect 1698 2827 1721 2847
rect 1741 2827 1748 2847
rect 1698 2797 1748 2827
rect 375 2748 425 2761
rect 593 2748 643 2761
rect 801 2748 851 2761
rect 1272 2739 1322 2755
rect 1490 2739 1540 2755
rect 1698 2739 1748 2755
rect 375 2620 425 2648
rect 375 2600 388 2620
rect 408 2600 425 2620
rect 375 2571 425 2600
rect 593 2623 643 2648
rect 593 2603 606 2623
rect 626 2603 643 2623
rect 593 2571 643 2603
rect 801 2621 851 2648
rect 801 2601 824 2621
rect 844 2601 851 2621
rect 801 2571 851 2601
rect 1173 2564 1223 2577
rect 1391 2564 1441 2577
rect 1599 2564 1649 2577
rect 375 2513 425 2529
rect 593 2513 643 2529
rect 801 2513 851 2529
rect 1173 2436 1223 2464
rect 1173 2416 1186 2436
rect 1206 2416 1223 2436
rect 1173 2387 1223 2416
rect 1391 2439 1441 2464
rect 1391 2419 1404 2439
rect 1424 2419 1441 2439
rect 1391 2387 1441 2419
rect 1599 2437 1649 2464
rect 1599 2417 1622 2437
rect 1642 2417 1649 2437
rect 1599 2387 1649 2417
rect 376 2336 426 2349
rect 594 2336 644 2349
rect 802 2336 852 2349
rect 1173 2329 1223 2345
rect 1391 2329 1441 2345
rect 1599 2329 1649 2345
rect 376 2208 426 2236
rect 376 2188 389 2208
rect 409 2188 426 2208
rect 376 2159 426 2188
rect 594 2211 644 2236
rect 594 2191 607 2211
rect 627 2191 644 2211
rect 594 2159 644 2191
rect 802 2209 852 2236
rect 802 2189 825 2209
rect 845 2189 852 2209
rect 802 2159 852 2189
rect 376 2101 426 2117
rect 594 2101 644 2117
rect 802 2101 852 2117
rect 1318 1954 1368 1967
rect 1536 1954 1586 1967
rect 1744 1954 1794 1967
rect 1318 1826 1368 1854
rect 1318 1806 1331 1826
rect 1351 1806 1368 1826
rect 1318 1777 1368 1806
rect 1536 1829 1586 1854
rect 1536 1809 1549 1829
rect 1569 1809 1586 1829
rect 1536 1777 1586 1809
rect 1744 1827 1794 1854
rect 1744 1807 1767 1827
rect 1787 1807 1794 1827
rect 1744 1777 1794 1807
rect 355 1730 405 1743
rect 573 1730 623 1743
rect 781 1730 831 1743
rect 1318 1719 1368 1735
rect 1536 1719 1586 1735
rect 1744 1719 1794 1735
rect 355 1602 405 1630
rect 355 1582 368 1602
rect 388 1582 405 1602
rect 355 1553 405 1582
rect 573 1605 623 1630
rect 573 1585 586 1605
rect 606 1585 623 1605
rect 573 1553 623 1585
rect 781 1603 831 1630
rect 781 1583 804 1603
rect 824 1583 831 1603
rect 781 1553 831 1583
rect 1153 1546 1203 1559
rect 1371 1546 1421 1559
rect 1579 1546 1629 1559
rect 355 1495 405 1511
rect 573 1495 623 1511
rect 781 1495 831 1511
rect 1153 1418 1203 1446
rect 1153 1398 1166 1418
rect 1186 1398 1203 1418
rect 1153 1369 1203 1398
rect 1371 1421 1421 1446
rect 1371 1401 1384 1421
rect 1404 1401 1421 1421
rect 1371 1369 1421 1401
rect 1579 1419 1629 1446
rect 1579 1399 1602 1419
rect 1622 1399 1629 1419
rect 1579 1369 1629 1399
rect 356 1318 406 1331
rect 574 1318 624 1331
rect 782 1318 832 1331
rect 1153 1311 1203 1327
rect 1371 1311 1421 1327
rect 1579 1311 1629 1327
rect 356 1190 406 1218
rect 356 1170 369 1190
rect 389 1170 406 1190
rect 356 1141 406 1170
rect 574 1193 624 1218
rect 574 1173 587 1193
rect 607 1173 624 1193
rect 574 1141 624 1173
rect 782 1191 832 1218
rect 782 1171 805 1191
rect 825 1171 832 1191
rect 782 1141 832 1171
rect 356 1083 406 1099
rect 574 1083 624 1099
rect 782 1083 832 1099
rect 1235 938 1285 951
rect 1453 938 1503 951
rect 1661 938 1711 951
rect 1235 810 1285 838
rect 1235 790 1248 810
rect 1268 790 1285 810
rect 1235 761 1285 790
rect 1453 813 1503 838
rect 1453 793 1466 813
rect 1486 793 1503 813
rect 1453 761 1503 793
rect 1661 811 1711 838
rect 1661 791 1684 811
rect 1704 791 1711 811
rect 1661 761 1711 791
rect 338 712 388 725
rect 556 712 606 725
rect 764 712 814 725
rect 1235 703 1285 719
rect 1453 703 1503 719
rect 1661 703 1711 719
rect 338 584 388 612
rect 338 564 351 584
rect 371 564 388 584
rect 338 535 388 564
rect 556 587 606 612
rect 556 567 569 587
rect 589 567 606 587
rect 556 535 606 567
rect 764 585 814 612
rect 764 565 787 585
rect 807 565 814 585
rect 764 535 814 565
rect 1136 528 1186 541
rect 1354 528 1404 541
rect 1562 528 1612 541
rect 338 477 388 493
rect 556 477 606 493
rect 764 477 814 493
rect 1136 400 1186 428
rect 1136 380 1149 400
rect 1169 380 1186 400
rect 1136 351 1186 380
rect 1354 403 1404 428
rect 1354 383 1367 403
rect 1387 383 1404 403
rect 1354 351 1404 383
rect 1562 401 1612 428
rect 1562 381 1585 401
rect 1605 381 1612 401
rect 1562 351 1612 381
rect 339 300 389 313
rect 557 300 607 313
rect 765 300 815 313
rect 1136 293 1186 309
rect 1354 293 1404 309
rect 1562 293 1612 309
rect 339 172 389 200
rect 339 152 352 172
rect 372 152 389 172
rect 339 123 389 152
rect 557 175 607 200
rect 557 155 570 175
rect 590 155 607 175
rect 557 123 607 155
rect 765 173 815 200
rect 765 153 788 173
rect 808 153 815 173
rect 765 123 815 153
rect 339 65 389 81
rect 557 65 607 81
rect 765 65 815 81
rect 1421 -84 1471 -71
rect 1639 -84 1689 -71
rect 1847 -84 1897 -71
rect 1421 -212 1471 -184
rect 1421 -232 1434 -212
rect 1454 -232 1471 -212
rect 1421 -261 1471 -232
rect 1639 -209 1689 -184
rect 1639 -229 1652 -209
rect 1672 -229 1689 -209
rect 1639 -261 1689 -229
rect 1847 -211 1897 -184
rect 1847 -231 1870 -211
rect 1890 -231 1897 -211
rect 1847 -261 1897 -231
rect 319 -306 369 -293
rect 537 -306 587 -293
rect 745 -306 795 -293
rect 1421 -319 1471 -303
rect 1639 -319 1689 -303
rect 1847 -319 1897 -303
rect 319 -434 369 -406
rect 319 -454 332 -434
rect 352 -454 369 -434
rect 319 -483 369 -454
rect 537 -431 587 -406
rect 537 -451 550 -431
rect 570 -451 587 -431
rect 537 -483 587 -451
rect 745 -433 795 -406
rect 745 -453 768 -433
rect 788 -453 795 -433
rect 745 -483 795 -453
rect 1117 -490 1167 -477
rect 1335 -490 1385 -477
rect 1543 -490 1593 -477
rect 319 -541 369 -525
rect 537 -541 587 -525
rect 745 -541 795 -525
rect 1117 -618 1167 -590
rect 1117 -638 1130 -618
rect 1150 -638 1167 -618
rect 1117 -667 1167 -638
rect 1335 -615 1385 -590
rect 1335 -635 1348 -615
rect 1368 -635 1385 -615
rect 1335 -667 1385 -635
rect 1543 -617 1593 -590
rect 1543 -637 1566 -617
rect 1586 -637 1593 -617
rect 1543 -667 1593 -637
rect 320 -718 370 -705
rect 538 -718 588 -705
rect 746 -718 796 -705
rect 1117 -725 1167 -709
rect 1335 -725 1385 -709
rect 1543 -725 1593 -709
rect 320 -846 370 -818
rect 320 -866 333 -846
rect 353 -866 370 -846
rect 320 -895 370 -866
rect 538 -843 588 -818
rect 538 -863 551 -843
rect 571 -863 588 -843
rect 538 -895 588 -863
rect 746 -845 796 -818
rect 746 -865 769 -845
rect 789 -865 796 -845
rect 746 -895 796 -865
rect 320 -953 370 -937
rect 538 -953 588 -937
rect 746 -953 796 -937
rect 1199 -1098 1249 -1085
rect 1417 -1098 1467 -1085
rect 1625 -1098 1675 -1085
rect 1199 -1226 1249 -1198
rect 1199 -1246 1212 -1226
rect 1232 -1246 1249 -1226
rect 1199 -1275 1249 -1246
rect 1417 -1223 1467 -1198
rect 1417 -1243 1430 -1223
rect 1450 -1243 1467 -1223
rect 1417 -1275 1467 -1243
rect 1625 -1225 1675 -1198
rect 1625 -1245 1648 -1225
rect 1668 -1245 1675 -1225
rect 1625 -1275 1675 -1245
rect 302 -1324 352 -1311
rect 520 -1324 570 -1311
rect 728 -1324 778 -1311
rect 1199 -1333 1249 -1317
rect 1417 -1333 1467 -1317
rect 1625 -1333 1675 -1317
rect 302 -1452 352 -1424
rect 302 -1472 315 -1452
rect 335 -1472 352 -1452
rect 302 -1501 352 -1472
rect 520 -1449 570 -1424
rect 520 -1469 533 -1449
rect 553 -1469 570 -1449
rect 520 -1501 570 -1469
rect 728 -1451 778 -1424
rect 728 -1471 751 -1451
rect 771 -1471 778 -1451
rect 728 -1501 778 -1471
rect 1100 -1508 1150 -1495
rect 1318 -1508 1368 -1495
rect 1526 -1508 1576 -1495
rect 302 -1559 352 -1543
rect 520 -1559 570 -1543
rect 728 -1559 778 -1543
rect 1100 -1636 1150 -1608
rect 1100 -1656 1113 -1636
rect 1133 -1656 1150 -1636
rect 1100 -1685 1150 -1656
rect 1318 -1633 1368 -1608
rect 1318 -1653 1331 -1633
rect 1351 -1653 1368 -1633
rect 1318 -1685 1368 -1653
rect 1526 -1635 1576 -1608
rect 1526 -1655 1549 -1635
rect 1569 -1655 1576 -1635
rect 1526 -1685 1576 -1655
rect 303 -1736 353 -1723
rect 521 -1736 571 -1723
rect 729 -1736 779 -1723
rect 1100 -1743 1150 -1727
rect 1318 -1743 1368 -1727
rect 1526 -1743 1576 -1727
rect 303 -1864 353 -1836
rect 303 -1884 316 -1864
rect 336 -1884 353 -1864
rect 303 -1913 353 -1884
rect 521 -1861 571 -1836
rect 521 -1881 534 -1861
rect 554 -1881 571 -1861
rect 521 -1913 571 -1881
rect 729 -1863 779 -1836
rect 729 -1883 752 -1863
rect 772 -1883 779 -1863
rect 729 -1913 779 -1883
rect 303 -1971 353 -1955
rect 521 -1971 571 -1955
rect 729 -1971 779 -1955
rect 1245 -2118 1295 -2105
rect 1463 -2118 1513 -2105
rect 1671 -2118 1721 -2105
rect 1245 -2246 1295 -2218
rect 1245 -2266 1258 -2246
rect 1278 -2266 1295 -2246
rect 1245 -2295 1295 -2266
rect 1463 -2243 1513 -2218
rect 1463 -2263 1476 -2243
rect 1496 -2263 1513 -2243
rect 1463 -2295 1513 -2263
rect 1671 -2245 1721 -2218
rect 1671 -2265 1694 -2245
rect 1714 -2265 1721 -2245
rect 1671 -2295 1721 -2265
rect 282 -2342 332 -2329
rect 500 -2342 550 -2329
rect 708 -2342 758 -2329
rect 1245 -2353 1295 -2337
rect 1463 -2353 1513 -2337
rect 1671 -2353 1721 -2337
rect 282 -2470 332 -2442
rect 282 -2490 295 -2470
rect 315 -2490 332 -2470
rect 282 -2519 332 -2490
rect 500 -2467 550 -2442
rect 500 -2487 513 -2467
rect 533 -2487 550 -2467
rect 500 -2519 550 -2487
rect 708 -2469 758 -2442
rect 708 -2489 731 -2469
rect 751 -2489 758 -2469
rect 708 -2519 758 -2489
rect 1080 -2526 1130 -2513
rect 1298 -2526 1348 -2513
rect 1506 -2526 1556 -2513
rect 282 -2577 332 -2561
rect 500 -2577 550 -2561
rect 708 -2577 758 -2561
rect 1080 -2654 1130 -2626
rect 1080 -2674 1093 -2654
rect 1113 -2674 1130 -2654
rect 1080 -2703 1130 -2674
rect 1298 -2651 1348 -2626
rect 1298 -2671 1311 -2651
rect 1331 -2671 1348 -2651
rect 1298 -2703 1348 -2671
rect 1506 -2653 1556 -2626
rect 1506 -2673 1529 -2653
rect 1549 -2673 1556 -2653
rect 1506 -2703 1556 -2673
rect 283 -2754 333 -2741
rect 501 -2754 551 -2741
rect 709 -2754 759 -2741
rect 1080 -2761 1130 -2745
rect 1298 -2761 1348 -2745
rect 1506 -2761 1556 -2745
rect 283 -2882 333 -2854
rect 283 -2902 296 -2882
rect 316 -2902 333 -2882
rect 283 -2931 333 -2902
rect 501 -2879 551 -2854
rect 501 -2899 514 -2879
rect 534 -2899 551 -2879
rect 501 -2931 551 -2899
rect 709 -2881 759 -2854
rect 709 -2901 732 -2881
rect 752 -2901 759 -2881
rect 709 -2931 759 -2901
rect 283 -2989 333 -2973
rect 501 -2989 551 -2973
rect 709 -2989 759 -2973
rect 1162 -3134 1212 -3121
rect 1380 -3134 1430 -3121
rect 1588 -3134 1638 -3121
rect 1162 -3262 1212 -3234
rect 1162 -3282 1175 -3262
rect 1195 -3282 1212 -3262
rect 1162 -3311 1212 -3282
rect 1380 -3259 1430 -3234
rect 1380 -3279 1393 -3259
rect 1413 -3279 1430 -3259
rect 1380 -3311 1430 -3279
rect 1588 -3261 1638 -3234
rect 1588 -3281 1611 -3261
rect 1631 -3281 1638 -3261
rect 1588 -3311 1638 -3281
rect 265 -3360 315 -3347
rect 483 -3360 533 -3347
rect 691 -3360 741 -3347
rect 1162 -3369 1212 -3353
rect 1380 -3369 1430 -3353
rect 1588 -3369 1638 -3353
rect 265 -3488 315 -3460
rect 265 -3508 278 -3488
rect 298 -3508 315 -3488
rect 265 -3537 315 -3508
rect 483 -3485 533 -3460
rect 483 -3505 496 -3485
rect 516 -3505 533 -3485
rect 483 -3537 533 -3505
rect 691 -3487 741 -3460
rect 691 -3507 714 -3487
rect 734 -3507 741 -3487
rect 691 -3537 741 -3507
rect 1063 -3544 1113 -3531
rect 1281 -3544 1331 -3531
rect 1489 -3544 1539 -3531
rect 265 -3595 315 -3579
rect 483 -3595 533 -3579
rect 691 -3595 741 -3579
rect 1063 -3672 1113 -3644
rect 1063 -3692 1076 -3672
rect 1096 -3692 1113 -3672
rect 1063 -3721 1113 -3692
rect 1281 -3669 1331 -3644
rect 1281 -3689 1294 -3669
rect 1314 -3689 1331 -3669
rect 1281 -3721 1331 -3689
rect 1489 -3671 1539 -3644
rect 1489 -3691 1512 -3671
rect 1532 -3691 1539 -3671
rect 1489 -3721 1539 -3691
rect 266 -3772 316 -3759
rect 484 -3772 534 -3759
rect 692 -3772 742 -3759
rect 1063 -3779 1113 -3763
rect 1281 -3779 1331 -3763
rect 1489 -3779 1539 -3763
rect 266 -3900 316 -3872
rect 266 -3920 279 -3900
rect 299 -3920 316 -3900
rect 266 -3949 316 -3920
rect 484 -3897 534 -3872
rect 484 -3917 497 -3897
rect 517 -3917 534 -3897
rect 484 -3949 534 -3917
rect 692 -3899 742 -3872
rect 692 -3919 715 -3899
rect 735 -3919 742 -3899
rect 692 -3949 742 -3919
rect 266 -4007 316 -3991
rect 484 -4007 534 -3991
rect 692 -4007 742 -3991
<< polycont >>
rect 405 3618 425 3638
rect 623 3621 643 3641
rect 841 3619 861 3639
rect 1203 3434 1223 3454
rect 1421 3437 1441 3457
rect 1639 3435 1659 3455
rect 406 3206 426 3226
rect 624 3209 644 3229
rect 842 3207 862 3227
rect 1285 2826 1305 2846
rect 1503 2829 1523 2849
rect 1721 2827 1741 2847
rect 388 2600 408 2620
rect 606 2603 626 2623
rect 824 2601 844 2621
rect 1186 2416 1206 2436
rect 1404 2419 1424 2439
rect 1622 2417 1642 2437
rect 389 2188 409 2208
rect 607 2191 627 2211
rect 825 2189 845 2209
rect 1331 1806 1351 1826
rect 1549 1809 1569 1829
rect 1767 1807 1787 1827
rect 368 1582 388 1602
rect 586 1585 606 1605
rect 804 1583 824 1603
rect 1166 1398 1186 1418
rect 1384 1401 1404 1421
rect 1602 1399 1622 1419
rect 369 1170 389 1190
rect 587 1173 607 1193
rect 805 1171 825 1191
rect 1248 790 1268 810
rect 1466 793 1486 813
rect 1684 791 1704 811
rect 351 564 371 584
rect 569 567 589 587
rect 787 565 807 585
rect 1149 380 1169 400
rect 1367 383 1387 403
rect 1585 381 1605 401
rect 352 152 372 172
rect 570 155 590 175
rect 788 153 808 173
rect 1434 -232 1454 -212
rect 1652 -229 1672 -209
rect 1870 -231 1890 -211
rect 332 -454 352 -434
rect 550 -451 570 -431
rect 768 -453 788 -433
rect 1130 -638 1150 -618
rect 1348 -635 1368 -615
rect 1566 -637 1586 -617
rect 333 -866 353 -846
rect 551 -863 571 -843
rect 769 -865 789 -845
rect 1212 -1246 1232 -1226
rect 1430 -1243 1450 -1223
rect 1648 -1245 1668 -1225
rect 315 -1472 335 -1452
rect 533 -1469 553 -1449
rect 751 -1471 771 -1451
rect 1113 -1656 1133 -1636
rect 1331 -1653 1351 -1633
rect 1549 -1655 1569 -1635
rect 316 -1884 336 -1864
rect 534 -1881 554 -1861
rect 752 -1883 772 -1863
rect 1258 -2266 1278 -2246
rect 1476 -2263 1496 -2243
rect 1694 -2265 1714 -2245
rect 295 -2490 315 -2470
rect 513 -2487 533 -2467
rect 731 -2489 751 -2469
rect 1093 -2674 1113 -2654
rect 1311 -2671 1331 -2651
rect 1529 -2673 1549 -2653
rect 296 -2902 316 -2882
rect 514 -2899 534 -2879
rect 732 -2901 752 -2881
rect 1175 -3282 1195 -3262
rect 1393 -3279 1413 -3259
rect 1611 -3281 1631 -3261
rect 278 -3508 298 -3488
rect 496 -3505 516 -3485
rect 714 -3507 734 -3487
rect 1076 -3692 1096 -3672
rect 1294 -3689 1314 -3669
rect 1512 -3691 1532 -3671
rect 279 -3920 299 -3900
rect 497 -3917 517 -3897
rect 715 -3919 735 -3899
<< ndiffres >>
rect 167 3988 228 4004
rect 72 3984 228 3988
rect 72 3966 190 3984
rect 208 3966 228 3984
rect 72 3945 228 3966
rect 72 3944 172 3945
rect 73 3908 115 3944
rect 73 3885 224 3908
rect 73 3870 188 3885
rect 167 3867 188 3870
rect 206 3867 224 3885
rect 167 3848 224 3867
rect 162 3664 223 3680
rect 67 3660 223 3664
rect 67 3642 185 3660
rect 203 3642 223 3660
rect 67 3621 223 3642
rect 67 3620 167 3621
rect 68 3584 110 3620
rect 68 3561 219 3584
rect 68 3546 183 3561
rect 162 3543 183 3546
rect 201 3543 219 3561
rect 162 3524 219 3543
rect 156 3481 217 3497
rect 61 3477 217 3481
rect 61 3459 179 3477
rect 197 3459 217 3477
rect 61 3438 217 3459
rect 61 3437 161 3438
rect 62 3401 104 3437
rect 62 3378 213 3401
rect 62 3363 177 3378
rect 156 3360 177 3363
rect 195 3360 213 3378
rect 156 3341 213 3360
rect 149 3263 210 3279
rect 54 3259 210 3263
rect 54 3241 172 3259
rect 190 3241 210 3259
rect 54 3220 210 3241
rect 54 3219 154 3220
rect 55 3183 97 3219
rect 55 3160 206 3183
rect 55 3145 170 3160
rect 149 3142 170 3145
rect 188 3142 206 3160
rect 149 3123 206 3142
rect 150 2970 211 2986
rect 55 2966 211 2970
rect 55 2948 173 2966
rect 191 2948 211 2966
rect 55 2927 211 2948
rect 55 2926 155 2927
rect 56 2890 98 2926
rect 56 2867 207 2890
rect 56 2852 171 2867
rect 150 2849 171 2852
rect 189 2849 207 2867
rect 150 2830 207 2849
rect 145 2646 206 2662
rect 50 2642 206 2646
rect 50 2624 168 2642
rect 186 2624 206 2642
rect 50 2603 206 2624
rect 50 2602 150 2603
rect 51 2566 93 2602
rect 51 2543 202 2566
rect 51 2528 166 2543
rect 145 2525 166 2528
rect 184 2525 202 2543
rect 145 2506 202 2525
rect 139 2463 200 2479
rect 44 2459 200 2463
rect 44 2441 162 2459
rect 180 2441 200 2459
rect 44 2420 200 2441
rect 44 2419 144 2420
rect 45 2383 87 2419
rect 45 2360 196 2383
rect 45 2345 160 2360
rect 139 2342 160 2345
rect 178 2342 196 2360
rect 139 2323 196 2342
rect 132 2245 193 2261
rect 37 2241 193 2245
rect 37 2223 155 2241
rect 173 2223 193 2241
rect 37 2202 193 2223
rect 37 2201 137 2202
rect 38 2165 80 2201
rect 38 2142 189 2165
rect 38 2127 153 2142
rect 132 2124 153 2127
rect 171 2124 189 2142
rect 132 2105 189 2124
rect 130 1952 191 1968
rect 35 1948 191 1952
rect 35 1930 153 1948
rect 171 1930 191 1948
rect 35 1909 191 1930
rect 35 1908 135 1909
rect 36 1872 78 1908
rect 36 1849 187 1872
rect 36 1834 151 1849
rect 130 1831 151 1834
rect 169 1831 187 1849
rect 130 1812 187 1831
rect 125 1628 186 1644
rect 30 1624 186 1628
rect 30 1606 148 1624
rect 166 1606 186 1624
rect 30 1585 186 1606
rect 30 1584 130 1585
rect 31 1548 73 1584
rect 31 1525 182 1548
rect 31 1510 146 1525
rect 125 1507 146 1510
rect 164 1507 182 1525
rect 125 1488 182 1507
rect 119 1445 180 1461
rect 24 1441 180 1445
rect 24 1423 142 1441
rect 160 1423 180 1441
rect 24 1402 180 1423
rect 24 1401 124 1402
rect 25 1365 67 1401
rect 25 1342 176 1365
rect 25 1327 140 1342
rect 119 1324 140 1327
rect 158 1324 176 1342
rect 119 1305 176 1324
rect 112 1227 173 1243
rect 17 1223 173 1227
rect 17 1205 135 1223
rect 153 1205 173 1223
rect 17 1184 173 1205
rect 17 1183 117 1184
rect 18 1147 60 1183
rect 18 1124 169 1147
rect 18 1109 133 1124
rect 112 1106 133 1109
rect 151 1106 169 1124
rect 112 1087 169 1106
rect 113 934 174 950
rect 18 930 174 934
rect 18 912 136 930
rect 154 912 174 930
rect 18 891 174 912
rect 18 890 118 891
rect 19 854 61 890
rect 19 831 170 854
rect 19 816 134 831
rect 113 813 134 816
rect 152 813 170 831
rect 113 794 170 813
rect 108 610 169 626
rect 13 606 169 610
rect 13 588 131 606
rect 149 588 169 606
rect 13 567 169 588
rect 13 566 113 567
rect 14 530 56 566
rect 14 507 165 530
rect 14 492 129 507
rect 108 489 129 492
rect 147 489 165 507
rect 108 470 165 489
rect 102 427 163 443
rect 7 423 163 427
rect 7 405 125 423
rect 143 405 163 423
rect 7 384 163 405
rect 7 383 107 384
rect 8 347 50 383
rect 8 324 159 347
rect 8 309 123 324
rect 102 306 123 309
rect 141 306 159 324
rect 102 287 159 306
rect 95 209 156 225
rect 0 205 156 209
rect 0 187 118 205
rect 136 187 156 205
rect 0 166 156 187
rect 0 165 100 166
rect 1 129 43 165
rect 1 106 152 129
rect 1 91 116 106
rect 95 88 116 91
rect 134 88 152 106
rect 95 69 152 88
rect 94 -84 155 -68
rect -1 -88 155 -84
rect -1 -106 117 -88
rect 135 -106 155 -88
rect -1 -127 155 -106
rect -1 -128 99 -127
rect 0 -164 42 -128
rect 0 -187 151 -164
rect 0 -202 115 -187
rect 94 -205 115 -202
rect 133 -205 151 -187
rect 94 -224 151 -205
rect 89 -408 150 -392
rect -6 -412 150 -408
rect -6 -430 112 -412
rect 130 -430 150 -412
rect -6 -451 150 -430
rect -6 -452 94 -451
rect -5 -488 37 -452
rect -5 -511 146 -488
rect -5 -526 110 -511
rect 89 -529 110 -526
rect 128 -529 146 -511
rect 89 -548 146 -529
rect 83 -591 144 -575
rect -12 -595 144 -591
rect -12 -613 106 -595
rect 124 -613 144 -595
rect -12 -634 144 -613
rect -12 -635 88 -634
rect -11 -671 31 -635
rect -11 -694 140 -671
rect -11 -709 104 -694
rect 83 -712 104 -709
rect 122 -712 140 -694
rect 83 -731 140 -712
rect 76 -809 137 -793
rect -19 -813 137 -809
rect -19 -831 99 -813
rect 117 -831 137 -813
rect -19 -852 137 -831
rect -19 -853 81 -852
rect -18 -889 24 -853
rect -18 -912 133 -889
rect -18 -927 97 -912
rect 76 -930 97 -927
rect 115 -930 133 -912
rect 76 -949 133 -930
rect 77 -1102 138 -1086
rect -18 -1106 138 -1102
rect -18 -1124 100 -1106
rect 118 -1124 138 -1106
rect -18 -1145 138 -1124
rect -18 -1146 82 -1145
rect -17 -1182 25 -1146
rect -17 -1205 134 -1182
rect -17 -1220 98 -1205
rect 77 -1223 98 -1220
rect 116 -1223 134 -1205
rect 77 -1242 134 -1223
rect 72 -1426 133 -1410
rect -23 -1430 133 -1426
rect -23 -1448 95 -1430
rect 113 -1448 133 -1430
rect -23 -1469 133 -1448
rect -23 -1470 77 -1469
rect -22 -1506 20 -1470
rect -22 -1529 129 -1506
rect -22 -1544 93 -1529
rect 72 -1547 93 -1544
rect 111 -1547 129 -1529
rect 72 -1566 129 -1547
rect 66 -1609 127 -1593
rect -29 -1613 127 -1609
rect -29 -1631 89 -1613
rect 107 -1631 127 -1613
rect -29 -1652 127 -1631
rect -29 -1653 71 -1652
rect -28 -1689 14 -1653
rect -28 -1712 123 -1689
rect -28 -1727 87 -1712
rect 66 -1730 87 -1727
rect 105 -1730 123 -1712
rect 66 -1749 123 -1730
rect 59 -1827 120 -1811
rect -36 -1831 120 -1827
rect -36 -1849 82 -1831
rect 100 -1849 120 -1831
rect -36 -1870 120 -1849
rect -36 -1871 64 -1870
rect -35 -1907 7 -1871
rect -35 -1930 116 -1907
rect -35 -1945 80 -1930
rect 59 -1948 80 -1945
rect 98 -1948 116 -1930
rect 59 -1967 116 -1948
rect 57 -2120 118 -2104
rect -38 -2124 118 -2120
rect -38 -2142 80 -2124
rect 98 -2142 118 -2124
rect -38 -2163 118 -2142
rect -38 -2164 62 -2163
rect -37 -2200 5 -2164
rect -37 -2223 114 -2200
rect -37 -2238 78 -2223
rect 57 -2241 78 -2238
rect 96 -2241 114 -2223
rect 57 -2260 114 -2241
rect 52 -2444 113 -2428
rect -43 -2448 113 -2444
rect -43 -2466 75 -2448
rect 93 -2466 113 -2448
rect -43 -2487 113 -2466
rect -43 -2488 57 -2487
rect -42 -2524 0 -2488
rect -42 -2547 109 -2524
rect -42 -2562 73 -2547
rect 52 -2565 73 -2562
rect 91 -2565 109 -2547
rect 52 -2584 109 -2565
rect 46 -2627 107 -2611
rect -49 -2631 107 -2627
rect -49 -2649 69 -2631
rect 87 -2649 107 -2631
rect -49 -2670 107 -2649
rect -49 -2671 51 -2670
rect -48 -2707 -6 -2671
rect -48 -2730 103 -2707
rect -48 -2745 67 -2730
rect 46 -2748 67 -2745
rect 85 -2748 103 -2730
rect 46 -2767 103 -2748
rect 39 -2845 100 -2829
rect -56 -2849 100 -2845
rect -56 -2867 62 -2849
rect 80 -2867 100 -2849
rect -56 -2888 100 -2867
rect -56 -2889 44 -2888
rect -55 -2925 -13 -2889
rect -55 -2948 96 -2925
rect -55 -2963 60 -2948
rect 39 -2966 60 -2963
rect 78 -2966 96 -2948
rect 39 -2985 96 -2966
rect 40 -3138 101 -3122
rect -55 -3142 101 -3138
rect -55 -3160 63 -3142
rect 81 -3160 101 -3142
rect -55 -3181 101 -3160
rect -55 -3182 45 -3181
rect -54 -3218 -12 -3182
rect -54 -3241 97 -3218
rect -54 -3256 61 -3241
rect 40 -3259 61 -3256
rect 79 -3259 97 -3241
rect 40 -3278 97 -3259
rect 35 -3462 96 -3446
rect -60 -3466 96 -3462
rect -60 -3484 58 -3466
rect 76 -3484 96 -3466
rect -60 -3505 96 -3484
rect -60 -3506 40 -3505
rect -59 -3542 -17 -3506
rect -59 -3565 92 -3542
rect -59 -3580 56 -3565
rect 35 -3583 56 -3580
rect 74 -3583 92 -3565
rect 35 -3602 92 -3583
rect 29 -3645 90 -3629
rect -66 -3649 90 -3645
rect -66 -3667 52 -3649
rect 70 -3667 90 -3649
rect -66 -3688 90 -3667
rect -66 -3689 34 -3688
rect -65 -3725 -23 -3689
rect -65 -3748 86 -3725
rect -65 -3763 50 -3748
rect 29 -3766 50 -3763
rect 68 -3766 86 -3748
rect 29 -3785 86 -3766
rect 22 -3863 83 -3847
rect -73 -3867 83 -3863
rect -73 -3885 45 -3867
rect 63 -3885 83 -3867
rect -73 -3906 83 -3885
rect -73 -3907 27 -3906
rect -72 -3943 -30 -3907
rect -72 -3966 79 -3943
rect -72 -3981 43 -3966
rect 22 -3984 43 -3981
rect 61 -3984 79 -3966
rect 22 -4003 79 -3984
<< locali >>
rect 180 3984 227 4100
rect 180 3966 190 3984
rect 208 3966 227 3984
rect 180 3962 227 3966
rect 181 3957 218 3962
rect 169 3895 221 3897
rect 167 3891 600 3895
rect 167 3885 606 3891
rect 167 3867 188 3885
rect 206 3867 606 3885
rect 167 3849 606 3867
rect 169 3660 221 3849
rect 567 3824 606 3849
rect 351 3799 538 3823
rect 567 3804 962 3824
rect 982 3804 985 3824
rect 567 3799 985 3804
rect 351 3728 388 3799
rect 567 3798 910 3799
rect 567 3795 606 3798
rect 872 3797 909 3798
rect 503 3738 534 3739
rect 351 3708 360 3728
rect 380 3708 388 3728
rect 351 3698 388 3708
rect 447 3728 534 3738
rect 447 3708 456 3728
rect 476 3708 534 3728
rect 447 3699 534 3708
rect 447 3698 484 3699
rect 169 3642 185 3660
rect 203 3642 221 3660
rect 503 3648 534 3699
rect 569 3728 606 3795
rect 721 3738 757 3739
rect 569 3708 578 3728
rect 598 3708 606 3728
rect 569 3698 606 3708
rect 665 3728 813 3738
rect 913 3735 1009 3737
rect 665 3708 674 3728
rect 694 3708 784 3728
rect 804 3708 813 3728
rect 665 3699 813 3708
rect 871 3728 1009 3735
rect 871 3708 880 3728
rect 900 3708 1009 3728
rect 871 3699 1009 3708
rect 665 3698 702 3699
rect 395 3645 436 3646
rect 169 3624 221 3642
rect 287 3638 436 3645
rect 287 3618 346 3638
rect 366 3618 405 3638
rect 425 3618 436 3638
rect 287 3610 436 3618
rect 503 3641 660 3648
rect 503 3621 623 3641
rect 643 3621 660 3641
rect 503 3611 660 3621
rect 503 3610 538 3611
rect 503 3589 534 3610
rect 721 3589 757 3699
rect 776 3698 813 3699
rect 872 3698 909 3699
rect 832 3639 922 3645
rect 832 3619 841 3639
rect 861 3637 922 3639
rect 861 3619 886 3637
rect 832 3617 886 3619
rect 906 3617 922 3637
rect 832 3611 922 3617
rect 346 3588 383 3589
rect 345 3579 383 3588
rect 173 3561 213 3571
rect 173 3543 183 3561
rect 201 3543 213 3561
rect 345 3559 354 3579
rect 374 3559 383 3579
rect 345 3551 383 3559
rect 449 3583 534 3589
rect 564 3588 601 3589
rect 449 3563 457 3583
rect 477 3563 534 3583
rect 449 3555 534 3563
rect 563 3579 601 3588
rect 563 3559 572 3579
rect 592 3559 601 3579
rect 449 3554 485 3555
rect 563 3551 601 3559
rect 667 3583 811 3589
rect 667 3563 675 3583
rect 695 3563 728 3583
rect 748 3563 783 3583
rect 803 3563 811 3583
rect 667 3555 811 3563
rect 667 3554 703 3555
rect 775 3554 811 3555
rect 877 3588 914 3589
rect 877 3587 915 3588
rect 877 3579 941 3587
rect 877 3559 886 3579
rect 906 3565 941 3579
rect 961 3565 964 3585
rect 906 3560 964 3565
rect 906 3559 941 3560
rect 173 3487 213 3543
rect 346 3522 383 3551
rect 347 3520 383 3522
rect 347 3498 538 3520
rect 564 3519 601 3551
rect 877 3547 941 3559
rect 981 3521 1008 3699
rect 840 3519 1008 3521
rect 564 3509 1008 3519
rect 1149 3615 1336 3639
rect 1367 3620 1760 3640
rect 1780 3620 1783 3640
rect 1367 3615 1783 3620
rect 1149 3544 1186 3615
rect 1367 3614 1708 3615
rect 1301 3554 1332 3555
rect 1149 3524 1158 3544
rect 1178 3524 1186 3544
rect 1149 3514 1186 3524
rect 1245 3544 1332 3554
rect 1245 3524 1254 3544
rect 1274 3524 1332 3544
rect 1245 3515 1332 3524
rect 1245 3514 1282 3515
rect 170 3482 213 3487
rect 561 3493 1008 3509
rect 561 3487 589 3493
rect 840 3492 1008 3493
rect 170 3479 320 3482
rect 561 3479 588 3487
rect 170 3477 588 3479
rect 170 3459 179 3477
rect 197 3459 588 3477
rect 1301 3464 1332 3515
rect 1367 3544 1404 3614
rect 1670 3613 1707 3614
rect 1519 3554 1555 3555
rect 1367 3524 1376 3544
rect 1396 3524 1404 3544
rect 1367 3514 1404 3524
rect 1463 3544 1611 3554
rect 1711 3551 1807 3553
rect 1463 3524 1472 3544
rect 1492 3524 1582 3544
rect 1602 3524 1611 3544
rect 1463 3515 1611 3524
rect 1669 3544 1807 3551
rect 1669 3524 1678 3544
rect 1698 3524 1807 3544
rect 1669 3515 1807 3524
rect 1463 3514 1500 3515
rect 1193 3461 1234 3462
rect 170 3456 588 3459
rect 170 3450 213 3456
rect 173 3447 213 3450
rect 1085 3454 1234 3461
rect 570 3438 610 3439
rect 281 3421 610 3438
rect 1085 3434 1144 3454
rect 1164 3434 1203 3454
rect 1223 3434 1234 3454
rect 1085 3426 1234 3434
rect 1301 3457 1458 3464
rect 1301 3437 1421 3457
rect 1441 3437 1458 3457
rect 1301 3427 1458 3437
rect 1301 3426 1336 3427
rect 165 3378 208 3389
rect 165 3360 177 3378
rect 195 3360 208 3378
rect 165 3334 208 3360
rect 281 3334 308 3421
rect 570 3412 610 3421
rect 165 3313 308 3334
rect 352 3386 386 3402
rect 570 3392 963 3412
rect 983 3392 986 3412
rect 1301 3405 1332 3426
rect 1519 3405 1555 3515
rect 1574 3514 1611 3515
rect 1670 3514 1707 3515
rect 1630 3455 1720 3461
rect 1630 3435 1639 3455
rect 1659 3453 1720 3455
rect 1659 3435 1684 3453
rect 1630 3433 1684 3435
rect 1704 3433 1720 3453
rect 1630 3427 1720 3433
rect 1144 3404 1181 3405
rect 570 3387 986 3392
rect 1143 3395 1181 3404
rect 570 3386 911 3387
rect 352 3316 389 3386
rect 504 3326 535 3327
rect 165 3311 302 3313
rect 165 3269 208 3311
rect 352 3296 361 3316
rect 381 3296 389 3316
rect 352 3286 389 3296
rect 448 3316 535 3326
rect 448 3296 457 3316
rect 477 3296 535 3316
rect 448 3287 535 3296
rect 448 3286 485 3287
rect 163 3259 208 3269
rect 163 3241 172 3259
rect 190 3241 208 3259
rect 163 3235 208 3241
rect 504 3236 535 3287
rect 570 3316 607 3386
rect 873 3385 910 3386
rect 1143 3375 1152 3395
rect 1172 3375 1181 3395
rect 1143 3367 1181 3375
rect 1247 3399 1332 3405
rect 1362 3404 1399 3405
rect 1247 3379 1255 3399
rect 1275 3379 1332 3399
rect 1247 3371 1332 3379
rect 1361 3395 1399 3404
rect 1361 3375 1370 3395
rect 1390 3375 1399 3395
rect 1247 3370 1283 3371
rect 1361 3367 1399 3375
rect 1465 3399 1609 3405
rect 1465 3379 1473 3399
rect 1493 3380 1525 3399
rect 1546 3380 1581 3399
rect 1493 3379 1581 3380
rect 1601 3379 1609 3399
rect 1465 3371 1609 3379
rect 1465 3370 1501 3371
rect 1573 3370 1609 3371
rect 1675 3404 1712 3405
rect 1675 3403 1713 3404
rect 1675 3395 1739 3403
rect 1675 3375 1684 3395
rect 1704 3381 1739 3395
rect 1759 3381 1762 3401
rect 1704 3376 1762 3381
rect 1704 3375 1739 3376
rect 1144 3338 1181 3367
rect 1145 3336 1181 3338
rect 722 3326 758 3327
rect 570 3296 579 3316
rect 599 3296 607 3316
rect 570 3286 607 3296
rect 666 3316 814 3326
rect 914 3323 1010 3325
rect 666 3296 675 3316
rect 695 3296 785 3316
rect 805 3296 814 3316
rect 666 3287 814 3296
rect 872 3316 1010 3323
rect 872 3296 881 3316
rect 901 3296 1010 3316
rect 1145 3314 1336 3336
rect 1362 3335 1399 3367
rect 1675 3363 1739 3375
rect 1779 3337 1806 3515
rect 1638 3335 1806 3337
rect 1362 3309 1806 3335
rect 872 3287 1010 3296
rect 666 3286 703 3287
rect 163 3232 200 3235
rect 396 3233 437 3234
rect 288 3226 437 3233
rect 288 3206 347 3226
rect 367 3206 406 3226
rect 426 3206 437 3226
rect 288 3198 437 3206
rect 504 3229 661 3236
rect 504 3209 624 3229
rect 644 3209 661 3229
rect 504 3199 661 3209
rect 504 3198 539 3199
rect 504 3177 535 3198
rect 722 3177 758 3287
rect 777 3286 814 3287
rect 873 3286 910 3287
rect 833 3227 923 3233
rect 833 3207 842 3227
rect 862 3225 923 3227
rect 862 3207 887 3225
rect 833 3205 887 3207
rect 907 3205 923 3225
rect 833 3199 923 3205
rect 347 3176 384 3177
rect 160 3168 197 3170
rect 160 3160 202 3168
rect 160 3142 170 3160
rect 188 3142 202 3160
rect 160 3133 202 3142
rect 346 3167 384 3176
rect 346 3147 355 3167
rect 375 3147 384 3167
rect 346 3139 384 3147
rect 450 3171 535 3177
rect 565 3176 602 3177
rect 450 3151 458 3171
rect 478 3151 535 3171
rect 450 3143 535 3151
rect 564 3167 602 3176
rect 564 3147 573 3167
rect 593 3147 602 3167
rect 450 3142 486 3143
rect 564 3139 602 3147
rect 668 3175 812 3177
rect 668 3171 720 3175
rect 668 3151 676 3171
rect 696 3155 720 3171
rect 740 3171 812 3175
rect 740 3155 784 3171
rect 696 3151 784 3155
rect 804 3151 812 3171
rect 668 3143 812 3151
rect 668 3142 704 3143
rect 776 3142 812 3143
rect 878 3176 915 3177
rect 878 3175 916 3176
rect 878 3167 942 3175
rect 878 3147 887 3167
rect 907 3153 942 3167
rect 962 3153 965 3173
rect 907 3148 965 3153
rect 907 3147 942 3148
rect 161 3108 202 3133
rect 347 3108 384 3139
rect 565 3108 602 3139
rect 878 3135 942 3147
rect 982 3109 1009 3287
rect 161 3081 210 3108
rect 346 3082 395 3108
rect 564 3107 645 3108
rect 841 3107 1009 3109
rect 564 3082 1009 3107
rect 565 3081 1009 3082
rect 163 3048 210 3081
rect 566 3048 606 3081
rect 841 3080 1009 3081
rect 1472 3085 1512 3309
rect 1638 3308 1806 3309
rect 1472 3063 1480 3085
rect 1504 3063 1512 3085
rect 1472 3055 1512 3063
rect 163 3009 606 3048
rect 163 2966 210 3009
rect 566 3004 606 3009
rect 1231 3007 1418 3031
rect 1449 3012 1842 3032
rect 1862 3012 1865 3032
rect 1449 3007 1865 3012
rect 163 2948 173 2966
rect 191 2948 210 2966
rect 163 2944 210 2948
rect 164 2939 201 2944
rect 1231 2936 1268 3007
rect 1449 3006 1790 3007
rect 1383 2946 1414 2947
rect 1231 2916 1240 2936
rect 1260 2916 1268 2936
rect 1231 2906 1268 2916
rect 1327 2936 1414 2946
rect 1327 2916 1336 2936
rect 1356 2916 1414 2936
rect 1327 2907 1414 2916
rect 1327 2906 1364 2907
rect 152 2877 204 2879
rect 150 2873 583 2877
rect 150 2867 589 2873
rect 150 2849 171 2867
rect 189 2849 589 2867
rect 1383 2856 1414 2907
rect 1449 2936 1486 3006
rect 1752 3005 1789 3006
rect 1601 2946 1637 2947
rect 1449 2916 1458 2936
rect 1478 2916 1486 2936
rect 1449 2906 1486 2916
rect 1545 2936 1693 2946
rect 1793 2943 1889 2945
rect 1545 2916 1554 2936
rect 1574 2916 1664 2936
rect 1684 2916 1693 2936
rect 1545 2907 1693 2916
rect 1751 2936 1889 2943
rect 1751 2916 1760 2936
rect 1780 2916 1889 2936
rect 1751 2907 1889 2916
rect 1545 2906 1582 2907
rect 1275 2853 1316 2854
rect 150 2831 589 2849
rect 152 2642 204 2831
rect 550 2806 589 2831
rect 1167 2846 1316 2853
rect 1167 2826 1226 2846
rect 1246 2826 1285 2846
rect 1305 2826 1316 2846
rect 1167 2818 1316 2826
rect 1383 2849 1540 2856
rect 1383 2829 1503 2849
rect 1523 2829 1540 2849
rect 1383 2819 1540 2829
rect 1383 2818 1418 2819
rect 334 2781 521 2805
rect 550 2786 945 2806
rect 965 2786 968 2806
rect 1383 2797 1414 2818
rect 1601 2797 1637 2907
rect 1656 2906 1693 2907
rect 1752 2906 1789 2907
rect 1712 2847 1802 2853
rect 1712 2827 1721 2847
rect 1741 2845 1802 2847
rect 1741 2827 1766 2845
rect 1712 2825 1766 2827
rect 1786 2825 1802 2845
rect 1712 2819 1802 2825
rect 1226 2796 1263 2797
rect 550 2781 968 2786
rect 1225 2787 1263 2796
rect 334 2710 371 2781
rect 550 2780 893 2781
rect 550 2777 589 2780
rect 855 2779 892 2780
rect 486 2720 517 2721
rect 334 2690 343 2710
rect 363 2690 371 2710
rect 334 2680 371 2690
rect 430 2710 517 2720
rect 430 2690 439 2710
rect 459 2690 517 2710
rect 430 2681 517 2690
rect 430 2680 467 2681
rect 152 2624 168 2642
rect 186 2624 204 2642
rect 486 2630 517 2681
rect 552 2710 589 2777
rect 1225 2767 1234 2787
rect 1254 2767 1263 2787
rect 1225 2759 1263 2767
rect 1329 2791 1414 2797
rect 1444 2796 1481 2797
rect 1329 2771 1337 2791
rect 1357 2771 1414 2791
rect 1329 2763 1414 2771
rect 1443 2787 1481 2796
rect 1443 2767 1452 2787
rect 1472 2767 1481 2787
rect 1329 2762 1365 2763
rect 1443 2759 1481 2767
rect 1547 2792 1691 2797
rect 1547 2791 1609 2792
rect 1547 2771 1555 2791
rect 1575 2773 1609 2791
rect 1630 2791 1691 2792
rect 1630 2773 1663 2791
rect 1575 2771 1663 2773
rect 1683 2771 1691 2791
rect 1547 2763 1691 2771
rect 1547 2762 1583 2763
rect 1655 2762 1691 2763
rect 1757 2796 1794 2797
rect 1757 2795 1795 2796
rect 1757 2787 1821 2795
rect 1757 2767 1766 2787
rect 1786 2773 1821 2787
rect 1841 2773 1844 2793
rect 1786 2768 1844 2773
rect 1786 2767 1821 2768
rect 1226 2730 1263 2759
rect 1227 2728 1263 2730
rect 704 2720 740 2721
rect 552 2690 561 2710
rect 581 2690 589 2710
rect 552 2680 589 2690
rect 648 2710 796 2720
rect 896 2717 992 2719
rect 648 2690 657 2710
rect 677 2690 767 2710
rect 787 2690 796 2710
rect 648 2681 796 2690
rect 854 2710 992 2717
rect 854 2690 863 2710
rect 883 2690 992 2710
rect 1227 2706 1418 2728
rect 1444 2727 1481 2759
rect 1757 2755 1821 2767
rect 1861 2729 1888 2907
rect 1720 2727 1888 2729
rect 1444 2713 1888 2727
rect 1444 2701 1891 2713
rect 1487 2699 1520 2701
rect 854 2681 992 2690
rect 648 2680 685 2681
rect 378 2627 419 2628
rect 152 2606 204 2624
rect 270 2620 419 2627
rect 270 2600 329 2620
rect 349 2600 388 2620
rect 408 2600 419 2620
rect 270 2592 419 2600
rect 486 2623 643 2630
rect 486 2603 606 2623
rect 626 2603 643 2623
rect 486 2593 643 2603
rect 486 2592 521 2593
rect 486 2571 517 2592
rect 704 2571 740 2681
rect 759 2680 796 2681
rect 855 2680 892 2681
rect 815 2621 905 2627
rect 815 2601 824 2621
rect 844 2619 905 2621
rect 844 2601 869 2619
rect 815 2599 869 2601
rect 889 2599 905 2619
rect 815 2593 905 2599
rect 329 2570 366 2571
rect 328 2561 366 2570
rect 156 2543 196 2553
rect 156 2525 166 2543
rect 184 2525 196 2543
rect 328 2541 337 2561
rect 357 2541 366 2561
rect 328 2533 366 2541
rect 432 2565 517 2571
rect 547 2570 584 2571
rect 432 2545 440 2565
rect 460 2545 517 2565
rect 432 2537 517 2545
rect 546 2561 584 2570
rect 546 2541 555 2561
rect 575 2541 584 2561
rect 432 2536 468 2537
rect 546 2533 584 2541
rect 650 2565 794 2571
rect 650 2545 658 2565
rect 678 2545 711 2565
rect 731 2545 766 2565
rect 786 2545 794 2565
rect 650 2537 794 2545
rect 650 2536 686 2537
rect 758 2536 794 2537
rect 860 2570 897 2571
rect 860 2569 898 2570
rect 860 2561 924 2569
rect 860 2541 869 2561
rect 889 2547 924 2561
rect 944 2547 947 2567
rect 889 2542 947 2547
rect 889 2541 924 2542
rect 156 2469 196 2525
rect 329 2504 366 2533
rect 330 2502 366 2504
rect 330 2480 521 2502
rect 547 2501 584 2533
rect 860 2529 924 2541
rect 964 2503 991 2681
rect 1849 2656 1891 2701
rect 823 2501 991 2503
rect 547 2491 991 2501
rect 1132 2597 1319 2621
rect 1350 2602 1743 2622
rect 1763 2602 1766 2622
rect 1350 2597 1766 2602
rect 1132 2526 1169 2597
rect 1350 2596 1691 2597
rect 1284 2536 1315 2537
rect 1132 2506 1141 2526
rect 1161 2506 1169 2526
rect 1132 2496 1169 2506
rect 1228 2526 1315 2536
rect 1228 2506 1237 2526
rect 1257 2506 1315 2526
rect 1228 2497 1315 2506
rect 1228 2496 1265 2497
rect 153 2464 196 2469
rect 544 2475 991 2491
rect 544 2469 572 2475
rect 823 2474 991 2475
rect 153 2461 303 2464
rect 544 2461 571 2469
rect 153 2459 571 2461
rect 153 2441 162 2459
rect 180 2441 571 2459
rect 1284 2446 1315 2497
rect 1350 2526 1387 2596
rect 1653 2595 1690 2596
rect 1502 2536 1538 2537
rect 1350 2506 1359 2526
rect 1379 2506 1387 2526
rect 1350 2496 1387 2506
rect 1446 2526 1594 2536
rect 1694 2533 1790 2535
rect 1446 2506 1455 2526
rect 1475 2506 1565 2526
rect 1585 2506 1594 2526
rect 1446 2497 1594 2506
rect 1652 2526 1790 2533
rect 1652 2506 1661 2526
rect 1681 2506 1790 2526
rect 1652 2497 1790 2506
rect 1446 2496 1483 2497
rect 1176 2443 1217 2444
rect 153 2438 571 2441
rect 153 2432 196 2438
rect 156 2429 196 2432
rect 1071 2436 1217 2443
rect 553 2420 593 2421
rect 264 2403 593 2420
rect 1071 2416 1127 2436
rect 1147 2416 1186 2436
rect 1206 2416 1217 2436
rect 1071 2408 1217 2416
rect 1284 2439 1441 2446
rect 1284 2419 1404 2439
rect 1424 2419 1441 2439
rect 1284 2409 1441 2419
rect 1284 2408 1319 2409
rect 148 2360 191 2371
rect 148 2342 160 2360
rect 178 2342 191 2360
rect 148 2316 191 2342
rect 264 2316 291 2403
rect 553 2394 593 2403
rect 148 2295 291 2316
rect 335 2368 369 2384
rect 553 2374 946 2394
rect 966 2374 969 2394
rect 1284 2387 1315 2408
rect 1502 2387 1538 2497
rect 1557 2496 1594 2497
rect 1653 2496 1690 2497
rect 1613 2437 1703 2443
rect 1613 2417 1622 2437
rect 1642 2435 1703 2437
rect 1642 2417 1667 2435
rect 1613 2415 1667 2417
rect 1687 2415 1703 2435
rect 1613 2409 1703 2415
rect 1127 2386 1164 2387
rect 553 2369 969 2374
rect 1126 2377 1164 2386
rect 553 2368 894 2369
rect 335 2298 372 2368
rect 487 2308 518 2309
rect 148 2293 285 2295
rect 148 2251 191 2293
rect 335 2278 344 2298
rect 364 2278 372 2298
rect 335 2268 372 2278
rect 431 2298 518 2308
rect 431 2278 440 2298
rect 460 2278 518 2298
rect 431 2269 518 2278
rect 431 2268 468 2269
rect 146 2241 191 2251
rect 146 2223 155 2241
rect 173 2223 191 2241
rect 146 2217 191 2223
rect 487 2218 518 2269
rect 553 2298 590 2368
rect 856 2367 893 2368
rect 1126 2357 1135 2377
rect 1155 2357 1164 2377
rect 1126 2349 1164 2357
rect 1230 2381 1315 2387
rect 1345 2386 1382 2387
rect 1230 2361 1238 2381
rect 1258 2361 1315 2381
rect 1230 2353 1315 2361
rect 1344 2377 1382 2386
rect 1344 2357 1353 2377
rect 1373 2357 1382 2377
rect 1230 2352 1266 2353
rect 1344 2349 1382 2357
rect 1448 2381 1592 2387
rect 1448 2361 1456 2381
rect 1476 2378 1564 2381
rect 1476 2361 1511 2378
rect 1448 2360 1511 2361
rect 1530 2361 1564 2378
rect 1584 2361 1592 2381
rect 1530 2360 1592 2361
rect 1448 2353 1592 2360
rect 1448 2352 1484 2353
rect 1556 2352 1592 2353
rect 1658 2386 1695 2387
rect 1658 2385 1696 2386
rect 1718 2385 1745 2389
rect 1658 2383 1745 2385
rect 1658 2377 1722 2383
rect 1658 2357 1667 2377
rect 1687 2363 1722 2377
rect 1742 2363 1745 2383
rect 1687 2358 1745 2363
rect 1687 2357 1722 2358
rect 1127 2320 1164 2349
rect 1128 2318 1164 2320
rect 705 2308 741 2309
rect 553 2278 562 2298
rect 582 2278 590 2298
rect 553 2268 590 2278
rect 649 2298 797 2308
rect 897 2305 993 2307
rect 649 2278 658 2298
rect 678 2278 768 2298
rect 788 2278 797 2298
rect 649 2269 797 2278
rect 855 2298 993 2305
rect 855 2278 864 2298
rect 884 2278 993 2298
rect 1128 2296 1319 2318
rect 1345 2317 1382 2349
rect 1658 2345 1722 2357
rect 1762 2319 1789 2497
rect 1621 2317 1789 2319
rect 1345 2291 1789 2317
rect 855 2269 993 2278
rect 649 2268 686 2269
rect 146 2214 183 2217
rect 379 2215 420 2216
rect 271 2208 420 2215
rect 271 2188 330 2208
rect 350 2188 389 2208
rect 409 2188 420 2208
rect 271 2180 420 2188
rect 487 2211 644 2218
rect 487 2191 607 2211
rect 627 2191 644 2211
rect 487 2181 644 2191
rect 487 2180 522 2181
rect 487 2159 518 2180
rect 705 2159 741 2269
rect 760 2268 797 2269
rect 856 2268 893 2269
rect 816 2209 906 2215
rect 816 2189 825 2209
rect 845 2207 906 2209
rect 845 2189 870 2207
rect 816 2187 870 2189
rect 890 2187 906 2207
rect 816 2181 906 2187
rect 330 2158 367 2159
rect 142 2150 180 2152
rect 142 2142 185 2150
rect 142 2124 153 2142
rect 171 2124 185 2142
rect 142 2097 185 2124
rect 329 2149 367 2158
rect 329 2129 338 2149
rect 358 2129 367 2149
rect 329 2121 367 2129
rect 433 2153 518 2159
rect 548 2158 585 2159
rect 433 2133 441 2153
rect 461 2133 518 2153
rect 433 2125 518 2133
rect 547 2149 585 2158
rect 547 2129 556 2149
rect 576 2129 585 2149
rect 433 2124 469 2125
rect 547 2121 585 2129
rect 651 2157 795 2159
rect 651 2153 703 2157
rect 651 2133 659 2153
rect 679 2137 703 2153
rect 723 2153 795 2157
rect 723 2137 767 2153
rect 679 2133 767 2137
rect 787 2133 795 2153
rect 651 2125 795 2133
rect 651 2124 687 2125
rect 759 2124 795 2125
rect 861 2158 898 2159
rect 861 2157 899 2158
rect 861 2149 925 2157
rect 861 2129 870 2149
rect 890 2135 925 2149
rect 945 2135 948 2155
rect 890 2130 948 2135
rect 890 2129 925 2130
rect 143 2090 185 2097
rect 330 2090 367 2121
rect 548 2090 585 2121
rect 861 2117 925 2129
rect 965 2091 992 2269
rect 143 2050 188 2090
rect 330 2065 475 2090
rect 548 2089 628 2090
rect 824 2089 992 2091
rect 548 2073 992 2089
rect 332 2064 475 2065
rect 547 2063 992 2073
rect 143 2029 190 2050
rect 547 2029 588 2063
rect 824 2062 992 2063
rect 1455 2067 1495 2291
rect 1621 2290 1789 2291
rect 1853 2323 1886 2656
rect 1853 2315 1890 2323
rect 1853 2296 1861 2315
rect 1882 2296 1890 2315
rect 1853 2290 1890 2296
rect 1455 2045 1463 2067
rect 1487 2045 1495 2067
rect 1455 2037 1495 2045
rect 143 1999 588 2029
rect 1626 2012 1691 2013
rect 143 1996 566 1999
rect 143 1948 190 1996
rect 143 1930 153 1948
rect 171 1930 190 1948
rect 143 1926 190 1930
rect 1277 1987 1464 2011
rect 1495 1992 1888 2012
rect 1908 1992 1911 2012
rect 1495 1987 1911 1992
rect 144 1921 181 1926
rect 1277 1916 1314 1987
rect 1495 1986 1836 1987
rect 1429 1926 1460 1927
rect 1277 1896 1286 1916
rect 1306 1896 1314 1916
rect 1277 1886 1314 1896
rect 1373 1916 1460 1926
rect 1373 1896 1382 1916
rect 1402 1896 1460 1916
rect 1373 1887 1460 1896
rect 1373 1886 1410 1887
rect 132 1859 184 1861
rect 130 1855 563 1859
rect 130 1849 569 1855
rect 130 1831 151 1849
rect 169 1831 569 1849
rect 1429 1836 1460 1887
rect 1495 1916 1532 1986
rect 1798 1985 1835 1986
rect 1647 1926 1683 1927
rect 1495 1896 1504 1916
rect 1524 1896 1532 1916
rect 1495 1886 1532 1896
rect 1591 1916 1739 1926
rect 1839 1923 1935 1925
rect 1591 1896 1600 1916
rect 1620 1896 1710 1916
rect 1730 1896 1739 1916
rect 1591 1887 1739 1896
rect 1797 1916 1935 1923
rect 1797 1896 1806 1916
rect 1826 1896 1935 1916
rect 1797 1887 1935 1896
rect 1591 1886 1628 1887
rect 1321 1833 1362 1834
rect 130 1813 569 1831
rect 132 1624 184 1813
rect 530 1788 569 1813
rect 1213 1826 1362 1833
rect 1213 1806 1272 1826
rect 1292 1806 1331 1826
rect 1351 1806 1362 1826
rect 1213 1798 1362 1806
rect 1429 1829 1586 1836
rect 1429 1809 1549 1829
rect 1569 1809 1586 1829
rect 1429 1799 1586 1809
rect 1429 1798 1464 1799
rect 314 1763 501 1787
rect 530 1768 925 1788
rect 945 1768 948 1788
rect 1429 1777 1460 1798
rect 1647 1777 1683 1887
rect 1702 1886 1739 1887
rect 1798 1886 1835 1887
rect 1758 1827 1848 1833
rect 1758 1807 1767 1827
rect 1787 1825 1848 1827
rect 1787 1807 1812 1825
rect 1758 1805 1812 1807
rect 1832 1805 1848 1825
rect 1758 1799 1848 1805
rect 1272 1776 1309 1777
rect 530 1763 948 1768
rect 1271 1767 1309 1776
rect 314 1692 351 1763
rect 530 1762 873 1763
rect 530 1759 569 1762
rect 835 1761 872 1762
rect 466 1702 497 1703
rect 314 1672 323 1692
rect 343 1672 351 1692
rect 314 1662 351 1672
rect 410 1692 497 1702
rect 410 1672 419 1692
rect 439 1672 497 1692
rect 410 1663 497 1672
rect 410 1662 447 1663
rect 132 1606 148 1624
rect 166 1606 184 1624
rect 466 1612 497 1663
rect 532 1692 569 1759
rect 1271 1747 1280 1767
rect 1300 1747 1309 1767
rect 1271 1739 1309 1747
rect 1375 1771 1460 1777
rect 1490 1776 1527 1777
rect 1375 1751 1383 1771
rect 1403 1751 1460 1771
rect 1375 1743 1460 1751
rect 1489 1767 1527 1776
rect 1489 1747 1498 1767
rect 1518 1747 1527 1767
rect 1375 1742 1411 1743
rect 1489 1739 1527 1747
rect 1593 1771 1737 1777
rect 1593 1751 1601 1771
rect 1621 1770 1709 1771
rect 1621 1752 1656 1770
rect 1674 1752 1709 1770
rect 1621 1751 1709 1752
rect 1729 1751 1737 1771
rect 1593 1743 1737 1751
rect 1593 1742 1629 1743
rect 1701 1742 1737 1743
rect 1803 1776 1840 1777
rect 1803 1775 1841 1776
rect 1803 1767 1867 1775
rect 1803 1747 1812 1767
rect 1832 1753 1867 1767
rect 1887 1753 1890 1773
rect 1832 1748 1890 1753
rect 1832 1747 1867 1748
rect 1272 1710 1309 1739
rect 1273 1708 1309 1710
rect 684 1702 720 1703
rect 532 1672 541 1692
rect 561 1672 569 1692
rect 532 1662 569 1672
rect 628 1692 776 1702
rect 876 1699 972 1701
rect 628 1672 637 1692
rect 657 1672 747 1692
rect 767 1672 776 1692
rect 628 1663 776 1672
rect 834 1692 972 1699
rect 834 1672 843 1692
rect 863 1672 972 1692
rect 1273 1686 1464 1708
rect 1490 1707 1527 1739
rect 1803 1735 1867 1747
rect 1907 1711 1934 1887
rect 1853 1709 1934 1711
rect 1766 1707 1934 1709
rect 1490 1681 1934 1707
rect 1600 1679 1640 1681
rect 1766 1680 1934 1681
rect 834 1663 972 1672
rect 1875 1678 1934 1680
rect 628 1662 665 1663
rect 358 1609 399 1610
rect 132 1588 184 1606
rect 250 1602 399 1609
rect 250 1582 309 1602
rect 329 1582 368 1602
rect 388 1582 399 1602
rect 250 1574 399 1582
rect 466 1605 623 1612
rect 466 1585 586 1605
rect 606 1585 623 1605
rect 466 1575 623 1585
rect 466 1574 501 1575
rect 466 1553 497 1574
rect 684 1553 720 1663
rect 739 1662 776 1663
rect 835 1662 872 1663
rect 795 1603 885 1609
rect 795 1583 804 1603
rect 824 1601 885 1603
rect 824 1583 849 1601
rect 795 1581 849 1583
rect 869 1581 885 1601
rect 795 1575 885 1581
rect 309 1552 346 1553
rect 308 1543 346 1552
rect 136 1525 176 1535
rect 136 1507 146 1525
rect 164 1507 176 1525
rect 308 1523 317 1543
rect 337 1523 346 1543
rect 308 1515 346 1523
rect 412 1547 497 1553
rect 527 1552 564 1553
rect 412 1527 420 1547
rect 440 1527 497 1547
rect 412 1519 497 1527
rect 526 1543 564 1552
rect 526 1523 535 1543
rect 555 1523 564 1543
rect 412 1518 448 1519
rect 526 1515 564 1523
rect 630 1547 774 1553
rect 630 1527 638 1547
rect 658 1527 691 1547
rect 711 1527 746 1547
rect 766 1527 774 1547
rect 630 1519 774 1527
rect 630 1518 666 1519
rect 738 1518 774 1519
rect 840 1552 877 1553
rect 840 1551 878 1552
rect 840 1543 904 1551
rect 840 1523 849 1543
rect 869 1529 904 1543
rect 924 1529 927 1549
rect 869 1524 927 1529
rect 869 1523 904 1524
rect 136 1451 176 1507
rect 309 1486 346 1515
rect 310 1484 346 1486
rect 310 1462 501 1484
rect 527 1483 564 1515
rect 840 1511 904 1523
rect 944 1485 971 1663
rect 1875 1660 1904 1678
rect 803 1483 971 1485
rect 527 1473 971 1483
rect 1112 1579 1299 1603
rect 1330 1584 1723 1604
rect 1743 1584 1746 1604
rect 1330 1579 1746 1584
rect 1112 1508 1149 1579
rect 1330 1578 1671 1579
rect 1264 1518 1295 1519
rect 1112 1488 1121 1508
rect 1141 1488 1149 1508
rect 1112 1478 1149 1488
rect 1208 1508 1295 1518
rect 1208 1488 1217 1508
rect 1237 1488 1295 1508
rect 1208 1479 1295 1488
rect 1208 1478 1245 1479
rect 133 1446 176 1451
rect 524 1457 971 1473
rect 524 1451 552 1457
rect 803 1456 971 1457
rect 133 1443 283 1446
rect 524 1443 551 1451
rect 133 1441 551 1443
rect 133 1423 142 1441
rect 160 1423 551 1441
rect 1264 1428 1295 1479
rect 1330 1508 1367 1578
rect 1633 1577 1670 1578
rect 1482 1518 1518 1519
rect 1330 1488 1339 1508
rect 1359 1488 1367 1508
rect 1330 1478 1367 1488
rect 1426 1508 1574 1518
rect 1674 1515 1770 1517
rect 1426 1488 1435 1508
rect 1455 1488 1545 1508
rect 1565 1488 1574 1508
rect 1426 1479 1574 1488
rect 1632 1508 1770 1515
rect 1632 1488 1641 1508
rect 1661 1488 1770 1508
rect 1632 1479 1770 1488
rect 1426 1478 1463 1479
rect 1156 1425 1197 1426
rect 133 1420 551 1423
rect 133 1414 176 1420
rect 136 1411 176 1414
rect 1048 1418 1197 1425
rect 533 1402 573 1403
rect 244 1385 573 1402
rect 1048 1398 1107 1418
rect 1127 1398 1166 1418
rect 1186 1398 1197 1418
rect 1048 1390 1197 1398
rect 1264 1421 1421 1428
rect 1264 1401 1384 1421
rect 1404 1401 1421 1421
rect 1264 1391 1421 1401
rect 1264 1390 1299 1391
rect 128 1342 171 1353
rect 128 1324 140 1342
rect 158 1324 171 1342
rect 128 1298 171 1324
rect 244 1298 271 1385
rect 533 1376 573 1385
rect 128 1277 271 1298
rect 315 1350 349 1366
rect 533 1356 926 1376
rect 946 1356 949 1376
rect 1264 1369 1295 1390
rect 1482 1369 1518 1479
rect 1537 1478 1574 1479
rect 1633 1478 1670 1479
rect 1593 1419 1683 1425
rect 1593 1399 1602 1419
rect 1622 1417 1683 1419
rect 1622 1399 1647 1417
rect 1593 1397 1647 1399
rect 1667 1397 1683 1417
rect 1593 1391 1683 1397
rect 1107 1368 1144 1369
rect 533 1351 949 1356
rect 1106 1359 1144 1368
rect 533 1350 874 1351
rect 315 1280 352 1350
rect 467 1290 498 1291
rect 128 1275 265 1277
rect 128 1233 171 1275
rect 315 1260 324 1280
rect 344 1260 352 1280
rect 315 1250 352 1260
rect 411 1280 498 1290
rect 411 1260 420 1280
rect 440 1260 498 1280
rect 411 1251 498 1260
rect 411 1250 448 1251
rect 126 1223 171 1233
rect 126 1205 135 1223
rect 153 1205 171 1223
rect 126 1199 171 1205
rect 467 1200 498 1251
rect 533 1280 570 1350
rect 836 1349 873 1350
rect 1106 1339 1115 1359
rect 1135 1339 1144 1359
rect 1106 1331 1144 1339
rect 1210 1363 1295 1369
rect 1325 1368 1362 1369
rect 1210 1343 1218 1363
rect 1238 1343 1295 1363
rect 1210 1335 1295 1343
rect 1324 1359 1362 1368
rect 1324 1339 1333 1359
rect 1353 1339 1362 1359
rect 1210 1334 1246 1335
rect 1324 1331 1362 1339
rect 1428 1363 1572 1369
rect 1428 1343 1436 1363
rect 1456 1344 1488 1363
rect 1509 1344 1544 1363
rect 1456 1343 1544 1344
rect 1564 1343 1572 1363
rect 1428 1335 1572 1343
rect 1428 1334 1464 1335
rect 1536 1334 1572 1335
rect 1638 1368 1675 1369
rect 1638 1367 1676 1368
rect 1638 1359 1702 1367
rect 1638 1339 1647 1359
rect 1667 1345 1702 1359
rect 1722 1345 1725 1365
rect 1667 1340 1725 1345
rect 1667 1339 1702 1340
rect 1107 1302 1144 1331
rect 1108 1300 1144 1302
rect 685 1290 721 1291
rect 533 1260 542 1280
rect 562 1260 570 1280
rect 533 1250 570 1260
rect 629 1280 777 1290
rect 877 1287 973 1289
rect 629 1260 638 1280
rect 658 1260 748 1280
rect 768 1260 777 1280
rect 629 1251 777 1260
rect 835 1280 973 1287
rect 835 1260 844 1280
rect 864 1260 973 1280
rect 1108 1278 1299 1300
rect 1325 1299 1362 1331
rect 1638 1327 1702 1339
rect 1742 1301 1769 1479
rect 1601 1299 1769 1301
rect 1325 1273 1769 1299
rect 835 1251 973 1260
rect 629 1250 666 1251
rect 126 1196 163 1199
rect 359 1197 400 1198
rect 251 1190 400 1197
rect 251 1170 310 1190
rect 330 1170 369 1190
rect 389 1170 400 1190
rect 251 1162 400 1170
rect 467 1193 624 1200
rect 467 1173 587 1193
rect 607 1173 624 1193
rect 467 1163 624 1173
rect 467 1162 502 1163
rect 467 1141 498 1162
rect 685 1141 721 1251
rect 740 1250 777 1251
rect 836 1250 873 1251
rect 796 1191 886 1197
rect 796 1171 805 1191
rect 825 1189 886 1191
rect 825 1171 850 1189
rect 796 1169 850 1171
rect 870 1169 886 1189
rect 796 1163 886 1169
rect 310 1140 347 1141
rect 123 1132 160 1134
rect 123 1124 165 1132
rect 123 1106 133 1124
rect 151 1106 165 1124
rect 123 1097 165 1106
rect 309 1131 347 1140
rect 309 1111 318 1131
rect 338 1111 347 1131
rect 309 1103 347 1111
rect 413 1135 498 1141
rect 528 1140 565 1141
rect 413 1115 421 1135
rect 441 1115 498 1135
rect 413 1107 498 1115
rect 527 1131 565 1140
rect 527 1111 536 1131
rect 556 1111 565 1131
rect 413 1106 449 1107
rect 527 1103 565 1111
rect 631 1139 775 1141
rect 631 1135 683 1139
rect 631 1115 639 1135
rect 659 1119 683 1135
rect 703 1135 775 1139
rect 703 1119 747 1135
rect 659 1115 747 1119
rect 767 1115 775 1135
rect 631 1107 775 1115
rect 631 1106 667 1107
rect 739 1106 775 1107
rect 841 1140 878 1141
rect 841 1139 879 1140
rect 841 1131 905 1139
rect 841 1111 850 1131
rect 870 1117 905 1131
rect 925 1117 928 1137
rect 870 1112 928 1117
rect 870 1111 905 1112
rect 124 1072 165 1097
rect 310 1072 347 1103
rect 528 1072 565 1103
rect 841 1099 905 1111
rect 945 1073 972 1251
rect 124 1045 173 1072
rect 309 1046 358 1072
rect 527 1071 608 1072
rect 804 1071 972 1073
rect 527 1046 972 1071
rect 528 1045 972 1046
rect 126 1012 173 1045
rect 529 1012 569 1045
rect 804 1044 972 1045
rect 1435 1049 1475 1273
rect 1601 1272 1769 1273
rect 1435 1027 1443 1049
rect 1467 1027 1475 1049
rect 1435 1019 1475 1027
rect 126 973 569 1012
rect 126 930 173 973
rect 529 968 569 973
rect 1194 971 1381 995
rect 1412 976 1805 996
rect 1825 976 1828 996
rect 1412 971 1828 976
rect 126 912 136 930
rect 154 912 173 930
rect 126 908 173 912
rect 127 903 164 908
rect 1194 900 1231 971
rect 1412 970 1753 971
rect 1346 910 1377 911
rect 1194 880 1203 900
rect 1223 880 1231 900
rect 1194 870 1231 880
rect 1290 900 1377 910
rect 1290 880 1299 900
rect 1319 880 1377 900
rect 1290 871 1377 880
rect 1290 870 1327 871
rect 115 841 167 843
rect 113 837 546 841
rect 113 831 552 837
rect 113 813 134 831
rect 152 813 552 831
rect 1346 820 1377 871
rect 1412 900 1449 970
rect 1715 969 1752 970
rect 1564 910 1600 911
rect 1412 880 1421 900
rect 1441 880 1449 900
rect 1412 870 1449 880
rect 1508 900 1656 910
rect 1756 907 1852 909
rect 1508 880 1517 900
rect 1537 880 1627 900
rect 1647 880 1656 900
rect 1508 871 1656 880
rect 1714 900 1852 907
rect 1714 880 1723 900
rect 1743 880 1852 900
rect 1714 871 1852 880
rect 1508 870 1545 871
rect 1238 817 1279 818
rect 113 795 552 813
rect 115 606 167 795
rect 513 770 552 795
rect 1130 810 1279 817
rect 1130 790 1189 810
rect 1209 790 1248 810
rect 1268 790 1279 810
rect 1130 782 1279 790
rect 1346 813 1503 820
rect 1346 793 1466 813
rect 1486 793 1503 813
rect 1346 783 1503 793
rect 1346 782 1381 783
rect 297 745 484 769
rect 513 750 908 770
rect 928 750 931 770
rect 1346 761 1377 782
rect 1564 761 1600 871
rect 1619 870 1656 871
rect 1715 870 1752 871
rect 1675 811 1765 817
rect 1675 791 1684 811
rect 1704 809 1765 811
rect 1704 791 1729 809
rect 1675 789 1729 791
rect 1749 789 1765 809
rect 1675 783 1765 789
rect 1189 760 1226 761
rect 513 745 931 750
rect 1188 751 1226 760
rect 297 674 334 745
rect 513 744 856 745
rect 513 741 552 744
rect 818 743 855 744
rect 449 684 480 685
rect 297 654 306 674
rect 326 654 334 674
rect 297 644 334 654
rect 393 674 480 684
rect 393 654 402 674
rect 422 654 480 674
rect 393 645 480 654
rect 393 644 430 645
rect 115 588 131 606
rect 149 588 167 606
rect 449 594 480 645
rect 515 674 552 741
rect 1188 731 1197 751
rect 1217 731 1226 751
rect 1188 723 1226 731
rect 1292 755 1377 761
rect 1407 760 1444 761
rect 1292 735 1300 755
rect 1320 735 1377 755
rect 1292 727 1377 735
rect 1406 751 1444 760
rect 1406 731 1415 751
rect 1435 731 1444 751
rect 1292 726 1328 727
rect 1406 723 1444 731
rect 1510 755 1654 761
rect 1510 735 1518 755
rect 1538 750 1626 755
rect 1538 735 1574 750
rect 1510 733 1574 735
rect 1593 735 1626 750
rect 1646 735 1654 755
rect 1593 733 1654 735
rect 1510 727 1654 733
rect 1510 726 1546 727
rect 1618 726 1654 727
rect 1720 760 1757 761
rect 1720 759 1758 760
rect 1720 751 1784 759
rect 1720 731 1729 751
rect 1749 737 1784 751
rect 1804 737 1807 757
rect 1749 732 1807 737
rect 1749 731 1784 732
rect 1189 694 1226 723
rect 1190 692 1226 694
rect 667 684 703 685
rect 515 654 524 674
rect 544 654 552 674
rect 515 644 552 654
rect 611 674 759 684
rect 859 681 955 683
rect 611 654 620 674
rect 640 654 730 674
rect 750 654 759 674
rect 611 645 759 654
rect 817 674 955 681
rect 817 654 826 674
rect 846 654 955 674
rect 1190 670 1381 692
rect 1407 691 1444 723
rect 1720 719 1784 731
rect 1824 693 1851 871
rect 1683 691 1851 693
rect 1407 677 1851 691
rect 1875 714 1903 1660
rect 1875 684 1920 714
rect 1407 665 1854 677
rect 1450 663 1483 665
rect 817 645 955 654
rect 611 644 648 645
rect 341 591 382 592
rect 115 570 167 588
rect 233 584 382 591
rect 233 564 292 584
rect 312 564 351 584
rect 371 564 382 584
rect 233 556 382 564
rect 449 587 606 594
rect 449 567 569 587
rect 589 567 606 587
rect 449 557 606 567
rect 449 556 484 557
rect 449 535 480 556
rect 667 535 703 645
rect 722 644 759 645
rect 818 644 855 645
rect 778 585 868 591
rect 778 565 787 585
rect 807 583 868 585
rect 807 565 832 583
rect 778 563 832 565
rect 852 563 868 583
rect 778 557 868 563
rect 292 534 329 535
rect 291 525 329 534
rect 119 507 159 517
rect 119 489 129 507
rect 147 489 159 507
rect 291 505 300 525
rect 320 505 329 525
rect 291 497 329 505
rect 395 529 480 535
rect 510 534 547 535
rect 395 509 403 529
rect 423 509 480 529
rect 395 501 480 509
rect 509 525 547 534
rect 509 505 518 525
rect 538 505 547 525
rect 395 500 431 501
rect 509 497 547 505
rect 613 529 757 535
rect 613 509 621 529
rect 641 509 674 529
rect 694 509 729 529
rect 749 509 757 529
rect 613 501 757 509
rect 613 500 649 501
rect 721 500 757 501
rect 823 534 860 535
rect 823 533 861 534
rect 823 525 887 533
rect 823 505 832 525
rect 852 511 887 525
rect 907 511 910 531
rect 852 506 910 511
rect 852 505 887 506
rect 119 433 159 489
rect 292 468 329 497
rect 293 466 329 468
rect 293 444 484 466
rect 510 465 547 497
rect 823 493 887 505
rect 927 467 954 645
rect 1812 620 1854 665
rect 1875 666 1886 684
rect 1908 666 1920 684
rect 1875 660 1920 666
rect 1876 659 1920 660
rect 786 465 954 467
rect 510 455 954 465
rect 1095 561 1282 585
rect 1313 566 1706 586
rect 1726 566 1729 586
rect 1313 561 1729 566
rect 1095 490 1132 561
rect 1313 560 1654 561
rect 1247 500 1278 501
rect 1095 470 1104 490
rect 1124 470 1132 490
rect 1095 460 1132 470
rect 1191 490 1278 500
rect 1191 470 1200 490
rect 1220 470 1278 490
rect 1191 461 1278 470
rect 1191 460 1228 461
rect 116 428 159 433
rect 507 439 954 455
rect 507 433 535 439
rect 786 438 954 439
rect 116 425 266 428
rect 507 425 534 433
rect 116 423 534 425
rect 116 405 125 423
rect 143 405 534 423
rect 1247 410 1278 461
rect 1313 490 1350 560
rect 1616 559 1653 560
rect 1465 500 1501 501
rect 1313 470 1322 490
rect 1342 470 1350 490
rect 1313 460 1350 470
rect 1409 490 1557 500
rect 1657 497 1753 499
rect 1409 470 1418 490
rect 1438 470 1528 490
rect 1548 470 1557 490
rect 1409 461 1557 470
rect 1615 490 1753 497
rect 1615 470 1624 490
rect 1644 470 1753 490
rect 1615 461 1753 470
rect 1409 460 1446 461
rect 1139 407 1180 408
rect 116 402 534 405
rect 116 396 159 402
rect 119 393 159 396
rect 1034 400 1180 407
rect 516 384 556 385
rect 227 367 556 384
rect 1034 380 1090 400
rect 1110 380 1149 400
rect 1169 380 1180 400
rect 1034 372 1180 380
rect 1247 403 1404 410
rect 1247 383 1367 403
rect 1387 383 1404 403
rect 1247 373 1404 383
rect 1247 372 1282 373
rect 111 324 154 335
rect 111 306 123 324
rect 141 306 154 324
rect 111 280 154 306
rect 227 280 254 367
rect 516 358 556 367
rect 111 259 254 280
rect 298 332 332 348
rect 516 338 909 358
rect 929 338 932 358
rect 1247 351 1278 372
rect 1465 351 1501 461
rect 1520 460 1557 461
rect 1616 460 1653 461
rect 1576 401 1666 407
rect 1576 381 1585 401
rect 1605 399 1666 401
rect 1605 381 1630 399
rect 1576 379 1630 381
rect 1650 379 1666 399
rect 1576 373 1666 379
rect 1090 350 1127 351
rect 516 333 932 338
rect 1089 341 1127 350
rect 516 332 857 333
rect 298 262 335 332
rect 450 272 481 273
rect 111 257 248 259
rect 111 215 154 257
rect 298 242 307 262
rect 327 242 335 262
rect 298 232 335 242
rect 394 262 481 272
rect 394 242 403 262
rect 423 242 481 262
rect 394 233 481 242
rect 394 232 431 233
rect 109 205 154 215
rect 109 187 118 205
rect 136 187 154 205
rect 109 181 154 187
rect 450 182 481 233
rect 516 262 553 332
rect 819 331 856 332
rect 1089 321 1098 341
rect 1118 321 1127 341
rect 1089 313 1127 321
rect 1193 345 1278 351
rect 1308 350 1345 351
rect 1193 325 1201 345
rect 1221 325 1278 345
rect 1193 317 1278 325
rect 1307 341 1345 350
rect 1307 321 1316 341
rect 1336 321 1345 341
rect 1193 316 1229 317
rect 1307 313 1345 321
rect 1411 345 1555 351
rect 1411 325 1419 345
rect 1439 342 1527 345
rect 1439 325 1474 342
rect 1411 324 1474 325
rect 1493 325 1527 342
rect 1547 325 1555 345
rect 1493 324 1555 325
rect 1411 317 1555 324
rect 1411 316 1447 317
rect 1519 316 1555 317
rect 1621 350 1658 351
rect 1621 349 1659 350
rect 1681 349 1708 353
rect 1621 347 1708 349
rect 1621 341 1685 347
rect 1621 321 1630 341
rect 1650 327 1685 341
rect 1705 327 1708 347
rect 1650 322 1708 327
rect 1650 321 1685 322
rect 1090 284 1127 313
rect 1091 282 1127 284
rect 668 272 704 273
rect 516 242 525 262
rect 545 242 553 262
rect 516 232 553 242
rect 612 262 760 272
rect 860 269 956 271
rect 612 242 621 262
rect 641 242 731 262
rect 751 242 760 262
rect 612 233 760 242
rect 818 262 956 269
rect 818 242 827 262
rect 847 242 956 262
rect 1091 260 1282 282
rect 1308 281 1345 313
rect 1621 309 1685 321
rect 1725 283 1752 461
rect 1584 281 1752 283
rect 1308 255 1752 281
rect 818 233 956 242
rect 612 232 649 233
rect 109 178 146 181
rect 342 179 383 180
rect 234 172 383 179
rect 234 152 293 172
rect 313 152 352 172
rect 372 152 383 172
rect 234 144 383 152
rect 450 175 607 182
rect 450 155 570 175
rect 590 155 607 175
rect 450 145 607 155
rect 450 144 485 145
rect 450 123 481 144
rect 668 123 704 233
rect 723 232 760 233
rect 819 232 856 233
rect 779 173 869 179
rect 779 153 788 173
rect 808 171 869 173
rect 808 153 833 171
rect 779 151 833 153
rect 853 151 869 171
rect 779 145 869 151
rect 293 122 330 123
rect 106 114 143 116
rect 106 106 148 114
rect 106 88 116 106
rect 134 88 148 106
rect 106 79 148 88
rect 292 113 330 122
rect 292 93 301 113
rect 321 93 330 113
rect 292 85 330 93
rect 396 117 481 123
rect 511 122 548 123
rect 396 97 404 117
rect 424 97 481 117
rect 396 89 481 97
rect 510 113 548 122
rect 510 93 519 113
rect 539 93 548 113
rect 396 88 432 89
rect 510 85 548 93
rect 614 121 758 123
rect 614 117 666 121
rect 614 97 622 117
rect 642 101 666 117
rect 686 117 758 121
rect 686 101 730 117
rect 642 97 730 101
rect 750 97 758 117
rect 614 89 758 97
rect 614 88 650 89
rect 722 88 758 89
rect 824 122 861 123
rect 824 121 862 122
rect 824 113 888 121
rect 824 93 833 113
rect 853 99 888 113
rect 908 99 911 119
rect 853 94 911 99
rect 853 93 888 94
rect 107 54 148 79
rect 293 54 330 85
rect 511 54 548 85
rect 824 81 888 93
rect 928 55 955 233
rect 107 20 150 54
rect 289 28 356 54
rect 511 53 591 54
rect 787 53 955 55
rect 511 27 955 53
rect 107 9 154 20
rect 511 10 546 27
rect 787 26 955 27
rect 1418 31 1458 255
rect 1584 254 1752 255
rect 1816 287 1849 620
rect 1816 279 1853 287
rect 1816 260 1824 279
rect 1845 260 1853 279
rect 1816 254 1853 260
rect 508 9 546 10
rect 107 -29 546 9
rect 1418 9 1426 31
rect 1450 9 1458 31
rect 1418 1 1458 9
rect 1729 -26 1794 -25
rect 107 -88 154 -29
rect 508 -30 546 -29
rect 107 -106 117 -88
rect 135 -106 154 -88
rect 107 -110 154 -106
rect 1380 -51 1567 -27
rect 1598 -46 1991 -26
rect 2011 -46 2014 -26
rect 1598 -51 2014 -46
rect 108 -115 145 -110
rect 1380 -122 1417 -51
rect 1598 -52 1939 -51
rect 1532 -112 1563 -111
rect 1380 -142 1389 -122
rect 1409 -142 1417 -122
rect 1380 -152 1417 -142
rect 1476 -122 1563 -112
rect 1476 -142 1485 -122
rect 1505 -142 1563 -122
rect 1476 -151 1563 -142
rect 1476 -152 1513 -151
rect 96 -177 148 -175
rect 94 -181 527 -177
rect 94 -187 533 -181
rect 94 -205 115 -187
rect 133 -205 533 -187
rect 1532 -202 1563 -151
rect 1598 -122 1635 -52
rect 1901 -53 1938 -52
rect 1750 -112 1786 -111
rect 1598 -142 1607 -122
rect 1627 -142 1635 -122
rect 1598 -152 1635 -142
rect 1694 -122 1842 -112
rect 1942 -115 2038 -113
rect 1694 -142 1703 -122
rect 1723 -142 1813 -122
rect 1833 -142 1842 -122
rect 1694 -151 1842 -142
rect 1900 -122 2038 -115
rect 1900 -142 1909 -122
rect 1929 -142 2038 -122
rect 1900 -151 2038 -142
rect 1694 -152 1731 -151
rect 1424 -205 1465 -204
rect 94 -223 533 -205
rect 96 -412 148 -223
rect 494 -248 533 -223
rect 1316 -212 1465 -205
rect 1316 -232 1375 -212
rect 1395 -232 1434 -212
rect 1454 -232 1465 -212
rect 1316 -240 1465 -232
rect 1532 -209 1689 -202
rect 1532 -229 1652 -209
rect 1672 -229 1689 -209
rect 1532 -239 1689 -229
rect 1532 -240 1567 -239
rect 278 -273 465 -249
rect 494 -268 889 -248
rect 909 -268 912 -248
rect 1532 -261 1563 -240
rect 1750 -261 1786 -151
rect 1805 -152 1842 -151
rect 1901 -152 1938 -151
rect 1861 -211 1951 -205
rect 1861 -231 1870 -211
rect 1890 -213 1951 -211
rect 1890 -231 1915 -213
rect 1861 -233 1915 -231
rect 1935 -233 1951 -213
rect 1861 -239 1951 -233
rect 1375 -262 1412 -261
rect 494 -273 912 -268
rect 1374 -271 1412 -262
rect 278 -344 315 -273
rect 494 -274 837 -273
rect 494 -277 533 -274
rect 799 -275 836 -274
rect 430 -334 461 -333
rect 278 -364 287 -344
rect 307 -364 315 -344
rect 278 -374 315 -364
rect 374 -344 461 -334
rect 374 -364 383 -344
rect 403 -364 461 -344
rect 374 -373 461 -364
rect 374 -374 411 -373
rect 96 -430 112 -412
rect 130 -430 148 -412
rect 430 -424 461 -373
rect 496 -344 533 -277
rect 1374 -291 1383 -271
rect 1403 -291 1412 -271
rect 1374 -299 1412 -291
rect 1478 -267 1563 -261
rect 1593 -262 1630 -261
rect 1478 -287 1486 -267
rect 1506 -287 1563 -267
rect 1478 -295 1563 -287
rect 1592 -271 1630 -262
rect 1592 -291 1601 -271
rect 1621 -291 1630 -271
rect 1478 -296 1514 -295
rect 1592 -299 1630 -291
rect 1696 -267 1840 -261
rect 1696 -287 1704 -267
rect 1724 -287 1812 -267
rect 1832 -287 1840 -267
rect 1696 -295 1840 -287
rect 1696 -296 1732 -295
rect 1804 -296 1840 -295
rect 1906 -262 1943 -261
rect 1906 -263 1944 -262
rect 1906 -271 1970 -263
rect 1906 -291 1915 -271
rect 1935 -285 1970 -271
rect 1990 -285 1993 -265
rect 1935 -290 1993 -285
rect 1935 -291 1970 -290
rect 1375 -328 1412 -299
rect 1376 -330 1412 -328
rect 648 -334 684 -333
rect 496 -364 505 -344
rect 525 -364 533 -344
rect 496 -374 533 -364
rect 592 -344 740 -334
rect 840 -337 936 -335
rect 592 -364 601 -344
rect 621 -364 711 -344
rect 731 -364 740 -344
rect 592 -373 740 -364
rect 798 -344 936 -337
rect 798 -364 807 -344
rect 827 -364 936 -344
rect 1376 -352 1567 -330
rect 1593 -331 1630 -299
rect 1906 -303 1970 -291
rect 2010 -329 2037 -151
rect 1869 -331 2037 -329
rect 1593 -357 2037 -331
rect 1703 -359 1743 -357
rect 1869 -358 2037 -357
rect 798 -373 936 -364
rect 1996 -363 2037 -358
rect 592 -374 629 -373
rect 322 -427 363 -426
rect 96 -448 148 -430
rect 214 -434 363 -427
rect 214 -454 273 -434
rect 293 -454 332 -434
rect 352 -454 363 -434
rect 214 -462 363 -454
rect 430 -431 587 -424
rect 430 -451 550 -431
rect 570 -451 587 -431
rect 430 -461 587 -451
rect 430 -462 465 -461
rect 430 -483 461 -462
rect 648 -483 684 -373
rect 703 -374 740 -373
rect 799 -374 836 -373
rect 759 -433 849 -427
rect 759 -453 768 -433
rect 788 -435 849 -433
rect 788 -453 813 -435
rect 759 -455 813 -453
rect 833 -455 849 -435
rect 759 -461 849 -455
rect 273 -484 310 -483
rect 272 -493 310 -484
rect 100 -511 140 -501
rect 100 -529 110 -511
rect 128 -529 140 -511
rect 272 -513 281 -493
rect 301 -513 310 -493
rect 272 -521 310 -513
rect 376 -489 461 -483
rect 491 -484 528 -483
rect 376 -509 384 -489
rect 404 -509 461 -489
rect 376 -517 461 -509
rect 490 -493 528 -484
rect 490 -513 499 -493
rect 519 -513 528 -493
rect 376 -518 412 -517
rect 490 -521 528 -513
rect 594 -489 738 -483
rect 594 -509 602 -489
rect 622 -509 655 -489
rect 675 -509 710 -489
rect 730 -509 738 -489
rect 594 -517 738 -509
rect 594 -518 630 -517
rect 702 -518 738 -517
rect 804 -484 841 -483
rect 804 -485 842 -484
rect 804 -493 868 -485
rect 804 -513 813 -493
rect 833 -507 868 -493
rect 888 -507 891 -487
rect 833 -512 891 -507
rect 833 -513 868 -512
rect 100 -585 140 -529
rect 273 -550 310 -521
rect 274 -552 310 -550
rect 274 -574 465 -552
rect 491 -553 528 -521
rect 804 -525 868 -513
rect 908 -551 935 -373
rect 767 -553 935 -551
rect 491 -563 935 -553
rect 1076 -457 1263 -433
rect 1294 -452 1687 -432
rect 1707 -452 1710 -432
rect 1294 -457 1710 -452
rect 1076 -528 1113 -457
rect 1294 -458 1635 -457
rect 1228 -518 1259 -517
rect 1076 -548 1085 -528
rect 1105 -548 1113 -528
rect 1076 -558 1113 -548
rect 1172 -528 1259 -518
rect 1172 -548 1181 -528
rect 1201 -548 1259 -528
rect 1172 -557 1259 -548
rect 1172 -558 1209 -557
rect 97 -590 140 -585
rect 488 -579 935 -563
rect 488 -585 516 -579
rect 767 -580 935 -579
rect 97 -593 247 -590
rect 488 -593 515 -585
rect 97 -595 515 -593
rect 97 -613 106 -595
rect 124 -613 515 -595
rect 1228 -608 1259 -557
rect 1294 -528 1331 -458
rect 1597 -459 1634 -458
rect 1446 -518 1482 -517
rect 1294 -548 1303 -528
rect 1323 -548 1331 -528
rect 1294 -558 1331 -548
rect 1390 -528 1538 -518
rect 1638 -521 1734 -519
rect 1390 -548 1399 -528
rect 1419 -548 1509 -528
rect 1529 -548 1538 -528
rect 1390 -557 1538 -548
rect 1596 -528 1734 -521
rect 1596 -548 1605 -528
rect 1625 -548 1734 -528
rect 1996 -545 2036 -363
rect 1596 -557 1734 -548
rect 1390 -558 1427 -557
rect 1120 -611 1161 -610
rect 97 -616 515 -613
rect 97 -622 140 -616
rect 100 -625 140 -622
rect 1012 -618 1161 -611
rect 497 -634 537 -633
rect 208 -651 537 -634
rect 1012 -638 1071 -618
rect 1091 -638 1130 -618
rect 1150 -638 1161 -618
rect 1012 -646 1161 -638
rect 1228 -615 1385 -608
rect 1228 -635 1348 -615
rect 1368 -635 1385 -615
rect 1228 -645 1385 -635
rect 1228 -646 1263 -645
rect 92 -694 135 -683
rect 92 -712 104 -694
rect 122 -712 135 -694
rect 92 -738 135 -712
rect 208 -738 235 -651
rect 497 -660 537 -651
rect 92 -759 235 -738
rect 279 -686 313 -670
rect 497 -680 890 -660
rect 910 -680 913 -660
rect 1228 -667 1259 -646
rect 1446 -667 1482 -557
rect 1501 -558 1538 -557
rect 1597 -558 1634 -557
rect 1557 -617 1647 -611
rect 1557 -637 1566 -617
rect 1586 -619 1647 -617
rect 1586 -637 1611 -619
rect 1557 -639 1611 -637
rect 1631 -639 1647 -619
rect 1557 -645 1647 -639
rect 1071 -668 1108 -667
rect 497 -685 913 -680
rect 1070 -677 1108 -668
rect 497 -686 838 -685
rect 279 -756 316 -686
rect 431 -746 462 -745
rect 92 -761 229 -759
rect 92 -803 135 -761
rect 279 -776 288 -756
rect 308 -776 316 -756
rect 279 -786 316 -776
rect 375 -756 462 -746
rect 375 -776 384 -756
rect 404 -776 462 -756
rect 375 -785 462 -776
rect 375 -786 412 -785
rect 90 -813 135 -803
rect 90 -831 99 -813
rect 117 -831 135 -813
rect 90 -837 135 -831
rect 431 -836 462 -785
rect 497 -756 534 -686
rect 800 -687 837 -686
rect 1070 -697 1079 -677
rect 1099 -697 1108 -677
rect 1070 -705 1108 -697
rect 1174 -673 1259 -667
rect 1289 -668 1326 -667
rect 1174 -693 1182 -673
rect 1202 -693 1259 -673
rect 1174 -701 1259 -693
rect 1288 -677 1326 -668
rect 1288 -697 1297 -677
rect 1317 -697 1326 -677
rect 1174 -702 1210 -701
rect 1288 -705 1326 -697
rect 1392 -673 1536 -667
rect 1392 -693 1400 -673
rect 1420 -692 1452 -673
rect 1473 -692 1508 -673
rect 1420 -693 1508 -692
rect 1528 -693 1536 -673
rect 1392 -701 1536 -693
rect 1392 -702 1428 -701
rect 1500 -702 1536 -701
rect 1602 -668 1639 -667
rect 1602 -669 1640 -668
rect 1602 -677 1666 -669
rect 1602 -697 1611 -677
rect 1631 -691 1666 -677
rect 1686 -691 1689 -671
rect 1631 -696 1689 -691
rect 1631 -697 1666 -696
rect 1071 -734 1108 -705
rect 1072 -736 1108 -734
rect 649 -746 685 -745
rect 497 -776 506 -756
rect 526 -776 534 -756
rect 497 -786 534 -776
rect 593 -756 741 -746
rect 841 -749 937 -747
rect 593 -776 602 -756
rect 622 -776 712 -756
rect 732 -776 741 -756
rect 593 -785 741 -776
rect 799 -756 937 -749
rect 799 -776 808 -756
rect 828 -776 937 -756
rect 1072 -758 1263 -736
rect 1289 -737 1326 -705
rect 1602 -709 1666 -697
rect 1706 -735 1733 -557
rect 1565 -737 1733 -735
rect 1289 -763 1733 -737
rect 799 -785 937 -776
rect 593 -786 630 -785
rect 90 -840 127 -837
rect 323 -839 364 -838
rect 215 -846 364 -839
rect 215 -866 274 -846
rect 294 -866 333 -846
rect 353 -866 364 -846
rect 215 -874 364 -866
rect 431 -843 588 -836
rect 431 -863 551 -843
rect 571 -863 588 -843
rect 431 -873 588 -863
rect 431 -874 466 -873
rect 431 -895 462 -874
rect 649 -895 685 -785
rect 704 -786 741 -785
rect 800 -786 837 -785
rect 760 -845 850 -839
rect 760 -865 769 -845
rect 789 -847 850 -845
rect 789 -865 814 -847
rect 760 -867 814 -865
rect 834 -867 850 -847
rect 760 -873 850 -867
rect 274 -896 311 -895
rect 87 -904 124 -902
rect 87 -912 129 -904
rect 87 -930 97 -912
rect 115 -930 129 -912
rect 87 -939 129 -930
rect 273 -905 311 -896
rect 273 -925 282 -905
rect 302 -925 311 -905
rect 273 -933 311 -925
rect 377 -901 462 -895
rect 492 -896 529 -895
rect 377 -921 385 -901
rect 405 -921 462 -901
rect 377 -929 462 -921
rect 491 -905 529 -896
rect 491 -925 500 -905
rect 520 -925 529 -905
rect 377 -930 413 -929
rect 491 -933 529 -925
rect 595 -897 739 -895
rect 595 -901 647 -897
rect 595 -921 603 -901
rect 623 -917 647 -901
rect 667 -901 739 -897
rect 667 -917 711 -901
rect 623 -921 711 -917
rect 731 -921 739 -901
rect 595 -929 739 -921
rect 595 -930 631 -929
rect 703 -930 739 -929
rect 805 -896 842 -895
rect 805 -897 843 -896
rect 805 -905 869 -897
rect 805 -925 814 -905
rect 834 -919 869 -905
rect 889 -919 892 -899
rect 834 -924 892 -919
rect 834 -925 869 -924
rect 88 -964 129 -939
rect 274 -964 311 -933
rect 492 -964 529 -933
rect 805 -937 869 -925
rect 909 -963 936 -785
rect 88 -991 137 -964
rect 273 -990 322 -964
rect 491 -965 572 -964
rect 768 -965 936 -963
rect 491 -990 936 -965
rect 492 -991 936 -990
rect 90 -1024 137 -991
rect 493 -1024 533 -991
rect 768 -992 936 -991
rect 1399 -987 1439 -763
rect 1565 -764 1733 -763
rect 1399 -1009 1407 -987
rect 1431 -1009 1439 -987
rect 1399 -1017 1439 -1009
rect 90 -1063 533 -1024
rect 90 -1106 137 -1063
rect 493 -1068 533 -1063
rect 1158 -1065 1345 -1041
rect 1376 -1060 1769 -1040
rect 1789 -1060 1792 -1040
rect 1376 -1065 1792 -1060
rect 90 -1124 100 -1106
rect 118 -1124 137 -1106
rect 90 -1128 137 -1124
rect 91 -1133 128 -1128
rect 1158 -1136 1195 -1065
rect 1376 -1066 1717 -1065
rect 1310 -1126 1341 -1125
rect 1158 -1156 1167 -1136
rect 1187 -1156 1195 -1136
rect 1158 -1166 1195 -1156
rect 1254 -1136 1341 -1126
rect 1254 -1156 1263 -1136
rect 1283 -1156 1341 -1136
rect 1254 -1165 1341 -1156
rect 1254 -1166 1291 -1165
rect 79 -1195 131 -1193
rect 77 -1199 510 -1195
rect 77 -1205 516 -1199
rect 77 -1223 98 -1205
rect 116 -1223 516 -1205
rect 1310 -1216 1341 -1165
rect 1376 -1136 1413 -1066
rect 1679 -1067 1716 -1066
rect 1528 -1126 1564 -1125
rect 1376 -1156 1385 -1136
rect 1405 -1156 1413 -1136
rect 1376 -1166 1413 -1156
rect 1472 -1136 1620 -1126
rect 1720 -1129 1816 -1127
rect 1472 -1156 1481 -1136
rect 1501 -1156 1591 -1136
rect 1611 -1156 1620 -1136
rect 1472 -1165 1620 -1156
rect 1678 -1136 1816 -1129
rect 1678 -1156 1687 -1136
rect 1707 -1156 1816 -1136
rect 1678 -1165 1816 -1156
rect 1472 -1166 1509 -1165
rect 1202 -1219 1243 -1218
rect 77 -1241 516 -1223
rect 79 -1430 131 -1241
rect 477 -1266 516 -1241
rect 1094 -1226 1243 -1219
rect 1094 -1246 1153 -1226
rect 1173 -1246 1212 -1226
rect 1232 -1246 1243 -1226
rect 1094 -1254 1243 -1246
rect 1310 -1223 1467 -1216
rect 1310 -1243 1430 -1223
rect 1450 -1243 1467 -1223
rect 1310 -1253 1467 -1243
rect 1310 -1254 1345 -1253
rect 261 -1291 448 -1267
rect 477 -1286 872 -1266
rect 892 -1286 895 -1266
rect 1310 -1275 1341 -1254
rect 1528 -1275 1564 -1165
rect 1583 -1166 1620 -1165
rect 1679 -1166 1716 -1165
rect 1639 -1225 1729 -1219
rect 1639 -1245 1648 -1225
rect 1668 -1227 1729 -1225
rect 1668 -1245 1693 -1227
rect 1639 -1247 1693 -1245
rect 1713 -1247 1729 -1227
rect 1639 -1253 1729 -1247
rect 1153 -1276 1190 -1275
rect 477 -1291 895 -1286
rect 1152 -1285 1190 -1276
rect 261 -1362 298 -1291
rect 477 -1292 820 -1291
rect 477 -1295 516 -1292
rect 782 -1293 819 -1292
rect 413 -1352 444 -1351
rect 261 -1382 270 -1362
rect 290 -1382 298 -1362
rect 261 -1392 298 -1382
rect 357 -1362 444 -1352
rect 357 -1382 366 -1362
rect 386 -1382 444 -1362
rect 357 -1391 444 -1382
rect 357 -1392 394 -1391
rect 79 -1448 95 -1430
rect 113 -1448 131 -1430
rect 413 -1442 444 -1391
rect 479 -1362 516 -1295
rect 1152 -1305 1161 -1285
rect 1181 -1305 1190 -1285
rect 1152 -1313 1190 -1305
rect 1256 -1281 1341 -1275
rect 1371 -1276 1408 -1275
rect 1256 -1301 1264 -1281
rect 1284 -1301 1341 -1281
rect 1256 -1309 1341 -1301
rect 1370 -1285 1408 -1276
rect 1370 -1305 1379 -1285
rect 1399 -1305 1408 -1285
rect 1256 -1310 1292 -1309
rect 1370 -1313 1408 -1305
rect 1474 -1280 1618 -1275
rect 1474 -1281 1536 -1280
rect 1474 -1301 1482 -1281
rect 1502 -1299 1536 -1281
rect 1557 -1281 1618 -1280
rect 1557 -1299 1590 -1281
rect 1502 -1301 1590 -1299
rect 1610 -1301 1618 -1281
rect 1474 -1309 1618 -1301
rect 1474 -1310 1510 -1309
rect 1582 -1310 1618 -1309
rect 1684 -1276 1721 -1275
rect 1684 -1277 1722 -1276
rect 1684 -1285 1748 -1277
rect 1684 -1305 1693 -1285
rect 1713 -1299 1748 -1285
rect 1768 -1299 1771 -1279
rect 1713 -1304 1771 -1299
rect 1713 -1305 1748 -1304
rect 1153 -1342 1190 -1313
rect 1154 -1344 1190 -1342
rect 631 -1352 667 -1351
rect 479 -1382 488 -1362
rect 508 -1382 516 -1362
rect 479 -1392 516 -1382
rect 575 -1362 723 -1352
rect 823 -1355 919 -1353
rect 575 -1382 584 -1362
rect 604 -1382 694 -1362
rect 714 -1382 723 -1362
rect 575 -1391 723 -1382
rect 781 -1362 919 -1355
rect 781 -1382 790 -1362
rect 810 -1382 919 -1362
rect 1154 -1366 1345 -1344
rect 1371 -1345 1408 -1313
rect 1684 -1317 1748 -1305
rect 1788 -1343 1815 -1165
rect 1647 -1345 1815 -1343
rect 1371 -1359 1815 -1345
rect 1371 -1371 1818 -1359
rect 1414 -1373 1447 -1371
rect 781 -1391 919 -1382
rect 575 -1392 612 -1391
rect 305 -1445 346 -1444
rect 79 -1466 131 -1448
rect 197 -1452 346 -1445
rect 197 -1472 256 -1452
rect 276 -1472 315 -1452
rect 335 -1472 346 -1452
rect 197 -1480 346 -1472
rect 413 -1449 570 -1442
rect 413 -1469 533 -1449
rect 553 -1469 570 -1449
rect 413 -1479 570 -1469
rect 413 -1480 448 -1479
rect 413 -1501 444 -1480
rect 631 -1501 667 -1391
rect 686 -1392 723 -1391
rect 782 -1392 819 -1391
rect 742 -1451 832 -1445
rect 742 -1471 751 -1451
rect 771 -1453 832 -1451
rect 771 -1471 796 -1453
rect 742 -1473 796 -1471
rect 816 -1473 832 -1453
rect 742 -1479 832 -1473
rect 256 -1502 293 -1501
rect 255 -1511 293 -1502
rect 83 -1529 123 -1519
rect 83 -1547 93 -1529
rect 111 -1547 123 -1529
rect 255 -1531 264 -1511
rect 284 -1531 293 -1511
rect 255 -1539 293 -1531
rect 359 -1507 444 -1501
rect 474 -1502 511 -1501
rect 359 -1527 367 -1507
rect 387 -1527 444 -1507
rect 359 -1535 444 -1527
rect 473 -1511 511 -1502
rect 473 -1531 482 -1511
rect 502 -1531 511 -1511
rect 359 -1536 395 -1535
rect 473 -1539 511 -1531
rect 577 -1507 721 -1501
rect 577 -1527 585 -1507
rect 605 -1527 638 -1507
rect 658 -1527 693 -1507
rect 713 -1527 721 -1507
rect 577 -1535 721 -1527
rect 577 -1536 613 -1535
rect 685 -1536 721 -1535
rect 787 -1502 824 -1501
rect 787 -1503 825 -1502
rect 787 -1511 851 -1503
rect 787 -1531 796 -1511
rect 816 -1525 851 -1511
rect 871 -1525 874 -1505
rect 816 -1530 874 -1525
rect 816 -1531 851 -1530
rect 83 -1603 123 -1547
rect 256 -1568 293 -1539
rect 257 -1570 293 -1568
rect 257 -1592 448 -1570
rect 474 -1571 511 -1539
rect 787 -1543 851 -1531
rect 891 -1569 918 -1391
rect 1776 -1416 1818 -1371
rect 750 -1571 918 -1569
rect 474 -1581 918 -1571
rect 1059 -1475 1246 -1451
rect 1277 -1470 1670 -1450
rect 1690 -1470 1693 -1450
rect 1277 -1475 1693 -1470
rect 1059 -1546 1096 -1475
rect 1277 -1476 1618 -1475
rect 1211 -1536 1242 -1535
rect 1059 -1566 1068 -1546
rect 1088 -1566 1096 -1546
rect 1059 -1576 1096 -1566
rect 1155 -1546 1242 -1536
rect 1155 -1566 1164 -1546
rect 1184 -1566 1242 -1546
rect 1155 -1575 1242 -1566
rect 1155 -1576 1192 -1575
rect 80 -1608 123 -1603
rect 471 -1597 918 -1581
rect 471 -1603 499 -1597
rect 750 -1598 918 -1597
rect 80 -1611 230 -1608
rect 471 -1611 498 -1603
rect 80 -1613 498 -1611
rect 80 -1631 89 -1613
rect 107 -1631 498 -1613
rect 1211 -1626 1242 -1575
rect 1277 -1546 1314 -1476
rect 1580 -1477 1617 -1476
rect 1429 -1536 1465 -1535
rect 1277 -1566 1286 -1546
rect 1306 -1566 1314 -1546
rect 1277 -1576 1314 -1566
rect 1373 -1546 1521 -1536
rect 1621 -1539 1717 -1537
rect 1373 -1566 1382 -1546
rect 1402 -1566 1492 -1546
rect 1512 -1566 1521 -1546
rect 1373 -1575 1521 -1566
rect 1579 -1546 1717 -1539
rect 1579 -1566 1588 -1546
rect 1608 -1566 1717 -1546
rect 1579 -1575 1717 -1566
rect 1373 -1576 1410 -1575
rect 1103 -1629 1144 -1628
rect 80 -1634 498 -1631
rect 80 -1640 123 -1634
rect 83 -1643 123 -1640
rect 998 -1636 1144 -1629
rect 480 -1652 520 -1651
rect 191 -1669 520 -1652
rect 998 -1656 1054 -1636
rect 1074 -1656 1113 -1636
rect 1133 -1656 1144 -1636
rect 998 -1664 1144 -1656
rect 1211 -1633 1368 -1626
rect 1211 -1653 1331 -1633
rect 1351 -1653 1368 -1633
rect 1211 -1663 1368 -1653
rect 1211 -1664 1246 -1663
rect 75 -1712 118 -1701
rect 75 -1730 87 -1712
rect 105 -1730 118 -1712
rect 75 -1756 118 -1730
rect 191 -1756 218 -1669
rect 480 -1678 520 -1669
rect 75 -1777 218 -1756
rect 262 -1704 296 -1688
rect 480 -1698 873 -1678
rect 893 -1698 896 -1678
rect 1211 -1685 1242 -1664
rect 1429 -1685 1465 -1575
rect 1484 -1576 1521 -1575
rect 1580 -1576 1617 -1575
rect 1540 -1635 1630 -1629
rect 1540 -1655 1549 -1635
rect 1569 -1637 1630 -1635
rect 1569 -1655 1594 -1637
rect 1540 -1657 1594 -1655
rect 1614 -1657 1630 -1637
rect 1540 -1663 1630 -1657
rect 1054 -1686 1091 -1685
rect 480 -1703 896 -1698
rect 1053 -1695 1091 -1686
rect 480 -1704 821 -1703
rect 262 -1774 299 -1704
rect 414 -1764 445 -1763
rect 75 -1779 212 -1777
rect 75 -1821 118 -1779
rect 262 -1794 271 -1774
rect 291 -1794 299 -1774
rect 262 -1804 299 -1794
rect 358 -1774 445 -1764
rect 358 -1794 367 -1774
rect 387 -1794 445 -1774
rect 358 -1803 445 -1794
rect 358 -1804 395 -1803
rect 73 -1831 118 -1821
rect 73 -1849 82 -1831
rect 100 -1849 118 -1831
rect 73 -1855 118 -1849
rect 414 -1854 445 -1803
rect 480 -1774 517 -1704
rect 783 -1705 820 -1704
rect 1053 -1715 1062 -1695
rect 1082 -1715 1091 -1695
rect 1053 -1723 1091 -1715
rect 1157 -1691 1242 -1685
rect 1272 -1686 1309 -1685
rect 1157 -1711 1165 -1691
rect 1185 -1711 1242 -1691
rect 1157 -1719 1242 -1711
rect 1271 -1695 1309 -1686
rect 1271 -1715 1280 -1695
rect 1300 -1715 1309 -1695
rect 1157 -1720 1193 -1719
rect 1271 -1723 1309 -1715
rect 1375 -1691 1519 -1685
rect 1375 -1711 1383 -1691
rect 1403 -1694 1491 -1691
rect 1403 -1711 1438 -1694
rect 1375 -1712 1438 -1711
rect 1457 -1711 1491 -1694
rect 1511 -1711 1519 -1691
rect 1457 -1712 1519 -1711
rect 1375 -1719 1519 -1712
rect 1375 -1720 1411 -1719
rect 1483 -1720 1519 -1719
rect 1585 -1686 1622 -1685
rect 1585 -1687 1623 -1686
rect 1645 -1687 1672 -1683
rect 1585 -1689 1672 -1687
rect 1585 -1695 1649 -1689
rect 1585 -1715 1594 -1695
rect 1614 -1709 1649 -1695
rect 1669 -1709 1672 -1689
rect 1614 -1714 1672 -1709
rect 1614 -1715 1649 -1714
rect 1054 -1752 1091 -1723
rect 1055 -1754 1091 -1752
rect 632 -1764 668 -1763
rect 480 -1794 489 -1774
rect 509 -1794 517 -1774
rect 480 -1804 517 -1794
rect 576 -1774 724 -1764
rect 824 -1767 920 -1765
rect 576 -1794 585 -1774
rect 605 -1794 695 -1774
rect 715 -1794 724 -1774
rect 576 -1803 724 -1794
rect 782 -1774 920 -1767
rect 782 -1794 791 -1774
rect 811 -1794 920 -1774
rect 1055 -1776 1246 -1754
rect 1272 -1755 1309 -1723
rect 1585 -1727 1649 -1715
rect 1689 -1753 1716 -1575
rect 1548 -1755 1716 -1753
rect 1272 -1781 1716 -1755
rect 782 -1803 920 -1794
rect 576 -1804 613 -1803
rect 73 -1858 110 -1855
rect 306 -1857 347 -1856
rect 198 -1864 347 -1857
rect 198 -1884 257 -1864
rect 277 -1884 316 -1864
rect 336 -1884 347 -1864
rect 198 -1892 347 -1884
rect 414 -1861 571 -1854
rect 414 -1881 534 -1861
rect 554 -1881 571 -1861
rect 414 -1891 571 -1881
rect 414 -1892 449 -1891
rect 414 -1913 445 -1892
rect 632 -1913 668 -1803
rect 687 -1804 724 -1803
rect 783 -1804 820 -1803
rect 743 -1863 833 -1857
rect 743 -1883 752 -1863
rect 772 -1865 833 -1863
rect 772 -1883 797 -1865
rect 743 -1885 797 -1883
rect 817 -1885 833 -1865
rect 743 -1891 833 -1885
rect 257 -1914 294 -1913
rect 69 -1922 107 -1920
rect 69 -1930 112 -1922
rect 69 -1948 80 -1930
rect 98 -1948 112 -1930
rect 69 -1975 112 -1948
rect 256 -1923 294 -1914
rect 256 -1943 265 -1923
rect 285 -1943 294 -1923
rect 256 -1951 294 -1943
rect 360 -1919 445 -1913
rect 475 -1914 512 -1913
rect 360 -1939 368 -1919
rect 388 -1939 445 -1919
rect 360 -1947 445 -1939
rect 474 -1923 512 -1914
rect 474 -1943 483 -1923
rect 503 -1943 512 -1923
rect 360 -1948 396 -1947
rect 474 -1951 512 -1943
rect 578 -1915 722 -1913
rect 578 -1919 630 -1915
rect 578 -1939 586 -1919
rect 606 -1935 630 -1919
rect 650 -1919 722 -1915
rect 650 -1935 694 -1919
rect 606 -1939 694 -1935
rect 714 -1939 722 -1919
rect 578 -1947 722 -1939
rect 578 -1948 614 -1947
rect 686 -1948 722 -1947
rect 788 -1914 825 -1913
rect 788 -1915 826 -1914
rect 788 -1923 852 -1915
rect 788 -1943 797 -1923
rect 817 -1937 852 -1923
rect 872 -1937 875 -1917
rect 817 -1942 875 -1937
rect 817 -1943 852 -1942
rect 70 -1982 112 -1975
rect 257 -1982 294 -1951
rect 475 -1982 512 -1951
rect 788 -1955 852 -1943
rect 892 -1981 919 -1803
rect 70 -2022 115 -1982
rect 257 -2007 402 -1982
rect 475 -1983 555 -1982
rect 751 -1983 919 -1981
rect 475 -1999 919 -1983
rect 259 -2008 402 -2007
rect 474 -2009 919 -1999
rect 70 -2043 117 -2022
rect 474 -2043 515 -2009
rect 751 -2010 919 -2009
rect 1382 -2005 1422 -1781
rect 1548 -1782 1716 -1781
rect 1780 -1749 1813 -1416
rect 1780 -1757 1817 -1749
rect 1780 -1776 1788 -1757
rect 1809 -1776 1817 -1757
rect 1780 -1782 1817 -1776
rect 1382 -2027 1390 -2005
rect 1414 -2027 1422 -2005
rect 1382 -2035 1422 -2027
rect 70 -2073 515 -2043
rect 1553 -2060 1618 -2059
rect 70 -2076 493 -2073
rect 70 -2124 117 -2076
rect 70 -2142 80 -2124
rect 98 -2142 117 -2124
rect 70 -2146 117 -2142
rect 1204 -2085 1391 -2061
rect 1422 -2080 1815 -2060
rect 1835 -2080 1838 -2060
rect 1422 -2085 1838 -2080
rect 71 -2151 108 -2146
rect 1204 -2156 1241 -2085
rect 1422 -2086 1763 -2085
rect 1356 -2146 1387 -2145
rect 1204 -2176 1213 -2156
rect 1233 -2176 1241 -2156
rect 1204 -2186 1241 -2176
rect 1300 -2156 1387 -2146
rect 1300 -2176 1309 -2156
rect 1329 -2176 1387 -2156
rect 1300 -2185 1387 -2176
rect 1300 -2186 1337 -2185
rect 59 -2213 111 -2211
rect 57 -2217 490 -2213
rect 57 -2223 496 -2217
rect 57 -2241 78 -2223
rect 96 -2241 496 -2223
rect 1356 -2236 1387 -2185
rect 1422 -2156 1459 -2086
rect 1725 -2087 1762 -2086
rect 1574 -2146 1610 -2145
rect 1422 -2176 1431 -2156
rect 1451 -2176 1459 -2156
rect 1422 -2186 1459 -2176
rect 1518 -2156 1666 -2146
rect 1766 -2149 1862 -2147
rect 1518 -2176 1527 -2156
rect 1547 -2176 1637 -2156
rect 1657 -2176 1666 -2156
rect 1518 -2185 1666 -2176
rect 1724 -2156 1862 -2149
rect 1724 -2176 1733 -2156
rect 1753 -2176 1862 -2156
rect 1724 -2185 1862 -2176
rect 1518 -2186 1555 -2185
rect 1248 -2239 1289 -2238
rect 57 -2259 496 -2241
rect 59 -2448 111 -2259
rect 457 -2284 496 -2259
rect 1140 -2246 1289 -2239
rect 1140 -2266 1199 -2246
rect 1219 -2266 1258 -2246
rect 1278 -2266 1289 -2246
rect 1140 -2274 1289 -2266
rect 1356 -2243 1513 -2236
rect 1356 -2263 1476 -2243
rect 1496 -2263 1513 -2243
rect 1356 -2273 1513 -2263
rect 1356 -2274 1391 -2273
rect 241 -2309 428 -2285
rect 457 -2304 852 -2284
rect 872 -2304 875 -2284
rect 1356 -2295 1387 -2274
rect 1574 -2295 1610 -2185
rect 1629 -2186 1666 -2185
rect 1725 -2186 1762 -2185
rect 1685 -2245 1775 -2239
rect 1685 -2265 1694 -2245
rect 1714 -2247 1775 -2245
rect 1714 -2265 1739 -2247
rect 1685 -2267 1739 -2265
rect 1759 -2267 1775 -2247
rect 1685 -2273 1775 -2267
rect 1199 -2296 1236 -2295
rect 457 -2309 875 -2304
rect 1198 -2305 1236 -2296
rect 241 -2380 278 -2309
rect 457 -2310 800 -2309
rect 457 -2313 496 -2310
rect 762 -2311 799 -2310
rect 393 -2370 424 -2369
rect 241 -2400 250 -2380
rect 270 -2400 278 -2380
rect 241 -2410 278 -2400
rect 337 -2380 424 -2370
rect 337 -2400 346 -2380
rect 366 -2400 424 -2380
rect 337 -2409 424 -2400
rect 337 -2410 374 -2409
rect 59 -2466 75 -2448
rect 93 -2466 111 -2448
rect 393 -2460 424 -2409
rect 459 -2380 496 -2313
rect 1198 -2325 1207 -2305
rect 1227 -2325 1236 -2305
rect 1198 -2333 1236 -2325
rect 1302 -2301 1387 -2295
rect 1417 -2296 1454 -2295
rect 1302 -2321 1310 -2301
rect 1330 -2321 1387 -2301
rect 1302 -2329 1387 -2321
rect 1416 -2305 1454 -2296
rect 1416 -2325 1425 -2305
rect 1445 -2325 1454 -2305
rect 1302 -2330 1338 -2329
rect 1416 -2333 1454 -2325
rect 1520 -2297 1664 -2295
rect 1520 -2301 1580 -2297
rect 1520 -2321 1528 -2301
rect 1548 -2319 1580 -2301
rect 1603 -2301 1664 -2297
rect 1603 -2319 1636 -2301
rect 1548 -2321 1636 -2319
rect 1656 -2321 1664 -2301
rect 1520 -2329 1664 -2321
rect 1520 -2330 1556 -2329
rect 1628 -2330 1664 -2329
rect 1730 -2296 1767 -2295
rect 1730 -2297 1768 -2296
rect 1730 -2305 1794 -2297
rect 1730 -2325 1739 -2305
rect 1759 -2319 1794 -2305
rect 1814 -2319 1817 -2299
rect 1759 -2324 1817 -2319
rect 1759 -2325 1794 -2324
rect 1199 -2362 1236 -2333
rect 1200 -2364 1236 -2362
rect 611 -2370 647 -2369
rect 459 -2400 468 -2380
rect 488 -2400 496 -2380
rect 459 -2410 496 -2400
rect 555 -2380 703 -2370
rect 803 -2373 899 -2371
rect 555 -2400 564 -2380
rect 584 -2400 674 -2380
rect 694 -2400 703 -2380
rect 555 -2409 703 -2400
rect 761 -2380 899 -2373
rect 761 -2400 770 -2380
rect 790 -2400 899 -2380
rect 1200 -2386 1391 -2364
rect 1417 -2365 1454 -2333
rect 1730 -2337 1794 -2325
rect 1417 -2366 1692 -2365
rect 1834 -2366 1861 -2185
rect 1417 -2391 1861 -2366
rect 1997 -2360 2036 -545
rect 1997 -2382 2004 -2360
rect 2028 -2382 2036 -2360
rect 1997 -2388 2036 -2382
rect 1527 -2393 1567 -2391
rect 1693 -2392 1861 -2391
rect 1795 -2393 1832 -2392
rect 761 -2409 899 -2400
rect 555 -2410 592 -2409
rect 285 -2463 326 -2462
rect 59 -2484 111 -2466
rect 177 -2470 326 -2463
rect 177 -2490 236 -2470
rect 256 -2490 295 -2470
rect 315 -2490 326 -2470
rect 177 -2498 326 -2490
rect 393 -2467 550 -2460
rect 393 -2487 513 -2467
rect 533 -2487 550 -2467
rect 393 -2497 550 -2487
rect 393 -2498 428 -2497
rect 393 -2519 424 -2498
rect 611 -2519 647 -2409
rect 666 -2410 703 -2409
rect 762 -2410 799 -2409
rect 722 -2469 812 -2463
rect 722 -2489 731 -2469
rect 751 -2471 812 -2469
rect 751 -2489 776 -2471
rect 722 -2491 776 -2489
rect 796 -2491 812 -2471
rect 722 -2497 812 -2491
rect 236 -2520 273 -2519
rect 235 -2529 273 -2520
rect 63 -2547 103 -2537
rect 63 -2565 73 -2547
rect 91 -2565 103 -2547
rect 235 -2549 244 -2529
rect 264 -2549 273 -2529
rect 235 -2557 273 -2549
rect 339 -2525 424 -2519
rect 454 -2520 491 -2519
rect 339 -2545 347 -2525
rect 367 -2545 424 -2525
rect 339 -2553 424 -2545
rect 453 -2529 491 -2520
rect 453 -2549 462 -2529
rect 482 -2549 491 -2529
rect 339 -2554 375 -2553
rect 453 -2557 491 -2549
rect 557 -2525 701 -2519
rect 557 -2545 565 -2525
rect 585 -2545 618 -2525
rect 638 -2545 673 -2525
rect 693 -2545 701 -2525
rect 557 -2553 701 -2545
rect 557 -2554 593 -2553
rect 665 -2554 701 -2553
rect 767 -2520 804 -2519
rect 767 -2521 805 -2520
rect 767 -2529 831 -2521
rect 767 -2549 776 -2529
rect 796 -2543 831 -2529
rect 851 -2543 854 -2523
rect 796 -2548 854 -2543
rect 796 -2549 831 -2548
rect 63 -2621 103 -2565
rect 236 -2586 273 -2557
rect 237 -2588 273 -2586
rect 237 -2610 428 -2588
rect 454 -2589 491 -2557
rect 767 -2561 831 -2549
rect 871 -2587 898 -2409
rect 730 -2589 898 -2587
rect 454 -2599 898 -2589
rect 1039 -2493 1226 -2469
rect 1257 -2488 1650 -2468
rect 1670 -2488 1673 -2468
rect 1257 -2493 1673 -2488
rect 1039 -2564 1076 -2493
rect 1257 -2494 1598 -2493
rect 1191 -2554 1222 -2553
rect 1039 -2584 1048 -2564
rect 1068 -2584 1076 -2564
rect 1039 -2594 1076 -2584
rect 1135 -2564 1222 -2554
rect 1135 -2584 1144 -2564
rect 1164 -2584 1222 -2564
rect 1135 -2593 1222 -2584
rect 1135 -2594 1172 -2593
rect 60 -2626 103 -2621
rect 451 -2615 898 -2599
rect 451 -2621 479 -2615
rect 730 -2616 898 -2615
rect 60 -2629 210 -2626
rect 451 -2629 478 -2621
rect 60 -2631 478 -2629
rect 60 -2649 69 -2631
rect 87 -2649 478 -2631
rect 1191 -2644 1222 -2593
rect 1257 -2564 1294 -2494
rect 1560 -2495 1597 -2494
rect 1798 -2552 1831 -2393
rect 1409 -2554 1445 -2553
rect 1257 -2584 1266 -2564
rect 1286 -2584 1294 -2564
rect 1257 -2594 1294 -2584
rect 1353 -2564 1501 -2554
rect 1601 -2557 1697 -2555
rect 1353 -2584 1362 -2564
rect 1382 -2584 1472 -2564
rect 1492 -2584 1501 -2564
rect 1353 -2593 1501 -2584
rect 1559 -2564 1697 -2557
rect 1559 -2584 1568 -2564
rect 1588 -2584 1697 -2564
rect 1798 -2556 1834 -2552
rect 1798 -2574 1807 -2556
rect 1829 -2574 1834 -2556
rect 1798 -2580 1834 -2574
rect 1559 -2593 1697 -2584
rect 1353 -2594 1390 -2593
rect 1083 -2647 1124 -2646
rect 60 -2652 478 -2649
rect 60 -2658 103 -2652
rect 63 -2661 103 -2658
rect 975 -2654 1124 -2647
rect 460 -2670 500 -2669
rect 171 -2687 500 -2670
rect 975 -2674 1034 -2654
rect 1054 -2674 1093 -2654
rect 1113 -2674 1124 -2654
rect 975 -2682 1124 -2674
rect 1191 -2651 1348 -2644
rect 1191 -2671 1311 -2651
rect 1331 -2671 1348 -2651
rect 1191 -2681 1348 -2671
rect 1191 -2682 1226 -2681
rect 55 -2730 98 -2719
rect 55 -2748 67 -2730
rect 85 -2748 98 -2730
rect 55 -2774 98 -2748
rect 171 -2774 198 -2687
rect 460 -2696 500 -2687
rect 55 -2795 198 -2774
rect 242 -2722 276 -2706
rect 460 -2716 853 -2696
rect 873 -2716 876 -2696
rect 1191 -2703 1222 -2682
rect 1409 -2703 1445 -2593
rect 1464 -2594 1501 -2593
rect 1560 -2594 1597 -2593
rect 1520 -2653 1610 -2647
rect 1520 -2673 1529 -2653
rect 1549 -2655 1610 -2653
rect 1549 -2673 1574 -2655
rect 1520 -2675 1574 -2673
rect 1594 -2675 1610 -2655
rect 1520 -2681 1610 -2675
rect 1034 -2704 1071 -2703
rect 460 -2721 876 -2716
rect 1033 -2713 1071 -2704
rect 460 -2722 801 -2721
rect 242 -2792 279 -2722
rect 394 -2782 425 -2781
rect 55 -2797 192 -2795
rect 55 -2839 98 -2797
rect 242 -2812 251 -2792
rect 271 -2812 279 -2792
rect 242 -2822 279 -2812
rect 338 -2792 425 -2782
rect 338 -2812 347 -2792
rect 367 -2812 425 -2792
rect 338 -2821 425 -2812
rect 338 -2822 375 -2821
rect 53 -2849 98 -2839
rect 53 -2867 62 -2849
rect 80 -2867 98 -2849
rect 53 -2873 98 -2867
rect 394 -2872 425 -2821
rect 460 -2792 497 -2722
rect 763 -2723 800 -2722
rect 1033 -2733 1042 -2713
rect 1062 -2733 1071 -2713
rect 1033 -2741 1071 -2733
rect 1137 -2709 1222 -2703
rect 1252 -2704 1289 -2703
rect 1137 -2729 1145 -2709
rect 1165 -2729 1222 -2709
rect 1137 -2737 1222 -2729
rect 1251 -2713 1289 -2704
rect 1251 -2733 1260 -2713
rect 1280 -2733 1289 -2713
rect 1137 -2738 1173 -2737
rect 1251 -2741 1289 -2733
rect 1355 -2709 1499 -2703
rect 1355 -2729 1363 -2709
rect 1383 -2728 1415 -2709
rect 1436 -2728 1471 -2709
rect 1383 -2729 1471 -2728
rect 1491 -2729 1499 -2709
rect 1355 -2737 1499 -2729
rect 1355 -2738 1391 -2737
rect 1463 -2738 1499 -2737
rect 1565 -2704 1602 -2703
rect 1565 -2705 1603 -2704
rect 1565 -2713 1629 -2705
rect 1565 -2733 1574 -2713
rect 1594 -2727 1629 -2713
rect 1649 -2727 1652 -2707
rect 1594 -2732 1652 -2727
rect 1594 -2733 1629 -2732
rect 1034 -2770 1071 -2741
rect 1035 -2772 1071 -2770
rect 612 -2782 648 -2781
rect 460 -2812 469 -2792
rect 489 -2812 497 -2792
rect 460 -2822 497 -2812
rect 556 -2792 704 -2782
rect 804 -2785 900 -2783
rect 556 -2812 565 -2792
rect 585 -2812 675 -2792
rect 695 -2812 704 -2792
rect 556 -2821 704 -2812
rect 762 -2792 900 -2785
rect 762 -2812 771 -2792
rect 791 -2812 900 -2792
rect 1035 -2794 1226 -2772
rect 1252 -2773 1289 -2741
rect 1565 -2745 1629 -2733
rect 1669 -2771 1696 -2593
rect 1528 -2773 1696 -2771
rect 1252 -2799 1696 -2773
rect 762 -2821 900 -2812
rect 556 -2822 593 -2821
rect 53 -2876 90 -2873
rect 286 -2875 327 -2874
rect 178 -2882 327 -2875
rect 178 -2902 237 -2882
rect 257 -2902 296 -2882
rect 316 -2902 327 -2882
rect 178 -2910 327 -2902
rect 394 -2879 551 -2872
rect 394 -2899 514 -2879
rect 534 -2899 551 -2879
rect 394 -2909 551 -2899
rect 394 -2910 429 -2909
rect 394 -2931 425 -2910
rect 612 -2931 648 -2821
rect 667 -2822 704 -2821
rect 763 -2822 800 -2821
rect 723 -2881 813 -2875
rect 723 -2901 732 -2881
rect 752 -2883 813 -2881
rect 752 -2901 777 -2883
rect 723 -2903 777 -2901
rect 797 -2903 813 -2883
rect 723 -2909 813 -2903
rect 237 -2932 274 -2931
rect 50 -2940 87 -2938
rect 50 -2948 92 -2940
rect 50 -2966 60 -2948
rect 78 -2966 92 -2948
rect 50 -2975 92 -2966
rect 236 -2941 274 -2932
rect 236 -2961 245 -2941
rect 265 -2961 274 -2941
rect 236 -2969 274 -2961
rect 340 -2937 425 -2931
rect 455 -2932 492 -2931
rect 340 -2957 348 -2937
rect 368 -2957 425 -2937
rect 340 -2965 425 -2957
rect 454 -2941 492 -2932
rect 454 -2961 463 -2941
rect 483 -2961 492 -2941
rect 340 -2966 376 -2965
rect 454 -2969 492 -2961
rect 558 -2933 702 -2931
rect 558 -2937 610 -2933
rect 558 -2957 566 -2937
rect 586 -2953 610 -2937
rect 630 -2937 702 -2933
rect 630 -2953 674 -2937
rect 586 -2957 674 -2953
rect 694 -2957 702 -2937
rect 558 -2965 702 -2957
rect 558 -2966 594 -2965
rect 666 -2966 702 -2965
rect 768 -2932 805 -2931
rect 768 -2933 806 -2932
rect 768 -2941 832 -2933
rect 768 -2961 777 -2941
rect 797 -2955 832 -2941
rect 852 -2955 855 -2935
rect 797 -2960 855 -2955
rect 797 -2961 832 -2960
rect 51 -3000 92 -2975
rect 237 -3000 274 -2969
rect 455 -3000 492 -2969
rect 768 -2973 832 -2961
rect 872 -2999 899 -2821
rect 51 -3027 100 -3000
rect 236 -3026 285 -3000
rect 454 -3001 535 -3000
rect 731 -3001 899 -2999
rect 454 -3026 899 -3001
rect 455 -3027 899 -3026
rect 53 -3060 100 -3027
rect 456 -3060 496 -3027
rect 731 -3028 899 -3027
rect 1362 -3023 1402 -2799
rect 1528 -2800 1696 -2799
rect 1362 -3045 1370 -3023
rect 1394 -3045 1402 -3023
rect 1362 -3053 1402 -3045
rect 53 -3099 496 -3060
rect 53 -3142 100 -3099
rect 456 -3104 496 -3099
rect 1121 -3101 1308 -3077
rect 1339 -3096 1732 -3076
rect 1752 -3096 1755 -3076
rect 1339 -3101 1755 -3096
rect 53 -3160 63 -3142
rect 81 -3160 100 -3142
rect 53 -3164 100 -3160
rect 54 -3169 91 -3164
rect 1121 -3172 1158 -3101
rect 1339 -3102 1680 -3101
rect 1273 -3162 1304 -3161
rect 1121 -3192 1130 -3172
rect 1150 -3192 1158 -3172
rect 1121 -3202 1158 -3192
rect 1217 -3172 1304 -3162
rect 1217 -3192 1226 -3172
rect 1246 -3192 1304 -3172
rect 1217 -3201 1304 -3192
rect 1217 -3202 1254 -3201
rect 42 -3231 94 -3229
rect 40 -3235 473 -3231
rect 40 -3241 479 -3235
rect 40 -3259 61 -3241
rect 79 -3259 479 -3241
rect 1273 -3252 1304 -3201
rect 1339 -3172 1376 -3102
rect 1642 -3103 1679 -3102
rect 1491 -3162 1527 -3161
rect 1339 -3192 1348 -3172
rect 1368 -3192 1376 -3172
rect 1339 -3202 1376 -3192
rect 1435 -3172 1583 -3162
rect 1683 -3165 1779 -3163
rect 1435 -3192 1444 -3172
rect 1464 -3192 1554 -3172
rect 1574 -3192 1583 -3172
rect 1435 -3201 1583 -3192
rect 1641 -3172 1779 -3165
rect 1641 -3192 1650 -3172
rect 1670 -3192 1779 -3172
rect 1641 -3201 1779 -3192
rect 1435 -3202 1472 -3201
rect 1165 -3255 1206 -3254
rect 40 -3277 479 -3259
rect 42 -3466 94 -3277
rect 440 -3302 479 -3277
rect 1057 -3262 1206 -3255
rect 1057 -3282 1116 -3262
rect 1136 -3282 1175 -3262
rect 1195 -3282 1206 -3262
rect 1057 -3290 1206 -3282
rect 1273 -3259 1430 -3252
rect 1273 -3279 1393 -3259
rect 1413 -3279 1430 -3259
rect 1273 -3289 1430 -3279
rect 1273 -3290 1308 -3289
rect 224 -3327 411 -3303
rect 440 -3322 835 -3302
rect 855 -3322 858 -3302
rect 1273 -3311 1304 -3290
rect 1491 -3311 1527 -3201
rect 1546 -3202 1583 -3201
rect 1642 -3202 1679 -3201
rect 1602 -3261 1692 -3255
rect 1602 -3281 1611 -3261
rect 1631 -3263 1692 -3261
rect 1631 -3281 1656 -3263
rect 1602 -3283 1656 -3281
rect 1676 -3283 1692 -3263
rect 1602 -3289 1692 -3283
rect 1116 -3312 1153 -3311
rect 440 -3327 858 -3322
rect 1115 -3321 1153 -3312
rect 224 -3398 261 -3327
rect 440 -3328 783 -3327
rect 440 -3331 479 -3328
rect 745 -3329 782 -3328
rect 376 -3388 407 -3387
rect 224 -3418 233 -3398
rect 253 -3418 261 -3398
rect 224 -3428 261 -3418
rect 320 -3398 407 -3388
rect 320 -3418 329 -3398
rect 349 -3418 407 -3398
rect 320 -3427 407 -3418
rect 320 -3428 357 -3427
rect 42 -3484 58 -3466
rect 76 -3484 94 -3466
rect 376 -3478 407 -3427
rect 442 -3398 479 -3331
rect 1115 -3341 1124 -3321
rect 1144 -3341 1153 -3321
rect 1115 -3349 1153 -3341
rect 1219 -3317 1304 -3311
rect 1334 -3312 1371 -3311
rect 1219 -3337 1227 -3317
rect 1247 -3337 1304 -3317
rect 1219 -3345 1304 -3337
rect 1333 -3321 1371 -3312
rect 1333 -3341 1342 -3321
rect 1362 -3341 1371 -3321
rect 1219 -3346 1255 -3345
rect 1333 -3349 1371 -3341
rect 1437 -3317 1581 -3311
rect 1437 -3337 1445 -3317
rect 1465 -3322 1553 -3317
rect 1465 -3337 1501 -3322
rect 1437 -3339 1501 -3337
rect 1520 -3337 1553 -3322
rect 1573 -3337 1581 -3317
rect 1520 -3339 1581 -3337
rect 1437 -3345 1581 -3339
rect 1437 -3346 1473 -3345
rect 1545 -3346 1581 -3345
rect 1647 -3312 1684 -3311
rect 1647 -3313 1685 -3312
rect 1647 -3321 1711 -3313
rect 1647 -3341 1656 -3321
rect 1676 -3335 1711 -3321
rect 1731 -3335 1734 -3315
rect 1676 -3340 1734 -3335
rect 1676 -3341 1711 -3340
rect 1116 -3378 1153 -3349
rect 1117 -3380 1153 -3378
rect 594 -3388 630 -3387
rect 442 -3418 451 -3398
rect 471 -3418 479 -3398
rect 442 -3428 479 -3418
rect 538 -3398 686 -3388
rect 786 -3391 882 -3389
rect 538 -3418 547 -3398
rect 567 -3418 657 -3398
rect 677 -3418 686 -3398
rect 538 -3427 686 -3418
rect 744 -3398 882 -3391
rect 744 -3418 753 -3398
rect 773 -3418 882 -3398
rect 1117 -3402 1308 -3380
rect 1334 -3381 1371 -3349
rect 1647 -3353 1711 -3341
rect 1751 -3379 1778 -3201
rect 1610 -3381 1778 -3379
rect 1334 -3395 1778 -3381
rect 1334 -3407 1781 -3395
rect 1377 -3409 1410 -3407
rect 744 -3427 882 -3418
rect 538 -3428 575 -3427
rect 268 -3481 309 -3480
rect 42 -3502 94 -3484
rect 160 -3488 309 -3481
rect 160 -3508 219 -3488
rect 239 -3508 278 -3488
rect 298 -3508 309 -3488
rect 160 -3516 309 -3508
rect 376 -3485 533 -3478
rect 376 -3505 496 -3485
rect 516 -3505 533 -3485
rect 376 -3515 533 -3505
rect 376 -3516 411 -3515
rect 376 -3537 407 -3516
rect 594 -3537 630 -3427
rect 649 -3428 686 -3427
rect 745 -3428 782 -3427
rect 705 -3487 795 -3481
rect 705 -3507 714 -3487
rect 734 -3489 795 -3487
rect 734 -3507 759 -3489
rect 705 -3509 759 -3507
rect 779 -3509 795 -3489
rect 705 -3515 795 -3509
rect 219 -3538 256 -3537
rect 218 -3547 256 -3538
rect 46 -3565 86 -3555
rect 46 -3583 56 -3565
rect 74 -3583 86 -3565
rect 218 -3567 227 -3547
rect 247 -3567 256 -3547
rect 218 -3575 256 -3567
rect 322 -3543 407 -3537
rect 437 -3538 474 -3537
rect 322 -3563 330 -3543
rect 350 -3563 407 -3543
rect 322 -3571 407 -3563
rect 436 -3547 474 -3538
rect 436 -3567 445 -3547
rect 465 -3567 474 -3547
rect 322 -3572 358 -3571
rect 436 -3575 474 -3567
rect 540 -3543 684 -3537
rect 540 -3563 548 -3543
rect 568 -3563 601 -3543
rect 621 -3563 656 -3543
rect 676 -3563 684 -3543
rect 540 -3571 684 -3563
rect 540 -3572 576 -3571
rect 648 -3572 684 -3571
rect 750 -3538 787 -3537
rect 750 -3539 788 -3538
rect 750 -3547 814 -3539
rect 750 -3567 759 -3547
rect 779 -3561 814 -3547
rect 834 -3561 837 -3541
rect 779 -3566 837 -3561
rect 779 -3567 814 -3566
rect 46 -3639 86 -3583
rect 219 -3604 256 -3575
rect 220 -3606 256 -3604
rect 220 -3628 411 -3606
rect 437 -3607 474 -3575
rect 750 -3579 814 -3567
rect 854 -3605 881 -3427
rect 1739 -3452 1781 -3407
rect 713 -3607 881 -3605
rect 437 -3617 881 -3607
rect 1022 -3511 1209 -3487
rect 1240 -3506 1633 -3486
rect 1653 -3506 1656 -3486
rect 1240 -3511 1656 -3506
rect 1022 -3582 1059 -3511
rect 1240 -3512 1581 -3511
rect 1174 -3572 1205 -3571
rect 1022 -3602 1031 -3582
rect 1051 -3602 1059 -3582
rect 1022 -3612 1059 -3602
rect 1118 -3582 1205 -3572
rect 1118 -3602 1127 -3582
rect 1147 -3602 1205 -3582
rect 1118 -3611 1205 -3602
rect 1118 -3612 1155 -3611
rect 43 -3644 86 -3639
rect 434 -3633 881 -3617
rect 434 -3639 462 -3633
rect 713 -3634 881 -3633
rect 43 -3647 193 -3644
rect 434 -3647 461 -3639
rect 43 -3649 461 -3647
rect 43 -3667 52 -3649
rect 70 -3667 461 -3649
rect 1174 -3662 1205 -3611
rect 1240 -3582 1277 -3512
rect 1543 -3513 1580 -3512
rect 1392 -3572 1428 -3571
rect 1240 -3602 1249 -3582
rect 1269 -3602 1277 -3582
rect 1240 -3612 1277 -3602
rect 1336 -3582 1484 -3572
rect 1584 -3575 1680 -3573
rect 1336 -3602 1345 -3582
rect 1365 -3602 1455 -3582
rect 1475 -3602 1484 -3582
rect 1336 -3611 1484 -3602
rect 1542 -3582 1680 -3575
rect 1542 -3602 1551 -3582
rect 1571 -3602 1680 -3582
rect 1542 -3611 1680 -3602
rect 1336 -3612 1373 -3611
rect 1066 -3665 1107 -3664
rect 43 -3670 461 -3667
rect 43 -3676 86 -3670
rect 46 -3679 86 -3676
rect 961 -3672 1107 -3665
rect 443 -3688 483 -3687
rect 154 -3705 483 -3688
rect 961 -3692 1017 -3672
rect 1037 -3692 1076 -3672
rect 1096 -3692 1107 -3672
rect 961 -3700 1107 -3692
rect 1174 -3669 1331 -3662
rect 1174 -3689 1294 -3669
rect 1314 -3689 1331 -3669
rect 1174 -3699 1331 -3689
rect 1174 -3700 1209 -3699
rect 38 -3748 81 -3737
rect 38 -3766 50 -3748
rect 68 -3766 81 -3748
rect 38 -3792 81 -3766
rect 154 -3792 181 -3705
rect 443 -3714 483 -3705
rect 38 -3813 181 -3792
rect 225 -3740 259 -3724
rect 443 -3734 836 -3714
rect 856 -3734 859 -3714
rect 1174 -3721 1205 -3700
rect 1392 -3721 1428 -3611
rect 1447 -3612 1484 -3611
rect 1543 -3612 1580 -3611
rect 1503 -3671 1593 -3665
rect 1503 -3691 1512 -3671
rect 1532 -3673 1593 -3671
rect 1532 -3691 1557 -3673
rect 1503 -3693 1557 -3691
rect 1577 -3693 1593 -3673
rect 1503 -3699 1593 -3693
rect 1017 -3722 1054 -3721
rect 443 -3739 859 -3734
rect 1016 -3731 1054 -3722
rect 443 -3740 784 -3739
rect 225 -3810 262 -3740
rect 377 -3800 408 -3799
rect 38 -3815 175 -3813
rect 38 -3857 81 -3815
rect 225 -3830 234 -3810
rect 254 -3830 262 -3810
rect 225 -3840 262 -3830
rect 321 -3810 408 -3800
rect 321 -3830 330 -3810
rect 350 -3830 408 -3810
rect 321 -3839 408 -3830
rect 321 -3840 358 -3839
rect 36 -3867 81 -3857
rect 36 -3885 45 -3867
rect 63 -3885 81 -3867
rect 36 -3891 81 -3885
rect 377 -3890 408 -3839
rect 443 -3810 480 -3740
rect 746 -3741 783 -3740
rect 1016 -3751 1025 -3731
rect 1045 -3751 1054 -3731
rect 1016 -3759 1054 -3751
rect 1120 -3727 1205 -3721
rect 1235 -3722 1272 -3721
rect 1120 -3747 1128 -3727
rect 1148 -3747 1205 -3727
rect 1120 -3755 1205 -3747
rect 1234 -3731 1272 -3722
rect 1234 -3751 1243 -3731
rect 1263 -3751 1272 -3731
rect 1120 -3756 1156 -3755
rect 1234 -3759 1272 -3751
rect 1338 -3727 1482 -3721
rect 1338 -3747 1346 -3727
rect 1366 -3730 1454 -3727
rect 1366 -3747 1401 -3730
rect 1338 -3748 1401 -3747
rect 1420 -3747 1454 -3730
rect 1474 -3747 1482 -3727
rect 1420 -3748 1482 -3747
rect 1338 -3755 1482 -3748
rect 1338 -3756 1374 -3755
rect 1446 -3756 1482 -3755
rect 1548 -3722 1585 -3721
rect 1548 -3723 1586 -3722
rect 1608 -3723 1635 -3719
rect 1548 -3725 1635 -3723
rect 1548 -3731 1612 -3725
rect 1548 -3751 1557 -3731
rect 1577 -3745 1612 -3731
rect 1632 -3745 1635 -3725
rect 1577 -3750 1635 -3745
rect 1577 -3751 1612 -3750
rect 1017 -3788 1054 -3759
rect 1018 -3790 1054 -3788
rect 595 -3800 631 -3799
rect 443 -3830 452 -3810
rect 472 -3830 480 -3810
rect 443 -3840 480 -3830
rect 539 -3810 687 -3800
rect 787 -3803 883 -3801
rect 539 -3830 548 -3810
rect 568 -3830 658 -3810
rect 678 -3830 687 -3810
rect 539 -3839 687 -3830
rect 745 -3810 883 -3803
rect 745 -3830 754 -3810
rect 774 -3830 883 -3810
rect 1018 -3812 1209 -3790
rect 1235 -3791 1272 -3759
rect 1548 -3763 1612 -3751
rect 1652 -3789 1679 -3611
rect 1511 -3791 1679 -3789
rect 1235 -3817 1679 -3791
rect 745 -3839 883 -3830
rect 539 -3840 576 -3839
rect 36 -3894 73 -3891
rect 269 -3893 310 -3892
rect 161 -3900 310 -3893
rect 161 -3920 220 -3900
rect 240 -3920 279 -3900
rect 299 -3920 310 -3900
rect 161 -3928 310 -3920
rect 377 -3897 534 -3890
rect 377 -3917 497 -3897
rect 517 -3917 534 -3897
rect 377 -3927 534 -3917
rect 377 -3928 412 -3927
rect 377 -3949 408 -3928
rect 595 -3949 631 -3839
rect 650 -3840 687 -3839
rect 746 -3840 783 -3839
rect 706 -3899 796 -3893
rect 706 -3919 715 -3899
rect 735 -3901 796 -3899
rect 735 -3919 760 -3901
rect 706 -3921 760 -3919
rect 780 -3921 796 -3901
rect 706 -3927 796 -3921
rect 220 -3950 257 -3949
rect 33 -3958 70 -3956
rect 33 -3966 75 -3958
rect 33 -3984 43 -3966
rect 61 -3984 75 -3966
rect 33 -3993 75 -3984
rect 219 -3959 257 -3950
rect 219 -3979 228 -3959
rect 248 -3979 257 -3959
rect 219 -3987 257 -3979
rect 323 -3955 408 -3949
rect 438 -3950 475 -3949
rect 323 -3975 331 -3955
rect 351 -3975 408 -3955
rect 323 -3983 408 -3975
rect 437 -3959 475 -3950
rect 437 -3979 446 -3959
rect 466 -3979 475 -3959
rect 323 -3984 359 -3983
rect 437 -3987 475 -3979
rect 541 -3951 685 -3949
rect 541 -3955 593 -3951
rect 541 -3975 549 -3955
rect 569 -3971 593 -3955
rect 613 -3955 685 -3951
rect 613 -3971 657 -3955
rect 569 -3975 657 -3971
rect 677 -3975 685 -3955
rect 541 -3983 685 -3975
rect 541 -3984 577 -3983
rect 649 -3984 685 -3983
rect 751 -3950 788 -3949
rect 751 -3951 789 -3950
rect 751 -3959 815 -3951
rect 751 -3979 760 -3959
rect 780 -3973 815 -3959
rect 835 -3973 838 -3953
rect 780 -3978 838 -3973
rect 780 -3979 815 -3978
rect 34 -4018 75 -3993
rect 220 -4018 257 -3987
rect 438 -4018 475 -3987
rect 751 -3991 815 -3979
rect 855 -4017 882 -3839
rect 34 -4019 518 -4018
rect 714 -4019 882 -4017
rect 34 -4044 882 -4019
rect 34 -4045 75 -4044
rect 438 -4045 882 -4044
rect 714 -4046 882 -4045
rect 1345 -4041 1385 -3817
rect 1511 -3818 1679 -3817
rect 1743 -3785 1776 -3452
rect 1743 -3793 1780 -3785
rect 1743 -3812 1751 -3793
rect 1772 -3812 1780 -3793
rect 1743 -3818 1780 -3812
rect 1345 -4063 1353 -4041
rect 1377 -4063 1385 -4041
rect 1345 -4071 1385 -4063
<< viali >>
rect 962 3804 982 3824
rect 346 3618 366 3638
rect 886 3617 906 3637
rect 728 3563 748 3583
rect 941 3565 961 3585
rect 1760 3620 1780 3640
rect 1144 3434 1164 3454
rect 963 3392 983 3412
rect 1684 3433 1704 3453
rect 1525 3380 1546 3399
rect 1739 3381 1759 3401
rect 347 3206 367 3226
rect 887 3205 907 3225
rect 720 3155 740 3175
rect 942 3153 962 3173
rect 1480 3063 1504 3085
rect 1842 3012 1862 3032
rect 1226 2826 1246 2846
rect 945 2786 965 2806
rect 1766 2825 1786 2845
rect 1609 2773 1630 2792
rect 1821 2773 1841 2793
rect 329 2600 349 2620
rect 869 2599 889 2619
rect 711 2545 731 2565
rect 924 2547 944 2567
rect 1743 2602 1763 2622
rect 1127 2416 1147 2436
rect 946 2374 966 2394
rect 1667 2415 1687 2435
rect 1511 2360 1530 2378
rect 1722 2363 1742 2383
rect 330 2188 350 2208
rect 870 2187 890 2207
rect 703 2137 723 2157
rect 925 2135 945 2155
rect 1861 2296 1882 2315
rect 1463 2045 1487 2067
rect 1888 1992 1908 2012
rect 1272 1806 1292 1826
rect 925 1768 945 1788
rect 1812 1805 1832 1825
rect 1656 1752 1674 1770
rect 1867 1753 1887 1773
rect 309 1582 329 1602
rect 849 1581 869 1601
rect 691 1527 711 1547
rect 904 1529 924 1549
rect 1723 1584 1743 1604
rect 1107 1398 1127 1418
rect 926 1356 946 1376
rect 1647 1397 1667 1417
rect 1488 1344 1509 1363
rect 1702 1345 1722 1365
rect 310 1170 330 1190
rect 850 1169 870 1189
rect 683 1119 703 1139
rect 905 1117 925 1137
rect 1443 1027 1467 1049
rect 1805 976 1825 996
rect 1189 790 1209 810
rect 908 750 928 770
rect 1729 789 1749 809
rect 1574 733 1593 750
rect 1784 737 1804 757
rect 292 564 312 584
rect 832 563 852 583
rect 674 509 694 529
rect 887 511 907 531
rect 1886 666 1908 684
rect 1706 566 1726 586
rect 1090 380 1110 400
rect 909 338 929 358
rect 1630 379 1650 399
rect 1474 324 1493 342
rect 1685 327 1705 347
rect 293 152 313 172
rect 833 151 853 171
rect 666 101 686 121
rect 888 99 908 119
rect 1824 260 1845 279
rect 1426 9 1450 31
rect 1991 -46 2011 -26
rect 1375 -232 1395 -212
rect 889 -268 909 -248
rect 1915 -233 1935 -213
rect 1970 -285 1990 -265
rect 273 -454 293 -434
rect 813 -455 833 -435
rect 655 -509 675 -489
rect 868 -507 888 -487
rect 1687 -452 1707 -432
rect 1071 -638 1091 -618
rect 890 -680 910 -660
rect 1611 -639 1631 -619
rect 1452 -692 1473 -673
rect 1666 -691 1686 -671
rect 274 -866 294 -846
rect 814 -867 834 -847
rect 647 -917 667 -897
rect 869 -919 889 -899
rect 1407 -1009 1431 -987
rect 1769 -1060 1789 -1040
rect 1153 -1246 1173 -1226
rect 872 -1286 892 -1266
rect 1693 -1247 1713 -1227
rect 1536 -1299 1557 -1280
rect 1748 -1299 1768 -1279
rect 256 -1472 276 -1452
rect 796 -1473 816 -1453
rect 638 -1527 658 -1507
rect 851 -1525 871 -1505
rect 1670 -1470 1690 -1450
rect 1054 -1656 1074 -1636
rect 873 -1698 893 -1678
rect 1594 -1657 1614 -1637
rect 1438 -1712 1457 -1694
rect 1649 -1709 1669 -1689
rect 257 -1884 277 -1864
rect 797 -1885 817 -1865
rect 630 -1935 650 -1915
rect 852 -1937 872 -1917
rect 1788 -1776 1809 -1757
rect 1390 -2027 1414 -2005
rect 1815 -2080 1835 -2060
rect 1199 -2266 1219 -2246
rect 852 -2304 872 -2284
rect 1739 -2267 1759 -2247
rect 1580 -2319 1603 -2297
rect 1794 -2319 1814 -2299
rect 2004 -2382 2028 -2360
rect 236 -2490 256 -2470
rect 776 -2491 796 -2471
rect 618 -2545 638 -2525
rect 831 -2543 851 -2523
rect 1650 -2488 1670 -2468
rect 1807 -2574 1829 -2556
rect 1034 -2674 1054 -2654
rect 853 -2716 873 -2696
rect 1574 -2675 1594 -2655
rect 1415 -2728 1436 -2709
rect 1629 -2727 1649 -2707
rect 237 -2902 257 -2882
rect 777 -2903 797 -2883
rect 610 -2953 630 -2933
rect 832 -2955 852 -2935
rect 1370 -3045 1394 -3023
rect 1732 -3096 1752 -3076
rect 1116 -3282 1136 -3262
rect 835 -3322 855 -3302
rect 1656 -3283 1676 -3263
rect 1501 -3339 1520 -3322
rect 1711 -3335 1731 -3315
rect 219 -3508 239 -3488
rect 759 -3509 779 -3489
rect 601 -3563 621 -3543
rect 814 -3561 834 -3541
rect 1633 -3506 1653 -3486
rect 1017 -3692 1037 -3672
rect 836 -3734 856 -3714
rect 1557 -3693 1577 -3673
rect 1401 -3748 1420 -3730
rect 1612 -3745 1632 -3725
rect 220 -3920 240 -3900
rect 760 -3921 780 -3901
rect 593 -3971 613 -3951
rect 815 -3973 835 -3953
rect 1751 -3812 1772 -3793
rect 1353 -4063 1377 -4041
<< metal1 >>
rect 958 3829 990 3830
rect 955 3824 990 3829
rect 955 3804 962 3824
rect 982 3804 990 3824
rect 955 3796 990 3804
rect 337 3638 922 3646
rect 337 3618 346 3638
rect 366 3637 922 3638
rect 366 3618 886 3637
rect 337 3617 886 3618
rect 906 3617 922 3637
rect 337 3611 922 3617
rect 956 3590 990 3796
rect 720 3583 755 3590
rect 720 3563 728 3583
rect 748 3563 755 3583
rect 720 3490 755 3563
rect 934 3585 990 3590
rect 934 3565 941 3585
rect 961 3565 990 3585
rect 934 3558 990 3565
rect 1025 3692 1055 3694
rect 1754 3692 1787 3693
rect 1025 3666 1788 3692
rect 934 3557 969 3558
rect 1025 3491 1055 3666
rect 1754 3645 1788 3666
rect 1753 3640 1788 3645
rect 1753 3620 1760 3640
rect 1780 3620 1788 3640
rect 1753 3612 1788 3620
rect 1020 3490 1055 3491
rect 719 3463 1055 3490
rect 1025 3462 1055 3463
rect 1135 3454 1720 3462
rect 1135 3434 1144 3454
rect 1164 3453 1720 3454
rect 1164 3434 1684 3453
rect 1135 3433 1684 3434
rect 1704 3433 1720 3453
rect 1135 3427 1720 3433
rect 959 3417 991 3418
rect 956 3412 991 3417
rect 956 3392 963 3412
rect 983 3392 991 3412
rect 1754 3406 1788 3612
rect 956 3384 991 3392
rect 338 3226 923 3234
rect 338 3206 347 3226
rect 367 3225 923 3226
rect 367 3206 887 3225
rect 338 3205 887 3206
rect 907 3205 923 3225
rect 338 3199 923 3205
rect 712 3175 751 3179
rect 957 3178 991 3384
rect 1520 3399 1555 3405
rect 1520 3380 1525 3399
rect 1546 3380 1555 3399
rect 1520 3371 1555 3380
rect 1732 3401 1788 3406
rect 1732 3381 1739 3401
rect 1759 3381 1788 3401
rect 1732 3374 1788 3381
rect 1732 3373 1767 3374
rect 1524 3303 1553 3371
rect 1524 3269 1870 3303
rect 712 3155 720 3175
rect 740 3155 751 3175
rect 712 3080 751 3155
rect 935 3173 991 3178
rect 935 3153 942 3173
rect 962 3153 991 3173
rect 935 3146 991 3153
rect 935 3145 970 3146
rect 1475 3085 1514 3098
rect 1475 3080 1480 3085
rect 712 3063 1480 3080
rect 1504 3080 1514 3085
rect 1504 3063 1515 3080
rect 712 3055 1515 3063
rect 714 3054 1000 3055
rect 1831 3032 1870 3269
rect 1831 3020 1842 3032
rect 1835 3012 1842 3020
rect 1862 3012 1870 3032
rect 1835 3004 1870 3012
rect 1217 2846 1802 2854
rect 1217 2826 1226 2846
rect 1246 2845 1802 2846
rect 1246 2826 1766 2845
rect 1217 2825 1766 2826
rect 1786 2825 1802 2845
rect 1217 2819 1802 2825
rect 941 2811 973 2812
rect 938 2806 973 2811
rect 938 2786 945 2806
rect 965 2786 973 2806
rect 1836 2798 1870 3004
rect 938 2778 973 2786
rect 320 2620 905 2628
rect 320 2600 329 2620
rect 349 2619 905 2620
rect 349 2600 869 2619
rect 320 2599 869 2600
rect 889 2599 905 2619
rect 320 2593 905 2599
rect 939 2572 973 2778
rect 1604 2792 1635 2798
rect 1604 2773 1609 2792
rect 1630 2773 1635 2792
rect 1604 2731 1635 2773
rect 1814 2793 1870 2798
rect 1814 2773 1821 2793
rect 1841 2773 1870 2793
rect 1814 2766 1870 2773
rect 1814 2765 1849 2766
rect 1604 2703 1943 2731
rect 703 2565 738 2572
rect 703 2545 711 2565
rect 731 2545 738 2565
rect 703 2472 738 2545
rect 917 2567 973 2572
rect 917 2547 924 2567
rect 944 2547 973 2567
rect 917 2540 973 2547
rect 1008 2674 1038 2676
rect 1737 2674 1770 2675
rect 1008 2648 1771 2674
rect 917 2539 952 2540
rect 1008 2473 1038 2648
rect 1737 2627 1771 2648
rect 1736 2622 1771 2627
rect 1736 2602 1743 2622
rect 1763 2602 1771 2622
rect 1736 2594 1771 2602
rect 1003 2472 1038 2473
rect 702 2445 1038 2472
rect 1008 2444 1038 2445
rect 1118 2436 1703 2444
rect 1118 2416 1127 2436
rect 1147 2435 1703 2436
rect 1147 2416 1667 2435
rect 1118 2415 1667 2416
rect 1687 2415 1703 2435
rect 1118 2409 1703 2415
rect 942 2399 974 2400
rect 939 2394 974 2399
rect 939 2374 946 2394
rect 966 2374 974 2394
rect 1737 2388 1771 2594
rect 939 2366 974 2374
rect 321 2208 906 2216
rect 321 2188 330 2208
rect 350 2207 906 2208
rect 350 2188 870 2207
rect 321 2187 870 2188
rect 890 2187 906 2207
rect 321 2181 906 2187
rect 695 2157 734 2161
rect 940 2160 974 2366
rect 1504 2378 1538 2386
rect 1504 2360 1511 2378
rect 1530 2360 1538 2378
rect 1504 2353 1538 2360
rect 1715 2383 1771 2388
rect 1715 2363 1722 2383
rect 1742 2363 1771 2383
rect 1715 2356 1771 2363
rect 1715 2355 1750 2356
rect 1508 2323 1537 2353
rect 1508 2315 1890 2323
rect 1508 2296 1861 2315
rect 1882 2296 1890 2315
rect 1508 2291 1890 2296
rect 695 2137 703 2157
rect 723 2137 734 2157
rect 695 2062 734 2137
rect 918 2155 974 2160
rect 918 2135 925 2155
rect 945 2135 974 2155
rect 918 2128 974 2135
rect 918 2127 953 2128
rect 1458 2067 1497 2080
rect 1458 2062 1463 2067
rect 695 2045 1463 2062
rect 1487 2062 1497 2067
rect 1487 2045 1498 2062
rect 695 2037 1498 2045
rect 697 2036 983 2037
rect 1914 2018 1943 2703
rect 1883 2015 1948 2018
rect 1881 2012 1948 2015
rect 1881 1992 1888 2012
rect 1908 1992 1948 2012
rect 1881 1985 1948 1992
rect 1881 1984 1916 1985
rect 1263 1826 1848 1834
rect 1263 1806 1272 1826
rect 1292 1825 1848 1826
rect 1292 1806 1812 1825
rect 1263 1805 1812 1806
rect 1832 1805 1848 1825
rect 1263 1799 1848 1805
rect 921 1793 953 1794
rect 918 1788 953 1793
rect 918 1768 925 1788
rect 945 1768 953 1788
rect 918 1760 953 1768
rect 300 1602 885 1610
rect 300 1582 309 1602
rect 329 1601 885 1602
rect 329 1582 849 1601
rect 300 1581 849 1582
rect 869 1581 885 1601
rect 300 1575 885 1581
rect 919 1554 953 1760
rect 1646 1770 1687 1781
rect 1882 1778 1916 1984
rect 1646 1752 1656 1770
rect 1674 1752 1687 1770
rect 1646 1744 1687 1752
rect 1860 1773 1916 1778
rect 1860 1753 1867 1773
rect 1887 1753 1916 1773
rect 1860 1746 1916 1753
rect 1860 1745 1895 1746
rect 1655 1714 1681 1744
rect 1655 1713 1993 1714
rect 1655 1677 2009 1713
rect 683 1547 718 1554
rect 683 1527 691 1547
rect 711 1527 718 1547
rect 683 1454 718 1527
rect 897 1549 953 1554
rect 897 1529 904 1549
rect 924 1529 953 1549
rect 897 1522 953 1529
rect 988 1656 1018 1658
rect 1717 1656 1750 1657
rect 988 1630 1751 1656
rect 897 1521 932 1522
rect 988 1455 1018 1630
rect 1717 1609 1751 1630
rect 1716 1604 1751 1609
rect 1716 1584 1723 1604
rect 1743 1584 1751 1604
rect 1716 1576 1751 1584
rect 983 1454 1018 1455
rect 682 1427 1018 1454
rect 988 1426 1018 1427
rect 1098 1418 1683 1426
rect 1098 1398 1107 1418
rect 1127 1417 1683 1418
rect 1127 1398 1647 1417
rect 1098 1397 1647 1398
rect 1667 1397 1683 1417
rect 1098 1391 1683 1397
rect 922 1381 954 1382
rect 919 1376 954 1381
rect 919 1356 926 1376
rect 946 1356 954 1376
rect 1717 1370 1751 1576
rect 919 1348 954 1356
rect 301 1190 886 1198
rect 301 1170 310 1190
rect 330 1189 886 1190
rect 330 1170 850 1189
rect 301 1169 850 1170
rect 870 1169 886 1189
rect 301 1163 886 1169
rect 675 1139 714 1143
rect 920 1142 954 1348
rect 1483 1363 1518 1369
rect 1483 1344 1488 1363
rect 1509 1344 1518 1363
rect 1483 1335 1518 1344
rect 1695 1365 1751 1370
rect 1695 1345 1702 1365
rect 1722 1345 1751 1365
rect 1695 1338 1751 1345
rect 1695 1337 1730 1338
rect 1487 1267 1516 1335
rect 1487 1233 1833 1267
rect 675 1119 683 1139
rect 703 1119 714 1139
rect 675 1044 714 1119
rect 898 1137 954 1142
rect 898 1117 905 1137
rect 925 1117 954 1137
rect 898 1110 954 1117
rect 898 1109 933 1110
rect 1438 1049 1477 1062
rect 1438 1044 1443 1049
rect 675 1027 1443 1044
rect 1467 1044 1477 1049
rect 1467 1027 1478 1044
rect 675 1019 1478 1027
rect 677 1018 963 1019
rect 1794 996 1833 1233
rect 1794 984 1805 996
rect 1798 976 1805 984
rect 1825 976 1833 996
rect 1798 968 1833 976
rect 1180 810 1765 818
rect 1180 790 1189 810
rect 1209 809 1765 810
rect 1209 790 1729 809
rect 1180 789 1729 790
rect 1749 789 1765 809
rect 1180 783 1765 789
rect 904 775 936 776
rect 901 770 936 775
rect 901 750 908 770
rect 928 750 936 770
rect 1799 762 1833 968
rect 901 742 936 750
rect 283 584 868 592
rect 283 564 292 584
rect 312 583 868 584
rect 312 564 832 583
rect 283 563 832 564
rect 852 563 868 583
rect 283 557 868 563
rect 902 536 936 742
rect 1565 750 1601 759
rect 1565 733 1574 750
rect 1593 733 1601 750
rect 1565 724 1601 733
rect 1777 757 1833 762
rect 1777 737 1784 757
rect 1804 737 1833 757
rect 1777 730 1833 737
rect 1777 729 1812 730
rect 1571 689 1597 724
rect 1879 689 1911 690
rect 1571 684 1911 689
rect 1571 666 1886 684
rect 1908 666 1911 684
rect 1571 661 1911 666
rect 1879 660 1911 661
rect 666 529 701 536
rect 666 509 674 529
rect 694 509 701 529
rect 666 436 701 509
rect 880 531 936 536
rect 880 511 887 531
rect 907 511 936 531
rect 880 504 936 511
rect 971 638 1001 640
rect 1700 638 1733 639
rect 971 612 1734 638
rect 880 503 915 504
rect 971 437 1001 612
rect 1700 591 1734 612
rect 1699 586 1734 591
rect 1699 566 1706 586
rect 1726 566 1734 586
rect 1699 558 1734 566
rect 966 436 1001 437
rect 665 409 1001 436
rect 971 408 1001 409
rect 1081 400 1666 408
rect 1081 380 1090 400
rect 1110 399 1666 400
rect 1110 380 1630 399
rect 1081 379 1630 380
rect 1650 379 1666 399
rect 1081 373 1666 379
rect 905 363 937 364
rect 902 358 937 363
rect 902 338 909 358
rect 929 338 937 358
rect 1700 352 1734 558
rect 902 330 937 338
rect 284 172 869 180
rect 284 152 293 172
rect 313 171 869 172
rect 313 152 833 171
rect 284 151 833 152
rect 853 151 869 171
rect 284 145 869 151
rect 658 121 697 125
rect 903 124 937 330
rect 1467 342 1501 350
rect 1467 324 1474 342
rect 1493 324 1501 342
rect 1467 317 1501 324
rect 1678 347 1734 352
rect 1678 327 1685 347
rect 1705 327 1734 347
rect 1678 320 1734 327
rect 1678 319 1713 320
rect 1471 287 1500 317
rect 1471 279 1853 287
rect 1471 260 1824 279
rect 1845 260 1853 279
rect 1471 255 1853 260
rect 658 101 666 121
rect 686 101 697 121
rect 658 26 697 101
rect 881 119 937 124
rect 881 99 888 119
rect 908 99 937 119
rect 881 92 937 99
rect 881 91 916 92
rect 1421 31 1460 44
rect 1421 26 1426 31
rect 658 9 1426 26
rect 1450 26 1460 31
rect 1450 9 1461 26
rect 658 1 1461 9
rect 660 0 946 1
rect 1982 -23 2009 1677
rect 1982 -26 2019 -23
rect 1982 -46 1991 -26
rect 2011 -46 2019 -26
rect 1982 -61 2019 -46
rect 1366 -212 1951 -204
rect 1366 -232 1375 -212
rect 1395 -213 1951 -212
rect 1395 -232 1915 -213
rect 1366 -233 1915 -232
rect 1935 -233 1951 -213
rect 1366 -239 1951 -233
rect 885 -243 917 -242
rect 882 -248 917 -243
rect 882 -268 889 -248
rect 909 -268 917 -248
rect 1985 -260 2019 -61
rect 882 -276 917 -268
rect 264 -434 849 -426
rect 264 -454 273 -434
rect 293 -435 849 -434
rect 293 -454 813 -435
rect 264 -455 813 -454
rect 833 -455 849 -435
rect 264 -461 849 -455
rect 883 -482 917 -276
rect 1963 -265 2019 -260
rect 1963 -285 1970 -265
rect 1990 -285 2019 -265
rect 1963 -292 2019 -285
rect 1963 -293 1998 -292
rect 647 -489 682 -482
rect 647 -509 655 -489
rect 675 -509 682 -489
rect 647 -582 682 -509
rect 861 -487 917 -482
rect 861 -507 868 -487
rect 888 -507 917 -487
rect 861 -514 917 -507
rect 952 -380 982 -378
rect 1681 -380 1714 -379
rect 952 -406 1715 -380
rect 861 -515 896 -514
rect 952 -581 982 -406
rect 1681 -427 1715 -406
rect 1680 -432 1715 -427
rect 1680 -452 1687 -432
rect 1707 -452 1715 -432
rect 1680 -460 1715 -452
rect 947 -582 982 -581
rect 646 -609 982 -582
rect 952 -610 982 -609
rect 1062 -618 1647 -610
rect 1062 -638 1071 -618
rect 1091 -619 1647 -618
rect 1091 -638 1611 -619
rect 1062 -639 1611 -638
rect 1631 -639 1647 -619
rect 1062 -645 1647 -639
rect 886 -655 918 -654
rect 883 -660 918 -655
rect 883 -680 890 -660
rect 910 -680 918 -660
rect 1681 -666 1715 -460
rect 883 -688 918 -680
rect 265 -846 850 -838
rect 265 -866 274 -846
rect 294 -847 850 -846
rect 294 -866 814 -847
rect 265 -867 814 -866
rect 834 -867 850 -847
rect 265 -873 850 -867
rect 639 -897 678 -893
rect 884 -894 918 -688
rect 1447 -673 1482 -667
rect 1447 -692 1452 -673
rect 1473 -692 1482 -673
rect 1447 -701 1482 -692
rect 1659 -671 1715 -666
rect 1659 -691 1666 -671
rect 1686 -691 1715 -671
rect 1659 -698 1715 -691
rect 1659 -699 1694 -698
rect 1451 -769 1480 -701
rect 1451 -803 1797 -769
rect 639 -917 647 -897
rect 667 -917 678 -897
rect 639 -992 678 -917
rect 862 -899 918 -894
rect 862 -919 869 -899
rect 889 -919 918 -899
rect 862 -926 918 -919
rect 862 -927 897 -926
rect 1402 -987 1441 -974
rect 1402 -992 1407 -987
rect 639 -1009 1407 -992
rect 1431 -992 1441 -987
rect 1431 -1009 1442 -992
rect 639 -1017 1442 -1009
rect 641 -1018 927 -1017
rect 1758 -1040 1797 -803
rect 1758 -1052 1769 -1040
rect 1762 -1060 1769 -1052
rect 1789 -1060 1797 -1040
rect 1762 -1068 1797 -1060
rect 1144 -1226 1729 -1218
rect 1144 -1246 1153 -1226
rect 1173 -1227 1729 -1226
rect 1173 -1246 1693 -1227
rect 1144 -1247 1693 -1246
rect 1713 -1247 1729 -1227
rect 1144 -1253 1729 -1247
rect 868 -1261 900 -1260
rect 865 -1266 900 -1261
rect 865 -1286 872 -1266
rect 892 -1286 900 -1266
rect 1763 -1274 1797 -1068
rect 865 -1294 900 -1286
rect 247 -1452 832 -1444
rect 247 -1472 256 -1452
rect 276 -1453 832 -1452
rect 276 -1472 796 -1453
rect 247 -1473 796 -1472
rect 816 -1473 832 -1453
rect 247 -1479 832 -1473
rect 866 -1500 900 -1294
rect 1531 -1280 1562 -1274
rect 1531 -1299 1536 -1280
rect 1557 -1299 1562 -1280
rect 1531 -1341 1562 -1299
rect 1741 -1279 1797 -1274
rect 1741 -1299 1748 -1279
rect 1768 -1299 1797 -1279
rect 1741 -1306 1797 -1299
rect 1741 -1307 1776 -1306
rect 1531 -1369 1870 -1341
rect 630 -1507 665 -1500
rect 630 -1527 638 -1507
rect 658 -1527 665 -1507
rect 630 -1600 665 -1527
rect 844 -1505 900 -1500
rect 844 -1525 851 -1505
rect 871 -1525 900 -1505
rect 844 -1532 900 -1525
rect 935 -1398 965 -1396
rect 1664 -1398 1697 -1397
rect 935 -1424 1698 -1398
rect 844 -1533 879 -1532
rect 935 -1599 965 -1424
rect 1664 -1445 1698 -1424
rect 1663 -1450 1698 -1445
rect 1663 -1470 1670 -1450
rect 1690 -1470 1698 -1450
rect 1663 -1478 1698 -1470
rect 930 -1600 965 -1599
rect 629 -1627 965 -1600
rect 935 -1628 965 -1627
rect 1045 -1636 1630 -1628
rect 1045 -1656 1054 -1636
rect 1074 -1637 1630 -1636
rect 1074 -1656 1594 -1637
rect 1045 -1657 1594 -1656
rect 1614 -1657 1630 -1637
rect 1045 -1663 1630 -1657
rect 869 -1673 901 -1672
rect 866 -1678 901 -1673
rect 866 -1698 873 -1678
rect 893 -1698 901 -1678
rect 1664 -1684 1698 -1478
rect 866 -1706 901 -1698
rect 248 -1864 833 -1856
rect 248 -1884 257 -1864
rect 277 -1865 833 -1864
rect 277 -1884 797 -1865
rect 248 -1885 797 -1884
rect 817 -1885 833 -1865
rect 248 -1891 833 -1885
rect 622 -1915 661 -1911
rect 867 -1912 901 -1706
rect 1431 -1694 1465 -1686
rect 1431 -1712 1438 -1694
rect 1457 -1712 1465 -1694
rect 1431 -1719 1465 -1712
rect 1642 -1689 1698 -1684
rect 1642 -1709 1649 -1689
rect 1669 -1709 1698 -1689
rect 1642 -1716 1698 -1709
rect 1642 -1717 1677 -1716
rect 1435 -1749 1464 -1719
rect 1435 -1757 1817 -1749
rect 1435 -1776 1788 -1757
rect 1809 -1776 1817 -1757
rect 1435 -1781 1817 -1776
rect 622 -1935 630 -1915
rect 650 -1935 661 -1915
rect 622 -2010 661 -1935
rect 845 -1917 901 -1912
rect 845 -1937 852 -1917
rect 872 -1937 901 -1917
rect 845 -1944 901 -1937
rect 845 -1945 880 -1944
rect 1385 -2005 1424 -1992
rect 1385 -2010 1390 -2005
rect 622 -2027 1390 -2010
rect 1414 -2010 1424 -2005
rect 1414 -2027 1425 -2010
rect 622 -2035 1425 -2027
rect 624 -2036 910 -2035
rect 1841 -2054 1870 -1369
rect 1810 -2057 1875 -2054
rect 1808 -2060 1875 -2057
rect 1808 -2080 1815 -2060
rect 1835 -2080 1875 -2060
rect 1808 -2087 1875 -2080
rect 1808 -2088 1843 -2087
rect 1190 -2246 1775 -2238
rect 1190 -2266 1199 -2246
rect 1219 -2247 1775 -2246
rect 1219 -2266 1739 -2247
rect 1190 -2267 1739 -2266
rect 1759 -2267 1775 -2247
rect 1190 -2273 1775 -2267
rect 848 -2279 880 -2278
rect 845 -2284 880 -2279
rect 845 -2304 852 -2284
rect 872 -2304 880 -2284
rect 845 -2312 880 -2304
rect 227 -2470 812 -2462
rect 227 -2490 236 -2470
rect 256 -2471 812 -2470
rect 256 -2490 776 -2471
rect 227 -2491 776 -2490
rect 796 -2491 812 -2471
rect 227 -2497 812 -2491
rect 846 -2518 880 -2312
rect 1575 -2297 1608 -2291
rect 1809 -2294 1843 -2088
rect 1575 -2319 1580 -2297
rect 1603 -2319 1608 -2297
rect 1575 -2328 1608 -2319
rect 1787 -2299 1843 -2294
rect 1787 -2319 1794 -2299
rect 1814 -2319 1843 -2299
rect 1787 -2326 1843 -2319
rect 1787 -2327 1822 -2326
rect 1577 -2359 1604 -2328
rect 1999 -2359 2038 -2347
rect 1577 -2360 2040 -2359
rect 1577 -2382 2004 -2360
rect 2028 -2382 2040 -2360
rect 1577 -2390 2040 -2382
rect 610 -2525 645 -2518
rect 610 -2545 618 -2525
rect 638 -2545 645 -2525
rect 610 -2618 645 -2545
rect 824 -2523 880 -2518
rect 824 -2543 831 -2523
rect 851 -2543 880 -2523
rect 824 -2550 880 -2543
rect 915 -2416 945 -2414
rect 1644 -2416 1677 -2415
rect 915 -2442 1678 -2416
rect 824 -2551 859 -2550
rect 915 -2617 945 -2442
rect 1644 -2463 1678 -2442
rect 1643 -2468 1678 -2463
rect 1643 -2488 1650 -2468
rect 1670 -2488 1678 -2468
rect 1643 -2496 1678 -2488
rect 910 -2618 945 -2617
rect 609 -2645 945 -2618
rect 915 -2646 945 -2645
rect 1025 -2654 1610 -2646
rect 1025 -2674 1034 -2654
rect 1054 -2655 1610 -2654
rect 1054 -2674 1574 -2655
rect 1025 -2675 1574 -2674
rect 1594 -2675 1610 -2655
rect 1025 -2681 1610 -2675
rect 849 -2691 881 -2690
rect 846 -2696 881 -2691
rect 846 -2716 853 -2696
rect 873 -2716 881 -2696
rect 1644 -2702 1678 -2496
rect 846 -2724 881 -2716
rect 228 -2882 813 -2874
rect 228 -2902 237 -2882
rect 257 -2883 813 -2882
rect 257 -2902 777 -2883
rect 228 -2903 777 -2902
rect 797 -2903 813 -2883
rect 228 -2909 813 -2903
rect 602 -2933 641 -2929
rect 847 -2930 881 -2724
rect 1410 -2709 1445 -2703
rect 1410 -2728 1415 -2709
rect 1436 -2728 1445 -2709
rect 1410 -2737 1445 -2728
rect 1622 -2707 1678 -2702
rect 1622 -2727 1629 -2707
rect 1649 -2727 1678 -2707
rect 1622 -2734 1678 -2727
rect 1800 -2556 1832 -2544
rect 1800 -2574 1807 -2556
rect 1829 -2574 1832 -2556
rect 1622 -2735 1657 -2734
rect 1414 -2805 1443 -2737
rect 1414 -2839 1760 -2805
rect 602 -2953 610 -2933
rect 630 -2953 641 -2933
rect 602 -3028 641 -2953
rect 825 -2935 881 -2930
rect 825 -2955 832 -2935
rect 852 -2955 881 -2935
rect 825 -2962 881 -2955
rect 825 -2963 860 -2962
rect 1365 -3023 1404 -3010
rect 1365 -3028 1370 -3023
rect 602 -3045 1370 -3028
rect 1394 -3028 1404 -3023
rect 1394 -3045 1405 -3028
rect 602 -3053 1405 -3045
rect 604 -3054 890 -3053
rect 1721 -3076 1760 -2839
rect 1721 -3088 1732 -3076
rect 1725 -3096 1732 -3088
rect 1752 -3096 1760 -3076
rect 1725 -3104 1760 -3096
rect 1107 -3262 1692 -3254
rect 1107 -3282 1116 -3262
rect 1136 -3263 1692 -3262
rect 1136 -3282 1656 -3263
rect 1107 -3283 1656 -3282
rect 1676 -3283 1692 -3263
rect 1107 -3289 1692 -3283
rect 831 -3297 863 -3296
rect 828 -3302 863 -3297
rect 828 -3322 835 -3302
rect 855 -3322 863 -3302
rect 1726 -3310 1760 -3104
rect 828 -3330 863 -3322
rect 210 -3488 795 -3480
rect 210 -3508 219 -3488
rect 239 -3489 795 -3488
rect 239 -3508 759 -3489
rect 210 -3509 759 -3508
rect 779 -3509 795 -3489
rect 210 -3515 795 -3509
rect 829 -3536 863 -3330
rect 1492 -3322 1528 -3313
rect 1492 -3339 1501 -3322
rect 1520 -3339 1528 -3322
rect 1492 -3348 1528 -3339
rect 1704 -3315 1760 -3310
rect 1704 -3335 1711 -3315
rect 1731 -3335 1760 -3315
rect 1704 -3342 1760 -3335
rect 1704 -3343 1739 -3342
rect 1498 -3383 1524 -3348
rect 1800 -3383 1832 -2574
rect 1498 -3411 1832 -3383
rect 593 -3543 628 -3536
rect 593 -3563 601 -3543
rect 621 -3563 628 -3543
rect 593 -3636 628 -3563
rect 807 -3541 863 -3536
rect 807 -3561 814 -3541
rect 834 -3561 863 -3541
rect 807 -3568 863 -3561
rect 898 -3434 928 -3432
rect 1627 -3434 1660 -3433
rect 898 -3460 1661 -3434
rect 807 -3569 842 -3568
rect 898 -3635 928 -3460
rect 1627 -3481 1661 -3460
rect 1626 -3486 1661 -3481
rect 1626 -3506 1633 -3486
rect 1653 -3506 1661 -3486
rect 1626 -3514 1661 -3506
rect 893 -3636 928 -3635
rect 592 -3663 928 -3636
rect 898 -3664 928 -3663
rect 1008 -3672 1593 -3664
rect 1008 -3692 1017 -3672
rect 1037 -3673 1593 -3672
rect 1037 -3692 1557 -3673
rect 1008 -3693 1557 -3692
rect 1577 -3693 1593 -3673
rect 1008 -3699 1593 -3693
rect 832 -3709 864 -3708
rect 829 -3714 864 -3709
rect 829 -3734 836 -3714
rect 856 -3734 864 -3714
rect 1627 -3720 1661 -3514
rect 829 -3742 864 -3734
rect 211 -3900 796 -3892
rect 211 -3920 220 -3900
rect 240 -3901 796 -3900
rect 240 -3920 760 -3901
rect 211 -3921 760 -3920
rect 780 -3921 796 -3901
rect 211 -3927 796 -3921
rect 585 -3951 624 -3947
rect 830 -3948 864 -3742
rect 1394 -3730 1428 -3722
rect 1394 -3748 1401 -3730
rect 1420 -3748 1428 -3730
rect 1394 -3755 1428 -3748
rect 1605 -3725 1661 -3720
rect 1605 -3745 1612 -3725
rect 1632 -3745 1661 -3725
rect 1605 -3752 1661 -3745
rect 1605 -3753 1640 -3752
rect 1398 -3785 1427 -3755
rect 1398 -3793 1780 -3785
rect 1398 -3812 1751 -3793
rect 1772 -3812 1780 -3793
rect 1398 -3817 1780 -3812
rect 585 -3971 593 -3951
rect 613 -3971 624 -3951
rect 585 -4046 624 -3971
rect 808 -3953 864 -3948
rect 808 -3973 815 -3953
rect 835 -3973 864 -3953
rect 808 -3980 864 -3973
rect 808 -3981 843 -3980
rect 1348 -4041 1387 -4028
rect 1348 -4046 1353 -4041
rect 585 -4063 1353 -4046
rect 1377 -4046 1387 -4041
rect 1377 -4063 1388 -4046
rect 585 -4071 1388 -4063
rect 587 -4072 873 -4071
<< labels >>
rlabel locali 300 3620 322 3635 1 d0
rlabel locali 354 3808 383 3814 1 vdd
rlabel locali 351 3509 380 3515 1 gnd
rlabel space 457 3527 486 3536 1 gnd
rlabel nwell 489 3785 512 3788 1 vdd
rlabel locali 301 3208 323 3223 1 d0
rlabel locali 355 3396 384 3402 1 vdd
rlabel locali 352 3097 381 3103 1 gnd
rlabel space 458 3115 487 3124 1 gnd
rlabel nwell 490 3373 513 3376 1 vdd
rlabel locali 191 4053 215 4083 1 vref
rlabel locali 283 2602 305 2617 1 d0
rlabel locali 337 2790 366 2796 1 vdd
rlabel locali 334 2491 363 2497 1 gnd
rlabel space 440 2509 469 2518 1 gnd
rlabel nwell 472 2767 495 2770 1 vdd
rlabel locali 284 2190 306 2205 1 d0
rlabel locali 338 2378 367 2384 1 vdd
rlabel locali 335 2079 364 2085 1 gnd
rlabel space 441 2097 470 2106 1 gnd
rlabel nwell 473 2355 496 2358 1 vdd
rlabel locali 1152 3624 1181 3630 1 vdd
rlabel locali 1149 3325 1178 3331 1 gnd
rlabel space 1255 3343 1284 3352 1 gnd
rlabel nwell 1287 3601 1310 3604 1 vdd
rlabel locali 1092 3432 1114 3449 1 d1
rlabel locali 1135 2606 1164 2612 1 vdd
rlabel locali 1132 2307 1161 2313 1 gnd
rlabel space 1238 2325 1267 2334 1 gnd
rlabel nwell 1270 2583 1293 2586 1 vdd
rlabel locali 1075 2414 1097 2431 1 d1
rlabel locali 1234 3016 1263 3022 1 vdd
rlabel locali 1231 2717 1260 2723 1 gnd
rlabel space 1337 2735 1366 2744 1 gnd
rlabel nwell 1369 2993 1392 2996 1 vdd
rlabel locali 1176 2824 1196 2848 1 d2
rlabel locali 263 1584 285 1599 1 d0
rlabel locali 317 1772 346 1778 1 vdd
rlabel locali 314 1473 343 1479 1 gnd
rlabel space 420 1491 449 1500 1 gnd
rlabel nwell 452 1749 475 1752 1 vdd
rlabel locali 264 1172 286 1187 1 d0
rlabel locali 318 1360 347 1366 1 vdd
rlabel locali 315 1061 344 1067 1 gnd
rlabel space 421 1079 450 1088 1 gnd
rlabel nwell 453 1337 476 1340 1 vdd
rlabel locali 246 566 268 581 1 d0
rlabel locali 300 754 329 760 1 vdd
rlabel locali 297 455 326 461 1 gnd
rlabel space 403 473 432 482 1 gnd
rlabel nwell 435 731 458 734 1 vdd
rlabel locali 247 154 269 169 1 d0
rlabel locali 301 342 330 348 1 vdd
rlabel locali 298 43 327 49 1 gnd
rlabel space 404 61 433 70 1 gnd
rlabel nwell 436 319 459 322 1 vdd
rlabel locali 1115 1588 1144 1594 1 vdd
rlabel locali 1112 1289 1141 1295 1 gnd
rlabel space 1218 1307 1247 1316 1 gnd
rlabel nwell 1250 1565 1273 1568 1 vdd
rlabel locali 1055 1396 1077 1413 1 d1
rlabel locali 1098 570 1127 576 1 vdd
rlabel locali 1095 271 1124 277 1 gnd
rlabel space 1201 289 1230 298 1 gnd
rlabel nwell 1233 547 1256 550 1 vdd
rlabel locali 1038 378 1060 395 1 d1
rlabel locali 1197 980 1226 986 1 vdd
rlabel locali 1194 681 1223 687 1 gnd
rlabel space 1300 699 1329 708 1 gnd
rlabel nwell 1332 957 1355 960 1 vdd
rlabel locali 1139 788 1159 812 1 d2
rlabel locali 1280 1996 1309 2002 1 vdd
rlabel locali 1277 1697 1306 1703 1 gnd
rlabel space 1383 1715 1412 1724 1 gnd
rlabel nwell 1415 1973 1438 1976 1 vdd
rlabel locali 1224 1810 1244 1823 1 d3
rlabel locali 227 -452 249 -437 1 d0
rlabel locali 281 -264 310 -258 1 vdd
rlabel locali 278 -563 307 -557 1 gnd
rlabel space 384 -545 413 -536 1 gnd
rlabel nwell 416 -287 439 -284 1 vdd
rlabel locali 228 -864 250 -849 1 d0
rlabel locali 282 -676 311 -670 1 vdd
rlabel locali 279 -975 308 -969 1 gnd
rlabel space 385 -957 414 -948 1 gnd
rlabel nwell 417 -699 440 -696 1 vdd
rlabel locali 210 -1470 232 -1455 1 d0
rlabel locali 264 -1282 293 -1276 1 vdd
rlabel locali 261 -1581 290 -1575 1 gnd
rlabel space 367 -1563 396 -1554 1 gnd
rlabel nwell 399 -1305 422 -1302 1 vdd
rlabel locali 211 -1882 233 -1867 1 d0
rlabel locali 265 -1694 294 -1688 1 vdd
rlabel locali 262 -1993 291 -1987 1 gnd
rlabel space 368 -1975 397 -1966 1 gnd
rlabel nwell 400 -1717 423 -1714 1 vdd
rlabel locali 1079 -448 1108 -442 1 vdd
rlabel locali 1076 -747 1105 -741 1 gnd
rlabel space 1182 -729 1211 -720 1 gnd
rlabel nwell 1214 -471 1237 -468 1 vdd
rlabel locali 1019 -640 1041 -623 1 d1
rlabel locali 1062 -1466 1091 -1460 1 vdd
rlabel locali 1059 -1765 1088 -1759 1 gnd
rlabel space 1165 -1747 1194 -1738 1 gnd
rlabel nwell 1197 -1489 1220 -1486 1 vdd
rlabel locali 1002 -1658 1024 -1641 1 d1
rlabel locali 1161 -1056 1190 -1050 1 vdd
rlabel locali 1158 -1355 1187 -1349 1 gnd
rlabel space 1264 -1337 1293 -1328 1 gnd
rlabel nwell 1296 -1079 1319 -1076 1 vdd
rlabel locali 1103 -1248 1123 -1224 1 d2
rlabel locali 190 -2488 212 -2473 1 d0
rlabel locali 244 -2300 273 -2294 1 vdd
rlabel locali 241 -2599 270 -2593 1 gnd
rlabel space 347 -2581 376 -2572 1 gnd
rlabel nwell 379 -2323 402 -2320 1 vdd
rlabel locali 191 -2900 213 -2885 1 d0
rlabel locali 245 -2712 274 -2706 1 vdd
rlabel locali 242 -3011 271 -3005 1 gnd
rlabel space 348 -2993 377 -2984 1 gnd
rlabel nwell 380 -2735 403 -2732 1 vdd
rlabel locali 173 -3506 195 -3491 1 d0
rlabel locali 227 -3318 256 -3312 1 vdd
rlabel locali 224 -3617 253 -3611 1 gnd
rlabel space 330 -3599 359 -3590 1 gnd
rlabel nwell 362 -3341 385 -3338 1 vdd
rlabel locali 174 -3918 196 -3903 1 d0
rlabel locali 228 -3730 257 -3724 1 vdd
rlabel locali 225 -4029 254 -4023 1 gnd
rlabel space 331 -4011 360 -4002 1 gnd
rlabel nwell 363 -3753 386 -3750 1 vdd
rlabel locali 40 -4030 68 -4012 1 gnd
rlabel locali 1042 -2484 1071 -2478 1 vdd
rlabel locali 1039 -2783 1068 -2777 1 gnd
rlabel space 1145 -2765 1174 -2756 1 gnd
rlabel nwell 1177 -2507 1200 -2504 1 vdd
rlabel locali 982 -2676 1004 -2659 1 d1
rlabel locali 1025 -3502 1054 -3496 1 vdd
rlabel locali 1022 -3801 1051 -3795 1 gnd
rlabel space 1128 -3783 1157 -3774 1 gnd
rlabel nwell 1160 -3525 1183 -3522 1 vdd
rlabel locali 965 -3694 987 -3677 1 d1
rlabel locali 1124 -3092 1153 -3086 1 vdd
rlabel locali 1121 -3391 1150 -3385 1 gnd
rlabel space 1227 -3373 1256 -3364 1 gnd
rlabel nwell 1259 -3115 1282 -3112 1 vdd
rlabel locali 1066 -3284 1086 -3260 1 d2
rlabel locali 1207 -2076 1236 -2070 1 vdd
rlabel locali 1204 -2375 1233 -2369 1 gnd
rlabel space 1310 -2357 1339 -2348 1 gnd
rlabel nwell 1342 -2099 1365 -2096 1 vdd
rlabel locali 1151 -2262 1171 -2249 1 d3
rlabel locali 1383 -42 1412 -36 1 vdd
rlabel locali 1380 -341 1409 -335 1 gnd
rlabel space 1486 -323 1515 -314 1 gnd
rlabel nwell 1518 -65 1541 -62 1 vdd
rlabel locali 1756 -195 1778 -180 1 vout
rlabel locali 1329 -232 1348 -215 1 d4
<< end >>

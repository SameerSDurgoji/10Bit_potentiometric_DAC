* SPICE3 file created from switchfinal.ext - technology: sky130A

.option scale=10000u

X0 a_1285_n167# d1 vout SUB sky130_fd_pr__nfet_01v8 w=42 l=50
X1 a_1161_n286# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=42 l=50
X2 vout a_1161_n286# a_1285_n167# vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X3 vout a_1161_n286# a_1280_n286# SUB sky130_fd_pr__nfet_01v8 w=42 l=50
X4 a_1280_n286# d1 vout vdd sky130_fd_pr__pfet_01v8 w=100 l=50
X5 a_1161_n286# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=100 l=50

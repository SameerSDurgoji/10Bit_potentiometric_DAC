* SPICE3 file created from 8bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_9437_6234# a_9219_6234# a_8956_6146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 a_4091_57# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2 a_4517_2569# a_4519_2862# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3 a_9365_1750# a_9147_1750# a_8876_1856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4 vdd d2 a_2793_5845# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5 a_1659_6433# a_1441_6433# a_1565_6552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6 a_1404_935# a_1186_935# a_606_1119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7 a_3401_4048# a_3654_4035# a_2599_4409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_2635_6445# d0 a_3437_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9 a_4970_1132# a_4752_1132# a_4495_1227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 a_13275_3806# a_13277_3905# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X11 a_660_4173# d1 a_1446_3500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 gnd d1 a_7276_7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_623_2137# a_405_2137# a_142_2049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X14 gnd d4 a_11312_4856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_13729_1763# a_13511_1763# a_13238_1770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_6864_4012# d1 a_6946_3404# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 a_12215_8145# a_12468_8132# a_11413_8506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_10218_5032# a_10000_5032# a_9420_5216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X19 a_679_5191# a_461_5191# a_204_5286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X20 a_7710_1419# a_7963_1406# a_6913_1191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X21 a_116_714# d0 a_607_707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X22 a_4555_4898# a_4562_5116# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X23 a_13802_5835# a_13584_5835# a_13311_5842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_12951_82# d6 a_8658_81# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X25 a_1322_3381# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X26 gnd d0 a_8000_3442# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_14381_6063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X28 a_8982_7347# d0 a_9457_7252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_3359_2601# a_3363_2424# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X30 a_14582_5045# a_14364_5045# a_13785_4817# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X31 a_7834_8310# a_7838_8133# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X32 a_5883_7585# d2 a_5929_6565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_153_2556# a_155_2849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X34 a_3397_4225# a_3654_4035# a_2599_4409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X35 a_9239_7252# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X36 a_16524_5516# a_16777_5503# a_15727_5288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X37 a_4879_8258# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 gnd d0 a_16759_4073# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 vdd d1 a_7276_7286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X40 a_4790_2756# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X41 a_168_3250# d0 a_643_3155# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X42 a_8911_3793# a_8913_3892# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X43 a_6864_4012# d1 a_6950_3227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X44 a_8930_4811# a_8932_4910# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X45 a_12211_8322# a_12468_8132# a_11413_8506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X46 a_8889_2257# a_8894_2581# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X47 a_13260_2887# d0 a_13749_2781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X48 a_425_3155# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X49 gnd d1 a_2875_5237# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X50 a_13340_7177# a_13346_7360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X51 a_6930_2209# a_7183_2196# a_6831_1799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 vdd d0 a_16795_6109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X53 a_9981_4014# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X54 a_13267_3105# d0 a_13748_3193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X55 a_5856_2493# a_5686_3394# a_5810_3513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X56 vdd d0 a_8000_3442# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X57 a_499_6815# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X58 a_3343_1171# a_3600_981# a_2545_1355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X59 a_13548_3799# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X60 a_16489_3068# a_16484_3657# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X61 a_13604_6853# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X62 a_13748_3193# d1 a_14546_3009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X63 a_7838_8133# a_7833_8722# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X64 a_14328_3009# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X65 a_7784_5079# a_8037_5066# a_6982_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X66 a_9474_8270# a_9256_8270# a_8993_8182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X67 vdd d0 a_16759_4073# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X68 vdd d3 a_15852_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X69 a_14670_6590# a_14500_7491# a_14624_7610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X70 a_4210_57# a_5966_144# a_6085_144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X71 gnd d0 a_12358_2024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_9129_1144# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X73 vdd d1 a_15944_3239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X74 a_4499_1844# a_4506_2062# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X75 a_660_4173# a_442_4173# a_179_4085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X76 a_13311_5842# a_13313_5941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X77 a_8883_2074# d0 a_9364_2162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X78 a_9202_5216# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_198_5103# a_204_5286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X80 gnd d0 a_3636_3429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X81 a_10187_3525# a_9981_4014# a_9401_4198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X82 a_2676_8304# a_2929_8291# a_2577_7894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X83 a_8976_7164# a_8982_7347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X84 a_3346_1406# a_3360_2189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X85 a_10109_2386# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X86 a_13765_4211# a_13547_4211# a_13290_4306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X87 a_10260_7597# a_10054_8086# a_9474_8270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X88 a_9347_1144# a_9129_1144# a_8872_1239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X89 a_215_6121# a_221_6304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X90 a_7780_5256# a_8037_5066# a_6982_5440# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X91 a_10228_2386# a_10026_1370# a_10145_960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_15723_5465# d0 a_16521_5281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 a_10182_6458# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 a_14551_3538# a_14345_4027# a_13766_3799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X95 a_9420_5216# a_9202_5216# a_8945_5311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X96 a_9437_6234# d1 a_10223_5561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X97 a_7820_7527# a_7834_8310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X98 a_6900_6048# a_7157_5858# a_6854_7068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X99 gnd d0 a_12450_7526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X100 a_16505_4498# a_16758_4485# a_15708_4270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_11235_6903# a_11488_6890# a_11059_4869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 gnd d0 a_3727_8107# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X103 vdd d0 a_12358_2024# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X104 a_8874_1757# a_8876_1856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X105 gnd a_16831_8557# a_15781_8342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X106 vdd d0 a_12414_5078# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X107 a_10400_6458# a_10182_6458# a_10306_6577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X108 a_8962_6329# a_8967_6653# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X109 gnd d1 a_2839_3201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 a_16506_4086# a_16501_4675# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X111 gnd d1 a_2856_4219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X112 a_7837_8545# a_8090_8532# a_7040_8317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X113 a_14691_2399# a_14473_2399# a_14592_2399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X114 gnd d1 a_2912_7273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X115 a_10462_156# d5 a_10561_156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X116 a_1602_131# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 a_8896_2874# d0 a_9385_2768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X118 a_2562_2373# d0 a_3364_2012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X119 a_4210_57# d6 a_4309_57# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X120 a_16489_3068# a_16742_3055# a_15687_3429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X121 a_5061_5810# a_4843_5810# a_4572_5916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X122 vdd d0 a_12450_7526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X123 a_6941_7907# a_7194_7894# a_6858_6891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X124 a_7765_4061# a_8018_4048# a_6963_4422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X125 a_16501_4675# a_16758_4485# a_15708_4270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X126 a_9240_6840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X127 a_4789_3168# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X128 a_6090_263# a_5908_4408# a_5950_2374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X129 vdd d4 a_6935_4844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X130 a_4862_7240# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X131 a_9130_732# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X132 a_2314_5021# d3 a_2421_2806# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X133 a_12177_6521# a_12194_7304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X134 a_14509_973# a_14291_973# a_13712_745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 a_12104_2449# a_12357_2436# a_11307_2221# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_11055_5046# d3 a_11158_3008# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 a_5929_6565# a_5759_7466# a_5878_7056# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X138 a_12160_5503# a_12413_5490# a_11363_5275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_7833_8722# a_8090_8532# a_7040_8317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X140 gnd d0 a_12395_4060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X141 a_243_7840# d0 a_734_7833# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X142 a_9166_3180# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X143 vdd d1 a_2912_7273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X144 a_7743_3632# a_7747_3455# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X145 a_4605_7335# d0 a_5080_7240# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X146 a_16485_3245# a_16742_3055# a_15687_3429# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X147 a_2500_3999# d1 a_2586_3214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X148 a_12215_8145# a_12210_8734# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X149 a_9402_3786# a_9184_3786# a_8911_3793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X150 a_15605_4037# a_15862_3847# a_15526_2844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X151 a_2536_6035# a_2793_5845# a_2490_7055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X152 a_6831_1799# d1 a_6926_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 a_4570_5817# a_4572_5916# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X154 a_15704_4447# d0 a_16502_4263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X155 a_9401_4198# a_9183_4198# a_8926_4293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X156 a_2545_1355# d0 a_3347_994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X157 a_3360_2189# a_3364_2012# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X158 a_5098_7846# d1 a_5883_7585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X159 a_7728_2025# a_7981_2012# a_6926_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X160 a_9927_960# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X161 a_12100_2626# a_12357_2436# a_11307_2221# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X162 a_5044_4792# d1 a_5841_5020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X163 a_11314_8096# d1 a_11400_7311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X164 a_4609_7952# a_4616_8170# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X165 a_4987_2150# d1 a_5773_1477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_5604_4002# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X167 a_14582_5045# d2 a_14665_6471# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X168 vdd d0 a_12395_4060# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X169 a_1487_2361# d3 a_1586_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X170 a_6982_5440# d0 a_7780_5256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X171 a_8949_5928# d0 a_9438_5822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X172 a_15645_5896# d1 a_15740_6483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 a_1659_6433# d4 a_1726_250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X174 a_1560_6433# a_1358_5417# a_1477_5007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X175 a_135_1831# d0 a_624_1725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X176 a_15704_4447# d0 a_16506_4086# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X177 a_12084_1196# a_12341_1006# a_11286_1380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X178 a_5732_2374# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X179 a_7724_2202# a_7981_2012# a_6926_2386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X180 a_3457_7102# a_3710_7089# a_2655_7463# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X181 a_3364_2012# a_3359_2601# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X182 a_13566_5229# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X183 a_11204_1988# a_11461_1798# a_11158_3008# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X184 a_7711_1007# a_7706_1596# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X185 a_11303_2398# d0 a_12101_2214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X186 a_8658_81# a_12832_82# a_10561_156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X187 a_5908_4408# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X188 a_14670_6590# d3 a_14764_6471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X189 a_6982_5440# d0 a_7784_5079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X190 a_10150_1489# a_9944_1978# a_9365_1750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X191 a_14546_6471# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X192 a_16538_6299# a_16795_6109# a_15740_6483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X193 a_13784_5229# a_13566_5229# a_13309_5324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X194 a_7784_5079# a_7779_5668# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X195 a_6854_7068# d2 a_6904_5871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X196 a_11327_3239# d0 a_12120_3644# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X197 a_6858_6891# a_7111_6878# a_6682_4857# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X198 a_11400_7311# d0 a_12193_7716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_3433_6261# a_3437_6084# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 a_10136_7478# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X201 a_7040_8317# d0 a_7833_8722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X202 a_2573_8071# a_2830_7881# a_2494_6878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X203 a_3379_3619# a_3383_3442# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X204 a_11303_2398# d0 a_12105_2037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X205 a_2549_1178# a_2802_1165# a_2463_1963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X206 a_14691_2399# d4 a_14831_288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X207 gnd d0 a_8074_7102# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X208 gnd d1 a_15944_3239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X209 vdd d0 a_3726_8519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X210 a_185_4268# a_189_4786# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X211 a_6858_6891# d2 a_6937_8084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X212 a_4519_2862# d0 a_5008_2756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X213 a_6946_3404# d0 a_7744_3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 gnd d0 a_12430_6508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_1726_250# d5 a_1820_131# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X216 a_13838_8283# d1 a_14624_7610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X217 a_14514_1502# a_14308_1991# a_13728_2175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X218 a_7036_8494# a_7293_8304# a_6941_7907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X219 a_11363_5275# a_11616_5262# a_11277_6060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X220 a_11327_3239# d0 a_12124_3467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X221 a_5805_2984# a_5587_2984# a_5008_2756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 a_3342_1583# a_3599_1393# a_2549_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X223 a_13284_4123# a_13290_4306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X224 a_11400_7311# d0 a_12197_7539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X225 a_7040_8317# d0 a_7837_8545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X226 vdd d0 a_3637_3017# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X227 a_2545_1355# a_2802_1165# a_2463_1963# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X228 a_228_6921# a_235_7139# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X229 gnd d0 a_12341_1006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X230 a_5677_8074# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X231 a_443_3761# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X232 a_5966_144# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X233 gnd d0 a_12414_5078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X234 a_2467_1786# d1 a_2562_2373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X235 a_644_2743# a_426_2743# a_153_2556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X236 a_8539_81# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X237 a_13766_3799# a_13548_3799# a_13275_3806# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X238 a_6946_3404# d0 a_7748_3043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X239 a_11359_5452# a_11616_5262# a_11277_6060# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X240 a_10255_7068# a_10037_7068# a_9457_7252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X241 a_5883_7585# a_5677_8074# a_5097_8258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X242 a_162_3067# a_168_3250# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X243 a_680_4779# d1 a_1477_5007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X244 a_13749_2781# a_13531_2781# a_13260_2887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X245 a_2490_7055# d2 a_2536_6035# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_13712_745# a_13494_745# a_13223_851# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X247 a_204_5286# d0 a_679_5191# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 a_3396_4637# a_3400_4460# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X249 a_11281_5883# d1 a_11376_6470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X250 a_3474_8120# a_3469_8709# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X251 a_13350_7977# a_13357_8195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X252 a_13253_2270# d0 a_13728_2175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X253 a_4843_5810# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X254 a_221_6304# d0 a_696_6209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X255 a_235_7139# a_241_7322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X256 a_4532_3263# a_4534_3781# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X257 vdd d0 a_16777_5503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X258 a_10327_2386# d4 a_10467_275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X259 a_9147_1750# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 a_16502_4263# a_16506_4086# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X261 a_5623_5020# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X262 a_10561_156# a_10343_156# a_10467_275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X263 a_2467_1786# d1 a_2566_2196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X264 a_15423_4882# a_15676_4869# a_14826_169# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X265 a_14463_5455# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X266 a_148_2232# a_153_2556# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X267 a_9220_5822# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X268 a_4605_7335# a_4607_7853# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X269 a_4769_2150# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X270 vdd d1 a_7166_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X271 a_1276_6025# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_5851_2374# d3 a_5950_2374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X273 vdd d2 a_11534_5870# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X274 a_14308_1991# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 a_1514_7043# d2 a_1565_6552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X276 a_13247_2087# a_13253_2270# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X277 a_11281_5883# d1 a_11380_6293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X278 a_1482_5536# a_1276_6025# a_696_6209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X279 a_15595_7093# d2 a_15645_5896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X280 a_3379_3619# a_3636_3429# a_2586_3214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X281 a_8986_7964# a_8993_8182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X282 a_16525_5104# a_16520_5693# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X283 a_14624_7610# d2 a_14670_6590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X284 a_6682_4857# d3 a_6854_7068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 vdd d0 a_16722_2037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X286 gnd d0 a_8090_8532# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X287 a_14587_5574# a_14381_6063# a_13802_5835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X288 a_8911_3793# d0 a_9402_3786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X289 a_661_3761# d1 a_1446_3500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X290 a_14831_288# a_14649_4433# a_14764_6471# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X291 a_9384_3180# a_9166_3180# a_8909_3275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X292 a_4807_3774# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X293 a_2494_6878# d2 a_2573_8071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X294 a_7711_1007# a_7964_994# a_6909_1368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X295 a_185_4268# d0 a_660_4173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_8883_2074# a_8889_2257# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X297 a_9458_6840# a_9240_6840# a_8969_6946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X298 a_5008_2756# a_4790_2756# a_4517_2569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X299 gnd d0 a_8001_3030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X300 a_4880_7846# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X301 a_9474_8270# d1 a_10260_7597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X302 a_16465_2227# a_16469_2050# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X303 a_1409_1464# d2 a_1487_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X304 vdd d0 a_16741_3467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X305 gnd d0 a_7963_1406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X306 a_2603_4232# d0 a_3400_4460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X307 a_515_8245# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X308 a_4590_6641# a_4592_6934# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X309 a_13748_3193# a_13530_3193# a_13267_3105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 a_3380_3207# a_3384_3030# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X311 a_5660_7056# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X312 a_16525_5104# a_16778_5091# a_15723_5465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X313 a_716_7227# a_498_7227# a_235_7139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X314 vdd d0 a_8090_8532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X315 a_8939_5128# d0 a_9420_5216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X316 a_5841_5020# d2 a_5924_6446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X317 a_11380_6293# d0 a_12173_6698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 a_13821_7265# a_13603_7265# a_13340_7177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X319 a_10223_5561# d2 a_10301_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X320 a_5097_8258# a_4879_8258# a_4616_8170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X321 a_13320_6159# a_13326_6342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X322 a_14418_8099# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X323 a_10301_6458# d3 a_10400_6458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X324 a_15654_1216# d0 a_16447_1621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 a_125_1031# d0 a_606_1119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X326 a_2504_3822# a_2757_3809# a_2421_2806# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X327 vdd d0 a_8001_3030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X328 a_8949_5928# a_8956_6146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X329 a_14597_2518# d3 a_14691_2399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X330 vdd d1 a_15961_4257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X331 gnd d2 a_7084_1786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X332 a_11286_1380# d0 a_12084_1196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X333 gnd d3 a_2674_2793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X334 vdd d1 a_16034_8329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X335 a_9219_6234# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_4506_2062# d0 a_4987_2150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X337 a_13294_4824# d0 a_13785_4817# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X338 vdd d0 a_12340_1418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X339 gnd d0 a_3709_7501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 a_2536_6035# d1 a_2622_5250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X341 a_1186_935# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X342 a_4570_5817# d0 a_5061_5810# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X343 gnd d0 a_3726_8519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X344 a_5929_6565# d3 a_6023_6446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X345 a_4770_1738# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X346 gnd d4 a_2571_4831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X347 vdd d0 a_12413_5490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X348 a_16464_2639# a_16721_2449# a_15671_2234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X349 a_243_7840# a_245_7939# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X350 a_4752_1132# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X351 a_7023_7299# a_7276_7286# a_6937_8084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X352 a_2314_5021# a_2571_4831# a_1721_131# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X353 a_9437_6234# a_9219_6234# a_8962_6329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X354 a_405_2137# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_12087_1431# a_12101_2214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X356 a_11059_4869# a_11312_4856# a_10462_156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X357 a_461_5191# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X358 a_13510_2175# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X359 a_12173_6698# a_12177_6521# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X360 a_15654_1216# d0 a_16451_1444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X361 a_13258_2594# a_13260_2887# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X362 vdd d2 a_7084_1786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X363 gnd d0 a_3637_3017# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X364 a_13584_5835# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_13346_7360# a_13348_7878# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X366 a_623_2137# a_405_2137# a_148_2232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X367 a_13729_1763# a_13511_1763# a_13240_1869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X368 gnd d1 a_2929_8291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X369 a_2582_3391# a_2839_3201# a_2500_3999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X370 a_14364_5045# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X371 a_697_5797# a_479_5797# a_208_5903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X372 a_1820_131# a_1602_131# a_1721_131# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X373 a_13802_5835# a_13584_5835# a_13313_5941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X374 vdd d2 a_15898_5883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X375 gnd d0 a_12451_7114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X376 a_14509_973# a_14291_973# a_13711_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X377 a_16506_4086# a_16759_4073# a_15704_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X378 a_8986_7964# d0 a_9475_7858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X379 a_8920_4110# d0 a_9401_4198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X380 a_7019_7476# a_7276_7286# a_6937_8084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X381 a_8976_7164# d0 a_9457_7252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X382 a_716_7227# d1 a_1514_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X383 a_16579_8158# a_16832_8145# a_15777_8519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X384 a_14582_5045# a_14364_5045# a_13784_5229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X385 a_5878_7056# d2 a_5929_6565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X386 a_15522_3021# d2 a_15572_1824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X387 vdd d4 a_15676_4869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X388 a_389_707# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X389 a_6941_7907# d1 a_7036_8494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X390 a_4879_8258# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X391 a_7838_8133# a_8091_8120# a_7036_8494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_5686_3394# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X393 a_7797_6274# a_7801_6097# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X394 a_162_3067# d0 a_643_3155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X395 vdd d2 a_2757_3809# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X396 a_2622_5250# d0 a_3415_5655# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 gnd d2 a_11498_3834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X398 gnd d2 a_11461_1798# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X399 a_14500_7491# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X400 a_3347_994# a_3600_981# a_2545_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_13275_3806# d0 a_13766_3799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X402 a_9256_8270# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X403 vdd d0 a_12451_7114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X404 a_16502_4263# a_16759_4073# a_15704_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X405 gnd d1 a_7166_1178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X406 a_2504_3822# d1 a_2603_4232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X407 a_2577_7894# d1 a_2676_8304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X408 a_16575_8335# a_16832_8145# a_15777_8519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X409 a_13749_2781# d1 a_14546_3009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X410 a_8658_81# d7 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X411 a_12160_5503# a_12174_6286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X412 a_15526_2844# d2 a_15605_4037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X413 a_12105_2037# a_12358_2024# a_11303_2398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X414 a_1519_7572# a_1313_8061# a_734_7833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X415 a_7834_8310# a_8091_8120# a_7036_8494# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X416 a_15671_2234# a_15924_2221# a_15572_1824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_5080_7240# a_4862_7240# a_4605_7335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X418 a_16579_8158# a_16574_8747# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X419 gnd d1 a_15980_5275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X420 a_3383_3442# a_3636_3429# a_2586_3214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X421 a_2622_5250# d0 a_3419_5478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X422 a_8872_1239# d0 a_9347_1144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X423 a_15691_3252# d0 a_16488_3480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X424 a_10017_6050# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X425 a_5773_1477# d2 a_5851_2374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X426 a_4210_57# a_5966_144# a_6090_263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X427 a_4482_826# a_4489_1044# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X428 a_10054_8086# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X429 a_9129_1144# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X430 a_660_4173# a_442_4173# a_185_4268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X431 a_9202_5216# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X432 gnd d0 a_16722_2037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X433 a_3415_5655# a_3419_5478# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X434 vdd d2 a_15862_3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X435 a_12101_2214# a_12358_2024# a_11303_2398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X436 a_3474_8120# a_3727_8107# a_2672_8481# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X437 a_1820_131# d6 a_4309_57# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X438 a_4987_2150# a_4769_2150# a_4512_2245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X439 a_12157_5268# a_12414_5078# a_11359_5452# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X440 a_11327_3239# a_11580_3226# a_11241_4024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 a_10182_6458# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X442 a_15667_2411# a_15924_2221# a_15572_1824# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X443 a_14551_3538# a_14345_4027# a_13765_4211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X444 a_12174_6286# a_12431_6096# a_11376_6470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X445 vdd d1 a_15980_5275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X446 a_14473_2399# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X447 a_5044_4792# a_4826_4792# a_4555_4898# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X448 a_6023_6446# a_5805_6446# a_5924_6446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X449 a_15568_2001# d1 a_15654_1216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X450 gnd d0 a_16741_3467# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X451 gnd d3 a_7038_2806# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X452 a_172_3867# a_179_4085# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X453 a_8945_5311# a_8947_5829# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X454 a_9364_2162# a_9146_2162# a_8883_2074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X455 a_2603_4232# d0 a_3396_4637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X456 a_11290_1203# d0 a_12087_1431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X457 a_2659_7286# d0 a_3452_7691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X458 a_14592_2399# a_14390_1383# a_14514_1502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X459 a_9964_2996# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X460 a_15599_6916# a_15852_6903# a_15423_4882# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X461 a_1721_131# d4 a_2314_5021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X462 gnd d0 a_8073_7514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X463 a_1602_131# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X464 a_8894_2581# d0 a_9385_2768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X465 a_11417_8329# d0 a_12210_8734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X466 a_11323_3416# a_11580_3226# a_11241_4024# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X467 a_5759_7466# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_2566_2196# a_2819_2183# a_2467_1786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X469 a_6090_263# a_5908_4408# a_6023_6446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X470 a_10467_275# a_10285_4420# a_10327_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X471 gnd d1 a_15961_4257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X472 a_228_6921# d0 a_717_6815# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X473 a_9130_732# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X474 gnd d1 a_16034_8329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X475 a_4549_4281# d0 a_5024_4186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 a_13333_6959# d0 a_13822_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X477 a_5929_6565# a_5759_7466# a_5883_7585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X478 a_9184_3786# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 gnd d0 a_12340_1418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 a_2536_6035# d1 a_2618_5427# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X481 a_4609_7952# d0 a_5098_7846# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X482 a_11396_7488# d0 a_12194_7304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X483 a_7036_8494# d0 a_7834_8310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X484 vdd d0 a_8073_7514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X485 a_9183_4198# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X486 vdd d3 a_11488_6890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X487 gnd d0 a_3617_1999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X488 a_6678_5034# d3 a_6785_2819# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X489 a_16468_2462# a_16721_2449# a_15671_2234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X490 a_11417_8329# d0 a_12214_8557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X491 a_4519_2862# a_4526_3080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X492 a_7747_3455# a_7761_4238# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X493 a_5080_7240# d1 a_5878_7056# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_16484_3657# a_16488_3480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X495 a_2562_2373# a_2819_2183# a_2467_1786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X496 a_7833_8722# a_7837_8545# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X497 a_1441_2971# a_1223_2971# a_643_3155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X498 vdd d0 a_3727_8107# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X499 gnd d1 a_2802_1165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X500 a_13547_4211# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 a_135_1831# a_142_2049# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X502 gnd d0 a_12431_6096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X503 a_15423_4882# d3 a_15599_6916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X504 a_1358_5417# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X505 vdd d2 a_7121_3822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X506 a_11158_3008# d2 a_11204_1988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X507 a_734_7833# a_516_7833# a_243_7840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X508 vdd d2 a_7194_7894# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X509 a_15605_4037# d1 a_15691_3252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X510 a_8947_5829# d0 a_9438_5822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X511 a_11396_7488# d0 a_12198_7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X512 a_7036_8494# d0 a_7838_8133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X513 a_5805_2984# a_5587_2984# a_5007_3168# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X514 a_1560_6433# a_1358_5417# a_1482_5536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X515 a_15641_6073# a_15898_5883# a_15595_7093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X516 a_15740_6483# d0 a_16538_6299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X517 a_5851_2374# a_5649_1358# a_5768_948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X518 a_4526_3080# a_4532_3263# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X519 a_133_1732# d0 a_624_1725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X520 vdd d1 a_2802_1165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X521 a_12120_3644# a_12124_3467# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X522 a_12198_7127# a_12193_7716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X523 a_14619_7081# a_14401_7081# a_13821_7265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X524 a_4495_1227# d0 a_4970_1132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X525 a_142_2049# a_148_2232# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X526 a_13566_5229# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X527 gnd d1 a_11653_7298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_606_1119# d1 a_1404_935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X529 a_4568_5299# d0 a_5043_5204# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X530 a_14665_6471# d3 a_14764_6471# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X531 a_1586_2361# a_1368_2361# a_1487_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X532 a_13221_752# a_13223_851# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X533 vdd d1 a_7256_6268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X534 a_2504_3822# d1 a_2599_4409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X535 vdd d0 a_16778_5091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X536 a_11204_1988# d1 a_11290_1203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X537 a_2573_8071# d1 a_2655_7463# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 a_16468_2462# a_16485_3245# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X539 a_16447_1621# a_16451_1444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X540 a_4497_1745# a_4499_1844# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X541 a_5550_948# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 a_10260_7597# d2 a_10306_6577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X543 a_7821_7115# a_8074_7102# a_7019_7476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X544 a_1240_3989# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X545 a_3416_5243# a_3420_5066# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X546 a_10136_7478# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X547 a_3469_8709# a_3726_8519# a_2676_8304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X548 a_4309_57# d7 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X549 a_2318_4844# d3 a_2494_6878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X550 a_15691_3252# d0 a_16484_3657# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_13346_7360# d0 a_13821_7265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 a_14308_1991# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X553 a_6085_144# d4 a_6682_4857# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X554 a_8939_5128# a_8945_5311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X555 a_5587_2984# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X556 a_5060_6222# a_4842_6222# a_4579_6134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_11307_2221# a_11560_2208# a_11208_1811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X558 a_3469_8709# a_3473_8532# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X559 a_252_8157# a_258_8340# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X560 a_4517_2569# d0 a_5008_2756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X561 a_3380_3207# a_3637_3017# a_2582_3391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X562 a_2467_1786# a_2720_1773# a_2417_2983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_2573_8071# d1 a_2659_7286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X564 vdd d2 a_11571_7906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X565 a_1721_131# d5 a_1820_131# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X566 a_3453_7279# a_3710_7089# a_2655_7463# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X567 a_1492_2480# a_1322_3381# a_1446_3500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X568 a_9474_8270# a_9256_8270# a_8999_8365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X569 a_15654_1216# a_15907_1203# a_15568_2001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 a_5024_4186# a_4806_4186# a_4543_4098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X571 a_12161_5091# a_12414_5078# a_11359_5452# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X572 gnd d0 a_3616_2411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X573 a_426_2743# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X574 a_5024_4186# d1 a_5810_3513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X575 gnd d0 a_8091_8120# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X576 a_13531_2781# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X577 a_7706_1596# a_7963_1406# a_6913_1191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X578 gnd d0 a_8053_6496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_5677_8074# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X580 a_5966_144# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X581 a_13530_3193# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X582 a_11055_5046# d3 a_11162_2831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X583 a_5878_7056# a_5660_7056# a_5081_6828# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X584 a_13838_8283# a_13620_8283# a_13357_8195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X585 a_644_2743# a_426_2743# a_155_2849# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X586 a_11290_1203# d0 a_12083_1608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_6930_2209# d0 a_7723_2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X588 a_2463_1963# a_2720_1773# a_2417_2983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X589 a_13253_2270# a_13258_2594# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X590 a_16520_5693# a_16777_5503# a_15727_5288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X591 gnd d0 a_7964_994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X592 a_208_5903# d0 a_697_5797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X593 a_13333_6959# a_13340_7177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X594 a_10228_2386# a_10026_1370# a_10150_1489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X595 a_4971_720# d1 a_5768_948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X596 vdd d0 a_3616_2411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X597 a_13247_2087# d0 a_13728_2175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X598 a_9438_5822# d1 a_10223_5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X599 a_215_6121# d0 a_696_6209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X600 a_15744_6306# d0 a_16537_6711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X601 vdd d0 a_8091_8120# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X602 a_6909_1368# a_7166_1178# a_6827_1976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X603 a_11277_6060# a_11534_5870# a_11231_7080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X604 a_8876_1856# d0 a_9365_1750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X605 a_10343_156# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 a_13221_752# a_16448_1209# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X607 a_11376_6470# d0 a_12174_6286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X608 a_6926_2386# a_7183_2196# a_6831_1799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X609 a_7706_1596# a_7710_1419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X610 a_4534_3781# a_4536_3880# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X611 a_12141_4485# a_12394_4472# a_11344_4257# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X612 vdd d0 a_12430_6508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X613 a_6930_2209# d0 a_7727_2437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X614 a_9220_5822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X615 a_4622_8353# a_3473_8532# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X616 a_1276_6025# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X617 a_9421_4804# a_9203_4804# a_8930_4811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X618 a_1477_5007# a_1259_5007# a_680_4779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X619 a_15744_6306# d0 a_16541_6534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X620 a_10327_2386# a_10109_2386# a_10233_2505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X621 a_191_4885# a_198_5103# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X622 a_11318_7919# a_11571_7906# a_11235_6903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X623 a_5773_1477# a_5567_1966# a_4987_2150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X624 a_16465_2227# a_16722_2037# a_15667_2411# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X625 a_12121_3232# a_12125_3055# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X626 vdd d4 a_11312_4856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X627 a_9384_3180# d1 a_10182_2996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X628 a_12137_4662# a_12394_4472# a_11344_4257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X629 a_2672_8481# a_2929_8291# a_2577_7894# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X630 a_15650_1393# d0 a_16452_1032# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X631 a_6967_4245# a_7220_4232# a_6868_3835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X632 a_7019_7476# d0 a_7817_7292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X633 a_15605_4037# d1 a_15687_3429# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_9166_3180# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X635 a_733_8245# d1 a_1519_7572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X636 a_8909_3275# a_8911_3793# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X637 a_15682_7932# a_15935_7919# a_15599_6916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X638 gnd d3 a_15779_2831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X639 a_14587_5574# a_14381_6063# a_13801_6247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X640 a_607_707# a_389_707# a_116_714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X641 a_4599_7152# d0 a_5080_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X642 a_1565_6552# a_1395_7453# a_1514_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X643 a_15723_5465# d0 a_16525_5104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X644 a_13277_3905# a_13284_4123# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X645 a_4970_1132# d1 a_5768_948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X646 a_4863_6828# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X647 a_16557_7729# a_16814_7539# a_15764_7324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X648 a_179_4085# d0 a_660_4173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X649 a_6854_7068# a_7111_6878# a_6682_4857# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X650 a_4482_826# d0 a_4971_720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X651 a_4579_6134# a_4585_6317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X652 a_498_7227# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_16448_1209# a_16452_1032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X654 a_5008_2756# a_4790_2756# a_4519_2862# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X655 vdd d1 a_2839_3201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X656 a_1404_935# d2 a_1487_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X657 a_13603_7265# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X658 a_6963_4422# a_7220_4232# a_6868_3835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X659 a_716_7227# a_498_7227# a_241_7322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X660 gnd d1 a_7256_6268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X661 gnd d0 a_16832_8145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 a_13821_7265# a_13603_7265# a_13346_7360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X663 a_11235_6903# d2 a_11318_7919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X664 a_10218_5032# d2 a_10301_6458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X665 a_2618_5427# d0 a_3416_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X666 a_2421_2806# a_2674_2793# a_2314_5021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X667 a_5097_8258# a_4879_8258# a_4622_8353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X668 a_3470_8297# a_3474_8120# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X669 a_3363_2424# a_3380_3207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X670 gnd d0 a_16704_1431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 a_14514_1502# d2 a_14592_2399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_15777_8519# a_16034_8329# a_15682_7932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X673 a_8932_4910# a_8939_5128# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X674 a_3456_7514# a_3709_7501# a_2659_7286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_4480_727# a_7707_1184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X676 a_3473_8532# a_3726_8519# a_2676_8304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X677 a_15781_8342# d0 gnd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X678 a_12156_5680# a_12413_5490# a_11363_5275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X679 a_9219_6234# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X680 a_8926_4293# a_8930_4811# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X681 a_8894_2581# a_8896_2874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X682 a_4842_6222# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X683 vdd d0 a_16832_8145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X684 a_5924_6446# d3 a_6023_6446# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X685 a_4770_1738# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X686 a_1544_4395# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X687 a_6827_1976# d1 a_6913_1191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X688 a_3384_3030# a_3637_3017# a_2582_3391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 a_2618_5427# d0 a_3420_5066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X690 a_11344_4257# a_11597_4244# a_11245_3847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X691 a_6831_1799# d1 a_6930_2209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X692 gnd d1 a_15924_2221# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X693 vdd d0 a_16704_1431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X694 a_405_2137# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X695 gnd d3 a_2747_6865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X696 a_11417_8329# a_11670_8316# a_11318_7919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X697 a_5550_948# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X698 a_13510_2175# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X699 a_606_1119# a_388_1119# a_125_1031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X700 a_11231_7080# d2 a_11277_6060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_479_5797# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X702 a_13711_1157# a_13493_1157# a_13230_1069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 a_13584_5835# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X704 a_13785_4817# a_13567_4817# a_13294_4824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X705 a_15645_5896# d1 a_15744_6306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X706 a_14649_4433# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X707 a_13348_7878# a_13350_7977# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X708 a_1820_131# a_1602_131# a_1726_250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X709 a_14364_5045# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X710 a_11380_6293# d0 a_12177_6521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X711 a_15419_5059# a_15676_4869# a_14826_169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X712 a_644_2743# d1 a_1441_2971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X713 a_11340_4434# a_11597_4244# a_11245_3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X714 a_8984_7865# d0 a_9475_7858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X715 a_7707_1184# a_7711_1007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X716 vdd d1 a_15924_2221# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X717 gnd d1 a_7293_8304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X718 a_717_6815# d1 a_1514_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X719 a_11413_8506# a_11670_8316# a_11318_7919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X720 a_14707_169# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X721 a_2500_3999# a_2757_3809# a_2421_2806# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X722 gnd d0 a_3599_1393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X723 a_2599_4409# d0 a_3397_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X724 a_389_707# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X725 a_258_8340# d0 a_733_8245# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X726 a_1446_3500# a_1240_3989# a_661_3761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X727 a_12832_82# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 a_1441_2971# a_1223_2971# a_644_2743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X729 a_13350_7977# d0 a_13839_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 a_6913_1191# a_7166_1178# a_6827_1976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X731 a_7800_6509# a_7817_7292# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X732 a_7760_4650# a_7764_4473# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X733 a_9964_2996# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X734 gnd d3 a_15852_6903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X735 a_13357_8195# d0 a_13838_8283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X736 a_6913_1191# d0 a_7706_1596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X737 a_13821_7265# d1 a_14619_7081# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 a_14597_2518# a_14427_3419# a_14546_3009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X739 a_1313_8061# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 a_206_5804# a_208_5903# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X741 a_6682_4857# d3 a_6858_6891# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X742 a_15419_5059# d3 a_15522_3021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X743 gnd d1 a_11543_1190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X744 a_9457_7252# a_9239_7252# a_8976_7164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X745 gnd d1 a_2819_2183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X746 a_2599_4409# d0 a_3401_4048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X747 a_13223_851# d0 a_13712_745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X748 a_15727_5288# d0 a_16520_5693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X749 a_1519_7572# a_1313_8061# a_733_8245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X750 gnd d1 a_2892_6255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_1565_6552# d3 a_1659_6433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X752 vdd d0 a_8074_7102# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X753 a_8866_1056# d0 a_9347_1144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X754 a_16469_2050# a_16722_2037# a_15667_2411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X755 a_9147_1750# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X756 a_5768_948# d2 a_5851_2374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X757 a_10150_1489# d2 a_10228_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X758 a_15682_7932# d1 a_15781_8342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X759 a_4769_2150# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X760 a_12174_6286# a_12178_6109# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X761 a_15650_1393# d0 a_16448_1209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X762 a_9927_960# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X763 a_5805_6446# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X764 a_9420_5216# d1 a_10218_5032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X765 a_4826_4792# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X766 a_4572_5916# a_4579_6134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X767 vdd d1 a_2819_2183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X768 a_14390_1383# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X769 a_6785_2819# a_7038_2806# a_6678_5034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X770 a_5924_6446# a_5722_5430# a_5841_5020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X771 vdd d0 a_12341_1006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X772 a_3419_5478# a_3433_6261# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X773 vdd d1 a_2892_6255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X774 gnd d0 a_3710_7089# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 a_16561_7552# a_16814_7539# a_15764_7324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_4585_6317# d0 a_5060_6222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X777 a_6023_6446# a_5805_6446# a_5929_6565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X778 a_4553_4799# a_4555_4898# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X779 vdd d2 a_11461_1798# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X780 a_4512_2245# a_4517_2569# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X781 a_7820_7527# a_8073_7514# a_7023_7299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_9364_2162# a_9146_2162# a_8889_2257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X783 a_1441_2971# d2 a_1492_2480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X784 a_8539_81# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X785 a_8947_5829# a_8949_5928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X786 a_10285_4420# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X787 gnd d3 a_7111_6878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X788 a_10223_5561# a_10017_6050# a_9438_5822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X789 a_15781_8342# a_16034_8329# a_15682_7932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X790 a_5759_7466# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X791 a_7816_7704# a_8073_7514# a_7023_7299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X792 a_3347_994# a_3342_1583# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X793 a_4543_4098# a_4549_4281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X794 a_15781_8342# d0 a_16574_8747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 a_226_6628# d0 a_717_6815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X796 a_3364_2012# a_3617_1999# a_2562_2373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X797 gnd d2 a_2830_7881# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X798 a_13331_6666# d0 a_13822_6853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X799 a_4599_7152# a_4605_7335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X800 a_4607_7853# d0 a_5098_7846# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X801 a_1223_2971# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X802 a_3470_8297# a_3727_8107# a_2672_8481# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X803 a_9385_2768# a_9167_2768# a_8894_2581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X804 a_1240_3989# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X805 a_6827_1976# d1 a_6909_1368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X806 a_15687_3429# d0 a_16485_3245# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X807 a_9401_4198# d1 a_10187_3525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X808 a_442_4173# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X809 a_16501_4675# a_16505_4498# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X810 a_5081_6828# d1 a_5878_7056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X811 a_10233_2505# a_10063_3406# a_10182_2996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X812 a_516_7833# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 a_13290_4306# d0 a_13765_4211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X814 a_5587_2984# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X815 a_16488_3480# a_16502_4263# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X816 a_13621_7871# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_13547_4211# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X818 a_8932_4910# d0 a_9421_4804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X819 a_16574_8747# gnd SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X820 a_1358_5417# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X821 a_11307_2221# d0 a_12100_2626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X822 a_13620_8283# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X823 a_14345_4027# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X824 a_11363_5275# d0 a_12156_5680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X825 a_10233_2505# d3 a_10327_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X826 a_734_7833# a_516_7833# a_245_7939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X827 a_14401_7081# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X828 a_7761_4238# a_7765_4061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X829 a_168_3250# a_170_3768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X830 gnd d1 a_15907_1203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X831 a_15687_3429# d0 a_16489_3068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X832 a_7707_1184# a_7964_994# a_6909_1368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X833 gnd d0 a_8054_6084# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X834 a_11400_7311# a_11653_7298# a_11314_8096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X835 a_5851_2374# a_5649_1358# a_5773_1477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X836 a_2490_7055# d2 a_2540_5858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X837 a_15526_2844# d2 a_15609_3860# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X838 a_1368_2361# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 a_4499_1844# d0 a_4988_1738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X840 a_6926_2386# d0 a_7724_2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 vdd d0 a_7963_1406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X842 a_15572_1824# a_15825_1811# a_15522_3021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X843 a_4489_1044# d0 a_4970_1132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X844 a_4555_4898# d0 a_5044_4792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 a_6999_6458# a_7256_6268# a_6904_5871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X846 a_13267_3105# a_13273_3288# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X847 a_12124_3467# a_12138_4250# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X848 a_4616_8170# a_4622_8353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X849 a_11307_2221# d0 a_12104_2449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X850 a_5773_1477# a_5567_1966# a_4988_1738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 a_16521_5281# a_16778_5091# a_15723_5465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X852 a_4562_5116# d0 a_5043_5204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X853 a_12210_8734# a_12214_8557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X854 a_14291_973# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X855 a_1586_2361# a_1368_2361# a_1492_2480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X856 a_9438_5822# a_9220_5822# a_8947_5829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 vdd d0 a_3617_1999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X858 a_7765_4061# a_7760_4650# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X859 a_1726_250# a_1544_4395# a_1586_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 vdd d0 a_8054_6084# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X861 a_5950_2374# a_5732_2374# a_5851_2374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X862 a_7023_7299# d0 a_7816_7704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 a_624_1725# a_406_1725# a_133_1732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X864 a_10255_7068# d2 a_10306_6577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X865 a_11286_1380# d0 a_12088_1019# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X866 a_12142_4073# a_12395_4060# a_11340_4434# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_6926_2386# d0 a_7728_2025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X868 vdd d3 a_2674_2793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X869 a_2655_7463# d0 a_3453_7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X870 a_4309_57# a_4091_57# a_4210_57# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X871 gnd d3 a_11415_2818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X872 a_2639_6268# a_2892_6255# a_2540_5858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 a_16561_7552# a_16575_8335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X874 a_11158_3008# d2 a_11208_1811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X875 a_16537_6711# a_16541_6534# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X876 vdd d0 a_3709_7501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X877 a_8909_3275# d0 a_9384_3180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X878 a_14764_6471# a_14546_6471# a_14665_6471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X879 a_13340_7177# d0 a_13821_7265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X880 a_8903_3092# a_8909_3275# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X881 a_5810_3513# d2 a_5856_2493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X882 a_16485_3245# a_16489_3068# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X883 a_1322_3381# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X884 a_8969_6946# d0 a_9458_6840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X885 a_15740_6483# d0 a_16542_6122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X886 a_5060_6222# a_4842_6222# a_4585_6317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X887 a_15682_7932# d1 a_15777_8519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X888 a_9256_8270# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X889 a_4806_4186# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X890 a_3363_2424# a_3616_2411# a_2566_2196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 a_131_1214# a_133_1732# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X892 a_7023_7299# d0 a_7820_7527# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X893 a_7800_6509# a_8053_6496# a_7003_6281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_155_2849# d0 a_644_2743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X895 a_12138_4250# a_12395_4060# a_11340_4434# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X896 vdd d1 a_11653_7298# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X897 a_15704_4447# a_15961_4257# a_15609_3860# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X898 a_7779_5668# a_7783_5491# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X899 a_2635_6445# a_2892_6255# a_2540_5858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X900 a_426_2743# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X901 a_9385_2768# d1 a_10182_2996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X902 a_5025_3774# d1 a_5810_3513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X903 a_2494_6878# d2 a_2577_7894# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X904 a_8913_3892# a_8920_4110# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X905 a_11162_2831# d2 a_11241_4024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X906 vdd d1 a_2929_8291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X907 a_13258_2594# d0 a_13749_2781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X908 a_6090_263# d5 a_4210_57# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X909 a_8969_6946# a_8976_7164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X910 gnd d2 a_15935_7919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X911 a_5878_7056# a_5660_7056# a_5080_7240# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X912 a_3359_2601# a_3616_2411# a_2566_2196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X913 a_16558_7317# a_16815_7127# a_15760_7501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X914 a_12138_4250# a_12142_4073# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X915 a_14624_7610# a_14418_8099# a_13839_7871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X916 a_13236_1252# d0 a_13711_1157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X917 a_11277_6060# d1 a_11359_5452# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X918 a_6941_7907# d1 a_7040_8317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X919 a_5081_6828# a_4863_6828# a_4590_6641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X920 vdd d0 a_16814_7539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X921 a_12194_7304# a_12198_7127# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X922 a_13309_5324# d0 a_13784_5229# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 a_3401_4048# a_3396_4637# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X924 a_661_3761# a_443_3761# a_170_3768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X925 a_10343_156# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X926 a_6963_4422# d0 a_7765_4061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X927 a_9203_4804# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X928 a_8866_1056# a_8872_1239# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X929 a_1259_5007# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X930 a_11303_2398# a_11560_2208# a_11208_1811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X931 a_4988_1738# a_4770_1738# a_4497_1745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X932 a_10109_2386# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X933 gnd d0 a_12377_3454# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X934 vdd d0 a_16721_2449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X935 a_9421_4804# a_9203_4804# a_8932_4910# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X936 a_11277_6060# d1 a_11363_5275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X937 a_7710_1419# a_7724_2202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X938 a_1477_5007# a_1259_5007# a_679_5191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X939 a_5567_1966# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X940 vdd d4 a_2571_4831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X941 a_643_3155# d1 a_1441_2971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 a_7796_6686# a_7800_6509# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X943 a_7764_4473# a_7780_5256# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X944 a_679_5191# a_461_5191# a_198_5103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_13728_2175# a_13510_2175# a_13247_2087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X946 a_4753_720# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X947 a_11055_5046# a_11312_4856# a_10462_156# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X948 a_696_6209# a_478_6209# a_215_6121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X949 a_13801_6247# a_13583_6247# a_13320_6159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X950 a_10467_275# a_10285_4420# a_10400_6458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X951 a_15526_2844# a_15779_2831# a_15419_5059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_1395_7453# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X953 a_16452_1032# a_16447_1621# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X954 a_14826_169# d4 a_15419_5059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X955 vdd d0 a_16705_1019# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X956 a_14691_2399# a_14473_2399# a_14597_2518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X957 a_13711_1157# d1 a_14509_973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X958 vdd d0 a_12377_3454# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X959 a_12951_82# a_14707_169# a_14826_169# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X960 a_734_7833# d1 a_1519_7572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X961 a_12211_8322# a_12215_8145# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X962 gnd d1 a_7203_3214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X963 a_607_707# a_389_707# a_118_813# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X964 a_1565_6552# a_1395_7453# a_1519_7572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X965 a_5856_2493# a_5686_3394# a_5805_2984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X966 gnd d0 a_3689_6483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X967 a_13273_3288# d0 a_13748_3193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_9457_7252# d1 a_10255_7068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X969 a_4863_6828# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X970 a_8999_8365# a_7837_8545# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X971 a_13548_3799# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X972 a_15727_5288# a_15980_5275# a_15641_6073# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 a_4562_5116# a_4568_5299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X974 a_2586_3214# d0 a_3383_3442# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X975 vdd d3 a_7038_2806# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X976 a_498_7227# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X977 a_12156_5680# a_12160_5503# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X978 a_7003_6281# a_7256_6268# a_6904_5871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X979 gnd d1 a_16017_7311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X980 a_2659_7286# d0 a_3456_7514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X981 a_13603_7265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X982 a_8857_739# a_12084_1196# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X983 vout a_8539_81# a_8658_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X984 a_10026_1370# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X985 vdd d2 a_11498_3834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X986 a_14670_6590# a_14500_7491# a_14619_7081# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X987 gnd d0 a_3600_981# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X988 a_7003_6281# d0 a_7796_6686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X989 a_16451_1444# a_16704_1431# a_15654_1216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X990 a_11059_4869# d3 a_11235_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X991 a_16538_6299# a_16542_6122# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X992 a_12105_2037# a_12100_2626# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X993 vdd d1 a_7203_3214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X994 a_16520_5693# a_16524_5516# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X995 gnd d1 a_11633_6280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X996 a_9402_3786# a_9184_3786# a_8913_3892# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X997 a_1446_3500# a_1240_3989# a_660_4173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X998 vdd d0 a_3689_6483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X999 a_15723_5465# a_15980_5275# a_15641_6073# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1000 a_6909_1368# d0 a_7707_1184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1001 vdd d1 a_16017_7311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1002 a_10260_7597# a_10054_8086# a_9475_7858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1003 a_1487_2361# a_1285_1345# a_1404_935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1004 a_696_6209# d1 a_1482_5536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1005 a_3456_7514# a_3470_8297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1006 a_13728_2175# d1 a_14514_1502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1007 a_7780_5256# a_7784_5079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1008 a_16447_1621# a_16704_1431# a_15654_1216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1009 a_2494_6878# a_2747_6865# a_2318_4844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 a_1586_2361# d4 a_1726_250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1011 a_388_1119# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1012 a_4842_6222# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1013 vdd d1 a_11633_6280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1014 a_6682_4857# a_6935_4844# a_6085_144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 a_9365_1750# d1 a_10150_1489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1016 a_10301_6458# a_10099_5442# a_10218_5032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1017 a_13493_1157# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1018 a_5043_5204# a_4825_5204# a_4562_5116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1019 a_5640_6038# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1020 a_8984_7865# a_8986_7964# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1021 a_13567_4817# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1022 gnd d1 a_11580_3226# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1023 a_4506_2062# a_4512_2245# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1024 a_606_1119# a_388_1119# a_131_1214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1025 a_10145_960# a_9927_960# a_9347_1144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1026 a_12141_4485# a_12157_5268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1027 vdd d0 a_12431_6096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1028 a_2421_2806# d2 a_2500_3999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1029 a_680_4779# a_462_4779# a_189_4786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 a_13711_1157# a_13493_1157# a_13236_1252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1031 a_15708_4270# a_15961_4257# a_15609_3860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1032 a_16562_7140# a_16557_7729# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1033 a_13785_4817# a_13567_4817# a_13296_4923# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1034 a_14649_4433# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1035 a_10187_3525# d2 a_10233_2505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1036 a_16562_7140# a_16815_7127# a_15760_7501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1037 a_15671_2234# d0 a_16468_2462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1038 a_8857_739# a_8859_838# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1039 a_6937_8084# d1 a_7019_7476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_1721_131# d4 a_2318_4844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1041 a_1223_2971# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1042 a_10462_156# d4 a_11055_5046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 vdd d1 a_11580_3226# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1044 gnd d0 a_16814_7539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1045 a_14707_169# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1046 a_4309_57# a_4091_57# a_1820_131# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1047 vdd d0 a_3653_4447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1048 a_252_8157# d0 a_733_8245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1049 a_14427_3419# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1050 a_13348_7878# d0 a_13839_7871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1051 a_11290_1203# a_11543_1190# a_11204_1988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1052 a_6963_4422# d0 a_7761_4238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1053 a_3437_6084# a_3690_6071# a_2635_6445# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1054 a_155_2849# a_162_3067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1055 a_9401_4198# a_9183_4198# a_8920_4110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1056 a_14597_2518# a_14427_3419# a_14551_3538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1057 a_6868_3835# a_7121_3822# a_6785_2819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1058 a_1313_8061# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1059 a_13839_7871# d1 a_14624_7610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1060 a_9475_7858# a_9257_7858# a_8984_7865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1061 a_6831_1799# a_7084_1786# a_6781_2996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1062 a_6937_8084# d1 a_7023_7299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1063 gnd d0 a_16721_2449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1064 a_15678_8109# a_15935_7919# a_15599_6916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1065 a_1514_7043# a_1296_7043# a_717_6815# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1066 a_9457_7252# a_9239_7252# a_8982_7347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1067 a_7817_7292# a_8074_7102# a_7019_7476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1068 a_15777_8519# d0 a_16575_8335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1069 gnd d0 a_7980_2424# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1070 a_13221_752# d0 a_13712_745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1071 a_8859_838# d0 a_9348_732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1072 a_8962_6329# d0 a_9437_6234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1073 a_8874_1757# d0 a_9365_1750# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1074 a_1560_6433# d3 a_1659_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1075 gnd d1 a_7183_2196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1076 a_607_707# d1 a_1404_935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1077 a_3433_6261# a_3690_6071# a_2635_6445# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1078 gnd d0 a_16705_1019# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 a_13766_3799# a_13548_3799# a_13277_3905# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1080 a_12157_5268# a_12161_5091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1081 a_226_6628# a_228_6921# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1082 a_5722_5430# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 a_148_2232# d0 a_623_2137# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1084 a_6827_1976# a_7084_1786# a_6781_2996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1085 a_13240_1869# a_13247_2087# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1086 a_13240_1869# d0 a_13729_1763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1087 gnd d2 a_7157_5858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1088 a_15777_8519# d0 a_16579_8158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1089 a_15650_1393# a_15907_1203# a_15568_2001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1090 gnd d1 a_15997_6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1091 a_5805_6446# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1092 a_9421_4804# d1 a_10218_5032# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1093 a_198_5103# d0 a_679_5191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1094 vdd d0 a_3600_981# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1095 a_13313_5941# d0 a_13802_5835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1096 a_7821_7115# a_7816_7704# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1097 vdd d0 a_7980_2424# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1098 vdd d0 a_8036_5478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1099 a_15572_1824# d1 a_15667_2411# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1100 a_16521_5281# a_16525_5104# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1101 a_7727_2437# a_7744_3220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1102 vdd d0 a_8053_6496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1103 a_4579_6134# d0 a_5060_6222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1104 a_2586_3214# d0 a_3379_3619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_13784_5229# d1 a_14582_5045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1106 a_7816_7704# a_7820_7527# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1107 a_4495_1227# a_4497_1745# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1108 a_5060_6222# d1 a_5846_5549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_1409_1464# a_1203_1953# a_623_2137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1110 vdd d0 a_7964_994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1111 a_11245_3847# a_11498_3834# a_11162_2831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1112 a_2672_8481# d0 a_3470_8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1113 a_8876_1856# a_8883_2074# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1114 gnd d2 a_15825_1811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1115 a_11241_4024# d1 a_11323_3416# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1116 a_11359_5452# d0 a_12161_5091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1117 a_15572_1824# d1 a_15671_2234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1118 gnd d0 a_3672_5465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1119 a_11376_6470# d0 a_12178_6109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1120 gnd d3 a_11488_6890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1121 a_4480_727# d0 a_4971_720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1122 a_4532_3263# d0 a_5007_3168# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1123 gnd d0 a_8017_4460# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1124 a_9167_2768# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_8999_8365# d0 a_9474_8270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1126 a_4592_6934# d0 a_5081_6828# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1127 a_14619_7081# d2 a_14670_6590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1128 a_12101_2214# a_12105_2037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1129 gnd d1 a_11560_2208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1130 a_15423_4882# d3 a_15595_7093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1131 a_258_8340# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1132 a_10063_3406# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1133 a_3437_6084# a_3432_6673# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1134 gnd d2 a_2720_1773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1135 a_9385_2768# a_9167_2768# a_8896_2874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1136 a_172_3867# d0 a_661_3761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1137 vdd d0 a_3710_7089# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1138 a_11241_4024# d1 a_11327_3239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1139 gnd d2 a_7194_7894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1140 a_9402_3786# d1 a_10187_3525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1141 a_13273_3288# a_13275_3806# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1142 a_442_4173# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1143 vdd d0 a_3672_5465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1144 a_10233_2505# a_10063_3406# a_10187_3525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1145 a_643_3155# a_425_3155# a_162_3067# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1146 a_13284_4123# d0 a_13765_4211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1147 a_9475_7858# d1 a_10260_7597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1148 a_516_7833# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1149 vdd d0 a_8017_4460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1150 a_6785_2819# d2 a_6864_4012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1151 a_4568_5299# a_4570_5817# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1152 a_13749_2781# a_13531_2781# a_13258_2594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1153 a_13621_7871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1154 a_6781_2996# d2 a_6827_1976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1155 a_717_6815# a_499_6815# a_226_6628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1156 a_13765_4211# d1 a_14551_3538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1157 a_8930_4811# d0 a_9421_4804# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1158 a_7019_7476# d0 a_7821_7115# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1159 a_13748_3193# a_13530_3193# a_13273_3288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1160 gnd d1 a_7239_5250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1161 a_13822_6853# a_13604_6853# a_13331_6666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1162 a_14345_4027# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1163 a_7801_6097# a_8054_6084# a_6999_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1164 a_5098_7846# a_4880_7846# a_4607_7853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1165 a_9348_732# a_9130_732# a_8857_739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1166 vdd d0 a_16831_8557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1167 vdd d2 a_2720_1773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1168 a_14546_3009# a_14328_3009# a_13749_2781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1169 a_15671_2234# d0 a_16464_2639# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1170 a_13326_6342# d0 a_13801_6247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1171 a_9146_2162# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1172 a_5567_1966# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1173 a_170_3768# a_172_3867# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1174 a_14592_2399# d3 a_14691_2399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1175 a_1368_2361# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1176 a_4497_1745# d0 a_4988_1738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1177 a_3360_2189# a_3617_1999# a_2562_2373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1178 gnd d0 a_3653_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1179 gnd d2 a_2793_5845# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 a_6781_2996# d2 a_6831_1799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1181 a_12104_2449# a_12121_3232# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1182 a_12193_7716# a_12197_7539# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1183 vdd d1 a_7239_5250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1184 vdd d0 a_16815_7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1185 a_7797_6274# a_8054_6084# a_6999_6458# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1186 a_6023_6446# d4 a_6090_263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1187 a_9438_5822# a_9220_5822# a_8949_5928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1188 a_221_6304# a_226_6628# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1189 a_13357_8195# a_13363_8378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1190 a_406_1725# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1191 gnd d0 a_12467_8544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1192 a_2417_2983# a_2674_2793# a_2314_5021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1193 a_13511_1763# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1194 a_4971_720# a_4753_720# a_4480_727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1195 a_11162_2831# a_11415_2818# a_11055_5046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 a_208_5903# a_215_6121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1197 a_1186_935# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1198 a_461_5191# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1199 a_5950_2374# a_5732_2374# a_5856_2493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1200 a_3452_7691# a_3709_7501# a_2659_7286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1201 a_13236_1252# a_13238_1770# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1202 a_5846_5549# a_5640_6038# a_5061_5810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1203 a_624_1725# a_406_1725# a_135_1831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1204 a_7747_3455# a_8000_3442# a_6950_3227# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1205 a_5841_5020# a_5623_5020# a_5044_4792# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1206 a_10037_7068# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1207 gnd d2 a_11571_7906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1208 a_11231_7080# a_11488_6890# a_11059_4869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1209 gnd d0 a_12378_3042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1210 a_8913_3892# d0 a_9402_3786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1211 a_14764_6471# a_14546_6471# a_14670_6590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1212 a_8920_4110# a_8926_4293# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1213 a_3342_1583# a_3346_1406# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1214 gnd d1 a_7220_4232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 vdd d0 a_12467_8544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1216 a_7817_7292# a_7821_7115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1217 a_11396_7488# a_11653_7298# a_11314_8096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1218 a_8993_8182# a_8999_8365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1219 vdd d3 a_15779_2831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1220 a_5007_3168# a_4789_3168# a_4526_3080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1221 a_2549_1178# d0 a_3342_1583# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1222 a_15744_6306# a_15997_6293# a_15645_5896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1223 a_16575_8335# a_16579_8158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1224 a_7743_3632# a_8000_3442# a_6950_3227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1225 a_12142_4073# a_12137_4662# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1226 a_10306_6577# a_10136_7478# a_10255_7068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1227 a_133_1732# a_135_1831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1228 a_4091_57# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1229 a_153_2556# d0 a_644_2743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1230 a_6937_8084# a_7194_7894# a_6858_6891# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1231 a_1482_5536# d2 a_1560_6433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1232 vdd d3 a_7111_6878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1233 a_2676_8304# d0 a_3473_8532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1234 vdd d0 a_12378_3042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1235 gnd d0 a_8036_5478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1236 a_7783_5491# a_7797_6274# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1237 a_14418_8099# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1238 a_5649_1358# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1239 a_14500_7491# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1240 a_10145_960# d2 a_10228_2386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1241 a_6085_144# d5 a_4210_57# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1242 vdd d1 a_7220_4232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1243 gnd d0 a_3690_6071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1244 a_11208_1811# d1 a_11303_2398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1245 vdd d1 a_7293_8304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1246 a_2582_3391# d0 a_3384_3030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1247 a_191_4885# d0 a_680_4779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_2417_2983# d2 a_2463_1963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 a_9944_1978# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1250 vdd d0 a_3599_1393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1251 a_16469_2050# a_16464_2639# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1252 a_13230_1069# d0 a_13711_1157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1253 a_5081_6828# a_4863_6828# a_4592_6934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1254 a_2655_7463# d0 a_3457_7102# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1255 a_9364_2162# d1 a_10150_1489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1256 a_5924_6446# a_5722_5430# a_5846_5549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1257 a_11359_5452# d0 a_12157_5268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1258 a_13303_5141# d0 a_13784_5229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1259 a_12832_82# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1260 a_6999_6458# d0 a_7797_6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1261 a_5810_3513# a_5604_4002# a_5025_3774# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1262 a_1441_6433# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_661_3761# a_443_3761# a_172_3867# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1264 a_12124_3467# a_12377_3454# a_11327_3239# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1265 a_6913_1191# d0 a_7710_1419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1266 a_9203_4804# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1267 a_1259_5007# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1268 a_6900_6048# d1 a_6982_5440# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1269 a_12197_7539# a_12450_7526# a_11400_7311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1270 vdd d0 a_3690_6071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1271 vdd d1 a_11543_1190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1272 a_478_6209# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1273 a_2417_2983# d2 a_2467_1786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1274 a_4988_1738# a_4770_1738# a_4499_1844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1275 a_8956_6146# a_8962_6329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1276 a_13583_6247# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1277 a_15727_5288# d0 a_16524_5516# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1278 a_10285_4420# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1279 a_697_5797# a_479_5797# a_206_5804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 gnd d1 a_11670_8316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1281 a_5768_948# a_5550_948# a_4970_1132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1282 a_6999_6458# d0 a_7801_6097# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1283 vdd d3 a_2747_6865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1284 a_13728_2175# a_13510_2175# a_13253_2270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1285 a_16448_1209# a_16705_1019# a_15650_1393# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1286 a_10223_5561# a_10017_6050# a_9437_6234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1287 a_696_6209# a_478_6209# a_221_6304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1288 a_14473_2399# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1289 a_13729_1763# d1 a_14514_1502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1290 a_9365_1750# a_9147_1750# a_8874_1757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1291 a_8926_4293# d0 a_9401_4198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1292 a_11231_7080# d2 a_11281_5883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1293 a_12120_3644# a_12377_3454# a_11327_3239# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1294 a_13801_6247# a_13583_6247# a_13326_6342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1295 a_5007_3168# d1 a_5805_2984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1296 a_6950_3227# a_7203_3214# a_6864_4012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1297 a_6900_6048# d1 a_6986_5263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1298 a_12193_7716# a_12450_7526# a_11400_7311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1299 a_3452_7691# a_3456_7514# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1300 a_1395_7453# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1301 a_11344_4257# d0 a_12137_4662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1302 gnd d4 a_6935_4844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1303 a_5686_3394# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1304 a_12951_82# a_14707_169# a_14831_288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1305 gnd d0 a_16831_8557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1306 a_6781_2996# a_7038_2806# a_6678_5034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1307 a_15764_7324# a_16017_7311# a_15678_8109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1308 vdd d1 a_11670_8316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1309 a_13277_3905# d0 a_13766_3799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1310 a_204_5286# a_206_5804# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1311 a_9458_6840# d1 a_10255_7068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1312 a_11235_6903# d2 a_11314_8096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1313 a_2463_1963# d1 a_2545_1355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1314 a_11323_3416# d0 a_12121_3232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1315 a_4536_3880# d0 a_5025_3774# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 a_2540_5858# a_2793_5845# a_2490_7055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1317 a_15667_2411# d0 a_16469_2050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1318 vdd d3 a_11415_2818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1319 a_6946_3404# a_7203_3214# a_6864_4012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1320 a_4543_4098# d0 a_5024_4186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1321 a_11380_6293# a_11633_6280# a_11281_5883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 a_7728_2025# a_7723_2614# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1323 a_10182_2996# a_9964_2996# a_9385_2768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1324 a_11344_4257# d0 a_12141_4485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1325 a_9184_3786# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1326 gnd d0 a_16815_7127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1327 a_6868_3835# d1 a_6963_4422# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 a_6858_6891# d2 a_6941_7907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1329 a_15599_6916# d2 a_15678_8109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1330 a_13331_6666# a_13333_6959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1331 a_7723_2614# a_7727_2437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1332 a_13290_4306# a_13294_4824# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1333 a_15760_7501# a_16017_7311# a_15678_8109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1334 a_15419_5059# d3 a_15526_2844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1335 a_10054_8086# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1336 a_1285_1345# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1337 a_16524_5516# a_16538_6299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1338 a_15764_7324# d0 a_16561_7552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1339 a_4592_6934# a_4599_7152# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1340 a_2463_1963# d1 a_2549_1178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1341 a_118_813# a_125_1031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1342 vout a_8539_81# a_4309_57# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1343 a_11323_3416# d0 a_12125_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1344 a_624_1725# d1 a_1409_1464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1345 a_116_714# a_118_813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1346 a_1487_2361# a_1285_1345# a_1409_1464# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1347 a_11376_6470# a_11633_6280# a_11281_5883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1348 a_3436_6496# a_3453_7279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1349 a_10099_5442# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1350 a_697_5797# d1 a_1482_5536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1351 a_4825_5204# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1352 a_6868_3835# d1 a_6967_4245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1353 gnd d0 a_7981_2012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1354 vdd d2 a_15935_7919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1355 a_5044_4792# a_4826_4792# a_4553_4799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1356 a_388_1119# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1357 a_462_4779# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_1409_1464# a_1203_1953# a_624_1725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1359 a_12088_1019# a_12083_1608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1360 a_10301_6458# a_10099_5442# a_10223_5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1361 a_13493_1157# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1362 a_189_4786# a_191_4885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1363 a_5043_5204# a_4825_5204# a_4568_5299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1364 a_2314_5021# d3 a_2417_2983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1365 a_5640_6038# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1366 a_8967_6653# a_8969_6946# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1367 a_14592_2399# a_14390_1383# a_14509_973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1368 a_13567_4817# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1369 a_13801_6247# d1 a_14587_5574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 a_12083_1608# a_12087_1431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1371 a_680_4779# a_462_4779# a_191_4885# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1372 a_14665_6471# a_14463_5455# a_14582_5045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1373 a_2676_8304# d0 a_3469_8709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1374 a_11363_5275# d0 a_12160_5503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1375 a_245_7939# a_252_8157# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1376 a_2500_3999# d1 a_2582_3391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1377 a_8903_3092# d0 a_9384_3180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1378 a_2577_7894# a_2830_7881# a_2494_6878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1379 vdd d0 a_7981_2012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1380 a_8967_6653# d0 a_9458_6840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1381 vdd d1 a_15907_1203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1382 a_10182_2996# d2 a_10233_2505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1383 a_3396_4637# a_3653_4447# a_2603_4232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1384 a_2582_3391# d0 a_3380_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1385 a_11245_3847# d1 a_11340_4434# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1386 a_14831_288# d5 a_12951_82# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 a_241_7322# d0 a_716_7227# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 a_11318_7919# d1 a_11413_8506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1389 a_14551_3538# d2 a_14597_2518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 a_12177_6521# a_12430_6508# a_11380_6293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1391 a_9183_4198# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1392 a_3383_3442# a_3397_4225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1393 a_14427_3419# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1394 a_3400_4460# a_3416_5243# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1395 a_4622_8353# d0 a_5097_8258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1396 a_5061_5810# a_4843_5810# a_4570_5817# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1397 a_9257_7858# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1398 a_4549_4281# a_4553_4799# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1399 a_9240_6840# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1400 a_1296_7043# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1401 a_15678_8109# d1 a_15760_7501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1402 a_14826_169# d4 a_15423_4882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1403 a_12088_1019# a_12341_1006# a_11286_1380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1404 gnd d0 a_3673_5053# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1405 a_4862_7240# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1406 vdd d2 a_2830_7881# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1407 a_11245_3847# d1 a_11344_4257# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1408 a_12161_5091# a_12156_5680# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1409 a_9475_7858# a_9257_7858# a_8986_7964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1410 a_5025_3774# a_4807_3774# a_4534_3781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1411 a_1514_7043# a_1296_7043# a_716_7227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1412 a_11318_7919# d1 a_11417_8329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1413 a_2421_2806# d2 a_2504_3822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1414 a_2618_5427# a_2875_5237# a_2536_6035# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1415 a_5024_4186# a_4806_4186# a_4549_4281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1416 a_733_8245# a_515_8245# a_252_8157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1417 a_16452_1032# a_16705_1019# a_15650_1393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1418 a_8857_739# d0 a_9348_732# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1419 a_13531_2781# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1420 a_8956_6146# d0 a_9437_6234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1421 a_13839_7871# a_13621_7871# a_13348_7878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1422 a_6904_5871# a_7157_5858# a_6854_7068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1423 a_15678_8109# d1 a_15764_7324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1424 a_13838_8283# a_13620_8283# a_13363_8378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1425 a_13494_745# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 vdd d0 a_3673_5053# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1427 a_14619_7081# a_14401_7081# a_13822_6853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1428 a_142_2049# d0 a_623_2137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1429 a_5043_5204# d1 a_5841_5020# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1430 a_13223_851# a_13230_1069# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1431 a_7779_5668# a_8036_5478# a_6986_5263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1432 vdd d0 a_8018_4048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1433 a_10000_5032# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1434 a_13238_1770# d0 a_13729_1763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1435 a_7796_6686# a_8053_6496# a_7003_6281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1436 gnd d2 a_11534_5870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1437 a_206_5804# d0 a_697_5797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1438 a_13311_5842# d0 a_13802_5835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1439 a_4753_720# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1440 a_116_714# a_3343_1171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1441 a_13712_745# d1 a_14509_973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1442 gnd d0 a_16795_6109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1443 a_1203_1953# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1444 a_4480_727# a_4482_826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1445 a_1659_6433# a_1441_6433# a_1560_6433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1446 a_15568_2001# a_15825_1811# a_15522_3021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1447 a_13785_4817# d1 a_14582_5045# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1448 a_15667_2411# d0 a_16465_2227# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1449 a_15595_7093# d2 a_15641_6073# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1450 a_7040_8317# a_7293_8304# a_6941_7907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1451 a_5061_5810# d1 a_5846_5549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1452 a_3346_1406# a_3599_1393# a_2549_1178# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1453 a_4970_1132# a_4752_1132# a_4489_1044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1454 a_16557_7729# a_16561_7552# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1455 a_4607_7853# a_4609_7952# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1456 a_1404_935# a_1186_935# a_607_707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1457 a_4585_6317# a_4590_6641# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1458 a_3397_4225# a_3401_4048# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1459 a_3419_5478# a_3672_5465# a_2622_5250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1460 gnd d0 a_3654_4035# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1461 a_10218_5032# a_10000_5032# a_9421_4804# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1462 a_118_813# d0 a_607_707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1463 a_7744_3220# a_7748_3043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1464 a_7764_4473# a_8017_4460# a_6967_4245# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1465 a_2599_4409# a_2856_4219# a_2504_3822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1466 a_14381_6063# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 a_15764_7324# d0 a_16557_7729# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1468 gnd d0 a_12468_8132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 a_4526_3080# d0 a_5007_3168# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1470 a_15609_3860# a_15862_3847# a_15526_2844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1471 a_9239_7252# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1472 a_1492_2480# a_1322_3381# a_1441_2971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1473 a_9167_2768# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1474 a_4590_6641# d0 a_5081_6828# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1475 a_10026_1370# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1476 a_4790_2756# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1477 a_7748_3043# a_8001_3030# a_6946_3404# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_3415_5655# a_3672_5465# a_2622_5250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1479 a_16484_3657# a_16741_3467# a_15691_3252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1480 vdd d0 a_3654_4035# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1481 a_10063_3406# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1482 a_425_3155# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1483 a_7760_4650# a_8017_4460# a_6967_4245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1484 gnd d0 a_16777_5503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1485 a_7748_3043# a_7743_3632# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1486 a_9981_4014# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1487 a_170_3768# d0 a_661_3761# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1488 a_2639_6268# d0 a_3432_6673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1489 a_13530_3193# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1490 a_499_6815# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1491 a_9944_1978# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1492 a_6986_5263# a_7239_5250# a_6900_6048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1493 a_13604_6853# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1494 vdd d0 a_12468_8132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1495 a_643_3155# a_425_3155# a_168_3250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1496 a_14328_3009# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1497 a_2562_2373# d0 a_3360_2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1498 a_11162_2831# d2 a_11245_3847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1499 a_717_6815# a_499_6815# a_228_6921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1500 a_13363_8378# a_12214_8557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1501 a_13766_3799# d1 a_14551_3538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1502 a_2545_1355# d0 a_3343_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1503 a_16541_6534# a_16558_7317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1504 a_13822_6853# a_13604_6853# a_13333_6959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1505 a_7744_3220# a_8001_3030# a_6946_3404# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1506 a_13309_5324# a_13311_5842# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1507 a_9348_732# a_9130_732# a_8859_838# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1508 a_2672_8481# d0 a_3474_8120# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1509 a_5098_7846# a_4880_7846# a_4609_7952# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1510 a_14546_3009# a_14328_3009# a_13748_3193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1511 gnd d0 a_8037_5066# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1512 a_3400_4460# a_3653_4447# a_2603_4232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1513 a_2639_6268# d0 a_3436_6496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1514 a_8889_2257# d0 a_9364_2162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1515 a_12083_1608# a_12340_1418# a_11290_1203# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1516 a_13320_6159# d0 a_13801_6247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1517 a_14509_973# d2 a_14592_2399# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1518 a_6854_7068# d2 a_6900_6048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1519 a_10187_3525# a_9981_4014# a_9402_3786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1520 a_9146_2162# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1521 a_6982_5440# a_7239_5250# a_6900_6048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1522 a_2318_4844# a_2571_4831# a_1721_131# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1523 a_13765_4211# a_13547_4211# a_13284_4123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1524 a_9347_1144# a_9129_1144# a_8866_1056# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1525 a_6986_5263# d0 a_7783_5491# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1526 a_12214_8557# a_12467_8544# a_11417_8329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1527 a_9420_5216# a_9202_5216# a_8939_5128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1528 a_8872_1239# a_8874_1757# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1529 a_4843_5810# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1530 a_7003_6281# d0 a_7800_6509# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1531 vdd d1 a_11560_2208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1532 gnd d0 a_16794_6521# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1533 a_10327_2386# a_10109_2386# a_10228_2386# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1534 a_5950_2374# d4 a_6090_263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1535 a_10400_6458# d4 a_10467_275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1536 a_406_1725# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1537 vdd d0 a_8037_5066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1538 a_12197_7539# a_12211_8322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1539 a_5623_5020# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_10400_6458# a_10182_6458# a_10301_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1541 a_13511_1763# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1542 vdd d2 a_7157_5858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1543 a_12125_3055# a_12378_3042# a_11323_3416# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1544 a_6909_1368# d0 a_7711_1007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1545 gnd d2 a_15898_5883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1546 a_11314_8096# d1 a_11396_7488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1547 gnd d0 a_16758_4485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1548 a_10467_275# d5 a_10561_156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1549 a_2622_5250# a_2875_5237# a_2536_6035# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1550 a_5846_5549# a_5640_6038# a_5060_6222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1551 a_12198_7127# a_12451_7114# a_11396_7488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1552 a_14291_973# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1553 a_15522_3021# d2 a_15568_2001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 a_10037_7068# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1555 a_13238_1770# a_13240_1869# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1556 a_6904_5871# d1 a_7003_6281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1557 a_12210_8734# a_12467_8544# a_11417_8329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1558 a_125_1031# a_131_1214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1559 vdd d0 a_16794_6521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1560 a_13326_6342# a_13331_6666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1561 a_15522_3021# a_15779_2831# a_15419_5059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1562 a_6967_4245# d0 a_7760_4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1563 a_13294_4824# a_13296_4923# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1564 a_4789_3168# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1565 gnd d0 a_16742_3055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1566 a_15595_7093# a_15852_6903# a_15423_4882# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1567 a_12121_3232# a_12378_3042# a_11323_3416# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1568 a_7783_5491# a_8036_5478# a_6986_5263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1569 a_11208_1811# a_11461_1798# a_11158_3008# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1570 gnd d0 a_8018_4048# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 vdd d0 a_16758_4485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1572 a_5007_3168# a_4789_3168# a_4532_3263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1573 a_245_7939# d0 a_734_7833# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1574 a_16558_7317# a_16562_7140# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1575 a_15687_3429# a_15944_3239# a_15605_4037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1576 a_12125_3055# a_12120_3644# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1577 a_3432_6673# a_3436_6496# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1578 a_12194_7304# a_12451_7114# a_11396_7488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1579 a_5008_2756# d1 a_5805_2984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1580 a_10306_6577# a_10136_7478# a_10260_7597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1581 a_11340_4434# d0 a_12138_4250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1582 a_1477_5007# d2 a_1560_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1583 gnd d0 a_12357_2436# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1584 a_16542_6122# a_16795_6109# a_15740_6483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1585 a_2540_5858# d1 a_2635_6445# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 a_11413_8506# d0 a_12211_8322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 gnd d0 a_12413_5490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1588 a_5768_948# a_5550_948# a_4971_720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1589 a_623_2137# d1 a_1409_1464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_9384_3180# a_9166_3180# a_8903_3092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1591 a_6967_4245# d0 a_7764_4473# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1592 a_5649_1358# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1593 a_5097_8258# d1 a_5883_7585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1594 a_13822_6853# d1 a_14619_7081# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1595 a_9458_6840# a_9240_6840# a_8967_6653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1596 vdd d0 a_16742_3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1597 a_5722_5430# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1598 a_2566_2196# d0 a_3359_2601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1599 a_5604_4002# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1600 a_189_4786# d0 a_680_4779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1601 a_14587_5574# d2 a_14665_6471# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1602 a_1492_2480# d3 a_1586_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1603 a_11340_4434# d0 a_12142_4073# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1604 a_2586_3214# a_2839_3201# a_2500_3999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1605 a_5846_5549# d2 a_5924_6446# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 vdd d0 a_12357_2436# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1607 a_2540_5858# d1 a_2639_6268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1608 a_15609_3860# d1 a_15708_4270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1609 a_2603_4232# a_2856_4219# a_2504_3822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1610 a_11413_8506# d0 a_12215_8145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1611 a_11286_1380# a_11543_1190# a_11204_1988# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1612 a_10182_2996# a_9964_2996# a_9384_3180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1613 a_1544_4395# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1614 a_1441_6433# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1615 a_2659_7286# a_2912_7273# a_2573_8071# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1616 a_5810_3513# a_5604_4002# a_5024_4186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1617 a_8982_7347# a_8984_7865# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1618 a_5732_2374# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1619 a_479_5797# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1620 a_2566_2196# d0 a_3363_2424# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1621 a_15760_7501# d0 a_16562_7140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1622 a_2490_7055# a_2747_6865# a_2318_4844# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1623 a_16488_3480# a_16741_3467# a_15691_3252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1624 a_5908_4408# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1625 a_478_6209# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1626 a_4512_2245# d0 a_4987_2150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1627 a_13583_6247# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1628 a_6678_5034# a_6935_4844# a_6085_144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1629 a_14546_6471# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1630 a_14390_1383# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1631 a_4572_5916# d0 a_5061_5810# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1632 a_13784_5229# a_13566_5229# a_13303_5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1633 a_7801_6097# a_7796_6686# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1634 a_3343_1171# a_3347_994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1635 a_4536_3880# a_4543_4098# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1636 a_2655_7463# a_2912_7273# a_2573_8071# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1637 vdd d1 a_7183_2196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1638 a_11208_1811# d1 a_11307_2221# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1639 gnd d0 a_12394_4472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1640 a_2577_7894# d1 a_2672_8481# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1641 a_8993_8182# d0 a_9474_8270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1642 vdd d1 a_15997_6293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1643 a_14764_6471# d4 a_14831_288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1644 a_13363_8378# d0 a_13838_8283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1645 a_11158_3008# a_11415_2818# a_11055_5046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1646 a_15708_4270# d0 a_16501_4675# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1647 a_12087_1431# a_12340_1418# a_11290_1203# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1648 a_11059_4869# d3 a_11231_7080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_7727_2437# a_7980_2424# a_6930_2209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1650 a_10462_156# d4 a_11059_4869# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1651 a_12137_4662# a_12141_4485# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1652 a_4489_1044# a_4495_1227# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1653 a_4534_3781# d0 a_5025_3774# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1654 vdd d0 a_12394_4472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1655 a_6986_5263# d0 a_7779_5668# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1656 a_16541_6534# a_16794_6521# a_15744_6306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 gnd d1 a_11616_5262# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1658 gnd d2 a_7121_3822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1659 a_12178_6109# a_12431_6096# a_11376_6470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1660 a_443_3761# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1661 a_6864_4012# a_7121_3822# a_6785_2819# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1662 a_15708_4270# d0 a_16505_4498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1663 a_1285_1345# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1664 a_15568_2001# d1 a_15650_1393# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1665 a_7723_2614# a_7980_2424# a_6930_2209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1666 a_15645_5896# a_15898_5883# a_15595_7093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1667 a_13260_2887# a_13267_3105# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1668 a_3384_3030# a_3379_3619# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1669 a_16505_4498# a_16521_5281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1670 a_10255_7068# a_10037_7068# a_9458_6840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1671 a_5883_7585# a_5677_8074# a_5098_7846# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1672 a_16464_2639# a_16468_2462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1673 a_15641_6073# d1 a_15723_5465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1674 a_679_5191# d1 a_1477_5007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1675 a_179_4085# a_185_4268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1676 a_13712_745# a_13494_745# a_13221_752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1677 a_4826_4792# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1678 a_6904_5871# d1 a_6999_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1679 a_1203_1953# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1680 a_10099_5442# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1681 a_16537_6711# a_16794_6521# a_15744_6306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1682 a_4825_5204# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1683 a_5080_7240# a_4862_7240# a_4599_7152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1684 a_10228_2386# d3 a_10327_2386# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1685 vdd d1 a_11616_5262# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1686 a_14401_7081# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1687 a_9348_732# d1 a_10145_960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1688 a_9347_1144# d1 a_10145_960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1689 a_10017_6050# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1690 a_4988_1738# d1 a_5773_1477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1691 vdd d1 a_2875_5237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1692 a_10561_156# a_10343_156# a_10462_156# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1693 a_462_4779# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1694 a_14463_5455# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1695 a_4971_720# a_4753_720# a_4482_826# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1696 a_5856_2493# d3 a_5950_2374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_1446_3500# d2 a_1492_2480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1698 a_15641_6073# d1 a_15727_5288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1699 a_3453_7279# a_3457_7102# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1700 a_15691_3252# a_15944_3239# a_15605_4037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1701 a_5841_5020# a_5623_5020# a_5043_5204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1702 a_12100_2626# a_12104_2449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1703 a_13802_5835# d1 a_14587_5574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1704 a_4553_4799# d0 a_5044_4792# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1705 a_1519_7572# d2 a_1565_6552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1706 a_12178_6109# a_12173_6698# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1707 a_8896_2874# a_8903_3092# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1708 gnd d4 a_15676_4869# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1709 a_14665_6471# a_14463_5455# a_14587_5574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1710 a_4987_2150# a_4769_2150# a_4506_2062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_6678_5034# d3 a_6781_2996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1712 a_1482_5536# a_1276_6025# a_697_5797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1713 a_14514_1502# a_14308_1991# a_13729_1763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1714 a_6950_3227# d0 a_7743_3632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_3436_6496# a_3689_6483# a_2639_6268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1716 a_2318_4844# d3 a_2490_7055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1717 a_1726_250# a_1544_4395# a_1659_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1718 gnd d1 a_11597_4244# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 a_6085_144# d4 a_6678_5034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1720 a_16542_6122# a_16537_6711# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1721 a_10150_1489# a_9944_1978# a_9364_2162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1722 vdd d0 a_3636_3429# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1723 a_16451_1444# a_16465_2227# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1724 a_3457_7102# a_3452_7691# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1725 a_14826_169# d5 a_12951_82# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1726 a_235_7139# d0 a_716_7227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1727 a_11241_4024# a_11498_3834# a_11162_2831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1728 vdd d2 a_15825_1811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1729 a_14546_3009# d2 a_14597_2518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1730 a_11314_8096# a_11571_7906# a_11235_6903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1731 a_15609_3860# d1 a_15704_4447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_3420_5066# a_3673_5053# a_2618_5427# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1733 a_14831_288# a_14649_4433# a_14691_2399# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1734 a_4616_8170# d0 a_5097_8258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1735 a_13296_4923# a_13303_5141# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1736 a_7724_2202# a_7728_2025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1737 a_5805_2984# d2 a_5856_2493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1738 a_9257_7858# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1739 a_4807_3774# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1740 a_6950_3227# d0 a_7747_3455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1741 a_3432_6673# a_3689_6483# a_2639_6268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1742 a_1296_7043# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1743 a_4880_7846# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 a_4806_4186# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1745 vdd d1 a_11597_4244# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1746 a_16574_8747# a_16831_8557# a_15781_8342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1747 a_15760_7501# d0 a_16558_7317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1748 a_515_8245# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1749 a_10561_156# d6 a_8658_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1750 a_5025_3774# a_4807_3774# a_4536_3880# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1751 vdd d1 a_2856_4219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1752 a_5660_7056# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1753 a_13620_8283# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1754 a_13230_1069# a_13236_1252# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1755 a_8945_5311# d0 a_9420_5216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1756 gnd d2 a_15862_3847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1757 a_8859_838# a_8866_1056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1758 a_3416_5243# a_3673_5053# a_2618_5427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1759 a_733_8245# a_515_8245# a_258_8340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1760 a_13303_5141# a_13309_5324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1761 a_13839_7871# a_13621_7871# a_13350_7977# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1762 a_6785_2819# d2 a_6868_3835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1763 a_7761_4238# a_8018_4048# a_6963_4422# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1764 gnd d0 a_16778_5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_10306_6577# d3 a_10400_6458# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_11204_1988# d1 a_11286_1380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_131_1214# d0 a_606_1119# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1768 a_2635_6445# d0 a_3433_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_11281_5883# a_11534_5870# a_11231_7080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1770 a_13494_745# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1771 a_2549_1178# d0 a_3346_1406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1772 a_12084_1196# a_12088_1019# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1773 a_14624_7610# a_14418_8099# a_13838_8283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1774 a_13296_4923# d0 a_13785_4817# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1775 a_15740_6483# a_15997_6293# a_15645_5896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1776 a_10000_5032# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1777 a_15599_6916# d2 a_15682_7932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1778 a_8658_81# a_12832_82# a_12951_82# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1779 a_241_7322# a_243_7840# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1780 gnd d2 a_2757_3809# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1781 a_12173_6698# a_12430_6508# a_11380_6293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1782 a_3420_5066# a_3415_5655# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1783 a_4752_1132# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1784 a_10145_960# a_9927_960# a_9348_732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1785 a_13313_5941# a_13320_6159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
C0 vdd gnd 4.85fF
C1 a_1721_131# a_1726_250# 5.60fF
C2 a_14826_169# a_14831_288# 5.60fF
C3 d0 gnd 9.63fF
C4 d2 gnd 2.53fF
C5 d0 vdd 3.61fF
C6 a_10462_156# a_10467_275# 5.60fF
C7 d1 gnd 5.06fF
C8 d1 vdd 2.14fF
C9 a_6085_144# a_6090_263# 5.60fF
C10 gnd SUB 55.31fF
C11 a_12951_82# SUB 3.15fF
C12 vdd SUB 238.89fF
C13 a_10561_156# SUB 3.77fF
C14 a_4210_57# SUB 3.15fF
C15 a_4309_57# SUB 5.69fF
C16 a_1820_131# SUB 3.77fF
C17 d5 SUB 2.25fF
C18 a_13221_752# SUB 5.34fF
C19 d0 SUB 78.42fF
C20 a_8857_739# SUB 5.34fF
C21 a_4480_727# SUB 5.34fF
C22 a_116_714# SUB 5.34fF
C23 a_13712_745# SUB 2.21fF
C24 d1 SUB 40.89fF
C25 a_13711_1157# SUB 2.30fF
C26 a_4971_720# SUB 2.21fF
C27 a_15650_1393# SUB 2.30fF
C28 a_9347_1144# SUB 2.30fF
C29 a_607_707# SUB 2.21fF
C30 a_11286_1380# SUB 2.30fF
C31 a_4970_1132# SUB 2.30fF
C32 a_6909_1368# SUB 2.30fF
C33 a_606_1119# SUB 2.30fF
C34 d2 SUB 18.36fF
C35 a_15654_1216# SUB 2.21fF
C36 a_2545_1355# SUB 2.30fF
C37 a_11290_1203# SUB 2.21fF
C38 a_6913_1191# SUB 2.21fF
C39 a_2549_1178# SUB 2.21fF
C40 a_13729_1763# SUB 2.21fF
C41 a_9365_1750# SUB 2.21fF
C42 a_13728_2175# SUB 2.30fF
C43 a_4988_1738# SUB 2.21fF
C44 a_624_1725# SUB 2.21fF
C45 a_15667_2411# SUB 2.30fF
C46 a_4987_2150# SUB 2.30fF
C47 a_11303_2398# SUB 2.30fF
C48 a_14592_2399# SUB 2.37fF
C49 a_623_2137# SUB 2.30fF
C50 a_6926_2386# SUB 2.30fF
C51 d3 SUB 11.41fF
C52 a_15671_2234# SUB 2.21fF
C53 a_10228_2386# SUB 2.37fF
C54 a_2562_2373# SUB 2.30fF
C55 a_11307_2221# SUB 2.21fF
C56 a_5851_2374# SUB 2.37fF
C57 a_6930_2209# SUB 2.21fF
C58 a_1487_2361# SUB 2.37fF
C59 a_2566_2196# SUB 2.21fF
C60 a_13749_2781# SUB 2.21fF
C61 a_9385_2768# SUB 2.21fF
C62 a_13748_3193# SUB 2.30fF
C63 a_5008_2756# SUB 2.21fF
C64 a_15687_3429# SUB 2.30fF
C65 a_9384_3180# SUB 2.30fF
C66 a_644_2743# SUB 2.21fF
C67 a_11323_3416# SUB 2.30fF
C68 a_5007_3168# SUB 2.30fF
C69 a_6946_3404# SUB 2.30fF
C70 a_643_3155# SUB 2.30fF
C71 a_15691_3252# SUB 2.21fF
C72 a_2582_3391# SUB 2.30fF
C73 a_11327_3239# SUB 2.21fF
C74 a_6950_3227# SUB 2.21fF
C75 a_2586_3214# SUB 2.21fF
C76 a_15526_2844# SUB 2.63fF
C77 a_11162_2831# SUB 2.63fF
C78 a_13766_3799# SUB 2.21fF
C79 a_6785_2819# SUB 2.63fF
C80 a_9402_3786# SUB 2.21fF
C81 a_2421_2806# SUB 2.63fF
C82 a_13765_4211# SUB 2.30fF
C83 a_5025_3774# SUB 2.21fF
C84 a_9401_4198# SUB 2.30fF
C85 a_661_3761# SUB 2.21fF
C86 a_15704_4447# SUB 2.30fF
C87 a_5024_4186# SUB 2.30fF
C88 a_11340_4434# SUB 2.30fF
C89 a_14691_2399# SUB 4.04fF
C90 a_14831_288# SUB 5.00fF
C91 a_660_4173# SUB 2.30fF
C92 a_6963_4422# SUB 2.30fF
C93 d4 SUB 5.48fF
C94 a_15708_4270# SUB 2.21fF
C95 a_10327_2386# SUB 4.04fF
C96 a_10467_275# SUB 5.00fF
C97 a_2599_4409# SUB 2.30fF
C98 a_11344_4257# SUB 2.21fF
C99 a_5950_2374# SUB 4.04fF
C100 a_6090_263# SUB 5.00fF
C101 a_6967_4245# SUB 2.21fF
C102 a_1586_2361# SUB 4.04fF
C103 a_1726_250# SUB 5.00fF
C104 a_2603_4232# SUB 2.21fF
C105 a_14826_169# SUB 5.75fF
C106 a_15419_5059# SUB 2.94fF
C107 a_10462_156# SUB 5.75fF
C108 a_11055_5046# SUB 2.94fF
C109 a_13785_4817# SUB 2.21fF
C110 a_6085_144# SUB 5.75fF
C111 a_6678_5034# SUB 2.94fF
C112 a_9421_4804# SUB 2.21fF
C113 a_1721_131# SUB 5.75fF
C114 a_2314_5021# SUB 2.94fF
C115 a_13784_5229# SUB 2.30fF
C116 a_5044_4792# SUB 2.21fF
C117 a_15723_5465# SUB 2.30fF
C118 a_9420_5216# SUB 2.30fF
C119 a_680_4779# SUB 2.21fF
C120 a_11359_5452# SUB 2.30fF
C121 a_5043_5204# SUB 2.30fF
C122 a_6982_5440# SUB 2.30fF
C123 a_679_5191# SUB 2.30fF
C124 a_15727_5288# SUB 2.21fF
C125 a_2618_5427# SUB 2.30fF
C126 a_11363_5275# SUB 2.21fF
C127 a_6986_5263# SUB 2.21fF
C128 a_2622_5250# SUB 2.21fF
C129 a_13802_5835# SUB 2.21fF
C130 a_9438_5822# SUB 2.21fF
C131 a_13801_6247# SUB 2.30fF
C132 a_9437_6234# SUB 2.30fF
C133 a_697_5797# SUB 2.21fF
C134 a_15740_6483# SUB 2.30fF
C135 a_5060_6222# SUB 2.30fF
C136 a_11376_6470# SUB 2.30fF
C137 a_14665_6471# SUB 2.63fF
C138 a_14764_6471# SUB 2.94fF
C139 a_696_6209# SUB 2.30fF
C140 a_6999_6458# SUB 2.30fF
C141 a_15744_6306# SUB 2.21fF
C142 a_10301_6458# SUB 2.63fF
C143 a_10400_6458# SUB 2.94fF
C144 a_2635_6445# SUB 2.30fF
C145 a_11380_6293# SUB 2.21fF
C146 a_5924_6446# SUB 2.63fF
C147 a_6023_6446# SUB 2.94fF
C148 a_7003_6281# SUB 2.21fF
C149 a_1560_6433# SUB 2.63fF
C150 a_1659_6433# SUB 2.94fF
C151 a_2639_6268# SUB 2.21fF
C152 a_15423_4882# SUB 4.03fF
C153 a_11059_4869# SUB 4.03fF
C154 a_13822_6853# SUB 2.21fF
C155 a_6682_4857# SUB 4.03fF
C156 a_9458_6840# SUB 2.21fF
C157 a_2318_4844# SUB 4.03fF
C158 a_13821_7265# SUB 2.30fF
C159 a_5081_6828# SUB 2.21fF
C160 a_15760_7501# SUB 2.30fF
C161 a_9457_7252# SUB 2.30fF
C162 a_717_6815# SUB 2.21fF
C163 a_11396_7488# SUB 2.30fF
C164 a_7019_7476# SUB 2.30fF
C165 a_716_7227# SUB 2.30fF
C166 a_15764_7324# SUB 2.21fF
C167 a_2655_7463# SUB 2.30fF
C168 a_11400_7311# SUB 2.21fF
C169 a_7023_7299# SUB 2.21fF
C170 a_2659_7286# SUB 2.21fF
C171 a_15599_6916# SUB 2.37fF
C172 a_11235_6903# SUB 2.37fF
C173 a_13839_7871# SUB 2.21fF
C174 a_6858_6891# SUB 2.37fF
C175 a_9475_7858# SUB 2.21fF
C176 a_2494_6878# SUB 2.37fF
C177 a_13838_8283# SUB 2.30fF
C178 a_9474_8270# SUB 2.30fF
C179 a_734_7833# SUB 2.21fF
C180 a_5097_8258# SUB 2.30fF
C181 a_733_8245# SUB 2.30fF
C182 a_15777_8519# SUB 2.30fF
C183 a_11413_8506# SUB 2.30fF
C184 a_7036_8494# SUB 2.30fF
C185 a_15781_8342# SUB 2.21fF
C186 a_2672_8481# SUB 2.30fF
C187 a_12214_8557# SUB 2.31fF
C188 a_11417_8329# SUB 2.21fF
C189 a_7837_8545# SUB 2.54fF
C190 a_7040_8317# SUB 2.21fF
C191 a_3473_8532# SUB 2.31fF
C192 a_2676_8304# SUB 2.21fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40ns 80ns)
Vd4 d4 0 pulse(0 1.8 0ns 0.1ns 0.1ns 80ns 160ns)
Vd5 d5 0 pulse(0 1.8 0ns 0.1ns 0.1ns 160ns 320ns)
Vd6 d6 0 pulse(0 1.8 0ns 0.1ns 0.1ns 320ns 640ns)
Vd7 d7 0 pulse(0 1.8 0ns 0.1ns 0.1ns 640ns 1280ns)


.tran 5ns 1280ns
.control
run
plot V(vout) 
.endc
.end

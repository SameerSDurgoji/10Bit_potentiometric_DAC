magic
tech sky130A
timestamp 1616088573
<< nwell >>
rect 291 1612 899 1762
rect 1089 1428 1697 1578
rect 292 1200 900 1350
rect 1171 820 1779 970
rect 274 594 882 744
rect 1072 410 1680 560
rect 275 182 883 332
rect 1217 -200 1825 -50
rect 254 -424 862 -274
rect 1052 -608 1660 -458
rect 255 -836 863 -686
rect 1134 -1216 1742 -1066
rect 237 -1442 845 -1292
rect 1035 -1626 1643 -1476
rect 238 -1854 846 -1704
<< nmos >>
rect 355 1511 405 1553
rect 573 1511 623 1553
rect 781 1511 831 1553
rect 1153 1327 1203 1369
rect 1371 1327 1421 1369
rect 1579 1327 1629 1369
rect 356 1099 406 1141
rect 574 1099 624 1141
rect 782 1099 832 1141
rect 1235 719 1285 761
rect 1453 719 1503 761
rect 1661 719 1711 761
rect 338 493 388 535
rect 556 493 606 535
rect 764 493 814 535
rect 1136 309 1186 351
rect 1354 309 1404 351
rect 1562 309 1612 351
rect 339 81 389 123
rect 557 81 607 123
rect 765 81 815 123
rect 1281 -301 1331 -259
rect 1499 -301 1549 -259
rect 1707 -301 1757 -259
rect 318 -525 368 -483
rect 536 -525 586 -483
rect 744 -525 794 -483
rect 1116 -709 1166 -667
rect 1334 -709 1384 -667
rect 1542 -709 1592 -667
rect 319 -937 369 -895
rect 537 -937 587 -895
rect 745 -937 795 -895
rect 1198 -1317 1248 -1275
rect 1416 -1317 1466 -1275
rect 1624 -1317 1674 -1275
rect 301 -1543 351 -1501
rect 519 -1543 569 -1501
rect 727 -1543 777 -1501
rect 1099 -1727 1149 -1685
rect 1317 -1727 1367 -1685
rect 1525 -1727 1575 -1685
rect 302 -1955 352 -1913
rect 520 -1955 570 -1913
rect 728 -1955 778 -1913
<< pmos >>
rect 355 1630 405 1730
rect 573 1630 623 1730
rect 781 1630 831 1730
rect 1153 1446 1203 1546
rect 1371 1446 1421 1546
rect 1579 1446 1629 1546
rect 356 1218 406 1318
rect 574 1218 624 1318
rect 782 1218 832 1318
rect 1235 838 1285 938
rect 1453 838 1503 938
rect 1661 838 1711 938
rect 338 612 388 712
rect 556 612 606 712
rect 764 612 814 712
rect 1136 428 1186 528
rect 1354 428 1404 528
rect 1562 428 1612 528
rect 339 200 389 300
rect 557 200 607 300
rect 765 200 815 300
rect 1281 -182 1331 -82
rect 1499 -182 1549 -82
rect 1707 -182 1757 -82
rect 318 -406 368 -306
rect 536 -406 586 -306
rect 744 -406 794 -306
rect 1116 -590 1166 -490
rect 1334 -590 1384 -490
rect 1542 -590 1592 -490
rect 319 -818 369 -718
rect 537 -818 587 -718
rect 745 -818 795 -718
rect 1198 -1198 1248 -1098
rect 1416 -1198 1466 -1098
rect 1624 -1198 1674 -1098
rect 301 -1424 351 -1324
rect 519 -1424 569 -1324
rect 727 -1424 777 -1324
rect 1099 -1608 1149 -1508
rect 1317 -1608 1367 -1508
rect 1525 -1608 1575 -1508
rect 302 -1836 352 -1736
rect 520 -1836 570 -1736
rect 728 -1836 778 -1736
<< ndiff >>
rect 306 1543 355 1553
rect 306 1523 317 1543
rect 337 1523 355 1543
rect 306 1511 355 1523
rect 405 1547 449 1553
rect 405 1527 420 1547
rect 440 1527 449 1547
rect 405 1511 449 1527
rect 524 1543 573 1553
rect 524 1523 535 1543
rect 555 1523 573 1543
rect 524 1511 573 1523
rect 623 1547 667 1553
rect 623 1527 638 1547
rect 658 1527 667 1547
rect 623 1511 667 1527
rect 737 1547 781 1553
rect 737 1527 746 1547
rect 766 1527 781 1547
rect 737 1511 781 1527
rect 831 1543 880 1553
rect 831 1523 849 1543
rect 869 1523 880 1543
rect 831 1511 880 1523
rect 1104 1359 1153 1369
rect 1104 1339 1115 1359
rect 1135 1339 1153 1359
rect 1104 1327 1153 1339
rect 1203 1363 1247 1369
rect 1203 1343 1218 1363
rect 1238 1343 1247 1363
rect 1203 1327 1247 1343
rect 1322 1359 1371 1369
rect 1322 1339 1333 1359
rect 1353 1339 1371 1359
rect 1322 1327 1371 1339
rect 1421 1363 1465 1369
rect 1421 1343 1436 1363
rect 1456 1343 1465 1363
rect 1421 1327 1465 1343
rect 1535 1363 1579 1369
rect 1535 1343 1544 1363
rect 1564 1343 1579 1363
rect 1535 1327 1579 1343
rect 1629 1359 1678 1369
rect 1629 1339 1647 1359
rect 1667 1339 1678 1359
rect 1629 1327 1678 1339
rect 307 1131 356 1141
rect 307 1111 318 1131
rect 338 1111 356 1131
rect 307 1099 356 1111
rect 406 1135 450 1141
rect 406 1115 421 1135
rect 441 1115 450 1135
rect 406 1099 450 1115
rect 525 1131 574 1141
rect 525 1111 536 1131
rect 556 1111 574 1131
rect 525 1099 574 1111
rect 624 1135 668 1141
rect 624 1115 639 1135
rect 659 1115 668 1135
rect 624 1099 668 1115
rect 738 1135 782 1141
rect 738 1115 747 1135
rect 767 1115 782 1135
rect 738 1099 782 1115
rect 832 1131 881 1141
rect 832 1111 850 1131
rect 870 1111 881 1131
rect 832 1099 881 1111
rect 1186 751 1235 761
rect 1186 731 1197 751
rect 1217 731 1235 751
rect 1186 719 1235 731
rect 1285 755 1329 761
rect 1285 735 1300 755
rect 1320 735 1329 755
rect 1285 719 1329 735
rect 1404 751 1453 761
rect 1404 731 1415 751
rect 1435 731 1453 751
rect 1404 719 1453 731
rect 1503 755 1547 761
rect 1503 735 1518 755
rect 1538 735 1547 755
rect 1503 719 1547 735
rect 1617 755 1661 761
rect 1617 735 1626 755
rect 1646 735 1661 755
rect 1617 719 1661 735
rect 1711 751 1760 761
rect 1711 731 1729 751
rect 1749 731 1760 751
rect 1711 719 1760 731
rect 289 525 338 535
rect 289 505 300 525
rect 320 505 338 525
rect 289 493 338 505
rect 388 529 432 535
rect 388 509 403 529
rect 423 509 432 529
rect 388 493 432 509
rect 507 525 556 535
rect 507 505 518 525
rect 538 505 556 525
rect 507 493 556 505
rect 606 529 650 535
rect 606 509 621 529
rect 641 509 650 529
rect 606 493 650 509
rect 720 529 764 535
rect 720 509 729 529
rect 749 509 764 529
rect 720 493 764 509
rect 814 525 863 535
rect 814 505 832 525
rect 852 505 863 525
rect 814 493 863 505
rect 1087 341 1136 351
rect 1087 321 1098 341
rect 1118 321 1136 341
rect 1087 309 1136 321
rect 1186 345 1230 351
rect 1186 325 1201 345
rect 1221 325 1230 345
rect 1186 309 1230 325
rect 1305 341 1354 351
rect 1305 321 1316 341
rect 1336 321 1354 341
rect 1305 309 1354 321
rect 1404 345 1448 351
rect 1404 325 1419 345
rect 1439 325 1448 345
rect 1404 309 1448 325
rect 1518 345 1562 351
rect 1518 325 1527 345
rect 1547 325 1562 345
rect 1518 309 1562 325
rect 1612 341 1661 351
rect 1612 321 1630 341
rect 1650 321 1661 341
rect 1612 309 1661 321
rect 290 113 339 123
rect 290 93 301 113
rect 321 93 339 113
rect 290 81 339 93
rect 389 117 433 123
rect 389 97 404 117
rect 424 97 433 117
rect 389 81 433 97
rect 508 113 557 123
rect 508 93 519 113
rect 539 93 557 113
rect 508 81 557 93
rect 607 117 651 123
rect 607 97 622 117
rect 642 97 651 117
rect 607 81 651 97
rect 721 117 765 123
rect 721 97 730 117
rect 750 97 765 117
rect 721 81 765 97
rect 815 113 864 123
rect 815 93 833 113
rect 853 93 864 113
rect 815 81 864 93
rect 1232 -269 1281 -259
rect 1232 -289 1243 -269
rect 1263 -289 1281 -269
rect 1232 -301 1281 -289
rect 1331 -265 1375 -259
rect 1331 -285 1346 -265
rect 1366 -285 1375 -265
rect 1331 -301 1375 -285
rect 1450 -269 1499 -259
rect 1450 -289 1461 -269
rect 1481 -289 1499 -269
rect 1450 -301 1499 -289
rect 1549 -265 1593 -259
rect 1549 -285 1564 -265
rect 1584 -285 1593 -265
rect 1549 -301 1593 -285
rect 1663 -265 1707 -259
rect 1663 -285 1672 -265
rect 1692 -285 1707 -265
rect 1663 -301 1707 -285
rect 1757 -269 1806 -259
rect 1757 -289 1775 -269
rect 1795 -289 1806 -269
rect 1757 -301 1806 -289
rect 269 -493 318 -483
rect 269 -513 280 -493
rect 300 -513 318 -493
rect 269 -525 318 -513
rect 368 -489 412 -483
rect 368 -509 383 -489
rect 403 -509 412 -489
rect 368 -525 412 -509
rect 487 -493 536 -483
rect 487 -513 498 -493
rect 518 -513 536 -493
rect 487 -525 536 -513
rect 586 -489 630 -483
rect 586 -509 601 -489
rect 621 -509 630 -489
rect 586 -525 630 -509
rect 700 -489 744 -483
rect 700 -509 709 -489
rect 729 -509 744 -489
rect 700 -525 744 -509
rect 794 -493 843 -483
rect 794 -513 812 -493
rect 832 -513 843 -493
rect 794 -525 843 -513
rect 1067 -677 1116 -667
rect 1067 -697 1078 -677
rect 1098 -697 1116 -677
rect 1067 -709 1116 -697
rect 1166 -673 1210 -667
rect 1166 -693 1181 -673
rect 1201 -693 1210 -673
rect 1166 -709 1210 -693
rect 1285 -677 1334 -667
rect 1285 -697 1296 -677
rect 1316 -697 1334 -677
rect 1285 -709 1334 -697
rect 1384 -673 1428 -667
rect 1384 -693 1399 -673
rect 1419 -693 1428 -673
rect 1384 -709 1428 -693
rect 1498 -673 1542 -667
rect 1498 -693 1507 -673
rect 1527 -693 1542 -673
rect 1498 -709 1542 -693
rect 1592 -677 1641 -667
rect 1592 -697 1610 -677
rect 1630 -697 1641 -677
rect 1592 -709 1641 -697
rect 270 -905 319 -895
rect 270 -925 281 -905
rect 301 -925 319 -905
rect 270 -937 319 -925
rect 369 -901 413 -895
rect 369 -921 384 -901
rect 404 -921 413 -901
rect 369 -937 413 -921
rect 488 -905 537 -895
rect 488 -925 499 -905
rect 519 -925 537 -905
rect 488 -937 537 -925
rect 587 -901 631 -895
rect 587 -921 602 -901
rect 622 -921 631 -901
rect 587 -937 631 -921
rect 701 -901 745 -895
rect 701 -921 710 -901
rect 730 -921 745 -901
rect 701 -937 745 -921
rect 795 -905 844 -895
rect 795 -925 813 -905
rect 833 -925 844 -905
rect 795 -937 844 -925
rect 1149 -1285 1198 -1275
rect 1149 -1305 1160 -1285
rect 1180 -1305 1198 -1285
rect 1149 -1317 1198 -1305
rect 1248 -1281 1292 -1275
rect 1248 -1301 1263 -1281
rect 1283 -1301 1292 -1281
rect 1248 -1317 1292 -1301
rect 1367 -1285 1416 -1275
rect 1367 -1305 1378 -1285
rect 1398 -1305 1416 -1285
rect 1367 -1317 1416 -1305
rect 1466 -1281 1510 -1275
rect 1466 -1301 1481 -1281
rect 1501 -1301 1510 -1281
rect 1466 -1317 1510 -1301
rect 1580 -1281 1624 -1275
rect 1580 -1301 1589 -1281
rect 1609 -1301 1624 -1281
rect 1580 -1317 1624 -1301
rect 1674 -1285 1723 -1275
rect 1674 -1305 1692 -1285
rect 1712 -1305 1723 -1285
rect 1674 -1317 1723 -1305
rect 252 -1511 301 -1501
rect 252 -1531 263 -1511
rect 283 -1531 301 -1511
rect 252 -1543 301 -1531
rect 351 -1507 395 -1501
rect 351 -1527 366 -1507
rect 386 -1527 395 -1507
rect 351 -1543 395 -1527
rect 470 -1511 519 -1501
rect 470 -1531 481 -1511
rect 501 -1531 519 -1511
rect 470 -1543 519 -1531
rect 569 -1507 613 -1501
rect 569 -1527 584 -1507
rect 604 -1527 613 -1507
rect 569 -1543 613 -1527
rect 683 -1507 727 -1501
rect 683 -1527 692 -1507
rect 712 -1527 727 -1507
rect 683 -1543 727 -1527
rect 777 -1511 826 -1501
rect 777 -1531 795 -1511
rect 815 -1531 826 -1511
rect 777 -1543 826 -1531
rect 1050 -1695 1099 -1685
rect 1050 -1715 1061 -1695
rect 1081 -1715 1099 -1695
rect 1050 -1727 1099 -1715
rect 1149 -1691 1193 -1685
rect 1149 -1711 1164 -1691
rect 1184 -1711 1193 -1691
rect 1149 -1727 1193 -1711
rect 1268 -1695 1317 -1685
rect 1268 -1715 1279 -1695
rect 1299 -1715 1317 -1695
rect 1268 -1727 1317 -1715
rect 1367 -1691 1411 -1685
rect 1367 -1711 1382 -1691
rect 1402 -1711 1411 -1691
rect 1367 -1727 1411 -1711
rect 1481 -1691 1525 -1685
rect 1481 -1711 1490 -1691
rect 1510 -1711 1525 -1691
rect 1481 -1727 1525 -1711
rect 1575 -1695 1624 -1685
rect 1575 -1715 1593 -1695
rect 1613 -1715 1624 -1695
rect 1575 -1727 1624 -1715
rect 253 -1923 302 -1913
rect 253 -1943 264 -1923
rect 284 -1943 302 -1923
rect 253 -1955 302 -1943
rect 352 -1919 396 -1913
rect 352 -1939 367 -1919
rect 387 -1939 396 -1919
rect 352 -1955 396 -1939
rect 471 -1923 520 -1913
rect 471 -1943 482 -1923
rect 502 -1943 520 -1923
rect 471 -1955 520 -1943
rect 570 -1919 614 -1913
rect 570 -1939 585 -1919
rect 605 -1939 614 -1919
rect 570 -1955 614 -1939
rect 684 -1919 728 -1913
rect 684 -1939 693 -1919
rect 713 -1939 728 -1919
rect 684 -1955 728 -1939
rect 778 -1923 827 -1913
rect 778 -1943 796 -1923
rect 816 -1943 827 -1923
rect 778 -1955 827 -1943
<< pdiff >>
rect 311 1692 355 1730
rect 311 1672 323 1692
rect 343 1672 355 1692
rect 311 1630 355 1672
rect 405 1692 447 1730
rect 405 1672 419 1692
rect 439 1672 447 1692
rect 405 1630 447 1672
rect 529 1692 573 1730
rect 529 1672 541 1692
rect 561 1672 573 1692
rect 529 1630 573 1672
rect 623 1692 665 1730
rect 623 1672 637 1692
rect 657 1672 665 1692
rect 623 1630 665 1672
rect 739 1692 781 1730
rect 739 1672 747 1692
rect 767 1672 781 1692
rect 739 1630 781 1672
rect 831 1699 876 1730
rect 831 1692 875 1699
rect 831 1672 843 1692
rect 863 1672 875 1692
rect 831 1630 875 1672
rect 1109 1508 1153 1546
rect 1109 1488 1121 1508
rect 1141 1488 1153 1508
rect 1109 1446 1153 1488
rect 1203 1508 1245 1546
rect 1203 1488 1217 1508
rect 1237 1488 1245 1508
rect 1203 1446 1245 1488
rect 1327 1508 1371 1546
rect 1327 1488 1339 1508
rect 1359 1488 1371 1508
rect 1327 1446 1371 1488
rect 1421 1508 1463 1546
rect 1421 1488 1435 1508
rect 1455 1488 1463 1508
rect 1421 1446 1463 1488
rect 1537 1508 1579 1546
rect 1537 1488 1545 1508
rect 1565 1488 1579 1508
rect 1537 1446 1579 1488
rect 1629 1515 1674 1546
rect 1629 1508 1673 1515
rect 1629 1488 1641 1508
rect 1661 1488 1673 1508
rect 1629 1446 1673 1488
rect 312 1280 356 1318
rect 312 1260 324 1280
rect 344 1260 356 1280
rect 312 1218 356 1260
rect 406 1280 448 1318
rect 406 1260 420 1280
rect 440 1260 448 1280
rect 406 1218 448 1260
rect 530 1280 574 1318
rect 530 1260 542 1280
rect 562 1260 574 1280
rect 530 1218 574 1260
rect 624 1280 666 1318
rect 624 1260 638 1280
rect 658 1260 666 1280
rect 624 1218 666 1260
rect 740 1280 782 1318
rect 740 1260 748 1280
rect 768 1260 782 1280
rect 740 1218 782 1260
rect 832 1287 877 1318
rect 832 1280 876 1287
rect 832 1260 844 1280
rect 864 1260 876 1280
rect 832 1218 876 1260
rect 1191 900 1235 938
rect 1191 880 1203 900
rect 1223 880 1235 900
rect 1191 838 1235 880
rect 1285 900 1327 938
rect 1285 880 1299 900
rect 1319 880 1327 900
rect 1285 838 1327 880
rect 1409 900 1453 938
rect 1409 880 1421 900
rect 1441 880 1453 900
rect 1409 838 1453 880
rect 1503 900 1545 938
rect 1503 880 1517 900
rect 1537 880 1545 900
rect 1503 838 1545 880
rect 1619 900 1661 938
rect 1619 880 1627 900
rect 1647 880 1661 900
rect 1619 838 1661 880
rect 1711 907 1756 938
rect 1711 900 1755 907
rect 1711 880 1723 900
rect 1743 880 1755 900
rect 1711 838 1755 880
rect 294 674 338 712
rect 294 654 306 674
rect 326 654 338 674
rect 294 612 338 654
rect 388 674 430 712
rect 388 654 402 674
rect 422 654 430 674
rect 388 612 430 654
rect 512 674 556 712
rect 512 654 524 674
rect 544 654 556 674
rect 512 612 556 654
rect 606 674 648 712
rect 606 654 620 674
rect 640 654 648 674
rect 606 612 648 654
rect 722 674 764 712
rect 722 654 730 674
rect 750 654 764 674
rect 722 612 764 654
rect 814 681 859 712
rect 814 674 858 681
rect 814 654 826 674
rect 846 654 858 674
rect 814 612 858 654
rect 1092 490 1136 528
rect 1092 470 1104 490
rect 1124 470 1136 490
rect 1092 428 1136 470
rect 1186 490 1228 528
rect 1186 470 1200 490
rect 1220 470 1228 490
rect 1186 428 1228 470
rect 1310 490 1354 528
rect 1310 470 1322 490
rect 1342 470 1354 490
rect 1310 428 1354 470
rect 1404 490 1446 528
rect 1404 470 1418 490
rect 1438 470 1446 490
rect 1404 428 1446 470
rect 1520 490 1562 528
rect 1520 470 1528 490
rect 1548 470 1562 490
rect 1520 428 1562 470
rect 1612 497 1657 528
rect 1612 490 1656 497
rect 1612 470 1624 490
rect 1644 470 1656 490
rect 1612 428 1656 470
rect 295 262 339 300
rect 295 242 307 262
rect 327 242 339 262
rect 295 200 339 242
rect 389 262 431 300
rect 389 242 403 262
rect 423 242 431 262
rect 389 200 431 242
rect 513 262 557 300
rect 513 242 525 262
rect 545 242 557 262
rect 513 200 557 242
rect 607 262 649 300
rect 607 242 621 262
rect 641 242 649 262
rect 607 200 649 242
rect 723 262 765 300
rect 723 242 731 262
rect 751 242 765 262
rect 723 200 765 242
rect 815 269 860 300
rect 815 262 859 269
rect 815 242 827 262
rect 847 242 859 262
rect 815 200 859 242
rect 1237 -120 1281 -82
rect 1237 -140 1249 -120
rect 1269 -140 1281 -120
rect 1237 -182 1281 -140
rect 1331 -120 1373 -82
rect 1331 -140 1345 -120
rect 1365 -140 1373 -120
rect 1331 -182 1373 -140
rect 1455 -120 1499 -82
rect 1455 -140 1467 -120
rect 1487 -140 1499 -120
rect 1455 -182 1499 -140
rect 1549 -120 1591 -82
rect 1549 -140 1563 -120
rect 1583 -140 1591 -120
rect 1549 -182 1591 -140
rect 1665 -120 1707 -82
rect 1665 -140 1673 -120
rect 1693 -140 1707 -120
rect 1665 -182 1707 -140
rect 1757 -113 1802 -82
rect 1757 -120 1801 -113
rect 1757 -140 1769 -120
rect 1789 -140 1801 -120
rect 1757 -182 1801 -140
rect 274 -344 318 -306
rect 274 -364 286 -344
rect 306 -364 318 -344
rect 274 -406 318 -364
rect 368 -344 410 -306
rect 368 -364 382 -344
rect 402 -364 410 -344
rect 368 -406 410 -364
rect 492 -344 536 -306
rect 492 -364 504 -344
rect 524 -364 536 -344
rect 492 -406 536 -364
rect 586 -344 628 -306
rect 586 -364 600 -344
rect 620 -364 628 -344
rect 586 -406 628 -364
rect 702 -344 744 -306
rect 702 -364 710 -344
rect 730 -364 744 -344
rect 702 -406 744 -364
rect 794 -337 839 -306
rect 794 -344 838 -337
rect 794 -364 806 -344
rect 826 -364 838 -344
rect 794 -406 838 -364
rect 1072 -528 1116 -490
rect 1072 -548 1084 -528
rect 1104 -548 1116 -528
rect 1072 -590 1116 -548
rect 1166 -528 1208 -490
rect 1166 -548 1180 -528
rect 1200 -548 1208 -528
rect 1166 -590 1208 -548
rect 1290 -528 1334 -490
rect 1290 -548 1302 -528
rect 1322 -548 1334 -528
rect 1290 -590 1334 -548
rect 1384 -528 1426 -490
rect 1384 -548 1398 -528
rect 1418 -548 1426 -528
rect 1384 -590 1426 -548
rect 1500 -528 1542 -490
rect 1500 -548 1508 -528
rect 1528 -548 1542 -528
rect 1500 -590 1542 -548
rect 1592 -521 1637 -490
rect 1592 -528 1636 -521
rect 1592 -548 1604 -528
rect 1624 -548 1636 -528
rect 1592 -590 1636 -548
rect 275 -756 319 -718
rect 275 -776 287 -756
rect 307 -776 319 -756
rect 275 -818 319 -776
rect 369 -756 411 -718
rect 369 -776 383 -756
rect 403 -776 411 -756
rect 369 -818 411 -776
rect 493 -756 537 -718
rect 493 -776 505 -756
rect 525 -776 537 -756
rect 493 -818 537 -776
rect 587 -756 629 -718
rect 587 -776 601 -756
rect 621 -776 629 -756
rect 587 -818 629 -776
rect 703 -756 745 -718
rect 703 -776 711 -756
rect 731 -776 745 -756
rect 703 -818 745 -776
rect 795 -749 840 -718
rect 795 -756 839 -749
rect 795 -776 807 -756
rect 827 -776 839 -756
rect 795 -818 839 -776
rect 1154 -1136 1198 -1098
rect 1154 -1156 1166 -1136
rect 1186 -1156 1198 -1136
rect 1154 -1198 1198 -1156
rect 1248 -1136 1290 -1098
rect 1248 -1156 1262 -1136
rect 1282 -1156 1290 -1136
rect 1248 -1198 1290 -1156
rect 1372 -1136 1416 -1098
rect 1372 -1156 1384 -1136
rect 1404 -1156 1416 -1136
rect 1372 -1198 1416 -1156
rect 1466 -1136 1508 -1098
rect 1466 -1156 1480 -1136
rect 1500 -1156 1508 -1136
rect 1466 -1198 1508 -1156
rect 1582 -1136 1624 -1098
rect 1582 -1156 1590 -1136
rect 1610 -1156 1624 -1136
rect 1582 -1198 1624 -1156
rect 1674 -1129 1719 -1098
rect 1674 -1136 1718 -1129
rect 1674 -1156 1686 -1136
rect 1706 -1156 1718 -1136
rect 1674 -1198 1718 -1156
rect 257 -1362 301 -1324
rect 257 -1382 269 -1362
rect 289 -1382 301 -1362
rect 257 -1424 301 -1382
rect 351 -1362 393 -1324
rect 351 -1382 365 -1362
rect 385 -1382 393 -1362
rect 351 -1424 393 -1382
rect 475 -1362 519 -1324
rect 475 -1382 487 -1362
rect 507 -1382 519 -1362
rect 475 -1424 519 -1382
rect 569 -1362 611 -1324
rect 569 -1382 583 -1362
rect 603 -1382 611 -1362
rect 569 -1424 611 -1382
rect 685 -1362 727 -1324
rect 685 -1382 693 -1362
rect 713 -1382 727 -1362
rect 685 -1424 727 -1382
rect 777 -1355 822 -1324
rect 777 -1362 821 -1355
rect 777 -1382 789 -1362
rect 809 -1382 821 -1362
rect 777 -1424 821 -1382
rect 1055 -1546 1099 -1508
rect 1055 -1566 1067 -1546
rect 1087 -1566 1099 -1546
rect 1055 -1608 1099 -1566
rect 1149 -1546 1191 -1508
rect 1149 -1566 1163 -1546
rect 1183 -1566 1191 -1546
rect 1149 -1608 1191 -1566
rect 1273 -1546 1317 -1508
rect 1273 -1566 1285 -1546
rect 1305 -1566 1317 -1546
rect 1273 -1608 1317 -1566
rect 1367 -1546 1409 -1508
rect 1367 -1566 1381 -1546
rect 1401 -1566 1409 -1546
rect 1367 -1608 1409 -1566
rect 1483 -1546 1525 -1508
rect 1483 -1566 1491 -1546
rect 1511 -1566 1525 -1546
rect 1483 -1608 1525 -1566
rect 1575 -1539 1620 -1508
rect 1575 -1546 1619 -1539
rect 1575 -1566 1587 -1546
rect 1607 -1566 1619 -1546
rect 1575 -1608 1619 -1566
rect 258 -1774 302 -1736
rect 258 -1794 270 -1774
rect 290 -1794 302 -1774
rect 258 -1836 302 -1794
rect 352 -1774 394 -1736
rect 352 -1794 366 -1774
rect 386 -1794 394 -1774
rect 352 -1836 394 -1794
rect 476 -1774 520 -1736
rect 476 -1794 488 -1774
rect 508 -1794 520 -1774
rect 476 -1836 520 -1794
rect 570 -1774 612 -1736
rect 570 -1794 584 -1774
rect 604 -1794 612 -1774
rect 570 -1836 612 -1794
rect 686 -1774 728 -1736
rect 686 -1794 694 -1774
rect 714 -1794 728 -1774
rect 686 -1836 728 -1794
rect 778 -1767 823 -1736
rect 778 -1774 822 -1767
rect 778 -1794 790 -1774
rect 810 -1794 822 -1774
rect 778 -1836 822 -1794
<< ndiffc >>
rect 153 1930 171 1948
rect 151 1831 169 1849
rect 148 1606 166 1624
rect 146 1507 164 1525
rect 317 1523 337 1543
rect 420 1527 440 1547
rect 535 1523 555 1543
rect 638 1527 658 1547
rect 746 1527 766 1547
rect 849 1523 869 1543
rect 142 1423 160 1441
rect 140 1324 158 1342
rect 1115 1339 1135 1359
rect 1218 1343 1238 1363
rect 1333 1339 1353 1359
rect 1436 1343 1456 1363
rect 1544 1343 1564 1363
rect 1647 1339 1667 1359
rect 135 1205 153 1223
rect 133 1106 151 1124
rect 318 1111 338 1131
rect 421 1115 441 1135
rect 536 1111 556 1131
rect 639 1115 659 1135
rect 747 1115 767 1135
rect 850 1111 870 1131
rect 136 912 154 930
rect 134 813 152 831
rect 1197 731 1217 751
rect 1300 735 1320 755
rect 1415 731 1435 751
rect 1518 735 1538 755
rect 1626 735 1646 755
rect 1729 731 1749 751
rect 131 588 149 606
rect 129 489 147 507
rect 300 505 320 525
rect 403 509 423 529
rect 518 505 538 525
rect 621 509 641 529
rect 729 509 749 529
rect 832 505 852 525
rect 125 405 143 423
rect 123 306 141 324
rect 1098 321 1118 341
rect 1201 325 1221 345
rect 1316 321 1336 341
rect 1419 325 1439 345
rect 1527 325 1547 345
rect 1630 321 1650 341
rect 118 187 136 205
rect 116 88 134 106
rect 301 93 321 113
rect 404 97 424 117
rect 519 93 539 113
rect 622 97 642 117
rect 730 97 750 117
rect 833 93 853 113
rect 116 -106 134 -88
rect 114 -205 132 -187
rect 1243 -289 1263 -269
rect 1346 -285 1366 -265
rect 1461 -289 1481 -269
rect 1564 -285 1584 -265
rect 1672 -285 1692 -265
rect 1775 -289 1795 -269
rect 111 -430 129 -412
rect 109 -529 127 -511
rect 280 -513 300 -493
rect 383 -509 403 -489
rect 498 -513 518 -493
rect 601 -509 621 -489
rect 709 -509 729 -489
rect 812 -513 832 -493
rect 105 -613 123 -595
rect 103 -712 121 -694
rect 1078 -697 1098 -677
rect 1181 -693 1201 -673
rect 1296 -697 1316 -677
rect 1399 -693 1419 -673
rect 1507 -693 1527 -673
rect 1610 -697 1630 -677
rect 98 -831 116 -813
rect 96 -930 114 -912
rect 281 -925 301 -905
rect 384 -921 404 -901
rect 499 -925 519 -905
rect 602 -921 622 -901
rect 710 -921 730 -901
rect 813 -925 833 -905
rect 99 -1124 117 -1106
rect 97 -1223 115 -1205
rect 1160 -1305 1180 -1285
rect 1263 -1301 1283 -1281
rect 1378 -1305 1398 -1285
rect 1481 -1301 1501 -1281
rect 1589 -1301 1609 -1281
rect 1692 -1305 1712 -1285
rect 94 -1448 112 -1430
rect 92 -1547 110 -1529
rect 263 -1531 283 -1511
rect 366 -1527 386 -1507
rect 481 -1531 501 -1511
rect 584 -1527 604 -1507
rect 692 -1527 712 -1507
rect 795 -1531 815 -1511
rect 88 -1631 106 -1613
rect 86 -1730 104 -1712
rect 1061 -1715 1081 -1695
rect 1164 -1711 1184 -1691
rect 1279 -1715 1299 -1695
rect 1382 -1711 1402 -1691
rect 1490 -1711 1510 -1691
rect 1593 -1715 1613 -1695
rect 81 -1849 99 -1831
rect 79 -1948 97 -1930
rect 264 -1943 284 -1923
rect 367 -1939 387 -1919
rect 482 -1943 502 -1923
rect 585 -1939 605 -1919
rect 693 -1939 713 -1919
rect 796 -1943 816 -1923
<< pdiffc >>
rect 323 1672 343 1692
rect 419 1672 439 1692
rect 541 1672 561 1692
rect 637 1672 657 1692
rect 747 1672 767 1692
rect 843 1672 863 1692
rect 1121 1488 1141 1508
rect 1217 1488 1237 1508
rect 1339 1488 1359 1508
rect 1435 1488 1455 1508
rect 1545 1488 1565 1508
rect 1641 1488 1661 1508
rect 324 1260 344 1280
rect 420 1260 440 1280
rect 542 1260 562 1280
rect 638 1260 658 1280
rect 748 1260 768 1280
rect 844 1260 864 1280
rect 1203 880 1223 900
rect 1299 880 1319 900
rect 1421 880 1441 900
rect 1517 880 1537 900
rect 1627 880 1647 900
rect 1723 880 1743 900
rect 306 654 326 674
rect 402 654 422 674
rect 524 654 544 674
rect 620 654 640 674
rect 730 654 750 674
rect 826 654 846 674
rect 1104 470 1124 490
rect 1200 470 1220 490
rect 1322 470 1342 490
rect 1418 470 1438 490
rect 1528 470 1548 490
rect 1624 470 1644 490
rect 307 242 327 262
rect 403 242 423 262
rect 525 242 545 262
rect 621 242 641 262
rect 731 242 751 262
rect 827 242 847 262
rect 1249 -140 1269 -120
rect 1345 -140 1365 -120
rect 1467 -140 1487 -120
rect 1563 -140 1583 -120
rect 1673 -140 1693 -120
rect 1769 -140 1789 -120
rect 286 -364 306 -344
rect 382 -364 402 -344
rect 504 -364 524 -344
rect 600 -364 620 -344
rect 710 -364 730 -344
rect 806 -364 826 -344
rect 1084 -548 1104 -528
rect 1180 -548 1200 -528
rect 1302 -548 1322 -528
rect 1398 -548 1418 -528
rect 1508 -548 1528 -528
rect 1604 -548 1624 -528
rect 287 -776 307 -756
rect 383 -776 403 -756
rect 505 -776 525 -756
rect 601 -776 621 -756
rect 711 -776 731 -756
rect 807 -776 827 -756
rect 1166 -1156 1186 -1136
rect 1262 -1156 1282 -1136
rect 1384 -1156 1404 -1136
rect 1480 -1156 1500 -1136
rect 1590 -1156 1610 -1136
rect 1686 -1156 1706 -1136
rect 269 -1382 289 -1362
rect 365 -1382 385 -1362
rect 487 -1382 507 -1362
rect 583 -1382 603 -1362
rect 693 -1382 713 -1362
rect 789 -1382 809 -1362
rect 1067 -1566 1087 -1546
rect 1163 -1566 1183 -1546
rect 1285 -1566 1305 -1546
rect 1381 -1566 1401 -1546
rect 1491 -1566 1511 -1546
rect 1587 -1566 1607 -1546
rect 270 -1794 290 -1774
rect 366 -1794 386 -1774
rect 488 -1794 508 -1774
rect 584 -1794 604 -1774
rect 694 -1794 714 -1774
rect 790 -1794 810 -1774
<< poly >>
rect 355 1730 405 1743
rect 573 1730 623 1743
rect 781 1730 831 1743
rect 355 1602 405 1630
rect 355 1582 368 1602
rect 388 1582 405 1602
rect 355 1553 405 1582
rect 573 1605 623 1630
rect 573 1585 586 1605
rect 606 1585 623 1605
rect 573 1553 623 1585
rect 781 1603 831 1630
rect 781 1583 804 1603
rect 824 1583 831 1603
rect 781 1553 831 1583
rect 1153 1546 1203 1559
rect 1371 1546 1421 1559
rect 1579 1546 1629 1559
rect 355 1495 405 1511
rect 573 1495 623 1511
rect 781 1495 831 1511
rect 1153 1418 1203 1446
rect 1153 1398 1166 1418
rect 1186 1398 1203 1418
rect 1153 1369 1203 1398
rect 1371 1421 1421 1446
rect 1371 1401 1384 1421
rect 1404 1401 1421 1421
rect 1371 1369 1421 1401
rect 1579 1419 1629 1446
rect 1579 1399 1602 1419
rect 1622 1399 1629 1419
rect 1579 1369 1629 1399
rect 356 1318 406 1331
rect 574 1318 624 1331
rect 782 1318 832 1331
rect 1153 1311 1203 1327
rect 1371 1311 1421 1327
rect 1579 1311 1629 1327
rect 356 1190 406 1218
rect 356 1170 369 1190
rect 389 1170 406 1190
rect 356 1141 406 1170
rect 574 1193 624 1218
rect 574 1173 587 1193
rect 607 1173 624 1193
rect 574 1141 624 1173
rect 782 1191 832 1218
rect 782 1171 805 1191
rect 825 1171 832 1191
rect 782 1141 832 1171
rect 356 1083 406 1099
rect 574 1083 624 1099
rect 782 1083 832 1099
rect 1235 938 1285 951
rect 1453 938 1503 951
rect 1661 938 1711 951
rect 1235 810 1285 838
rect 1235 790 1248 810
rect 1268 790 1285 810
rect 1235 761 1285 790
rect 1453 813 1503 838
rect 1453 793 1466 813
rect 1486 793 1503 813
rect 1453 761 1503 793
rect 1661 811 1711 838
rect 1661 791 1684 811
rect 1704 791 1711 811
rect 1661 761 1711 791
rect 338 712 388 725
rect 556 712 606 725
rect 764 712 814 725
rect 1235 703 1285 719
rect 1453 703 1503 719
rect 1661 703 1711 719
rect 338 584 388 612
rect 338 564 351 584
rect 371 564 388 584
rect 338 535 388 564
rect 556 587 606 612
rect 556 567 569 587
rect 589 567 606 587
rect 556 535 606 567
rect 764 585 814 612
rect 764 565 787 585
rect 807 565 814 585
rect 764 535 814 565
rect 1136 528 1186 541
rect 1354 528 1404 541
rect 1562 528 1612 541
rect 338 477 388 493
rect 556 477 606 493
rect 764 477 814 493
rect 1136 400 1186 428
rect 1136 380 1149 400
rect 1169 380 1186 400
rect 1136 351 1186 380
rect 1354 403 1404 428
rect 1354 383 1367 403
rect 1387 383 1404 403
rect 1354 351 1404 383
rect 1562 401 1612 428
rect 1562 381 1585 401
rect 1605 381 1612 401
rect 1562 351 1612 381
rect 339 300 389 313
rect 557 300 607 313
rect 765 300 815 313
rect 1136 293 1186 309
rect 1354 293 1404 309
rect 1562 293 1612 309
rect 339 172 389 200
rect 339 152 352 172
rect 372 152 389 172
rect 339 123 389 152
rect 557 175 607 200
rect 557 155 570 175
rect 590 155 607 175
rect 557 123 607 155
rect 765 173 815 200
rect 765 153 788 173
rect 808 153 815 173
rect 765 123 815 153
rect 339 65 389 81
rect 557 65 607 81
rect 765 65 815 81
rect 1281 -82 1331 -69
rect 1499 -82 1549 -69
rect 1707 -82 1757 -69
rect 1281 -210 1331 -182
rect 1281 -230 1294 -210
rect 1314 -230 1331 -210
rect 1281 -259 1331 -230
rect 1499 -207 1549 -182
rect 1499 -227 1512 -207
rect 1532 -227 1549 -207
rect 1499 -259 1549 -227
rect 1707 -209 1757 -182
rect 1707 -229 1730 -209
rect 1750 -229 1757 -209
rect 1707 -259 1757 -229
rect 318 -306 368 -293
rect 536 -306 586 -293
rect 744 -306 794 -293
rect 1281 -317 1331 -301
rect 1499 -317 1549 -301
rect 1707 -317 1757 -301
rect 318 -434 368 -406
rect 318 -454 331 -434
rect 351 -454 368 -434
rect 318 -483 368 -454
rect 536 -431 586 -406
rect 536 -451 549 -431
rect 569 -451 586 -431
rect 536 -483 586 -451
rect 744 -433 794 -406
rect 744 -453 767 -433
rect 787 -453 794 -433
rect 744 -483 794 -453
rect 1116 -490 1166 -477
rect 1334 -490 1384 -477
rect 1542 -490 1592 -477
rect 318 -541 368 -525
rect 536 -541 586 -525
rect 744 -541 794 -525
rect 1116 -618 1166 -590
rect 1116 -638 1129 -618
rect 1149 -638 1166 -618
rect 1116 -667 1166 -638
rect 1334 -615 1384 -590
rect 1334 -635 1347 -615
rect 1367 -635 1384 -615
rect 1334 -667 1384 -635
rect 1542 -617 1592 -590
rect 1542 -637 1565 -617
rect 1585 -637 1592 -617
rect 1542 -667 1592 -637
rect 319 -718 369 -705
rect 537 -718 587 -705
rect 745 -718 795 -705
rect 1116 -725 1166 -709
rect 1334 -725 1384 -709
rect 1542 -725 1592 -709
rect 319 -846 369 -818
rect 319 -866 332 -846
rect 352 -866 369 -846
rect 319 -895 369 -866
rect 537 -843 587 -818
rect 537 -863 550 -843
rect 570 -863 587 -843
rect 537 -895 587 -863
rect 745 -845 795 -818
rect 745 -865 768 -845
rect 788 -865 795 -845
rect 745 -895 795 -865
rect 319 -953 369 -937
rect 537 -953 587 -937
rect 745 -953 795 -937
rect 1198 -1098 1248 -1085
rect 1416 -1098 1466 -1085
rect 1624 -1098 1674 -1085
rect 1198 -1226 1248 -1198
rect 1198 -1246 1211 -1226
rect 1231 -1246 1248 -1226
rect 1198 -1275 1248 -1246
rect 1416 -1223 1466 -1198
rect 1416 -1243 1429 -1223
rect 1449 -1243 1466 -1223
rect 1416 -1275 1466 -1243
rect 1624 -1225 1674 -1198
rect 1624 -1245 1647 -1225
rect 1667 -1245 1674 -1225
rect 1624 -1275 1674 -1245
rect 301 -1324 351 -1311
rect 519 -1324 569 -1311
rect 727 -1324 777 -1311
rect 1198 -1333 1248 -1317
rect 1416 -1333 1466 -1317
rect 1624 -1333 1674 -1317
rect 301 -1452 351 -1424
rect 301 -1472 314 -1452
rect 334 -1472 351 -1452
rect 301 -1501 351 -1472
rect 519 -1449 569 -1424
rect 519 -1469 532 -1449
rect 552 -1469 569 -1449
rect 519 -1501 569 -1469
rect 727 -1451 777 -1424
rect 727 -1471 750 -1451
rect 770 -1471 777 -1451
rect 727 -1501 777 -1471
rect 1099 -1508 1149 -1495
rect 1317 -1508 1367 -1495
rect 1525 -1508 1575 -1495
rect 301 -1559 351 -1543
rect 519 -1559 569 -1543
rect 727 -1559 777 -1543
rect 1099 -1636 1149 -1608
rect 1099 -1656 1112 -1636
rect 1132 -1656 1149 -1636
rect 1099 -1685 1149 -1656
rect 1317 -1633 1367 -1608
rect 1317 -1653 1330 -1633
rect 1350 -1653 1367 -1633
rect 1317 -1685 1367 -1653
rect 1525 -1635 1575 -1608
rect 1525 -1655 1548 -1635
rect 1568 -1655 1575 -1635
rect 1525 -1685 1575 -1655
rect 302 -1736 352 -1723
rect 520 -1736 570 -1723
rect 728 -1736 778 -1723
rect 1099 -1743 1149 -1727
rect 1317 -1743 1367 -1727
rect 1525 -1743 1575 -1727
rect 302 -1864 352 -1836
rect 302 -1884 315 -1864
rect 335 -1884 352 -1864
rect 302 -1913 352 -1884
rect 520 -1861 570 -1836
rect 520 -1881 533 -1861
rect 553 -1881 570 -1861
rect 520 -1913 570 -1881
rect 728 -1863 778 -1836
rect 728 -1883 751 -1863
rect 771 -1883 778 -1863
rect 728 -1913 778 -1883
rect 302 -1971 352 -1955
rect 520 -1971 570 -1955
rect 728 -1971 778 -1955
<< polycont >>
rect 368 1582 388 1602
rect 586 1585 606 1605
rect 804 1583 824 1603
rect 1166 1398 1186 1418
rect 1384 1401 1404 1421
rect 1602 1399 1622 1419
rect 369 1170 389 1190
rect 587 1173 607 1193
rect 805 1171 825 1191
rect 1248 790 1268 810
rect 1466 793 1486 813
rect 1684 791 1704 811
rect 351 564 371 584
rect 569 567 589 587
rect 787 565 807 585
rect 1149 380 1169 400
rect 1367 383 1387 403
rect 1585 381 1605 401
rect 352 152 372 172
rect 570 155 590 175
rect 788 153 808 173
rect 1294 -230 1314 -210
rect 1512 -227 1532 -207
rect 1730 -229 1750 -209
rect 331 -454 351 -434
rect 549 -451 569 -431
rect 767 -453 787 -433
rect 1129 -638 1149 -618
rect 1347 -635 1367 -615
rect 1565 -637 1585 -617
rect 332 -866 352 -846
rect 550 -863 570 -843
rect 768 -865 788 -845
rect 1211 -1246 1231 -1226
rect 1429 -1243 1449 -1223
rect 1647 -1245 1667 -1225
rect 314 -1472 334 -1452
rect 532 -1469 552 -1449
rect 750 -1471 770 -1451
rect 1112 -1656 1132 -1636
rect 1330 -1653 1350 -1633
rect 1548 -1655 1568 -1635
rect 315 -1884 335 -1864
rect 533 -1881 553 -1861
rect 751 -1883 771 -1863
<< ndiffres >>
rect 130 1952 191 1968
rect 35 1948 191 1952
rect 35 1930 153 1948
rect 171 1930 191 1948
rect 35 1909 191 1930
rect 35 1908 135 1909
rect 36 1872 78 1908
rect 36 1849 187 1872
rect 36 1834 151 1849
rect 130 1831 151 1834
rect 169 1831 187 1849
rect 130 1812 187 1831
rect 125 1628 186 1644
rect 30 1624 186 1628
rect 30 1606 148 1624
rect 166 1606 186 1624
rect 30 1585 186 1606
rect 30 1584 130 1585
rect 31 1548 73 1584
rect 31 1525 182 1548
rect 31 1510 146 1525
rect 125 1507 146 1510
rect 164 1507 182 1525
rect 125 1488 182 1507
rect 119 1445 180 1461
rect 24 1441 180 1445
rect 24 1423 142 1441
rect 160 1423 180 1441
rect 24 1402 180 1423
rect 24 1401 124 1402
rect 25 1365 67 1401
rect 25 1342 176 1365
rect 25 1327 140 1342
rect 119 1324 140 1327
rect 158 1324 176 1342
rect 119 1305 176 1324
rect 112 1227 173 1243
rect 17 1223 173 1227
rect 17 1205 135 1223
rect 153 1205 173 1223
rect 17 1184 173 1205
rect 17 1183 117 1184
rect 18 1147 60 1183
rect 18 1124 169 1147
rect 18 1109 133 1124
rect 112 1106 133 1109
rect 151 1106 169 1124
rect 112 1087 169 1106
rect 113 934 174 950
rect 18 930 174 934
rect 18 912 136 930
rect 154 912 174 930
rect 18 891 174 912
rect 18 890 118 891
rect 19 854 61 890
rect 19 831 170 854
rect 19 816 134 831
rect 113 813 134 816
rect 152 813 170 831
rect 113 794 170 813
rect 108 610 169 626
rect 13 606 169 610
rect 13 588 131 606
rect 149 588 169 606
rect 13 567 169 588
rect 13 566 113 567
rect 14 530 56 566
rect 14 507 165 530
rect 14 492 129 507
rect 108 489 129 492
rect 147 489 165 507
rect 108 470 165 489
rect 102 427 163 443
rect 7 423 163 427
rect 7 405 125 423
rect 143 405 163 423
rect 7 384 163 405
rect 7 383 107 384
rect 8 347 50 383
rect 8 324 159 347
rect 8 309 123 324
rect 102 306 123 309
rect 141 306 159 324
rect 102 287 159 306
rect 95 209 156 225
rect 0 205 156 209
rect 0 187 118 205
rect 136 187 156 205
rect 0 166 156 187
rect 0 165 100 166
rect 1 129 43 165
rect 1 106 152 129
rect 1 91 116 106
rect 95 88 116 91
rect 134 88 152 106
rect 95 69 152 88
rect 93 -84 154 -68
rect -2 -88 154 -84
rect -2 -106 116 -88
rect 134 -106 154 -88
rect -2 -127 154 -106
rect -2 -128 98 -127
rect -1 -164 41 -128
rect -1 -187 150 -164
rect -1 -202 114 -187
rect 93 -205 114 -202
rect 132 -205 150 -187
rect 93 -224 150 -205
rect 88 -408 149 -392
rect -7 -412 149 -408
rect -7 -430 111 -412
rect 129 -430 149 -412
rect -7 -451 149 -430
rect -7 -452 93 -451
rect -6 -488 36 -452
rect -6 -511 145 -488
rect -6 -526 109 -511
rect 88 -529 109 -526
rect 127 -529 145 -511
rect 88 -548 145 -529
rect 82 -591 143 -575
rect -13 -595 143 -591
rect -13 -613 105 -595
rect 123 -613 143 -595
rect -13 -634 143 -613
rect -13 -635 87 -634
rect -12 -671 30 -635
rect -12 -694 139 -671
rect -12 -709 103 -694
rect 82 -712 103 -709
rect 121 -712 139 -694
rect 82 -731 139 -712
rect 75 -809 136 -793
rect -20 -813 136 -809
rect -20 -831 98 -813
rect 116 -831 136 -813
rect -20 -852 136 -831
rect -20 -853 80 -852
rect -19 -889 23 -853
rect -19 -912 132 -889
rect -19 -927 96 -912
rect 75 -930 96 -927
rect 114 -930 132 -912
rect 75 -949 132 -930
rect 76 -1102 137 -1086
rect -19 -1106 137 -1102
rect -19 -1124 99 -1106
rect 117 -1124 137 -1106
rect -19 -1145 137 -1124
rect -19 -1146 81 -1145
rect -18 -1182 24 -1146
rect -18 -1205 133 -1182
rect -18 -1220 97 -1205
rect 76 -1223 97 -1220
rect 115 -1223 133 -1205
rect 76 -1242 133 -1223
rect 71 -1426 132 -1410
rect -24 -1430 132 -1426
rect -24 -1448 94 -1430
rect 112 -1448 132 -1430
rect -24 -1469 132 -1448
rect -24 -1470 76 -1469
rect -23 -1506 19 -1470
rect -23 -1529 128 -1506
rect -23 -1544 92 -1529
rect 71 -1547 92 -1544
rect 110 -1547 128 -1529
rect 71 -1566 128 -1547
rect 65 -1609 126 -1593
rect -30 -1613 126 -1609
rect -30 -1631 88 -1613
rect 106 -1631 126 -1613
rect -30 -1652 126 -1631
rect -30 -1653 70 -1652
rect -29 -1689 13 -1653
rect -29 -1712 122 -1689
rect -29 -1727 86 -1712
rect 65 -1730 86 -1727
rect 104 -1730 122 -1712
rect 65 -1749 122 -1730
rect 58 -1827 119 -1811
rect -37 -1831 119 -1827
rect -37 -1849 81 -1831
rect 99 -1849 119 -1831
rect -37 -1870 119 -1849
rect -37 -1871 63 -1870
rect -36 -1907 6 -1871
rect -36 -1930 115 -1907
rect -36 -1945 79 -1930
rect 58 -1948 79 -1945
rect 97 -1948 115 -1930
rect 58 -1967 115 -1948
<< locali >>
rect 143 1948 190 2064
rect 143 1930 153 1948
rect 171 1930 190 1948
rect 143 1926 190 1930
rect 144 1921 181 1926
rect 132 1859 184 1861
rect 130 1855 563 1859
rect 130 1849 569 1855
rect 130 1831 151 1849
rect 169 1831 569 1849
rect 130 1813 569 1831
rect 132 1624 184 1813
rect 530 1788 569 1813
rect 314 1763 501 1787
rect 530 1768 925 1788
rect 945 1768 948 1788
rect 530 1763 948 1768
rect 314 1692 351 1763
rect 530 1762 873 1763
rect 530 1759 569 1762
rect 835 1761 872 1762
rect 466 1702 497 1703
rect 314 1672 323 1692
rect 343 1672 351 1692
rect 314 1662 351 1672
rect 410 1692 497 1702
rect 410 1672 419 1692
rect 439 1672 497 1692
rect 410 1663 497 1672
rect 410 1662 447 1663
rect 132 1606 148 1624
rect 166 1606 184 1624
rect 466 1612 497 1663
rect 532 1692 569 1759
rect 684 1702 720 1703
rect 532 1672 541 1692
rect 561 1672 569 1692
rect 532 1662 569 1672
rect 628 1692 776 1702
rect 876 1699 972 1701
rect 628 1672 637 1692
rect 657 1672 747 1692
rect 767 1672 776 1692
rect 628 1663 776 1672
rect 834 1692 972 1699
rect 834 1672 843 1692
rect 863 1672 972 1692
rect 834 1663 972 1672
rect 628 1662 665 1663
rect 358 1609 399 1610
rect 132 1588 184 1606
rect 250 1602 399 1609
rect 250 1582 309 1602
rect 329 1582 368 1602
rect 388 1582 399 1602
rect 250 1574 399 1582
rect 466 1605 623 1612
rect 466 1585 586 1605
rect 606 1585 623 1605
rect 466 1575 623 1585
rect 466 1574 501 1575
rect 466 1553 497 1574
rect 684 1553 720 1663
rect 739 1662 776 1663
rect 835 1662 872 1663
rect 795 1603 885 1609
rect 795 1583 804 1603
rect 824 1601 885 1603
rect 824 1583 849 1601
rect 795 1581 849 1583
rect 869 1581 885 1601
rect 795 1575 885 1581
rect 309 1552 346 1553
rect 308 1543 346 1552
rect 136 1525 176 1535
rect 136 1507 146 1525
rect 164 1507 176 1525
rect 308 1523 317 1543
rect 337 1523 346 1543
rect 308 1515 346 1523
rect 412 1547 497 1553
rect 527 1552 564 1553
rect 412 1527 420 1547
rect 440 1527 497 1547
rect 412 1519 497 1527
rect 526 1543 564 1552
rect 526 1523 535 1543
rect 555 1523 564 1543
rect 412 1518 448 1519
rect 526 1515 564 1523
rect 630 1547 774 1553
rect 630 1527 638 1547
rect 658 1527 691 1547
rect 711 1527 746 1547
rect 766 1527 774 1547
rect 630 1519 774 1527
rect 630 1518 666 1519
rect 738 1518 774 1519
rect 840 1552 877 1553
rect 840 1551 878 1552
rect 840 1543 904 1551
rect 840 1523 849 1543
rect 869 1529 904 1543
rect 924 1529 927 1549
rect 869 1524 927 1529
rect 869 1523 904 1524
rect 136 1451 176 1507
rect 309 1486 346 1515
rect 310 1484 346 1486
rect 310 1462 501 1484
rect 527 1483 564 1515
rect 840 1511 904 1523
rect 944 1485 971 1663
rect 803 1483 971 1485
rect 527 1473 971 1483
rect 1112 1579 1299 1603
rect 1330 1584 1723 1604
rect 1743 1584 1746 1604
rect 1330 1579 1746 1584
rect 1112 1508 1149 1579
rect 1330 1578 1671 1579
rect 1264 1518 1295 1519
rect 1112 1488 1121 1508
rect 1141 1488 1149 1508
rect 1112 1478 1149 1488
rect 1208 1508 1295 1518
rect 1208 1488 1217 1508
rect 1237 1488 1295 1508
rect 1208 1479 1295 1488
rect 1208 1478 1245 1479
rect 133 1446 176 1451
rect 524 1457 971 1473
rect 524 1451 552 1457
rect 803 1456 971 1457
rect 133 1443 283 1446
rect 524 1443 551 1451
rect 133 1441 551 1443
rect 133 1423 142 1441
rect 160 1423 551 1441
rect 1264 1428 1295 1479
rect 1330 1508 1367 1578
rect 1633 1577 1670 1578
rect 1482 1518 1518 1519
rect 1330 1488 1339 1508
rect 1359 1488 1367 1508
rect 1330 1478 1367 1488
rect 1426 1508 1574 1518
rect 1674 1515 1770 1517
rect 1426 1488 1435 1508
rect 1455 1488 1545 1508
rect 1565 1488 1574 1508
rect 1426 1479 1574 1488
rect 1632 1508 1770 1515
rect 1632 1488 1641 1508
rect 1661 1488 1770 1508
rect 1632 1479 1770 1488
rect 1426 1478 1463 1479
rect 1156 1425 1197 1426
rect 133 1420 551 1423
rect 133 1414 176 1420
rect 136 1411 176 1414
rect 1048 1418 1197 1425
rect 533 1402 573 1403
rect 244 1385 573 1402
rect 1048 1398 1107 1418
rect 1127 1398 1166 1418
rect 1186 1398 1197 1418
rect 1048 1390 1197 1398
rect 1264 1421 1421 1428
rect 1264 1401 1384 1421
rect 1404 1401 1421 1421
rect 1264 1391 1421 1401
rect 1264 1390 1299 1391
rect 128 1342 171 1353
rect 128 1324 140 1342
rect 158 1324 171 1342
rect 128 1298 171 1324
rect 244 1298 271 1385
rect 533 1376 573 1385
rect 128 1277 271 1298
rect 315 1350 349 1366
rect 533 1356 926 1376
rect 946 1356 949 1376
rect 1264 1369 1295 1390
rect 1482 1369 1518 1479
rect 1537 1478 1574 1479
rect 1633 1478 1670 1479
rect 1593 1419 1683 1425
rect 1593 1399 1602 1419
rect 1622 1417 1683 1419
rect 1622 1399 1647 1417
rect 1593 1397 1647 1399
rect 1667 1397 1683 1417
rect 1593 1391 1683 1397
rect 1107 1368 1144 1369
rect 533 1351 949 1356
rect 1106 1359 1144 1368
rect 533 1350 874 1351
rect 315 1280 352 1350
rect 467 1290 498 1291
rect 128 1275 265 1277
rect 128 1233 171 1275
rect 315 1260 324 1280
rect 344 1260 352 1280
rect 315 1250 352 1260
rect 411 1280 498 1290
rect 411 1260 420 1280
rect 440 1260 498 1280
rect 411 1251 498 1260
rect 411 1250 448 1251
rect 126 1223 171 1233
rect 126 1205 135 1223
rect 153 1205 171 1223
rect 126 1199 171 1205
rect 467 1200 498 1251
rect 533 1280 570 1350
rect 836 1349 873 1350
rect 1106 1339 1115 1359
rect 1135 1339 1144 1359
rect 1106 1331 1144 1339
rect 1210 1363 1295 1369
rect 1325 1368 1362 1369
rect 1210 1343 1218 1363
rect 1238 1343 1295 1363
rect 1210 1335 1295 1343
rect 1324 1359 1362 1368
rect 1324 1339 1333 1359
rect 1353 1339 1362 1359
rect 1210 1334 1246 1335
rect 1324 1331 1362 1339
rect 1428 1363 1572 1369
rect 1428 1343 1436 1363
rect 1456 1344 1488 1363
rect 1509 1344 1544 1363
rect 1456 1343 1544 1344
rect 1564 1343 1572 1363
rect 1428 1335 1572 1343
rect 1428 1334 1464 1335
rect 1536 1334 1572 1335
rect 1638 1368 1675 1369
rect 1638 1367 1676 1368
rect 1638 1359 1702 1367
rect 1638 1339 1647 1359
rect 1667 1345 1702 1359
rect 1722 1345 1725 1365
rect 1667 1340 1725 1345
rect 1667 1339 1702 1340
rect 1107 1302 1144 1331
rect 1108 1300 1144 1302
rect 685 1290 721 1291
rect 533 1260 542 1280
rect 562 1260 570 1280
rect 533 1250 570 1260
rect 629 1280 777 1290
rect 877 1287 973 1289
rect 629 1260 638 1280
rect 658 1260 748 1280
rect 768 1260 777 1280
rect 629 1251 777 1260
rect 835 1280 973 1287
rect 835 1260 844 1280
rect 864 1260 973 1280
rect 1108 1278 1299 1300
rect 1325 1299 1362 1331
rect 1638 1327 1702 1339
rect 1742 1301 1769 1479
rect 1601 1299 1769 1301
rect 1325 1273 1769 1299
rect 835 1251 973 1260
rect 629 1250 666 1251
rect 126 1196 163 1199
rect 359 1197 400 1198
rect 251 1190 400 1197
rect 251 1170 310 1190
rect 330 1170 369 1190
rect 389 1170 400 1190
rect 251 1162 400 1170
rect 467 1193 624 1200
rect 467 1173 587 1193
rect 607 1173 624 1193
rect 467 1163 624 1173
rect 467 1162 502 1163
rect 467 1141 498 1162
rect 685 1141 721 1251
rect 740 1250 777 1251
rect 836 1250 873 1251
rect 796 1191 886 1197
rect 796 1171 805 1191
rect 825 1189 886 1191
rect 825 1171 850 1189
rect 796 1169 850 1171
rect 870 1169 886 1189
rect 796 1163 886 1169
rect 310 1140 347 1141
rect 123 1132 160 1134
rect 123 1124 165 1132
rect 123 1106 133 1124
rect 151 1106 165 1124
rect 123 1097 165 1106
rect 309 1131 347 1140
rect 309 1111 318 1131
rect 338 1111 347 1131
rect 309 1103 347 1111
rect 413 1135 498 1141
rect 528 1140 565 1141
rect 413 1115 421 1135
rect 441 1115 498 1135
rect 413 1107 498 1115
rect 527 1131 565 1140
rect 527 1111 536 1131
rect 556 1111 565 1131
rect 413 1106 449 1107
rect 527 1103 565 1111
rect 631 1139 775 1141
rect 631 1135 683 1139
rect 631 1115 639 1135
rect 659 1119 683 1135
rect 703 1135 775 1139
rect 703 1119 747 1135
rect 659 1115 747 1119
rect 767 1115 775 1135
rect 631 1107 775 1115
rect 631 1106 667 1107
rect 739 1106 775 1107
rect 841 1140 878 1141
rect 841 1139 879 1140
rect 841 1131 905 1139
rect 841 1111 850 1131
rect 870 1117 905 1131
rect 925 1117 928 1137
rect 870 1112 928 1117
rect 870 1111 905 1112
rect 124 1072 165 1097
rect 310 1072 347 1103
rect 528 1072 565 1103
rect 841 1099 905 1111
rect 945 1073 972 1251
rect 124 1045 173 1072
rect 309 1046 358 1072
rect 527 1071 608 1072
rect 804 1071 972 1073
rect 527 1046 972 1071
rect 528 1045 972 1046
rect 126 1012 173 1045
rect 529 1012 569 1045
rect 804 1044 972 1045
rect 1435 1049 1475 1273
rect 1601 1272 1769 1273
rect 1435 1027 1443 1049
rect 1467 1027 1475 1049
rect 1435 1019 1475 1027
rect 126 973 569 1012
rect 126 930 173 973
rect 529 968 569 973
rect 1194 971 1381 995
rect 1412 976 1805 996
rect 1825 976 1828 996
rect 1412 971 1828 976
rect 126 912 136 930
rect 154 912 173 930
rect 126 908 173 912
rect 127 903 164 908
rect 1194 900 1231 971
rect 1412 970 1753 971
rect 1346 910 1377 911
rect 1194 880 1203 900
rect 1223 880 1231 900
rect 1194 870 1231 880
rect 1290 900 1377 910
rect 1290 880 1299 900
rect 1319 880 1377 900
rect 1290 871 1377 880
rect 1290 870 1327 871
rect 115 841 167 843
rect 113 837 546 841
rect 113 831 552 837
rect 113 813 134 831
rect 152 813 552 831
rect 1346 820 1377 871
rect 1412 900 1449 970
rect 1715 969 1752 970
rect 1564 910 1600 911
rect 1412 880 1421 900
rect 1441 880 1449 900
rect 1412 870 1449 880
rect 1508 900 1656 910
rect 1756 907 1852 909
rect 1508 880 1517 900
rect 1537 880 1627 900
rect 1647 880 1656 900
rect 1508 871 1656 880
rect 1714 900 1852 907
rect 1714 880 1723 900
rect 1743 880 1852 900
rect 1714 871 1852 880
rect 1508 870 1545 871
rect 1238 817 1279 818
rect 113 795 552 813
rect 115 606 167 795
rect 513 770 552 795
rect 1130 810 1279 817
rect 1130 790 1189 810
rect 1209 790 1248 810
rect 1268 790 1279 810
rect 1130 782 1279 790
rect 1346 813 1503 820
rect 1346 793 1466 813
rect 1486 793 1503 813
rect 1346 783 1503 793
rect 1346 782 1381 783
rect 297 745 484 769
rect 513 750 908 770
rect 928 750 931 770
rect 1346 761 1377 782
rect 1564 761 1600 871
rect 1619 870 1656 871
rect 1715 870 1752 871
rect 1675 811 1765 817
rect 1675 791 1684 811
rect 1704 809 1765 811
rect 1704 791 1729 809
rect 1675 789 1729 791
rect 1749 789 1765 809
rect 1675 783 1765 789
rect 1189 760 1226 761
rect 513 745 931 750
rect 1188 751 1226 760
rect 297 674 334 745
rect 513 744 856 745
rect 513 741 552 744
rect 818 743 855 744
rect 449 684 480 685
rect 297 654 306 674
rect 326 654 334 674
rect 297 644 334 654
rect 393 674 480 684
rect 393 654 402 674
rect 422 654 480 674
rect 393 645 480 654
rect 393 644 430 645
rect 115 588 131 606
rect 149 588 167 606
rect 449 594 480 645
rect 515 674 552 741
rect 1188 731 1197 751
rect 1217 731 1226 751
rect 1188 723 1226 731
rect 1292 755 1377 761
rect 1407 760 1444 761
rect 1292 735 1300 755
rect 1320 735 1377 755
rect 1292 727 1377 735
rect 1406 751 1444 760
rect 1406 731 1415 751
rect 1435 731 1444 751
rect 1292 726 1328 727
rect 1406 723 1444 731
rect 1510 756 1654 761
rect 1510 755 1572 756
rect 1510 735 1518 755
rect 1538 737 1572 755
rect 1593 755 1654 756
rect 1593 737 1626 755
rect 1538 735 1626 737
rect 1646 735 1654 755
rect 1510 727 1654 735
rect 1510 726 1546 727
rect 1618 726 1654 727
rect 1720 760 1757 761
rect 1720 759 1758 760
rect 1720 751 1784 759
rect 1720 731 1729 751
rect 1749 737 1784 751
rect 1804 737 1807 757
rect 1749 732 1807 737
rect 1749 731 1784 732
rect 1189 694 1226 723
rect 1190 692 1226 694
rect 667 684 703 685
rect 515 654 524 674
rect 544 654 552 674
rect 515 644 552 654
rect 611 674 759 684
rect 859 681 955 683
rect 611 654 620 674
rect 640 654 730 674
rect 750 654 759 674
rect 611 645 759 654
rect 817 674 955 681
rect 817 654 826 674
rect 846 654 955 674
rect 1190 670 1381 692
rect 1407 691 1444 723
rect 1720 719 1784 731
rect 1824 693 1851 871
rect 1683 691 1851 693
rect 1407 677 1851 691
rect 1407 665 1854 677
rect 1450 663 1483 665
rect 817 645 955 654
rect 611 644 648 645
rect 341 591 382 592
rect 115 570 167 588
rect 233 584 382 591
rect 233 564 292 584
rect 312 564 351 584
rect 371 564 382 584
rect 233 556 382 564
rect 449 587 606 594
rect 449 567 569 587
rect 589 567 606 587
rect 449 557 606 567
rect 449 556 484 557
rect 449 535 480 556
rect 667 535 703 645
rect 722 644 759 645
rect 818 644 855 645
rect 778 585 868 591
rect 778 565 787 585
rect 807 583 868 585
rect 807 565 832 583
rect 778 563 832 565
rect 852 563 868 583
rect 778 557 868 563
rect 292 534 329 535
rect 291 525 329 534
rect 119 507 159 517
rect 119 489 129 507
rect 147 489 159 507
rect 291 505 300 525
rect 320 505 329 525
rect 291 497 329 505
rect 395 529 480 535
rect 510 534 547 535
rect 395 509 403 529
rect 423 509 480 529
rect 395 501 480 509
rect 509 525 547 534
rect 509 505 518 525
rect 538 505 547 525
rect 395 500 431 501
rect 509 497 547 505
rect 613 529 757 535
rect 613 509 621 529
rect 641 509 674 529
rect 694 509 729 529
rect 749 509 757 529
rect 613 501 757 509
rect 613 500 649 501
rect 721 500 757 501
rect 823 534 860 535
rect 823 533 861 534
rect 823 525 887 533
rect 823 505 832 525
rect 852 511 887 525
rect 907 511 910 531
rect 852 506 910 511
rect 852 505 887 506
rect 119 433 159 489
rect 292 468 329 497
rect 293 466 329 468
rect 293 444 484 466
rect 510 465 547 497
rect 823 493 887 505
rect 927 467 954 645
rect 1812 620 1854 665
rect 786 465 954 467
rect 510 455 954 465
rect 1095 561 1282 585
rect 1313 566 1706 586
rect 1726 566 1729 586
rect 1313 561 1729 566
rect 1095 490 1132 561
rect 1313 560 1654 561
rect 1247 500 1278 501
rect 1095 470 1104 490
rect 1124 470 1132 490
rect 1095 460 1132 470
rect 1191 490 1278 500
rect 1191 470 1200 490
rect 1220 470 1278 490
rect 1191 461 1278 470
rect 1191 460 1228 461
rect 116 428 159 433
rect 507 439 954 455
rect 507 433 535 439
rect 786 438 954 439
rect 116 425 266 428
rect 507 425 534 433
rect 116 423 534 425
rect 116 405 125 423
rect 143 405 534 423
rect 1247 410 1278 461
rect 1313 490 1350 560
rect 1616 559 1653 560
rect 1465 500 1501 501
rect 1313 470 1322 490
rect 1342 470 1350 490
rect 1313 460 1350 470
rect 1409 490 1557 500
rect 1657 497 1753 499
rect 1409 470 1418 490
rect 1438 470 1528 490
rect 1548 470 1557 490
rect 1409 461 1557 470
rect 1615 490 1753 497
rect 1615 470 1624 490
rect 1644 470 1753 490
rect 1615 461 1753 470
rect 1409 460 1446 461
rect 1139 407 1180 408
rect 116 402 534 405
rect 116 396 159 402
rect 119 393 159 396
rect 1034 400 1180 407
rect 516 384 556 385
rect 227 367 556 384
rect 1034 380 1090 400
rect 1110 380 1149 400
rect 1169 380 1180 400
rect 1034 372 1180 380
rect 1247 403 1404 410
rect 1247 383 1367 403
rect 1387 383 1404 403
rect 1247 373 1404 383
rect 1247 372 1282 373
rect 111 324 154 335
rect 111 306 123 324
rect 141 306 154 324
rect 111 280 154 306
rect 227 280 254 367
rect 516 358 556 367
rect 111 259 254 280
rect 298 332 332 348
rect 516 338 909 358
rect 929 338 932 358
rect 1247 351 1278 372
rect 1465 351 1501 461
rect 1520 460 1557 461
rect 1616 460 1653 461
rect 1576 401 1666 407
rect 1576 381 1585 401
rect 1605 399 1666 401
rect 1605 381 1630 399
rect 1576 379 1630 381
rect 1650 379 1666 399
rect 1576 373 1666 379
rect 1090 350 1127 351
rect 516 333 932 338
rect 1089 341 1127 350
rect 516 332 857 333
rect 298 262 335 332
rect 450 272 481 273
rect 111 257 248 259
rect 111 215 154 257
rect 298 242 307 262
rect 327 242 335 262
rect 298 232 335 242
rect 394 262 481 272
rect 394 242 403 262
rect 423 242 481 262
rect 394 233 481 242
rect 394 232 431 233
rect 109 205 154 215
rect 109 187 118 205
rect 136 187 154 205
rect 109 181 154 187
rect 450 182 481 233
rect 516 262 553 332
rect 819 331 856 332
rect 1089 321 1098 341
rect 1118 321 1127 341
rect 1089 313 1127 321
rect 1193 345 1278 351
rect 1308 350 1345 351
rect 1193 325 1201 345
rect 1221 325 1278 345
rect 1193 317 1278 325
rect 1307 341 1345 350
rect 1307 321 1316 341
rect 1336 321 1345 341
rect 1193 316 1229 317
rect 1307 313 1345 321
rect 1411 345 1555 351
rect 1411 325 1419 345
rect 1439 342 1527 345
rect 1439 325 1474 342
rect 1411 324 1474 325
rect 1493 325 1527 342
rect 1547 325 1555 345
rect 1493 324 1555 325
rect 1411 317 1555 324
rect 1411 316 1447 317
rect 1519 316 1555 317
rect 1621 350 1658 351
rect 1621 349 1659 350
rect 1681 349 1708 353
rect 1621 347 1708 349
rect 1621 341 1685 347
rect 1621 321 1630 341
rect 1650 327 1685 341
rect 1705 327 1708 347
rect 1650 322 1708 327
rect 1650 321 1685 322
rect 1090 284 1127 313
rect 1091 282 1127 284
rect 668 272 704 273
rect 516 242 525 262
rect 545 242 553 262
rect 516 232 553 242
rect 612 262 760 272
rect 860 269 956 271
rect 612 242 621 262
rect 641 242 731 262
rect 751 242 760 262
rect 612 233 760 242
rect 818 262 956 269
rect 818 242 827 262
rect 847 242 956 262
rect 1091 260 1282 282
rect 1308 281 1345 313
rect 1621 309 1685 321
rect 1725 283 1752 461
rect 1584 281 1752 283
rect 1308 255 1752 281
rect 818 233 956 242
rect 612 232 649 233
rect 109 178 146 181
rect 342 179 383 180
rect 234 172 383 179
rect 234 152 293 172
rect 313 152 352 172
rect 372 152 383 172
rect 234 144 383 152
rect 450 175 607 182
rect 450 155 570 175
rect 590 155 607 175
rect 450 145 607 155
rect 450 144 485 145
rect 450 123 481 144
rect 668 123 704 233
rect 723 232 760 233
rect 819 232 856 233
rect 779 173 869 179
rect 779 153 788 173
rect 808 171 869 173
rect 808 153 833 171
rect 779 151 833 153
rect 853 151 869 171
rect 779 145 869 151
rect 293 122 330 123
rect 105 114 143 116
rect 105 106 148 114
rect 105 88 116 106
rect 134 88 148 106
rect 105 61 148 88
rect 292 113 330 122
rect 292 93 301 113
rect 321 93 330 113
rect 292 85 330 93
rect 396 117 481 123
rect 511 122 548 123
rect 396 97 404 117
rect 424 97 481 117
rect 396 89 481 97
rect 510 113 548 122
rect 510 93 519 113
rect 539 93 548 113
rect 396 88 432 89
rect 510 85 548 93
rect 614 121 758 123
rect 614 117 666 121
rect 614 97 622 117
rect 642 101 666 117
rect 686 117 758 121
rect 686 101 730 117
rect 642 97 730 101
rect 750 97 758 117
rect 614 89 758 97
rect 614 88 650 89
rect 722 88 758 89
rect 824 122 861 123
rect 824 121 862 122
rect 824 113 888 121
rect 824 93 833 113
rect 853 99 888 113
rect 908 99 911 119
rect 853 94 911 99
rect 853 93 888 94
rect 106 54 148 61
rect 293 54 330 85
rect 511 54 548 85
rect 824 81 888 93
rect 928 55 955 233
rect 106 14 151 54
rect 293 29 438 54
rect 511 53 591 54
rect 787 53 955 55
rect 511 37 955 53
rect 295 28 438 29
rect 510 27 955 37
rect 106 -7 153 14
rect 510 -7 551 27
rect 787 26 955 27
rect 1418 31 1458 255
rect 1584 254 1752 255
rect 1816 287 1849 620
rect 1816 279 1853 287
rect 1816 260 1824 279
rect 1845 260 1853 279
rect 1816 254 1853 260
rect 1418 9 1426 31
rect 1450 9 1458 31
rect 1418 1 1458 9
rect 106 -37 551 -7
rect 1589 -24 1654 -23
rect 106 -40 529 -37
rect 106 -88 153 -40
rect 106 -106 116 -88
rect 134 -106 153 -88
rect 106 -110 153 -106
rect 1240 -49 1427 -25
rect 1458 -44 1851 -24
rect 1871 -44 1874 -24
rect 1458 -49 1874 -44
rect 107 -115 144 -110
rect 1240 -120 1277 -49
rect 1458 -50 1799 -49
rect 1392 -110 1423 -109
rect 1240 -140 1249 -120
rect 1269 -140 1277 -120
rect 1240 -150 1277 -140
rect 1336 -120 1423 -110
rect 1336 -140 1345 -120
rect 1365 -140 1423 -120
rect 1336 -149 1423 -140
rect 1336 -150 1373 -149
rect 95 -177 147 -175
rect 93 -181 526 -177
rect 93 -187 532 -181
rect 93 -205 114 -187
rect 132 -205 532 -187
rect 1392 -200 1423 -149
rect 1458 -120 1495 -50
rect 1761 -51 1798 -50
rect 1610 -110 1646 -109
rect 1458 -140 1467 -120
rect 1487 -140 1495 -120
rect 1458 -150 1495 -140
rect 1554 -120 1702 -110
rect 1802 -113 1898 -111
rect 1554 -140 1563 -120
rect 1583 -140 1673 -120
rect 1693 -140 1702 -120
rect 1554 -149 1702 -140
rect 1760 -120 1898 -113
rect 1760 -140 1769 -120
rect 1789 -140 1898 -120
rect 1760 -149 1898 -140
rect 1554 -150 1591 -149
rect 1284 -203 1325 -202
rect 93 -223 532 -205
rect 95 -412 147 -223
rect 493 -248 532 -223
rect 1176 -210 1325 -203
rect 1176 -230 1235 -210
rect 1255 -230 1294 -210
rect 1314 -230 1325 -210
rect 1176 -238 1325 -230
rect 1392 -207 1549 -200
rect 1392 -227 1512 -207
rect 1532 -227 1549 -207
rect 1392 -237 1549 -227
rect 1392 -238 1427 -237
rect 277 -273 464 -249
rect 493 -268 888 -248
rect 908 -268 911 -248
rect 1392 -259 1423 -238
rect 1610 -259 1646 -149
rect 1665 -150 1702 -149
rect 1761 -150 1798 -149
rect 1721 -209 1811 -203
rect 1721 -229 1730 -209
rect 1750 -211 1811 -209
rect 1750 -229 1775 -211
rect 1721 -231 1775 -229
rect 1795 -231 1811 -211
rect 1721 -237 1811 -231
rect 1235 -260 1272 -259
rect 493 -273 911 -268
rect 1234 -269 1272 -260
rect 277 -344 314 -273
rect 493 -274 836 -273
rect 493 -277 532 -274
rect 798 -275 835 -274
rect 429 -334 460 -333
rect 277 -364 286 -344
rect 306 -364 314 -344
rect 277 -374 314 -364
rect 373 -344 460 -334
rect 373 -364 382 -344
rect 402 -364 460 -344
rect 373 -373 460 -364
rect 373 -374 410 -373
rect 95 -430 111 -412
rect 129 -430 147 -412
rect 429 -424 460 -373
rect 495 -344 532 -277
rect 1234 -289 1243 -269
rect 1263 -289 1272 -269
rect 1234 -297 1272 -289
rect 1338 -265 1423 -259
rect 1453 -260 1490 -259
rect 1338 -285 1346 -265
rect 1366 -285 1423 -265
rect 1338 -293 1423 -285
rect 1452 -269 1490 -260
rect 1452 -289 1461 -269
rect 1481 -289 1490 -269
rect 1338 -294 1374 -293
rect 1452 -297 1490 -289
rect 1556 -265 1700 -259
rect 1556 -285 1564 -265
rect 1584 -285 1672 -265
rect 1692 -285 1700 -265
rect 1556 -293 1700 -285
rect 1556 -294 1592 -293
rect 1664 -294 1700 -293
rect 1766 -260 1803 -259
rect 1766 -261 1804 -260
rect 1766 -269 1830 -261
rect 1766 -289 1775 -269
rect 1795 -283 1830 -269
rect 1850 -283 1853 -263
rect 1795 -288 1853 -283
rect 1795 -289 1830 -288
rect 1235 -326 1272 -297
rect 1236 -328 1272 -326
rect 647 -334 683 -333
rect 495 -364 504 -344
rect 524 -364 532 -344
rect 495 -374 532 -364
rect 591 -344 739 -334
rect 839 -337 935 -335
rect 591 -364 600 -344
rect 620 -364 710 -344
rect 730 -364 739 -344
rect 591 -373 739 -364
rect 797 -344 935 -337
rect 797 -364 806 -344
rect 826 -364 935 -344
rect 1236 -350 1427 -328
rect 1453 -329 1490 -297
rect 1766 -301 1830 -289
rect 1870 -327 1897 -149
rect 1729 -329 1897 -327
rect 1453 -331 1897 -329
rect 1453 -349 1843 -331
rect 1865 -349 1897 -331
rect 1453 -355 1897 -349
rect 1563 -357 1603 -355
rect 1729 -356 1897 -355
rect 797 -373 935 -364
rect 591 -374 628 -373
rect 321 -427 362 -426
rect 95 -448 147 -430
rect 213 -434 362 -427
rect 213 -454 272 -434
rect 292 -454 331 -434
rect 351 -454 362 -434
rect 213 -462 362 -454
rect 429 -431 586 -424
rect 429 -451 549 -431
rect 569 -451 586 -431
rect 429 -461 586 -451
rect 429 -462 464 -461
rect 429 -483 460 -462
rect 647 -483 683 -373
rect 702 -374 739 -373
rect 798 -374 835 -373
rect 758 -433 848 -427
rect 758 -453 767 -433
rect 787 -435 848 -433
rect 787 -453 812 -435
rect 758 -455 812 -453
rect 832 -455 848 -435
rect 758 -461 848 -455
rect 272 -484 309 -483
rect 271 -493 309 -484
rect 99 -511 139 -501
rect 99 -529 109 -511
rect 127 -529 139 -511
rect 271 -513 280 -493
rect 300 -513 309 -493
rect 271 -521 309 -513
rect 375 -489 460 -483
rect 490 -484 527 -483
rect 375 -509 383 -489
rect 403 -509 460 -489
rect 375 -517 460 -509
rect 489 -493 527 -484
rect 489 -513 498 -493
rect 518 -513 527 -493
rect 375 -518 411 -517
rect 489 -521 527 -513
rect 593 -489 737 -483
rect 593 -509 601 -489
rect 621 -509 654 -489
rect 674 -509 709 -489
rect 729 -509 737 -489
rect 593 -517 737 -509
rect 593 -518 629 -517
rect 701 -518 737 -517
rect 803 -484 840 -483
rect 803 -485 841 -484
rect 803 -493 867 -485
rect 803 -513 812 -493
rect 832 -507 867 -493
rect 887 -507 890 -487
rect 832 -512 890 -507
rect 832 -513 867 -512
rect 99 -585 139 -529
rect 272 -550 309 -521
rect 273 -552 309 -550
rect 273 -574 464 -552
rect 490 -553 527 -521
rect 803 -525 867 -513
rect 907 -551 934 -373
rect 766 -553 934 -551
rect 490 -563 934 -553
rect 1075 -457 1262 -433
rect 1293 -452 1686 -432
rect 1706 -452 1709 -432
rect 1293 -457 1709 -452
rect 1075 -528 1112 -457
rect 1293 -458 1634 -457
rect 1227 -518 1258 -517
rect 1075 -548 1084 -528
rect 1104 -548 1112 -528
rect 1075 -558 1112 -548
rect 1171 -528 1258 -518
rect 1171 -548 1180 -528
rect 1200 -548 1258 -528
rect 1171 -557 1258 -548
rect 1171 -558 1208 -557
rect 96 -590 139 -585
rect 487 -579 934 -563
rect 487 -585 515 -579
rect 766 -580 934 -579
rect 96 -593 246 -590
rect 487 -593 514 -585
rect 96 -595 514 -593
rect 96 -613 105 -595
rect 123 -613 514 -595
rect 1227 -608 1258 -557
rect 1293 -528 1330 -458
rect 1596 -459 1633 -458
rect 1445 -518 1481 -517
rect 1293 -548 1302 -528
rect 1322 -548 1330 -528
rect 1293 -558 1330 -548
rect 1389 -528 1537 -518
rect 1637 -521 1733 -519
rect 1389 -548 1398 -528
rect 1418 -548 1508 -528
rect 1528 -548 1537 -528
rect 1389 -557 1537 -548
rect 1595 -528 1733 -521
rect 1595 -548 1604 -528
rect 1624 -548 1733 -528
rect 1595 -557 1733 -548
rect 1389 -558 1426 -557
rect 1119 -611 1160 -610
rect 96 -616 514 -613
rect 96 -622 139 -616
rect 99 -625 139 -622
rect 1011 -618 1160 -611
rect 496 -634 536 -633
rect 207 -651 536 -634
rect 1011 -638 1070 -618
rect 1090 -638 1129 -618
rect 1149 -638 1160 -618
rect 1011 -646 1160 -638
rect 1227 -615 1384 -608
rect 1227 -635 1347 -615
rect 1367 -635 1384 -615
rect 1227 -645 1384 -635
rect 1227 -646 1262 -645
rect 91 -694 134 -683
rect 91 -712 103 -694
rect 121 -712 134 -694
rect 91 -738 134 -712
rect 207 -738 234 -651
rect 496 -660 536 -651
rect 91 -759 234 -738
rect 278 -686 312 -670
rect 496 -680 889 -660
rect 909 -680 912 -660
rect 1227 -667 1258 -646
rect 1445 -667 1481 -557
rect 1500 -558 1537 -557
rect 1596 -558 1633 -557
rect 1556 -617 1646 -611
rect 1556 -637 1565 -617
rect 1585 -619 1646 -617
rect 1585 -637 1610 -619
rect 1556 -639 1610 -637
rect 1630 -639 1646 -619
rect 1556 -645 1646 -639
rect 1070 -668 1107 -667
rect 496 -685 912 -680
rect 1069 -677 1107 -668
rect 496 -686 837 -685
rect 278 -756 315 -686
rect 430 -746 461 -745
rect 91 -761 228 -759
rect 91 -803 134 -761
rect 278 -776 287 -756
rect 307 -776 315 -756
rect 278 -786 315 -776
rect 374 -756 461 -746
rect 374 -776 383 -756
rect 403 -776 461 -756
rect 374 -785 461 -776
rect 374 -786 411 -785
rect 89 -813 134 -803
rect 89 -831 98 -813
rect 116 -831 134 -813
rect 89 -837 134 -831
rect 430 -836 461 -785
rect 496 -756 533 -686
rect 799 -687 836 -686
rect 1069 -697 1078 -677
rect 1098 -697 1107 -677
rect 1069 -705 1107 -697
rect 1173 -673 1258 -667
rect 1288 -668 1325 -667
rect 1173 -693 1181 -673
rect 1201 -693 1258 -673
rect 1173 -701 1258 -693
rect 1287 -677 1325 -668
rect 1287 -697 1296 -677
rect 1316 -697 1325 -677
rect 1173 -702 1209 -701
rect 1287 -705 1325 -697
rect 1391 -673 1535 -667
rect 1391 -693 1399 -673
rect 1419 -692 1451 -673
rect 1472 -692 1507 -673
rect 1419 -693 1507 -692
rect 1527 -693 1535 -673
rect 1391 -701 1535 -693
rect 1391 -702 1427 -701
rect 1499 -702 1535 -701
rect 1601 -668 1638 -667
rect 1601 -669 1639 -668
rect 1601 -677 1665 -669
rect 1601 -697 1610 -677
rect 1630 -691 1665 -677
rect 1685 -691 1688 -671
rect 1630 -696 1688 -691
rect 1630 -697 1665 -696
rect 1070 -734 1107 -705
rect 1071 -736 1107 -734
rect 648 -746 684 -745
rect 496 -776 505 -756
rect 525 -776 533 -756
rect 496 -786 533 -776
rect 592 -756 740 -746
rect 840 -749 936 -747
rect 592 -776 601 -756
rect 621 -776 711 -756
rect 731 -776 740 -756
rect 592 -785 740 -776
rect 798 -756 936 -749
rect 798 -776 807 -756
rect 827 -776 936 -756
rect 1071 -758 1262 -736
rect 1288 -737 1325 -705
rect 1601 -709 1665 -697
rect 1705 -735 1732 -557
rect 1564 -737 1732 -735
rect 1288 -763 1732 -737
rect 798 -785 936 -776
rect 592 -786 629 -785
rect 89 -840 126 -837
rect 322 -839 363 -838
rect 214 -846 363 -839
rect 214 -866 273 -846
rect 293 -866 332 -846
rect 352 -866 363 -846
rect 214 -874 363 -866
rect 430 -843 587 -836
rect 430 -863 550 -843
rect 570 -863 587 -843
rect 430 -873 587 -863
rect 430 -874 465 -873
rect 430 -895 461 -874
rect 648 -895 684 -785
rect 703 -786 740 -785
rect 799 -786 836 -785
rect 759 -845 849 -839
rect 759 -865 768 -845
rect 788 -847 849 -845
rect 788 -865 813 -847
rect 759 -867 813 -865
rect 833 -867 849 -847
rect 759 -873 849 -867
rect 273 -896 310 -895
rect 86 -904 123 -902
rect 86 -912 128 -904
rect 86 -930 96 -912
rect 114 -930 128 -912
rect 86 -939 128 -930
rect 272 -905 310 -896
rect 272 -925 281 -905
rect 301 -925 310 -905
rect 272 -933 310 -925
rect 376 -901 461 -895
rect 491 -896 528 -895
rect 376 -921 384 -901
rect 404 -921 461 -901
rect 376 -929 461 -921
rect 490 -905 528 -896
rect 490 -925 499 -905
rect 519 -925 528 -905
rect 376 -930 412 -929
rect 490 -933 528 -925
rect 594 -897 738 -895
rect 594 -901 646 -897
rect 594 -921 602 -901
rect 622 -917 646 -901
rect 666 -901 738 -897
rect 666 -917 710 -901
rect 622 -921 710 -917
rect 730 -921 738 -901
rect 594 -929 738 -921
rect 594 -930 630 -929
rect 702 -930 738 -929
rect 804 -896 841 -895
rect 804 -897 842 -896
rect 804 -905 868 -897
rect 804 -925 813 -905
rect 833 -919 868 -905
rect 888 -919 891 -899
rect 833 -924 891 -919
rect 833 -925 868 -924
rect 87 -964 128 -939
rect 273 -964 310 -933
rect 491 -964 528 -933
rect 804 -937 868 -925
rect 908 -963 935 -785
rect 87 -991 136 -964
rect 272 -990 321 -964
rect 490 -965 571 -964
rect 767 -965 935 -963
rect 490 -990 935 -965
rect 491 -991 935 -990
rect 89 -1024 136 -991
rect 492 -1024 532 -991
rect 767 -992 935 -991
rect 1398 -987 1438 -763
rect 1564 -764 1732 -763
rect 1398 -1009 1406 -987
rect 1430 -1009 1438 -987
rect 1398 -1017 1438 -1009
rect 89 -1063 532 -1024
rect 89 -1106 136 -1063
rect 492 -1068 532 -1063
rect 1157 -1065 1344 -1041
rect 1375 -1060 1768 -1040
rect 1788 -1060 1791 -1040
rect 1375 -1065 1791 -1060
rect 89 -1124 99 -1106
rect 117 -1124 136 -1106
rect 89 -1128 136 -1124
rect 90 -1133 127 -1128
rect 1157 -1136 1194 -1065
rect 1375 -1066 1716 -1065
rect 1309 -1126 1340 -1125
rect 1157 -1156 1166 -1136
rect 1186 -1156 1194 -1136
rect 1157 -1166 1194 -1156
rect 1253 -1136 1340 -1126
rect 1253 -1156 1262 -1136
rect 1282 -1156 1340 -1136
rect 1253 -1165 1340 -1156
rect 1253 -1166 1290 -1165
rect 78 -1195 130 -1193
rect 76 -1199 509 -1195
rect 76 -1205 515 -1199
rect 76 -1223 97 -1205
rect 115 -1223 515 -1205
rect 1309 -1216 1340 -1165
rect 1375 -1136 1412 -1066
rect 1678 -1067 1715 -1066
rect 1527 -1126 1563 -1125
rect 1375 -1156 1384 -1136
rect 1404 -1156 1412 -1136
rect 1375 -1166 1412 -1156
rect 1471 -1136 1619 -1126
rect 1719 -1129 1815 -1127
rect 1471 -1156 1480 -1136
rect 1500 -1156 1590 -1136
rect 1610 -1156 1619 -1136
rect 1471 -1165 1619 -1156
rect 1677 -1136 1815 -1129
rect 1677 -1156 1686 -1136
rect 1706 -1156 1815 -1136
rect 1677 -1165 1815 -1156
rect 1471 -1166 1508 -1165
rect 1201 -1219 1242 -1218
rect 76 -1241 515 -1223
rect 78 -1430 130 -1241
rect 476 -1266 515 -1241
rect 1093 -1226 1242 -1219
rect 1093 -1246 1152 -1226
rect 1172 -1246 1211 -1226
rect 1231 -1246 1242 -1226
rect 1093 -1254 1242 -1246
rect 1309 -1223 1466 -1216
rect 1309 -1243 1429 -1223
rect 1449 -1243 1466 -1223
rect 1309 -1253 1466 -1243
rect 1309 -1254 1344 -1253
rect 260 -1291 447 -1267
rect 476 -1286 871 -1266
rect 891 -1286 894 -1266
rect 1309 -1275 1340 -1254
rect 1527 -1275 1563 -1165
rect 1582 -1166 1619 -1165
rect 1678 -1166 1715 -1165
rect 1638 -1225 1728 -1219
rect 1638 -1245 1647 -1225
rect 1667 -1227 1728 -1225
rect 1667 -1245 1692 -1227
rect 1638 -1247 1692 -1245
rect 1712 -1247 1728 -1227
rect 1638 -1253 1728 -1247
rect 1152 -1276 1189 -1275
rect 476 -1291 894 -1286
rect 1151 -1285 1189 -1276
rect 260 -1362 297 -1291
rect 476 -1292 819 -1291
rect 476 -1295 515 -1292
rect 781 -1293 818 -1292
rect 412 -1352 443 -1351
rect 260 -1382 269 -1362
rect 289 -1382 297 -1362
rect 260 -1392 297 -1382
rect 356 -1362 443 -1352
rect 356 -1382 365 -1362
rect 385 -1382 443 -1362
rect 356 -1391 443 -1382
rect 356 -1392 393 -1391
rect 78 -1448 94 -1430
rect 112 -1448 130 -1430
rect 412 -1442 443 -1391
rect 478 -1362 515 -1295
rect 1151 -1305 1160 -1285
rect 1180 -1305 1189 -1285
rect 1151 -1313 1189 -1305
rect 1255 -1281 1340 -1275
rect 1370 -1276 1407 -1275
rect 1255 -1301 1263 -1281
rect 1283 -1301 1340 -1281
rect 1255 -1309 1340 -1301
rect 1369 -1285 1407 -1276
rect 1369 -1305 1378 -1285
rect 1398 -1305 1407 -1285
rect 1255 -1310 1291 -1309
rect 1369 -1313 1407 -1305
rect 1473 -1281 1617 -1275
rect 1473 -1301 1481 -1281
rect 1501 -1286 1589 -1281
rect 1501 -1301 1537 -1286
rect 1473 -1303 1537 -1301
rect 1556 -1301 1589 -1286
rect 1609 -1301 1617 -1281
rect 1556 -1303 1617 -1301
rect 1473 -1309 1617 -1303
rect 1473 -1310 1509 -1309
rect 1581 -1310 1617 -1309
rect 1683 -1276 1720 -1275
rect 1683 -1277 1721 -1276
rect 1683 -1285 1747 -1277
rect 1683 -1305 1692 -1285
rect 1712 -1299 1747 -1285
rect 1767 -1299 1770 -1279
rect 1712 -1304 1770 -1299
rect 1712 -1305 1747 -1304
rect 1152 -1342 1189 -1313
rect 1153 -1344 1189 -1342
rect 630 -1352 666 -1351
rect 478 -1382 487 -1362
rect 507 -1382 515 -1362
rect 478 -1392 515 -1382
rect 574 -1362 722 -1352
rect 822 -1355 918 -1353
rect 574 -1382 583 -1362
rect 603 -1382 693 -1362
rect 713 -1382 722 -1362
rect 574 -1391 722 -1382
rect 780 -1362 918 -1355
rect 780 -1382 789 -1362
rect 809 -1382 918 -1362
rect 1153 -1366 1344 -1344
rect 1370 -1345 1407 -1313
rect 1683 -1317 1747 -1305
rect 1787 -1343 1814 -1165
rect 1646 -1345 1814 -1343
rect 1370 -1359 1814 -1345
rect 1370 -1371 1817 -1359
rect 1413 -1373 1446 -1371
rect 780 -1391 918 -1382
rect 574 -1392 611 -1391
rect 304 -1445 345 -1444
rect 78 -1466 130 -1448
rect 196 -1452 345 -1445
rect 196 -1472 255 -1452
rect 275 -1472 314 -1452
rect 334 -1472 345 -1452
rect 196 -1480 345 -1472
rect 412 -1449 569 -1442
rect 412 -1469 532 -1449
rect 552 -1469 569 -1449
rect 412 -1479 569 -1469
rect 412 -1480 447 -1479
rect 412 -1501 443 -1480
rect 630 -1501 666 -1391
rect 685 -1392 722 -1391
rect 781 -1392 818 -1391
rect 741 -1451 831 -1445
rect 741 -1471 750 -1451
rect 770 -1453 831 -1451
rect 770 -1471 795 -1453
rect 741 -1473 795 -1471
rect 815 -1473 831 -1453
rect 741 -1479 831 -1473
rect 255 -1502 292 -1501
rect 254 -1511 292 -1502
rect 82 -1529 122 -1519
rect 82 -1547 92 -1529
rect 110 -1547 122 -1529
rect 254 -1531 263 -1511
rect 283 -1531 292 -1511
rect 254 -1539 292 -1531
rect 358 -1507 443 -1501
rect 473 -1502 510 -1501
rect 358 -1527 366 -1507
rect 386 -1527 443 -1507
rect 358 -1535 443 -1527
rect 472 -1511 510 -1502
rect 472 -1531 481 -1511
rect 501 -1531 510 -1511
rect 358 -1536 394 -1535
rect 472 -1539 510 -1531
rect 576 -1507 720 -1501
rect 576 -1527 584 -1507
rect 604 -1527 637 -1507
rect 657 -1527 692 -1507
rect 712 -1527 720 -1507
rect 576 -1535 720 -1527
rect 576 -1536 612 -1535
rect 684 -1536 720 -1535
rect 786 -1502 823 -1501
rect 786 -1503 824 -1502
rect 786 -1511 850 -1503
rect 786 -1531 795 -1511
rect 815 -1525 850 -1511
rect 870 -1525 873 -1505
rect 815 -1530 873 -1525
rect 815 -1531 850 -1530
rect 82 -1603 122 -1547
rect 255 -1568 292 -1539
rect 256 -1570 292 -1568
rect 256 -1592 447 -1570
rect 473 -1571 510 -1539
rect 786 -1543 850 -1531
rect 890 -1569 917 -1391
rect 1775 -1416 1817 -1371
rect 749 -1571 917 -1569
rect 473 -1581 917 -1571
rect 1058 -1475 1245 -1451
rect 1276 -1470 1669 -1450
rect 1689 -1470 1692 -1450
rect 1276 -1475 1692 -1470
rect 1058 -1546 1095 -1475
rect 1276 -1476 1617 -1475
rect 1210 -1536 1241 -1535
rect 1058 -1566 1067 -1546
rect 1087 -1566 1095 -1546
rect 1058 -1576 1095 -1566
rect 1154 -1546 1241 -1536
rect 1154 -1566 1163 -1546
rect 1183 -1566 1241 -1546
rect 1154 -1575 1241 -1566
rect 1154 -1576 1191 -1575
rect 79 -1608 122 -1603
rect 470 -1597 917 -1581
rect 470 -1603 498 -1597
rect 749 -1598 917 -1597
rect 79 -1611 229 -1608
rect 470 -1611 497 -1603
rect 79 -1613 497 -1611
rect 79 -1631 88 -1613
rect 106 -1631 497 -1613
rect 1210 -1626 1241 -1575
rect 1276 -1546 1313 -1476
rect 1579 -1477 1616 -1476
rect 1428 -1536 1464 -1535
rect 1276 -1566 1285 -1546
rect 1305 -1566 1313 -1546
rect 1276 -1576 1313 -1566
rect 1372 -1546 1520 -1536
rect 1620 -1539 1716 -1537
rect 1372 -1566 1381 -1546
rect 1401 -1566 1491 -1546
rect 1511 -1566 1520 -1546
rect 1372 -1575 1520 -1566
rect 1578 -1546 1716 -1539
rect 1578 -1566 1587 -1546
rect 1607 -1566 1716 -1546
rect 1578 -1575 1716 -1566
rect 1372 -1576 1409 -1575
rect 1102 -1629 1143 -1628
rect 79 -1634 497 -1631
rect 79 -1640 122 -1634
rect 82 -1643 122 -1640
rect 997 -1636 1143 -1629
rect 479 -1652 519 -1651
rect 190 -1669 519 -1652
rect 997 -1656 1053 -1636
rect 1073 -1656 1112 -1636
rect 1132 -1656 1143 -1636
rect 997 -1664 1143 -1656
rect 1210 -1633 1367 -1626
rect 1210 -1653 1330 -1633
rect 1350 -1653 1367 -1633
rect 1210 -1663 1367 -1653
rect 1210 -1664 1245 -1663
rect 74 -1712 117 -1701
rect 74 -1730 86 -1712
rect 104 -1730 117 -1712
rect 74 -1756 117 -1730
rect 190 -1756 217 -1669
rect 479 -1678 519 -1669
rect 74 -1777 217 -1756
rect 261 -1704 295 -1688
rect 479 -1698 872 -1678
rect 892 -1698 895 -1678
rect 1210 -1685 1241 -1664
rect 1428 -1685 1464 -1575
rect 1483 -1576 1520 -1575
rect 1579 -1576 1616 -1575
rect 1539 -1635 1629 -1629
rect 1539 -1655 1548 -1635
rect 1568 -1637 1629 -1635
rect 1568 -1655 1593 -1637
rect 1539 -1657 1593 -1655
rect 1613 -1657 1629 -1637
rect 1539 -1663 1629 -1657
rect 1053 -1686 1090 -1685
rect 479 -1703 895 -1698
rect 1052 -1695 1090 -1686
rect 479 -1704 820 -1703
rect 261 -1774 298 -1704
rect 413 -1764 444 -1763
rect 74 -1779 211 -1777
rect 74 -1821 117 -1779
rect 261 -1794 270 -1774
rect 290 -1794 298 -1774
rect 261 -1804 298 -1794
rect 357 -1774 444 -1764
rect 357 -1794 366 -1774
rect 386 -1794 444 -1774
rect 357 -1803 444 -1794
rect 357 -1804 394 -1803
rect 72 -1831 117 -1821
rect 72 -1849 81 -1831
rect 99 -1849 117 -1831
rect 72 -1855 117 -1849
rect 413 -1854 444 -1803
rect 479 -1774 516 -1704
rect 782 -1705 819 -1704
rect 1052 -1715 1061 -1695
rect 1081 -1715 1090 -1695
rect 1052 -1723 1090 -1715
rect 1156 -1691 1241 -1685
rect 1271 -1686 1308 -1685
rect 1156 -1711 1164 -1691
rect 1184 -1711 1241 -1691
rect 1156 -1719 1241 -1711
rect 1270 -1695 1308 -1686
rect 1270 -1715 1279 -1695
rect 1299 -1715 1308 -1695
rect 1156 -1720 1192 -1719
rect 1270 -1723 1308 -1715
rect 1374 -1691 1518 -1685
rect 1374 -1711 1382 -1691
rect 1402 -1694 1490 -1691
rect 1402 -1711 1437 -1694
rect 1374 -1712 1437 -1711
rect 1456 -1711 1490 -1694
rect 1510 -1711 1518 -1691
rect 1456 -1712 1518 -1711
rect 1374 -1719 1518 -1712
rect 1374 -1720 1410 -1719
rect 1482 -1720 1518 -1719
rect 1584 -1686 1621 -1685
rect 1584 -1687 1622 -1686
rect 1644 -1687 1671 -1683
rect 1584 -1689 1671 -1687
rect 1584 -1695 1648 -1689
rect 1584 -1715 1593 -1695
rect 1613 -1709 1648 -1695
rect 1668 -1709 1671 -1689
rect 1613 -1714 1671 -1709
rect 1613 -1715 1648 -1714
rect 1053 -1752 1090 -1723
rect 1054 -1754 1090 -1752
rect 631 -1764 667 -1763
rect 479 -1794 488 -1774
rect 508 -1794 516 -1774
rect 479 -1804 516 -1794
rect 575 -1774 723 -1764
rect 823 -1767 919 -1765
rect 575 -1794 584 -1774
rect 604 -1794 694 -1774
rect 714 -1794 723 -1774
rect 575 -1803 723 -1794
rect 781 -1774 919 -1767
rect 781 -1794 790 -1774
rect 810 -1794 919 -1774
rect 1054 -1776 1245 -1754
rect 1271 -1755 1308 -1723
rect 1584 -1727 1648 -1715
rect 1688 -1753 1715 -1575
rect 1547 -1755 1715 -1753
rect 1271 -1781 1715 -1755
rect 781 -1803 919 -1794
rect 575 -1804 612 -1803
rect 72 -1858 109 -1855
rect 305 -1857 346 -1856
rect 197 -1864 346 -1857
rect 197 -1884 256 -1864
rect 276 -1884 315 -1864
rect 335 -1884 346 -1864
rect 197 -1892 346 -1884
rect 413 -1861 570 -1854
rect 413 -1881 533 -1861
rect 553 -1881 570 -1861
rect 413 -1891 570 -1881
rect 413 -1892 448 -1891
rect 413 -1913 444 -1892
rect 631 -1913 667 -1803
rect 686 -1804 723 -1803
rect 782 -1804 819 -1803
rect 742 -1863 832 -1857
rect 742 -1883 751 -1863
rect 771 -1865 832 -1863
rect 771 -1883 796 -1865
rect 742 -1885 796 -1883
rect 816 -1885 832 -1865
rect 742 -1891 832 -1885
rect 256 -1914 293 -1913
rect 69 -1922 106 -1920
rect 69 -1930 111 -1922
rect 69 -1948 79 -1930
rect 97 -1948 111 -1930
rect 69 -1957 111 -1948
rect 255 -1923 293 -1914
rect 255 -1943 264 -1923
rect 284 -1943 293 -1923
rect 255 -1951 293 -1943
rect 359 -1919 444 -1913
rect 474 -1914 511 -1913
rect 359 -1939 367 -1919
rect 387 -1939 444 -1919
rect 359 -1947 444 -1939
rect 473 -1923 511 -1914
rect 473 -1943 482 -1923
rect 502 -1943 511 -1923
rect 359 -1948 395 -1947
rect 473 -1951 511 -1943
rect 577 -1915 721 -1913
rect 577 -1919 629 -1915
rect 577 -1939 585 -1919
rect 605 -1935 629 -1919
rect 649 -1919 721 -1915
rect 649 -1935 693 -1919
rect 605 -1939 693 -1935
rect 713 -1939 721 -1919
rect 577 -1947 721 -1939
rect 577 -1948 613 -1947
rect 685 -1948 721 -1947
rect 787 -1914 824 -1913
rect 787 -1915 825 -1914
rect 787 -1923 851 -1915
rect 787 -1943 796 -1923
rect 816 -1937 851 -1923
rect 871 -1937 874 -1917
rect 816 -1942 874 -1937
rect 816 -1943 851 -1942
rect 70 -1982 111 -1957
rect 256 -1982 293 -1951
rect 474 -1982 511 -1951
rect 787 -1955 851 -1943
rect 891 -1981 918 -1803
rect 70 -1983 554 -1982
rect 750 -1983 918 -1981
rect 70 -2008 918 -1983
rect 70 -2009 111 -2008
rect 474 -2009 918 -2008
rect 750 -2010 918 -2009
rect 1381 -2005 1421 -1781
rect 1547 -1782 1715 -1781
rect 1779 -1749 1812 -1416
rect 1779 -1757 1816 -1749
rect 1779 -1776 1787 -1757
rect 1808 -1776 1816 -1757
rect 1779 -1782 1816 -1776
rect 1381 -2027 1389 -2005
rect 1413 -2027 1421 -2005
rect 1381 -2035 1421 -2027
<< viali >>
rect 925 1768 945 1788
rect 309 1582 329 1602
rect 849 1581 869 1601
rect 691 1527 711 1547
rect 904 1529 924 1549
rect 1723 1584 1743 1604
rect 1107 1398 1127 1418
rect 926 1356 946 1376
rect 1647 1397 1667 1417
rect 1488 1344 1509 1363
rect 1702 1345 1722 1365
rect 310 1170 330 1190
rect 850 1169 870 1189
rect 683 1119 703 1139
rect 905 1117 925 1137
rect 1443 1027 1467 1049
rect 1805 976 1825 996
rect 1189 790 1209 810
rect 908 750 928 770
rect 1729 789 1749 809
rect 1572 737 1593 756
rect 1784 737 1804 757
rect 292 564 312 584
rect 832 563 852 583
rect 674 509 694 529
rect 887 511 907 531
rect 1706 566 1726 586
rect 1090 380 1110 400
rect 909 338 929 358
rect 1630 379 1650 399
rect 1474 324 1493 342
rect 1685 327 1705 347
rect 293 152 313 172
rect 833 151 853 171
rect 666 101 686 121
rect 888 99 908 119
rect 1824 260 1845 279
rect 1426 9 1450 31
rect 1851 -44 1871 -24
rect 1235 -230 1255 -210
rect 888 -268 908 -248
rect 1775 -231 1795 -211
rect 1830 -283 1850 -263
rect 1843 -349 1865 -331
rect 272 -454 292 -434
rect 812 -455 832 -435
rect 654 -509 674 -489
rect 867 -507 887 -487
rect 1686 -452 1706 -432
rect 1070 -638 1090 -618
rect 889 -680 909 -660
rect 1610 -639 1630 -619
rect 1451 -692 1472 -673
rect 1665 -691 1685 -671
rect 273 -866 293 -846
rect 813 -867 833 -847
rect 646 -917 666 -897
rect 868 -919 888 -899
rect 1406 -1009 1430 -987
rect 1768 -1060 1788 -1040
rect 1152 -1246 1172 -1226
rect 871 -1286 891 -1266
rect 1692 -1247 1712 -1227
rect 1537 -1303 1556 -1286
rect 1747 -1299 1767 -1279
rect 255 -1472 275 -1452
rect 795 -1473 815 -1453
rect 637 -1527 657 -1507
rect 850 -1525 870 -1505
rect 1669 -1470 1689 -1450
rect 1053 -1656 1073 -1636
rect 872 -1698 892 -1678
rect 1593 -1657 1613 -1637
rect 1437 -1712 1456 -1694
rect 1648 -1709 1668 -1689
rect 256 -1884 276 -1864
rect 796 -1885 816 -1865
rect 629 -1935 649 -1915
rect 851 -1937 871 -1917
rect 1787 -1776 1808 -1757
rect 1389 -2027 1413 -2005
<< metal1 >>
rect 921 1793 953 1794
rect 918 1788 953 1793
rect 918 1768 925 1788
rect 945 1768 953 1788
rect 918 1760 953 1768
rect 300 1602 885 1610
rect 300 1582 309 1602
rect 329 1601 885 1602
rect 329 1582 849 1601
rect 300 1581 849 1582
rect 869 1581 885 1601
rect 300 1575 885 1581
rect 919 1554 953 1760
rect 683 1547 718 1554
rect 683 1527 691 1547
rect 711 1527 718 1547
rect 683 1454 718 1527
rect 897 1549 953 1554
rect 897 1529 904 1549
rect 924 1529 953 1549
rect 897 1522 953 1529
rect 988 1656 1018 1658
rect 1717 1656 1750 1657
rect 988 1630 1751 1656
rect 897 1521 932 1522
rect 988 1455 1018 1630
rect 1717 1609 1751 1630
rect 1716 1604 1751 1609
rect 1716 1584 1723 1604
rect 1743 1584 1751 1604
rect 1716 1576 1751 1584
rect 983 1454 1018 1455
rect 682 1427 1018 1454
rect 988 1426 1018 1427
rect 1098 1418 1683 1426
rect 1098 1398 1107 1418
rect 1127 1417 1683 1418
rect 1127 1398 1647 1417
rect 1098 1397 1647 1398
rect 1667 1397 1683 1417
rect 1098 1391 1683 1397
rect 922 1381 954 1382
rect 919 1376 954 1381
rect 919 1356 926 1376
rect 946 1356 954 1376
rect 1717 1370 1751 1576
rect 919 1348 954 1356
rect 301 1190 886 1198
rect 301 1170 310 1190
rect 330 1189 886 1190
rect 330 1170 850 1189
rect 301 1169 850 1170
rect 870 1169 886 1189
rect 301 1163 886 1169
rect 675 1139 714 1143
rect 920 1142 954 1348
rect 1483 1363 1518 1369
rect 1483 1344 1488 1363
rect 1509 1344 1518 1363
rect 1483 1335 1518 1344
rect 1695 1365 1751 1370
rect 1695 1345 1702 1365
rect 1722 1345 1751 1365
rect 1695 1338 1751 1345
rect 1695 1337 1730 1338
rect 1487 1267 1516 1335
rect 1487 1233 1833 1267
rect 675 1119 683 1139
rect 703 1119 714 1139
rect 675 1044 714 1119
rect 898 1137 954 1142
rect 898 1117 905 1137
rect 925 1117 954 1137
rect 898 1110 954 1117
rect 898 1109 933 1110
rect 1438 1049 1477 1062
rect 1438 1044 1443 1049
rect 675 1027 1443 1044
rect 1467 1044 1477 1049
rect 1467 1027 1478 1044
rect 675 1019 1478 1027
rect 677 1018 963 1019
rect 1794 996 1833 1233
rect 1794 984 1805 996
rect 1798 976 1805 984
rect 1825 976 1833 996
rect 1798 968 1833 976
rect 1180 810 1765 818
rect 1180 790 1189 810
rect 1209 809 1765 810
rect 1209 790 1729 809
rect 1180 789 1729 790
rect 1749 789 1765 809
rect 1180 783 1765 789
rect 904 775 936 776
rect 901 770 936 775
rect 901 750 908 770
rect 928 750 936 770
rect 1799 762 1833 968
rect 901 742 936 750
rect 283 584 868 592
rect 283 564 292 584
rect 312 583 868 584
rect 312 564 832 583
rect 283 563 832 564
rect 852 563 868 583
rect 283 557 868 563
rect 902 536 936 742
rect 1567 756 1598 762
rect 1567 737 1572 756
rect 1593 737 1598 756
rect 1567 695 1598 737
rect 1777 757 1833 762
rect 1777 737 1784 757
rect 1804 737 1833 757
rect 1777 730 1833 737
rect 1777 729 1812 730
rect 1567 667 1906 695
rect 666 529 701 536
rect 666 509 674 529
rect 694 509 701 529
rect 666 436 701 509
rect 880 531 936 536
rect 880 511 887 531
rect 907 511 936 531
rect 880 504 936 511
rect 971 638 1001 640
rect 1700 638 1733 639
rect 971 612 1734 638
rect 880 503 915 504
rect 971 437 1001 612
rect 1700 591 1734 612
rect 1699 586 1734 591
rect 1699 566 1706 586
rect 1726 566 1734 586
rect 1699 558 1734 566
rect 966 436 1001 437
rect 665 409 1001 436
rect 971 408 1001 409
rect 1081 400 1666 408
rect 1081 380 1090 400
rect 1110 399 1666 400
rect 1110 380 1630 399
rect 1081 379 1630 380
rect 1650 379 1666 399
rect 1081 373 1666 379
rect 905 363 937 364
rect 902 358 937 363
rect 902 338 909 358
rect 929 338 937 358
rect 1700 352 1734 558
rect 902 330 937 338
rect 284 172 869 180
rect 284 152 293 172
rect 313 171 869 172
rect 313 152 833 171
rect 284 151 833 152
rect 853 151 869 171
rect 284 145 869 151
rect 658 121 697 125
rect 903 124 937 330
rect 1467 342 1501 350
rect 1467 324 1474 342
rect 1493 324 1501 342
rect 1467 317 1501 324
rect 1678 347 1734 352
rect 1678 327 1685 347
rect 1705 327 1734 347
rect 1678 320 1734 327
rect 1678 319 1713 320
rect 1471 287 1500 317
rect 1471 279 1853 287
rect 1471 260 1824 279
rect 1845 260 1853 279
rect 1471 255 1853 260
rect 658 101 666 121
rect 686 101 697 121
rect 658 26 697 101
rect 881 119 937 124
rect 881 99 888 119
rect 908 99 937 119
rect 881 92 937 99
rect 881 91 916 92
rect 1421 31 1460 44
rect 1421 26 1426 31
rect 658 9 1426 26
rect 1450 26 1460 31
rect 1450 9 1461 26
rect 658 1 1461 9
rect 660 0 946 1
rect 1877 -18 1906 667
rect 1846 -21 1911 -18
rect 1844 -24 1911 -21
rect 1844 -44 1851 -24
rect 1871 -44 1911 -24
rect 1844 -51 1911 -44
rect 1844 -52 1879 -51
rect 1226 -210 1811 -202
rect 1226 -230 1235 -210
rect 1255 -211 1811 -210
rect 1255 -230 1775 -211
rect 1226 -231 1775 -230
rect 1795 -231 1811 -211
rect 1226 -237 1811 -231
rect 884 -243 916 -242
rect 881 -248 916 -243
rect 881 -268 888 -248
rect 908 -268 916 -248
rect 1845 -258 1879 -52
rect 881 -276 916 -268
rect 263 -434 848 -426
rect 263 -454 272 -434
rect 292 -435 848 -434
rect 292 -454 812 -435
rect 263 -455 812 -454
rect 832 -455 848 -435
rect 263 -461 848 -455
rect 882 -482 916 -276
rect 1823 -263 1879 -258
rect 1823 -283 1830 -263
rect 1850 -283 1879 -263
rect 1823 -290 1879 -283
rect 1823 -291 1858 -290
rect 1836 -331 1868 -325
rect 1836 -349 1843 -331
rect 1865 -349 1868 -331
rect 646 -489 681 -482
rect 646 -509 654 -489
rect 674 -509 681 -489
rect 646 -582 681 -509
rect 860 -487 916 -482
rect 860 -507 867 -487
rect 887 -507 916 -487
rect 860 -514 916 -507
rect 951 -380 981 -378
rect 1680 -380 1713 -379
rect 951 -406 1714 -380
rect 860 -515 895 -514
rect 951 -581 981 -406
rect 1680 -427 1714 -406
rect 1679 -432 1714 -427
rect 1679 -452 1686 -432
rect 1706 -452 1714 -432
rect 1679 -460 1714 -452
rect 946 -582 981 -581
rect 645 -609 981 -582
rect 951 -610 981 -609
rect 1061 -618 1646 -610
rect 1061 -638 1070 -618
rect 1090 -619 1646 -618
rect 1090 -638 1610 -619
rect 1061 -639 1610 -638
rect 1630 -639 1646 -619
rect 1061 -645 1646 -639
rect 885 -655 917 -654
rect 882 -660 917 -655
rect 882 -680 889 -660
rect 909 -680 917 -660
rect 1680 -666 1714 -460
rect 882 -688 917 -680
rect 264 -846 849 -838
rect 264 -866 273 -846
rect 293 -847 849 -846
rect 293 -866 813 -847
rect 264 -867 813 -866
rect 833 -867 849 -847
rect 264 -873 849 -867
rect 638 -897 677 -893
rect 883 -894 917 -688
rect 1446 -673 1481 -667
rect 1446 -692 1451 -673
rect 1472 -692 1481 -673
rect 1446 -701 1481 -692
rect 1658 -671 1714 -666
rect 1658 -691 1665 -671
rect 1685 -691 1714 -671
rect 1658 -698 1714 -691
rect 1658 -699 1693 -698
rect 1450 -769 1479 -701
rect 1450 -803 1796 -769
rect 638 -917 646 -897
rect 666 -917 677 -897
rect 638 -992 677 -917
rect 861 -899 917 -894
rect 861 -919 868 -899
rect 888 -919 917 -899
rect 861 -926 917 -919
rect 861 -927 896 -926
rect 1401 -987 1440 -974
rect 1401 -992 1406 -987
rect 638 -1009 1406 -992
rect 1430 -992 1440 -987
rect 1430 -1009 1441 -992
rect 638 -1017 1441 -1009
rect 640 -1018 926 -1017
rect 1757 -1040 1796 -803
rect 1757 -1052 1768 -1040
rect 1761 -1060 1768 -1052
rect 1788 -1060 1796 -1040
rect 1761 -1068 1796 -1060
rect 1143 -1226 1728 -1218
rect 1143 -1246 1152 -1226
rect 1172 -1227 1728 -1226
rect 1172 -1246 1692 -1227
rect 1143 -1247 1692 -1246
rect 1712 -1247 1728 -1227
rect 1143 -1253 1728 -1247
rect 867 -1261 899 -1260
rect 864 -1266 899 -1261
rect 864 -1286 871 -1266
rect 891 -1286 899 -1266
rect 1762 -1274 1796 -1068
rect 864 -1294 899 -1286
rect 246 -1452 831 -1444
rect 246 -1472 255 -1452
rect 275 -1453 831 -1452
rect 275 -1472 795 -1453
rect 246 -1473 795 -1472
rect 815 -1473 831 -1453
rect 246 -1479 831 -1473
rect 865 -1500 899 -1294
rect 1528 -1286 1564 -1277
rect 1528 -1303 1537 -1286
rect 1556 -1303 1564 -1286
rect 1528 -1312 1564 -1303
rect 1740 -1279 1796 -1274
rect 1740 -1299 1747 -1279
rect 1767 -1299 1796 -1279
rect 1740 -1306 1796 -1299
rect 1740 -1307 1775 -1306
rect 1534 -1347 1560 -1312
rect 1836 -1347 1868 -349
rect 1534 -1375 1868 -1347
rect 629 -1507 664 -1500
rect 629 -1527 637 -1507
rect 657 -1527 664 -1507
rect 629 -1600 664 -1527
rect 843 -1505 899 -1500
rect 843 -1525 850 -1505
rect 870 -1525 899 -1505
rect 843 -1532 899 -1525
rect 934 -1398 964 -1396
rect 1663 -1398 1696 -1397
rect 934 -1424 1697 -1398
rect 843 -1533 878 -1532
rect 934 -1599 964 -1424
rect 1663 -1445 1697 -1424
rect 1662 -1450 1697 -1445
rect 1662 -1470 1669 -1450
rect 1689 -1470 1697 -1450
rect 1662 -1478 1697 -1470
rect 929 -1600 964 -1599
rect 628 -1627 964 -1600
rect 934 -1628 964 -1627
rect 1044 -1636 1629 -1628
rect 1044 -1656 1053 -1636
rect 1073 -1637 1629 -1636
rect 1073 -1656 1593 -1637
rect 1044 -1657 1593 -1656
rect 1613 -1657 1629 -1637
rect 1044 -1663 1629 -1657
rect 868 -1673 900 -1672
rect 865 -1678 900 -1673
rect 865 -1698 872 -1678
rect 892 -1698 900 -1678
rect 1663 -1684 1697 -1478
rect 865 -1706 900 -1698
rect 247 -1864 832 -1856
rect 247 -1884 256 -1864
rect 276 -1865 832 -1864
rect 276 -1884 796 -1865
rect 247 -1885 796 -1884
rect 816 -1885 832 -1865
rect 247 -1891 832 -1885
rect 621 -1915 660 -1911
rect 866 -1912 900 -1706
rect 1430 -1694 1464 -1686
rect 1430 -1712 1437 -1694
rect 1456 -1712 1464 -1694
rect 1430 -1719 1464 -1712
rect 1641 -1689 1697 -1684
rect 1641 -1709 1648 -1689
rect 1668 -1709 1697 -1689
rect 1641 -1716 1697 -1709
rect 1641 -1717 1676 -1716
rect 1434 -1749 1463 -1719
rect 1434 -1757 1816 -1749
rect 1434 -1776 1787 -1757
rect 1808 -1776 1816 -1757
rect 1434 -1781 1816 -1776
rect 621 -1935 629 -1915
rect 649 -1935 660 -1915
rect 621 -2010 660 -1935
rect 844 -1917 900 -1912
rect 844 -1937 851 -1917
rect 871 -1937 900 -1917
rect 844 -1944 900 -1937
rect 844 -1945 879 -1944
rect 1384 -2005 1423 -1992
rect 1384 -2010 1389 -2005
rect 621 -2027 1389 -2010
rect 1413 -2010 1423 -2005
rect 1413 -2027 1424 -2010
rect 621 -2035 1424 -2027
rect 623 -2036 909 -2035
<< labels >>
rlabel locali 263 1584 285 1599 1 d0
rlabel locali 317 1772 346 1778 1 vdd
rlabel locali 314 1473 343 1479 1 gnd
rlabel space 420 1491 449 1500 1 gnd
rlabel nwell 452 1749 475 1752 1 vdd
rlabel locali 264 1172 286 1187 1 d0
rlabel locali 318 1360 347 1366 1 vdd
rlabel locali 315 1061 344 1067 1 gnd
rlabel space 421 1079 450 1088 1 gnd
rlabel nwell 453 1337 476 1340 1 vdd
rlabel locali 154 2017 178 2047 1 vref
rlabel locali 246 566 268 581 1 d0
rlabel locali 300 754 329 760 1 vdd
rlabel locali 297 455 326 461 1 gnd
rlabel space 403 473 432 482 1 gnd
rlabel nwell 435 731 458 734 1 vdd
rlabel locali 247 154 269 169 1 d0
rlabel locali 301 342 330 348 1 vdd
rlabel locali 298 43 327 49 1 gnd
rlabel space 404 61 433 70 1 gnd
rlabel nwell 436 319 459 322 1 vdd
rlabel locali 1115 1588 1144 1594 1 vdd
rlabel locali 1112 1289 1141 1295 1 gnd
rlabel space 1218 1307 1247 1316 1 gnd
rlabel nwell 1250 1565 1273 1568 1 vdd
rlabel locali 1055 1396 1077 1413 1 d1
rlabel locali 1098 570 1127 576 1 vdd
rlabel locali 1095 271 1124 277 1 gnd
rlabel space 1201 289 1230 298 1 gnd
rlabel nwell 1233 547 1256 550 1 vdd
rlabel locali 1038 378 1060 395 1 d1
rlabel locali 1197 980 1226 986 1 vdd
rlabel locali 1194 681 1223 687 1 gnd
rlabel space 1300 699 1329 708 1 gnd
rlabel nwell 1332 957 1355 960 1 vdd
rlabel locali 1139 788 1159 812 1 d2
rlabel locali 226 -452 248 -437 1 d0
rlabel locali 280 -264 309 -258 1 vdd
rlabel locali 277 -563 306 -557 1 gnd
rlabel space 383 -545 412 -536 1 gnd
rlabel nwell 415 -287 438 -284 1 vdd
rlabel locali 227 -864 249 -849 1 d0
rlabel locali 281 -676 310 -670 1 vdd
rlabel locali 278 -975 307 -969 1 gnd
rlabel space 384 -957 413 -948 1 gnd
rlabel nwell 416 -699 439 -696 1 vdd
rlabel locali 209 -1470 231 -1455 1 d0
rlabel locali 263 -1282 292 -1276 1 vdd
rlabel locali 260 -1581 289 -1575 1 gnd
rlabel space 366 -1563 395 -1554 1 gnd
rlabel nwell 398 -1305 421 -1302 1 vdd
rlabel locali 210 -1882 232 -1867 1 d0
rlabel locali 264 -1694 293 -1688 1 vdd
rlabel locali 261 -1993 290 -1987 1 gnd
rlabel space 367 -1975 396 -1966 1 gnd
rlabel nwell 399 -1717 422 -1714 1 vdd
rlabel locali 76 -1994 104 -1976 1 gnd
rlabel locali 1078 -448 1107 -442 1 vdd
rlabel locali 1075 -747 1104 -741 1 gnd
rlabel space 1181 -729 1210 -720 1 gnd
rlabel nwell 1213 -471 1236 -468 1 vdd
rlabel locali 1018 -640 1040 -623 1 d1
rlabel locali 1061 -1466 1090 -1460 1 vdd
rlabel locali 1058 -1765 1087 -1759 1 gnd
rlabel space 1164 -1747 1193 -1738 1 gnd
rlabel nwell 1196 -1489 1219 -1486 1 vdd
rlabel locali 1001 -1658 1023 -1641 1 d1
rlabel locali 1160 -1056 1189 -1050 1 vdd
rlabel locali 1157 -1355 1186 -1349 1 gnd
rlabel space 1263 -1337 1292 -1328 1 gnd
rlabel nwell 1295 -1079 1318 -1076 1 vdd
rlabel locali 1102 -1248 1122 -1224 1 d2
rlabel locali 1243 -40 1272 -34 1 vdd
rlabel locali 1240 -339 1269 -333 1 gnd
rlabel space 1346 -321 1375 -312 1 gnd
rlabel nwell 1378 -63 1401 -60 1 vdd
rlabel locali 1616 -193 1638 -178 1 vout
rlabel locali 1187 -226 1207 -213 1 d3
<< end >>

magic
tech sky130A
timestamp 1616084917
<< nwell >>
rect 185 -1 793 149
rect 1047 -185 1655 -35
rect 186 -413 794 -263
<< nmos >>
rect 249 -102 299 -60
rect 467 -102 517 -60
rect 675 -102 725 -60
rect 1111 -286 1161 -244
rect 1329 -286 1379 -244
rect 1537 -286 1587 -244
rect 250 -514 300 -472
rect 468 -514 518 -472
rect 676 -514 726 -472
<< pmos >>
rect 249 17 299 117
rect 467 17 517 117
rect 675 17 725 117
rect 1111 -167 1161 -67
rect 1329 -167 1379 -67
rect 1537 -167 1587 -67
rect 250 -395 300 -295
rect 468 -395 518 -295
rect 676 -395 726 -295
<< ndiff >>
rect 200 -70 249 -60
rect 200 -90 211 -70
rect 231 -90 249 -70
rect 200 -102 249 -90
rect 299 -66 343 -60
rect 299 -86 314 -66
rect 334 -86 343 -66
rect 299 -102 343 -86
rect 418 -70 467 -60
rect 418 -90 429 -70
rect 449 -90 467 -70
rect 418 -102 467 -90
rect 517 -66 561 -60
rect 517 -86 532 -66
rect 552 -86 561 -66
rect 517 -102 561 -86
rect 631 -66 675 -60
rect 631 -86 640 -66
rect 660 -86 675 -66
rect 631 -102 675 -86
rect 725 -70 774 -60
rect 725 -90 743 -70
rect 763 -90 774 -70
rect 725 -102 774 -90
rect 1062 -254 1111 -244
rect 1062 -274 1073 -254
rect 1093 -274 1111 -254
rect 1062 -286 1111 -274
rect 1161 -250 1205 -244
rect 1161 -270 1176 -250
rect 1196 -270 1205 -250
rect 1161 -286 1205 -270
rect 1280 -254 1329 -244
rect 1280 -274 1291 -254
rect 1311 -274 1329 -254
rect 1280 -286 1329 -274
rect 1379 -250 1423 -244
rect 1379 -270 1394 -250
rect 1414 -270 1423 -250
rect 1379 -286 1423 -270
rect 1493 -250 1537 -244
rect 1493 -270 1502 -250
rect 1522 -270 1537 -250
rect 1493 -286 1537 -270
rect 1587 -254 1636 -244
rect 1587 -274 1605 -254
rect 1625 -274 1636 -254
rect 1587 -286 1636 -274
rect 201 -482 250 -472
rect 201 -502 212 -482
rect 232 -502 250 -482
rect 201 -514 250 -502
rect 300 -478 344 -472
rect 300 -498 315 -478
rect 335 -498 344 -478
rect 300 -514 344 -498
rect 419 -482 468 -472
rect 419 -502 430 -482
rect 450 -502 468 -482
rect 419 -514 468 -502
rect 518 -478 562 -472
rect 518 -498 533 -478
rect 553 -498 562 -478
rect 518 -514 562 -498
rect 632 -478 676 -472
rect 632 -498 641 -478
rect 661 -498 676 -478
rect 632 -514 676 -498
rect 726 -482 775 -472
rect 726 -502 744 -482
rect 764 -502 775 -482
rect 726 -514 775 -502
<< pdiff >>
rect 205 79 249 117
rect 205 59 217 79
rect 237 59 249 79
rect 205 17 249 59
rect 299 79 341 117
rect 299 59 313 79
rect 333 59 341 79
rect 299 17 341 59
rect 423 79 467 117
rect 423 59 435 79
rect 455 59 467 79
rect 423 17 467 59
rect 517 79 559 117
rect 517 59 531 79
rect 551 59 559 79
rect 517 17 559 59
rect 633 79 675 117
rect 633 59 641 79
rect 661 59 675 79
rect 633 17 675 59
rect 725 86 770 117
rect 725 79 769 86
rect 725 59 737 79
rect 757 59 769 79
rect 725 17 769 59
rect 1067 -105 1111 -67
rect 1067 -125 1079 -105
rect 1099 -125 1111 -105
rect 1067 -167 1111 -125
rect 1161 -105 1203 -67
rect 1161 -125 1175 -105
rect 1195 -125 1203 -105
rect 1161 -167 1203 -125
rect 1285 -105 1329 -67
rect 1285 -125 1297 -105
rect 1317 -125 1329 -105
rect 1285 -167 1329 -125
rect 1379 -105 1421 -67
rect 1379 -125 1393 -105
rect 1413 -125 1421 -105
rect 1379 -167 1421 -125
rect 1495 -105 1537 -67
rect 1495 -125 1503 -105
rect 1523 -125 1537 -105
rect 1495 -167 1537 -125
rect 1587 -98 1632 -67
rect 1587 -105 1631 -98
rect 1587 -125 1599 -105
rect 1619 -125 1631 -105
rect 1587 -167 1631 -125
rect 206 -333 250 -295
rect 206 -353 218 -333
rect 238 -353 250 -333
rect 206 -395 250 -353
rect 300 -333 342 -295
rect 300 -353 314 -333
rect 334 -353 342 -333
rect 300 -395 342 -353
rect 424 -333 468 -295
rect 424 -353 436 -333
rect 456 -353 468 -333
rect 424 -395 468 -353
rect 518 -333 560 -295
rect 518 -353 532 -333
rect 552 -353 560 -333
rect 518 -395 560 -353
rect 634 -333 676 -295
rect 634 -353 642 -333
rect 662 -353 676 -333
rect 634 -395 676 -353
rect 726 -326 771 -295
rect 726 -333 770 -326
rect 726 -353 738 -333
rect 758 -353 770 -333
rect 726 -395 770 -353
<< ndiffc >>
rect 47 317 65 335
rect 45 218 63 236
rect 42 -7 60 11
rect 40 -106 58 -88
rect 211 -90 231 -70
rect 314 -86 334 -66
rect 429 -90 449 -70
rect 532 -86 552 -66
rect 640 -86 660 -66
rect 743 -90 763 -70
rect 36 -190 54 -172
rect 34 -289 52 -271
rect 1073 -274 1093 -254
rect 1176 -270 1196 -250
rect 1291 -274 1311 -254
rect 1394 -270 1414 -250
rect 1502 -270 1522 -250
rect 1605 -274 1625 -254
rect 29 -408 47 -390
rect 27 -507 45 -489
rect 212 -502 232 -482
rect 315 -498 335 -478
rect 430 -502 450 -482
rect 533 -498 553 -478
rect 641 -498 661 -478
rect 744 -502 764 -482
<< pdiffc >>
rect 217 59 237 79
rect 313 59 333 79
rect 435 59 455 79
rect 531 59 551 79
rect 641 59 661 79
rect 737 59 757 79
rect 1079 -125 1099 -105
rect 1175 -125 1195 -105
rect 1297 -125 1317 -105
rect 1393 -125 1413 -105
rect 1503 -125 1523 -105
rect 1599 -125 1619 -105
rect 218 -353 238 -333
rect 314 -353 334 -333
rect 436 -353 456 -333
rect 532 -353 552 -333
rect 642 -353 662 -333
rect 738 -353 758 -333
<< poly >>
rect 249 117 299 130
rect 467 117 517 130
rect 675 117 725 130
rect 249 -11 299 17
rect 249 -31 262 -11
rect 282 -31 299 -11
rect 249 -60 299 -31
rect 467 -8 517 17
rect 467 -28 480 -8
rect 500 -28 517 -8
rect 467 -60 517 -28
rect 675 -10 725 17
rect 675 -30 698 -10
rect 718 -30 725 -10
rect 675 -60 725 -30
rect 1111 -67 1161 -54
rect 1329 -67 1379 -54
rect 1537 -67 1587 -54
rect 249 -118 299 -102
rect 467 -118 517 -102
rect 675 -118 725 -102
rect 1111 -195 1161 -167
rect 1111 -215 1124 -195
rect 1144 -215 1161 -195
rect 1111 -244 1161 -215
rect 1329 -192 1379 -167
rect 1329 -212 1342 -192
rect 1362 -212 1379 -192
rect 1329 -244 1379 -212
rect 1537 -194 1587 -167
rect 1537 -214 1560 -194
rect 1580 -214 1587 -194
rect 1537 -244 1587 -214
rect 250 -295 300 -282
rect 468 -295 518 -282
rect 676 -295 726 -282
rect 1111 -302 1161 -286
rect 1329 -302 1379 -286
rect 1537 -302 1587 -286
rect 250 -423 300 -395
rect 250 -443 263 -423
rect 283 -443 300 -423
rect 250 -472 300 -443
rect 468 -420 518 -395
rect 468 -440 481 -420
rect 501 -440 518 -420
rect 468 -472 518 -440
rect 676 -422 726 -395
rect 676 -442 699 -422
rect 719 -442 726 -422
rect 676 -472 726 -442
rect 250 -530 300 -514
rect 468 -530 518 -514
rect 676 -530 726 -514
<< polycont >>
rect 262 -31 282 -11
rect 480 -28 500 -8
rect 698 -30 718 -10
rect 1124 -215 1144 -195
rect 1342 -212 1362 -192
rect 1560 -214 1580 -194
rect 263 -443 283 -423
rect 481 -440 501 -420
rect 699 -442 719 -422
<< ndiffres >>
rect 24 339 85 355
rect -71 335 85 339
rect -71 317 47 335
rect 65 317 85 335
rect -71 296 85 317
rect -71 295 29 296
rect -70 259 -28 295
rect -70 236 81 259
rect -70 221 45 236
rect 24 218 45 221
rect 63 218 81 236
rect 24 199 81 218
rect 19 15 80 31
rect -76 11 80 15
rect -76 -7 42 11
rect 60 -7 80 11
rect -76 -28 80 -7
rect -76 -29 24 -28
rect -75 -65 -33 -29
rect -75 -88 76 -65
rect -75 -103 40 -88
rect 19 -106 40 -103
rect 58 -106 76 -88
rect 19 -125 76 -106
rect 13 -168 74 -152
rect -82 -172 74 -168
rect -82 -190 36 -172
rect 54 -190 74 -172
rect -82 -211 74 -190
rect -82 -212 18 -211
rect -81 -248 -39 -212
rect -81 -271 70 -248
rect -81 -286 34 -271
rect 13 -289 34 -286
rect 52 -289 70 -271
rect 13 -308 70 -289
rect 6 -386 67 -370
rect -89 -390 67 -386
rect -89 -408 29 -390
rect 47 -408 67 -390
rect -89 -429 67 -408
rect -89 -430 11 -429
rect -88 -466 -46 -430
rect -88 -489 63 -466
rect -88 -504 27 -489
rect 6 -507 27 -504
rect 45 -507 63 -489
rect 6 -526 63 -507
<< locali >>
rect 37 335 84 451
rect 37 317 47 335
rect 65 317 84 335
rect 37 313 84 317
rect 38 308 75 313
rect 26 246 78 248
rect 24 242 457 246
rect 24 236 463 242
rect 24 218 45 236
rect 63 218 463 236
rect 24 200 463 218
rect 26 11 78 200
rect 424 175 463 200
rect 208 150 395 174
rect 424 155 819 175
rect 839 155 842 175
rect 424 150 842 155
rect 208 79 245 150
rect 424 149 767 150
rect 424 146 463 149
rect 729 148 766 149
rect 360 89 391 90
rect 208 59 217 79
rect 237 59 245 79
rect 208 49 245 59
rect 304 79 391 89
rect 304 59 313 79
rect 333 59 391 79
rect 304 50 391 59
rect 304 49 341 50
rect 26 -7 42 11
rect 60 -7 78 11
rect 360 -1 391 50
rect 426 79 463 146
rect 578 89 614 90
rect 426 59 435 79
rect 455 59 463 79
rect 426 49 463 59
rect 522 79 670 89
rect 770 86 866 88
rect 522 59 531 79
rect 551 59 641 79
rect 661 59 670 79
rect 522 50 670 59
rect 728 79 866 86
rect 728 59 737 79
rect 757 59 866 79
rect 728 50 866 59
rect 522 49 559 50
rect 252 -4 293 -3
rect 26 -25 78 -7
rect 144 -11 293 -4
rect 144 -31 203 -11
rect 223 -31 262 -11
rect 282 -31 293 -11
rect 144 -39 293 -31
rect 360 -8 517 -1
rect 360 -28 480 -8
rect 500 -28 517 -8
rect 360 -38 517 -28
rect 360 -39 395 -38
rect 360 -60 391 -39
rect 578 -60 614 50
rect 633 49 670 50
rect 729 49 766 50
rect 689 -10 779 -4
rect 689 -30 698 -10
rect 718 -12 779 -10
rect 718 -30 743 -12
rect 689 -32 743 -30
rect 763 -32 779 -12
rect 689 -38 779 -32
rect 203 -61 240 -60
rect 202 -70 240 -61
rect 30 -88 70 -78
rect 30 -106 40 -88
rect 58 -106 70 -88
rect 202 -90 211 -70
rect 231 -90 240 -70
rect 202 -98 240 -90
rect 306 -66 391 -60
rect 421 -61 458 -60
rect 306 -86 314 -66
rect 334 -86 391 -66
rect 306 -94 391 -86
rect 420 -70 458 -61
rect 420 -90 429 -70
rect 449 -90 458 -70
rect 306 -95 342 -94
rect 420 -98 458 -90
rect 524 -66 668 -60
rect 524 -86 532 -66
rect 552 -86 585 -66
rect 605 -86 640 -66
rect 660 -86 668 -66
rect 524 -94 668 -86
rect 524 -95 560 -94
rect 632 -95 668 -94
rect 734 -61 771 -60
rect 734 -62 772 -61
rect 734 -70 798 -62
rect 734 -90 743 -70
rect 763 -84 798 -70
rect 818 -84 821 -64
rect 763 -89 821 -84
rect 763 -90 798 -89
rect 30 -162 70 -106
rect 203 -127 240 -98
rect 204 -129 240 -127
rect 204 -151 395 -129
rect 421 -130 458 -98
rect 734 -102 798 -90
rect 838 -128 865 50
rect 697 -130 865 -128
rect 421 -140 865 -130
rect 1070 -34 1257 -10
rect 1288 -29 1681 -9
rect 1701 -29 1704 -9
rect 1288 -34 1704 -29
rect 1070 -105 1107 -34
rect 1288 -35 1629 -34
rect 1222 -95 1253 -94
rect 1070 -125 1079 -105
rect 1099 -125 1107 -105
rect 1070 -135 1107 -125
rect 1166 -105 1253 -95
rect 1166 -125 1175 -105
rect 1195 -125 1253 -105
rect 1166 -134 1253 -125
rect 1166 -135 1203 -134
rect 27 -167 70 -162
rect 418 -156 865 -140
rect 418 -162 446 -156
rect 697 -157 865 -156
rect 27 -170 177 -167
rect 418 -170 445 -162
rect 27 -172 445 -170
rect 27 -190 36 -172
rect 54 -190 445 -172
rect 1222 -185 1253 -134
rect 1288 -105 1325 -35
rect 1591 -36 1628 -35
rect 1440 -95 1476 -94
rect 1288 -125 1297 -105
rect 1317 -125 1325 -105
rect 1288 -135 1325 -125
rect 1384 -105 1532 -95
rect 1632 -98 1728 -96
rect 1384 -125 1393 -105
rect 1413 -125 1503 -105
rect 1523 -125 1532 -105
rect 1384 -134 1532 -125
rect 1590 -105 1728 -98
rect 1590 -125 1599 -105
rect 1619 -125 1728 -105
rect 1590 -134 1728 -125
rect 1384 -135 1421 -134
rect 1114 -188 1155 -187
rect 27 -193 445 -190
rect 27 -199 70 -193
rect 30 -202 70 -199
rect 1006 -195 1155 -188
rect 427 -211 467 -210
rect 138 -228 467 -211
rect 1006 -215 1065 -195
rect 1085 -215 1124 -195
rect 1144 -215 1155 -195
rect 1006 -223 1155 -215
rect 1222 -192 1379 -185
rect 1222 -212 1342 -192
rect 1362 -212 1379 -192
rect 1222 -222 1379 -212
rect 1222 -223 1257 -222
rect 22 -271 65 -260
rect 22 -289 34 -271
rect 52 -289 65 -271
rect 22 -315 65 -289
rect 138 -315 165 -228
rect 427 -237 467 -228
rect 22 -336 165 -315
rect 209 -263 243 -247
rect 427 -257 820 -237
rect 840 -257 843 -237
rect 1222 -244 1253 -223
rect 1440 -244 1476 -134
rect 1495 -135 1532 -134
rect 1591 -135 1628 -134
rect 1551 -194 1641 -188
rect 1551 -214 1560 -194
rect 1580 -196 1641 -194
rect 1580 -214 1605 -196
rect 1551 -216 1605 -214
rect 1625 -216 1641 -196
rect 1551 -222 1641 -216
rect 1065 -245 1102 -244
rect 427 -262 843 -257
rect 1064 -254 1102 -245
rect 427 -263 768 -262
rect 209 -333 246 -263
rect 361 -323 392 -322
rect 22 -338 159 -336
rect 22 -380 65 -338
rect 209 -353 218 -333
rect 238 -353 246 -333
rect 209 -363 246 -353
rect 305 -333 392 -323
rect 305 -353 314 -333
rect 334 -353 392 -333
rect 305 -362 392 -353
rect 305 -363 342 -362
rect 20 -390 65 -380
rect 20 -408 29 -390
rect 47 -408 65 -390
rect 20 -414 65 -408
rect 361 -413 392 -362
rect 427 -333 464 -263
rect 730 -264 767 -263
rect 1064 -274 1073 -254
rect 1093 -274 1102 -254
rect 1064 -282 1102 -274
rect 1168 -250 1253 -244
rect 1283 -245 1320 -244
rect 1168 -270 1176 -250
rect 1196 -270 1253 -250
rect 1168 -278 1253 -270
rect 1282 -254 1320 -245
rect 1282 -274 1291 -254
rect 1311 -274 1320 -254
rect 1168 -279 1204 -278
rect 1282 -282 1320 -274
rect 1386 -250 1530 -244
rect 1386 -270 1394 -250
rect 1414 -270 1502 -250
rect 1522 -270 1530 -250
rect 1386 -278 1530 -270
rect 1386 -279 1422 -278
rect 1494 -279 1530 -278
rect 1596 -245 1633 -244
rect 1596 -246 1634 -245
rect 1596 -254 1660 -246
rect 1596 -274 1605 -254
rect 1625 -268 1660 -254
rect 1680 -268 1683 -248
rect 1625 -273 1683 -268
rect 1625 -274 1660 -273
rect 1065 -311 1102 -282
rect 1066 -313 1102 -311
rect 579 -323 615 -322
rect 427 -353 436 -333
rect 456 -353 464 -333
rect 427 -363 464 -353
rect 523 -333 671 -323
rect 771 -326 867 -324
rect 523 -353 532 -333
rect 552 -353 642 -333
rect 662 -353 671 -333
rect 523 -362 671 -353
rect 729 -333 867 -326
rect 729 -353 738 -333
rect 758 -353 867 -333
rect 1066 -335 1257 -313
rect 1283 -314 1320 -282
rect 1596 -286 1660 -274
rect 1700 -312 1727 -134
rect 1559 -314 1727 -312
rect 1283 -340 1727 -314
rect 729 -362 867 -353
rect 523 -363 560 -362
rect 20 -417 57 -414
rect 253 -416 294 -415
rect 145 -423 294 -416
rect 145 -443 204 -423
rect 224 -443 263 -423
rect 283 -443 294 -423
rect 145 -451 294 -443
rect 361 -420 518 -413
rect 361 -440 481 -420
rect 501 -440 518 -420
rect 361 -450 518 -440
rect 361 -451 396 -450
rect 361 -472 392 -451
rect 579 -472 615 -362
rect 634 -363 671 -362
rect 730 -363 767 -362
rect 690 -422 780 -416
rect 690 -442 699 -422
rect 719 -424 780 -422
rect 719 -442 744 -424
rect 690 -444 744 -442
rect 764 -444 780 -424
rect 690 -450 780 -444
rect 204 -473 241 -472
rect 17 -481 54 -479
rect 17 -489 59 -481
rect 17 -507 27 -489
rect 45 -507 59 -489
rect 17 -516 59 -507
rect 203 -482 241 -473
rect 203 -502 212 -482
rect 232 -502 241 -482
rect 203 -510 241 -502
rect 307 -478 392 -472
rect 422 -473 459 -472
rect 307 -498 315 -478
rect 335 -498 392 -478
rect 307 -506 392 -498
rect 421 -482 459 -473
rect 421 -502 430 -482
rect 450 -502 459 -482
rect 307 -507 343 -506
rect 421 -510 459 -502
rect 525 -474 669 -472
rect 525 -478 577 -474
rect 525 -498 533 -478
rect 553 -494 577 -478
rect 597 -478 669 -474
rect 597 -494 641 -478
rect 553 -498 641 -494
rect 661 -498 669 -478
rect 525 -506 669 -498
rect 525 -507 561 -506
rect 633 -507 669 -506
rect 735 -473 772 -472
rect 735 -474 773 -473
rect 735 -482 799 -474
rect 735 -502 744 -482
rect 764 -496 799 -482
rect 819 -496 822 -476
rect 764 -501 822 -496
rect 764 -502 799 -501
rect 18 -541 59 -516
rect 204 -541 241 -510
rect 422 -541 459 -510
rect 735 -514 799 -502
rect 839 -540 866 -362
rect 18 -542 502 -541
rect 698 -542 866 -540
rect 18 -567 866 -542
rect 18 -568 59 -567
rect 422 -568 866 -567
rect 698 -569 866 -568
rect 1393 -564 1433 -340
rect 1559 -341 1727 -340
rect 1393 -586 1401 -564
rect 1425 -586 1433 -564
rect 1393 -594 1433 -586
<< viali >>
rect 819 155 839 175
rect 203 -31 223 -11
rect 743 -32 763 -12
rect 585 -86 605 -66
rect 798 -84 818 -64
rect 1681 -29 1701 -9
rect 1065 -215 1085 -195
rect 820 -257 840 -237
rect 1605 -216 1625 -196
rect 1660 -268 1680 -248
rect 204 -443 224 -423
rect 744 -444 764 -424
rect 577 -494 597 -474
rect 799 -496 819 -476
rect 1401 -586 1425 -564
<< metal1 >>
rect 815 180 847 181
rect 812 175 847 180
rect 812 155 819 175
rect 839 155 847 175
rect 812 147 847 155
rect 194 -11 779 -3
rect 194 -31 203 -11
rect 223 -12 779 -11
rect 223 -31 743 -12
rect 194 -32 743 -31
rect 763 -32 779 -12
rect 194 -38 779 -32
rect 813 -59 847 147
rect 577 -66 612 -59
rect 577 -86 585 -66
rect 605 -86 612 -66
rect 577 -159 612 -86
rect 791 -64 847 -59
rect 791 -84 798 -64
rect 818 -84 847 -64
rect 791 -91 847 -84
rect 882 43 912 45
rect 1675 43 1708 44
rect 882 17 1709 43
rect 791 -92 826 -91
rect 882 -158 912 17
rect 1675 -4 1709 17
rect 1674 -9 1709 -4
rect 1674 -29 1681 -9
rect 1701 -29 1709 -9
rect 1674 -37 1709 -29
rect 877 -159 912 -158
rect 576 -186 912 -159
rect 882 -187 912 -186
rect 1056 -195 1641 -187
rect 1056 -215 1065 -195
rect 1085 -196 1641 -195
rect 1085 -215 1605 -196
rect 1056 -216 1605 -215
rect 1625 -216 1641 -196
rect 1056 -222 1641 -216
rect 816 -232 848 -231
rect 813 -237 848 -232
rect 813 -257 820 -237
rect 840 -257 848 -237
rect 1675 -243 1709 -37
rect 813 -265 848 -257
rect 195 -423 780 -415
rect 195 -443 204 -423
rect 224 -424 780 -423
rect 224 -443 744 -424
rect 195 -444 744 -443
rect 764 -444 780 -424
rect 195 -450 780 -444
rect 569 -474 608 -470
rect 814 -471 848 -265
rect 1653 -248 1709 -243
rect 1653 -268 1660 -248
rect 1680 -268 1709 -248
rect 1653 -275 1709 -268
rect 1653 -276 1688 -275
rect 569 -494 577 -474
rect 597 -494 608 -474
rect 569 -569 608 -494
rect 792 -476 848 -471
rect 792 -496 799 -476
rect 819 -496 848 -476
rect 792 -503 848 -496
rect 792 -504 827 -503
rect 1396 -564 1435 -551
rect 1396 -569 1401 -564
rect 569 -586 1401 -569
rect 1425 -569 1435 -564
rect 1425 -586 1436 -569
rect 569 -594 1436 -586
rect 571 -595 857 -594
<< labels >>
rlabel locali 157 -29 179 -14 1 d0
rlabel locali 211 159 240 165 1 vdd
rlabel locali 208 -140 237 -134 1 gnd
rlabel space 314 -122 343 -113 1 gnd
rlabel nwell 346 136 369 139 1 vdd
rlabel locali 158 -441 180 -426 1 d0
rlabel locali 212 -253 241 -247 1 vdd
rlabel locali 209 -552 238 -546 1 gnd
rlabel space 315 -534 344 -525 1 gnd
rlabel nwell 347 -276 370 -273 1 vdd
rlabel locali 1073 -25 1102 -19 1 vdd
rlabel locali 1070 -324 1099 -318 1 gnd
rlabel space 1176 -306 1205 -297 1 gnd
rlabel nwell 1208 -48 1231 -45 1 vdd
rlabel locali 1446 -178 1468 -163 1 vout
rlabel locali 1442 -333 1481 -330 1 vrefl
rlabel locali 1440 -21 1479 -18 1 vrefh
rlabel locali 1013 -217 1035 -200 1 d1
rlabel locali 48 404 72 434 1 vref
rlabel locali 24 -553 52 -535 1 gnd
<< end >>

magic
tech sky130A
timestamp 1616132309
<< nwell >>
rect 3450 8615 4058 8765
rect 7814 8628 8422 8778
rect 12191 8640 12799 8790
rect 16555 8653 17163 8803
rect 401 8461 1009 8611
rect 1199 8277 1807 8427
rect 2653 8387 3261 8537
rect 4765 8474 5373 8624
rect 3451 8203 4059 8353
rect 5563 8290 6171 8440
rect 7017 8400 7625 8550
rect 9142 8486 9750 8636
rect 7815 8216 8423 8366
rect 9940 8302 10548 8452
rect 11394 8412 12002 8562
rect 13506 8499 14114 8649
rect 20821 8627 21429 8777
rect 25185 8640 25793 8790
rect 29562 8652 30170 8802
rect 33926 8665 34534 8815
rect 12192 8228 12800 8378
rect 14304 8315 14912 8465
rect 15758 8425 16366 8575
rect 17772 8473 18380 8623
rect 16556 8241 17164 8391
rect 18570 8289 19178 8439
rect 20024 8399 20632 8549
rect 22136 8486 22744 8636
rect 402 8049 1010 8199
rect 2554 7977 3162 8127
rect 4766 8062 5374 8212
rect 6918 7990 7526 8140
rect 9143 8074 9751 8224
rect 11295 8002 11903 8152
rect 13507 8087 14115 8237
rect 20822 8215 21430 8365
rect 22934 8302 23542 8452
rect 24388 8412 24996 8562
rect 26513 8498 27121 8648
rect 25186 8228 25794 8378
rect 27311 8314 27919 8464
rect 28765 8424 29373 8574
rect 30877 8511 31485 8661
rect 29563 8240 30171 8390
rect 31675 8327 32283 8477
rect 33129 8437 33737 8587
rect 33927 8253 34535 8403
rect 15659 8015 16267 8165
rect 17773 8061 18381 8211
rect 19925 7989 20533 8139
rect 22137 8074 22745 8224
rect 24289 8002 24897 8152
rect 26514 8086 27122 8236
rect 28666 8014 29274 8164
rect 30878 8099 31486 8249
rect 33030 8027 33638 8177
rect 1281 7669 1889 7819
rect 3433 7597 4041 7747
rect 5645 7682 6253 7832
rect 7797 7610 8405 7760
rect 10022 7694 10630 7844
rect 12174 7622 12782 7772
rect 14386 7707 14994 7857
rect 16538 7635 17146 7785
rect 18652 7681 19260 7831
rect 384 7443 992 7593
rect 1182 7259 1790 7409
rect 2636 7369 3244 7519
rect 4748 7456 5356 7606
rect 3434 7185 4042 7335
rect 5546 7272 6154 7422
rect 7000 7382 7608 7532
rect 9125 7468 9733 7618
rect 7798 7198 8406 7348
rect 9923 7284 10531 7434
rect 11377 7394 11985 7544
rect 13489 7481 14097 7631
rect 20804 7609 21412 7759
rect 23016 7694 23624 7844
rect 25168 7622 25776 7772
rect 27393 7706 28001 7856
rect 29545 7634 30153 7784
rect 31757 7719 32365 7869
rect 33909 7647 34517 7797
rect 12175 7210 12783 7360
rect 14287 7297 14895 7447
rect 15741 7407 16349 7557
rect 17755 7455 18363 7605
rect 16539 7223 17147 7373
rect 18553 7271 19161 7421
rect 20007 7381 20615 7531
rect 22119 7468 22727 7618
rect 385 7031 993 7181
rect 2471 6961 3079 7111
rect 4749 7044 5357 7194
rect 6835 6974 7443 7124
rect 9126 7056 9734 7206
rect 11212 6986 11820 7136
rect 13490 7069 14098 7219
rect 20805 7197 21413 7347
rect 22917 7284 23525 7434
rect 24371 7394 24979 7544
rect 26496 7480 27104 7630
rect 25169 7210 25777 7360
rect 27294 7296 27902 7446
rect 28748 7406 29356 7556
rect 30860 7493 31468 7643
rect 29546 7222 30154 7372
rect 31658 7309 32266 7459
rect 33112 7419 33720 7569
rect 33910 7235 34518 7385
rect 15576 6999 16184 7149
rect 17756 7043 18364 7193
rect 19842 6973 20450 7123
rect 22120 7056 22728 7206
rect 24206 6986 24814 7136
rect 26497 7068 27105 7218
rect 28583 6998 29191 7148
rect 30861 7081 31469 7231
rect 32947 7011 33555 7161
rect 1327 6649 1935 6799
rect 3413 6579 4021 6729
rect 5691 6662 6299 6812
rect 7777 6592 8385 6742
rect 10068 6674 10676 6824
rect 12154 6604 12762 6754
rect 14432 6687 15040 6837
rect 16518 6617 17126 6767
rect 18698 6661 19306 6811
rect 364 6425 972 6575
rect 1162 6241 1770 6391
rect 2616 6351 3224 6501
rect 4728 6438 5336 6588
rect 3414 6167 4022 6317
rect 5526 6254 6134 6404
rect 6980 6364 7588 6514
rect 9105 6450 9713 6600
rect 7778 6180 8386 6330
rect 9903 6266 10511 6416
rect 11357 6376 11965 6526
rect 13469 6463 14077 6613
rect 20784 6591 21392 6741
rect 23062 6674 23670 6824
rect 25148 6604 25756 6754
rect 27439 6686 28047 6836
rect 29525 6616 30133 6766
rect 31803 6699 32411 6849
rect 33889 6629 34497 6779
rect 12155 6192 12763 6342
rect 14267 6279 14875 6429
rect 15721 6389 16329 6539
rect 17735 6437 18343 6587
rect 16519 6205 17127 6355
rect 18533 6253 19141 6403
rect 19987 6363 20595 6513
rect 22099 6450 22707 6600
rect 365 6013 973 6163
rect 2517 5941 3125 6091
rect 4729 6026 5337 6176
rect 6881 5954 7489 6104
rect 9106 6038 9714 6188
rect 11258 5966 11866 6116
rect 13470 6051 14078 6201
rect 20785 6179 21393 6329
rect 22897 6266 23505 6416
rect 24351 6376 24959 6526
rect 26476 6462 27084 6612
rect 25149 6192 25757 6342
rect 27274 6278 27882 6428
rect 28728 6388 29336 6538
rect 30840 6475 31448 6625
rect 29526 6204 30134 6354
rect 31638 6291 32246 6441
rect 33092 6401 33700 6551
rect 33890 6217 34498 6367
rect 15622 5979 16230 6129
rect 17736 6025 18344 6175
rect 19888 5953 20496 6103
rect 22100 6038 22708 6188
rect 24252 5966 24860 6116
rect 26477 6050 27085 6200
rect 28629 5978 29237 6128
rect 30841 6063 31449 6213
rect 32993 5991 33601 6141
rect 1244 5633 1852 5783
rect 3396 5561 4004 5711
rect 5608 5646 6216 5796
rect 7760 5574 8368 5724
rect 9985 5658 10593 5808
rect 12137 5586 12745 5736
rect 14349 5671 14957 5821
rect 16501 5599 17109 5749
rect 18615 5645 19223 5795
rect 347 5407 955 5557
rect 1145 5223 1753 5373
rect 2599 5333 3207 5483
rect 4711 5420 5319 5570
rect 3397 5149 4005 5299
rect 5509 5236 6117 5386
rect 6963 5346 7571 5496
rect 9088 5432 9696 5582
rect 7761 5162 8369 5312
rect 9886 5248 10494 5398
rect 11340 5358 11948 5508
rect 13452 5445 14060 5595
rect 20767 5573 21375 5723
rect 22979 5658 23587 5808
rect 25131 5586 25739 5736
rect 27356 5670 27964 5820
rect 29508 5598 30116 5748
rect 31720 5683 32328 5833
rect 33872 5611 34480 5761
rect 12138 5174 12746 5324
rect 14250 5261 14858 5411
rect 15704 5371 16312 5521
rect 17718 5419 18326 5569
rect 16502 5187 17110 5337
rect 18516 5235 19124 5385
rect 19970 5345 20578 5495
rect 22082 5432 22690 5582
rect 348 4995 956 5145
rect 2295 4927 2903 5077
rect 4712 5008 5320 5158
rect 6659 4940 7267 5090
rect 9089 5020 9697 5170
rect 11036 4952 11644 5102
rect 13453 5033 14061 5183
rect 20768 5161 21376 5311
rect 22880 5248 23488 5398
rect 24334 5358 24942 5508
rect 26459 5444 27067 5594
rect 25132 5174 25740 5324
rect 27257 5260 27865 5410
rect 28711 5370 29319 5520
rect 30823 5457 31431 5607
rect 29509 5186 30117 5336
rect 31621 5273 32229 5423
rect 33075 5383 33683 5533
rect 33873 5199 34481 5349
rect 15400 4965 16008 5115
rect 17719 5007 18327 5157
rect 19666 4939 20274 5089
rect 22083 5020 22691 5170
rect 24030 4952 24638 5102
rect 26460 5032 27068 5182
rect 28407 4964 29015 5114
rect 30824 5045 31432 5195
rect 32771 4977 33379 5127
rect 1430 4611 2038 4761
rect 3377 4543 3985 4693
rect 5794 4624 6402 4774
rect 7741 4556 8349 4706
rect 10171 4636 10779 4786
rect 12118 4568 12726 4718
rect 14535 4649 15143 4799
rect 16482 4581 17090 4731
rect 18801 4623 19409 4773
rect 328 4389 936 4539
rect 1126 4205 1734 4355
rect 2580 4315 3188 4465
rect 4692 4402 5300 4552
rect 3378 4131 3986 4281
rect 5490 4218 6098 4368
rect 6944 4328 7552 4478
rect 9069 4414 9677 4564
rect 7742 4144 8350 4294
rect 9867 4230 10475 4380
rect 11321 4340 11929 4490
rect 13433 4427 14041 4577
rect 20748 4555 21356 4705
rect 23165 4636 23773 4786
rect 25112 4568 25720 4718
rect 27542 4648 28150 4798
rect 29489 4580 30097 4730
rect 31906 4661 32514 4811
rect 33853 4593 34461 4743
rect 12119 4156 12727 4306
rect 14231 4243 14839 4393
rect 15685 4353 16293 4503
rect 17699 4401 18307 4551
rect 16483 4169 17091 4319
rect 18497 4217 19105 4367
rect 19951 4327 20559 4477
rect 22063 4414 22671 4564
rect 329 3977 937 4127
rect 2481 3905 3089 4055
rect 4693 3990 5301 4140
rect 6845 3918 7453 4068
rect 9070 4002 9678 4152
rect 11222 3930 11830 4080
rect 13434 4015 14042 4165
rect 20749 4143 21357 4293
rect 22861 4230 23469 4380
rect 24315 4340 24923 4490
rect 26440 4426 27048 4576
rect 25113 4156 25721 4306
rect 27238 4242 27846 4392
rect 28692 4352 29300 4502
rect 30804 4439 31412 4589
rect 29490 4168 30098 4318
rect 31602 4255 32210 4405
rect 33056 4365 33664 4515
rect 33854 4181 34462 4331
rect 15586 3943 16194 4093
rect 17700 3989 18308 4139
rect 19852 3917 20460 4067
rect 22064 4002 22672 4152
rect 24216 3930 24824 4080
rect 26441 4014 27049 4164
rect 28593 3942 29201 4092
rect 30805 4027 31413 4177
rect 32957 3955 33565 4105
rect 1208 3597 1816 3747
rect 3360 3525 3968 3675
rect 5572 3610 6180 3760
rect 7724 3538 8332 3688
rect 9949 3622 10557 3772
rect 12101 3550 12709 3700
rect 14313 3635 14921 3785
rect 16465 3563 17073 3713
rect 18579 3609 19187 3759
rect 311 3371 919 3521
rect 1109 3187 1717 3337
rect 2563 3297 3171 3447
rect 4675 3384 5283 3534
rect 3361 3113 3969 3263
rect 5473 3200 6081 3350
rect 6927 3310 7535 3460
rect 9052 3396 9660 3546
rect 7725 3126 8333 3276
rect 9850 3212 10458 3362
rect 11304 3322 11912 3472
rect 13416 3409 14024 3559
rect 20731 3537 21339 3687
rect 22943 3622 23551 3772
rect 25095 3550 25703 3700
rect 27320 3634 27928 3784
rect 29472 3562 30080 3712
rect 31684 3647 32292 3797
rect 33836 3575 34444 3725
rect 12102 3138 12710 3288
rect 14214 3225 14822 3375
rect 15668 3335 16276 3485
rect 17682 3383 18290 3533
rect 16466 3151 17074 3301
rect 18480 3199 19088 3349
rect 19934 3309 20542 3459
rect 22046 3396 22654 3546
rect 312 2959 920 3109
rect 2398 2889 3006 3039
rect 4676 2972 5284 3122
rect 6762 2902 7370 3052
rect 9053 2984 9661 3134
rect 11139 2914 11747 3064
rect 13417 2997 14025 3147
rect 20732 3125 21340 3275
rect 22844 3212 23452 3362
rect 24298 3322 24906 3472
rect 26423 3408 27031 3558
rect 25096 3138 25704 3288
rect 27221 3224 27829 3374
rect 28675 3334 29283 3484
rect 30787 3421 31395 3571
rect 29473 3150 30081 3300
rect 31585 3237 32193 3387
rect 33039 3347 33647 3497
rect 33837 3163 34445 3313
rect 15503 2927 16111 3077
rect 17683 2971 18291 3121
rect 19769 2901 20377 3051
rect 22047 2984 22655 3134
rect 24133 2914 24741 3064
rect 26424 2996 27032 3146
rect 28510 2926 29118 3076
rect 30788 3009 31396 3159
rect 32874 2939 33482 3089
rect 1254 2577 1862 2727
rect 3340 2507 3948 2657
rect 5618 2590 6226 2740
rect 7704 2520 8312 2670
rect 9995 2602 10603 2752
rect 12081 2532 12689 2682
rect 14359 2615 14967 2765
rect 16445 2545 17053 2695
rect 18625 2589 19233 2739
rect 291 2353 899 2503
rect 1089 2169 1697 2319
rect 2543 2279 3151 2429
rect 4655 2366 5263 2516
rect 3341 2095 3949 2245
rect 5453 2182 6061 2332
rect 6907 2292 7515 2442
rect 9032 2378 9640 2528
rect 7705 2108 8313 2258
rect 9830 2194 10438 2344
rect 11284 2304 11892 2454
rect 13396 2391 14004 2541
rect 20711 2519 21319 2669
rect 22989 2602 23597 2752
rect 25075 2532 25683 2682
rect 27366 2614 27974 2764
rect 29452 2544 30060 2694
rect 31730 2627 32338 2777
rect 33816 2557 34424 2707
rect 12082 2120 12690 2270
rect 14194 2207 14802 2357
rect 15648 2317 16256 2467
rect 17662 2365 18270 2515
rect 16446 2133 17054 2283
rect 18460 2181 19068 2331
rect 19914 2291 20522 2441
rect 22026 2378 22634 2528
rect 292 1941 900 2091
rect 2444 1869 3052 2019
rect 4656 1954 5264 2104
rect 6808 1882 7416 2032
rect 9033 1966 9641 2116
rect 11185 1894 11793 2044
rect 13397 1979 14005 2129
rect 20712 2107 21320 2257
rect 22824 2194 23432 2344
rect 24278 2304 24886 2454
rect 26403 2390 27011 2540
rect 25076 2120 25684 2270
rect 27201 2206 27809 2356
rect 28655 2316 29263 2466
rect 30767 2403 31375 2553
rect 29453 2132 30061 2282
rect 31565 2219 32173 2369
rect 33019 2329 33627 2479
rect 33817 2145 34425 2295
rect 15549 1907 16157 2057
rect 17663 1953 18271 2103
rect 19815 1881 20423 2031
rect 22027 1966 22635 2116
rect 24179 1894 24787 2044
rect 26404 1978 27012 2128
rect 28556 1906 29164 2056
rect 30768 1991 31376 2141
rect 32920 1919 33528 2069
rect 1171 1561 1779 1711
rect 3323 1489 3931 1639
rect 5535 1574 6143 1724
rect 7687 1502 8295 1652
rect 9912 1586 10520 1736
rect 12064 1514 12672 1664
rect 14276 1599 14884 1749
rect 16428 1527 17036 1677
rect 18542 1573 19150 1723
rect 274 1335 882 1485
rect 1072 1151 1680 1301
rect 2526 1261 3134 1411
rect 4638 1348 5246 1498
rect 3324 1077 3932 1227
rect 5436 1164 6044 1314
rect 6890 1274 7498 1424
rect 9015 1360 9623 1510
rect 7688 1090 8296 1240
rect 9813 1176 10421 1326
rect 11267 1286 11875 1436
rect 13379 1373 13987 1523
rect 20694 1501 21302 1651
rect 22906 1586 23514 1736
rect 25058 1514 25666 1664
rect 27283 1598 27891 1748
rect 29435 1526 30043 1676
rect 31647 1611 32255 1761
rect 33799 1539 34407 1689
rect 12065 1102 12673 1252
rect 14177 1189 14785 1339
rect 15631 1299 16239 1449
rect 17645 1347 18253 1497
rect 16429 1115 17037 1265
rect 18443 1163 19051 1313
rect 19897 1273 20505 1423
rect 22009 1360 22617 1510
rect 275 923 883 1073
rect 4639 936 5247 1086
rect 9016 948 9624 1098
rect 13380 961 13988 1111
rect 20695 1089 21303 1239
rect 22807 1176 23415 1326
rect 24261 1286 24869 1436
rect 26386 1372 26994 1522
rect 25059 1102 25667 1252
rect 27184 1188 27792 1338
rect 28638 1298 29246 1448
rect 30750 1385 31358 1535
rect 29436 1114 30044 1264
rect 31548 1201 32156 1351
rect 33002 1311 33610 1461
rect 33800 1127 34408 1277
rect 17646 935 18254 1085
rect 22010 948 22618 1098
rect 26387 960 26995 1110
rect 30751 973 31359 1123
rect 1488 347 2096 497
rect 3977 273 4585 423
rect 5852 360 6460 510
rect 8425 297 9033 447
rect 10229 372 10837 522
rect 12718 298 13326 448
rect 14593 385 15201 535
rect 16915 234 17523 384
rect 18859 359 19467 509
rect 21348 285 21956 435
rect 23223 372 23831 522
rect 25796 309 26404 459
rect 27600 384 28208 534
rect 30089 310 30697 460
rect 31964 397 32572 547
<< nmos >>
rect 3518 8824 3568 8866
rect 3726 8824 3776 8866
rect 3944 8824 3994 8866
rect 7882 8837 7932 8879
rect 8090 8837 8140 8879
rect 8308 8837 8358 8879
rect 12259 8849 12309 8891
rect 12467 8849 12517 8891
rect 12685 8849 12735 8891
rect 2721 8596 2771 8638
rect 2929 8596 2979 8638
rect 3147 8596 3197 8638
rect 16623 8862 16673 8904
rect 16831 8862 16881 8904
rect 17049 8862 17099 8904
rect 7085 8609 7135 8651
rect 7293 8609 7343 8651
rect 7511 8609 7561 8651
rect 20889 8836 20939 8878
rect 21097 8836 21147 8878
rect 21315 8836 21365 8878
rect 11462 8621 11512 8663
rect 11670 8621 11720 8663
rect 11888 8621 11938 8663
rect 25253 8849 25303 8891
rect 25461 8849 25511 8891
rect 25679 8849 25729 8891
rect 15826 8634 15876 8676
rect 16034 8634 16084 8676
rect 16252 8634 16302 8676
rect 29630 8861 29680 8903
rect 29838 8861 29888 8903
rect 30056 8861 30106 8903
rect 465 8360 515 8402
rect 683 8360 733 8402
rect 891 8360 941 8402
rect 3519 8412 3569 8454
rect 3727 8412 3777 8454
rect 3945 8412 3995 8454
rect 4829 8373 4879 8415
rect 5047 8373 5097 8415
rect 5255 8373 5305 8415
rect 7883 8425 7933 8467
rect 8091 8425 8141 8467
rect 8309 8425 8359 8467
rect 20092 8608 20142 8650
rect 20300 8608 20350 8650
rect 20518 8608 20568 8650
rect 33994 8874 34044 8916
rect 34202 8874 34252 8916
rect 34420 8874 34470 8916
rect 24456 8621 24506 8663
rect 24664 8621 24714 8663
rect 24882 8621 24932 8663
rect 28833 8633 28883 8675
rect 29041 8633 29091 8675
rect 29259 8633 29309 8675
rect 33197 8646 33247 8688
rect 33405 8646 33455 8688
rect 33623 8646 33673 8688
rect 9206 8385 9256 8427
rect 9424 8385 9474 8427
rect 9632 8385 9682 8427
rect 12260 8437 12310 8479
rect 12468 8437 12518 8479
rect 12686 8437 12736 8479
rect 1263 8176 1313 8218
rect 1481 8176 1531 8218
rect 1689 8176 1739 8218
rect 2622 8186 2672 8228
rect 2830 8186 2880 8228
rect 3048 8186 3098 8228
rect 13570 8398 13620 8440
rect 13788 8398 13838 8440
rect 13996 8398 14046 8440
rect 16624 8450 16674 8492
rect 16832 8450 16882 8492
rect 17050 8450 17100 8492
rect 5627 8189 5677 8231
rect 5845 8189 5895 8231
rect 6053 8189 6103 8231
rect 6986 8199 7036 8241
rect 7194 8199 7244 8241
rect 7412 8199 7462 8241
rect 10004 8201 10054 8243
rect 10222 8201 10272 8243
rect 10430 8201 10480 8243
rect 11363 8211 11413 8253
rect 11571 8211 11621 8253
rect 11789 8211 11839 8253
rect 17836 8372 17886 8414
rect 18054 8372 18104 8414
rect 18262 8372 18312 8414
rect 20890 8424 20940 8466
rect 21098 8424 21148 8466
rect 21316 8424 21366 8466
rect 22200 8385 22250 8427
rect 22418 8385 22468 8427
rect 22626 8385 22676 8427
rect 25254 8437 25304 8479
rect 25462 8437 25512 8479
rect 25680 8437 25730 8479
rect 466 7948 516 7990
rect 684 7948 734 7990
rect 892 7948 942 7990
rect 14368 8214 14418 8256
rect 14586 8214 14636 8256
rect 14794 8214 14844 8256
rect 15727 8224 15777 8266
rect 15935 8224 15985 8266
rect 16153 8224 16203 8266
rect 26577 8397 26627 8439
rect 26795 8397 26845 8439
rect 27003 8397 27053 8439
rect 29631 8449 29681 8491
rect 29839 8449 29889 8491
rect 30057 8449 30107 8491
rect 4830 7961 4880 8003
rect 5048 7961 5098 8003
rect 5256 7961 5306 8003
rect 18634 8188 18684 8230
rect 18852 8188 18902 8230
rect 19060 8188 19110 8230
rect 19993 8198 20043 8240
rect 20201 8198 20251 8240
rect 20419 8198 20469 8240
rect 30941 8410 30991 8452
rect 31159 8410 31209 8452
rect 31367 8410 31417 8452
rect 33995 8462 34045 8504
rect 34203 8462 34253 8504
rect 34421 8462 34471 8504
rect 9207 7973 9257 8015
rect 9425 7973 9475 8015
rect 9633 7973 9683 8015
rect 22998 8201 23048 8243
rect 23216 8201 23266 8243
rect 23424 8201 23474 8243
rect 24357 8211 24407 8253
rect 24565 8211 24615 8253
rect 24783 8211 24833 8253
rect 13571 7986 13621 8028
rect 13789 7986 13839 8028
rect 13997 7986 14047 8028
rect 27375 8213 27425 8255
rect 27593 8213 27643 8255
rect 27801 8213 27851 8255
rect 28734 8223 28784 8265
rect 28942 8223 28992 8265
rect 29160 8223 29210 8265
rect 17837 7960 17887 8002
rect 18055 7960 18105 8002
rect 18263 7960 18313 8002
rect 31739 8226 31789 8268
rect 31957 8226 32007 8268
rect 32165 8226 32215 8268
rect 33098 8236 33148 8278
rect 33306 8236 33356 8278
rect 33524 8236 33574 8278
rect 22201 7973 22251 8015
rect 22419 7973 22469 8015
rect 22627 7973 22677 8015
rect 26578 7985 26628 8027
rect 26796 7985 26846 8027
rect 27004 7985 27054 8027
rect 30942 7998 30992 8040
rect 31160 7998 31210 8040
rect 31368 7998 31418 8040
rect 3501 7806 3551 7848
rect 3709 7806 3759 7848
rect 3927 7806 3977 7848
rect 7865 7819 7915 7861
rect 8073 7819 8123 7861
rect 8291 7819 8341 7861
rect 12242 7831 12292 7873
rect 12450 7831 12500 7873
rect 12668 7831 12718 7873
rect 1345 7568 1395 7610
rect 1563 7568 1613 7610
rect 1771 7568 1821 7610
rect 2704 7578 2754 7620
rect 2912 7578 2962 7620
rect 3130 7578 3180 7620
rect 16606 7844 16656 7886
rect 16814 7844 16864 7886
rect 17032 7844 17082 7886
rect 5709 7581 5759 7623
rect 5927 7581 5977 7623
rect 6135 7581 6185 7623
rect 7068 7591 7118 7633
rect 7276 7591 7326 7633
rect 7494 7591 7544 7633
rect 20872 7818 20922 7860
rect 21080 7818 21130 7860
rect 21298 7818 21348 7860
rect 10086 7593 10136 7635
rect 10304 7593 10354 7635
rect 10512 7593 10562 7635
rect 11445 7603 11495 7645
rect 11653 7603 11703 7645
rect 11871 7603 11921 7645
rect 25236 7831 25286 7873
rect 25444 7831 25494 7873
rect 25662 7831 25712 7873
rect 448 7342 498 7384
rect 666 7342 716 7384
rect 874 7342 924 7384
rect 3502 7394 3552 7436
rect 3710 7394 3760 7436
rect 3928 7394 3978 7436
rect 14450 7606 14500 7648
rect 14668 7606 14718 7648
rect 14876 7606 14926 7648
rect 15809 7616 15859 7658
rect 16017 7616 16067 7658
rect 16235 7616 16285 7658
rect 29613 7843 29663 7885
rect 29821 7843 29871 7885
rect 30039 7843 30089 7885
rect 4812 7355 4862 7397
rect 5030 7355 5080 7397
rect 5238 7355 5288 7397
rect 7866 7407 7916 7449
rect 8074 7407 8124 7449
rect 8292 7407 8342 7449
rect 18716 7580 18766 7622
rect 18934 7580 18984 7622
rect 19142 7580 19192 7622
rect 20075 7590 20125 7632
rect 20283 7590 20333 7632
rect 20501 7590 20551 7632
rect 33977 7856 34027 7898
rect 34185 7856 34235 7898
rect 34403 7856 34453 7898
rect 9189 7367 9239 7409
rect 9407 7367 9457 7409
rect 9615 7367 9665 7409
rect 12243 7419 12293 7461
rect 12451 7419 12501 7461
rect 12669 7419 12719 7461
rect 1246 7158 1296 7200
rect 1464 7158 1514 7200
rect 1672 7158 1722 7200
rect 2539 7170 2589 7212
rect 2747 7170 2797 7212
rect 2965 7170 3015 7212
rect 13553 7380 13603 7422
rect 13771 7380 13821 7422
rect 13979 7380 14029 7422
rect 16607 7432 16657 7474
rect 16815 7432 16865 7474
rect 17033 7432 17083 7474
rect 23080 7593 23130 7635
rect 23298 7593 23348 7635
rect 23506 7593 23556 7635
rect 24439 7603 24489 7645
rect 24647 7603 24697 7645
rect 24865 7603 24915 7645
rect 5610 7171 5660 7213
rect 5828 7171 5878 7213
rect 6036 7171 6086 7213
rect 6903 7183 6953 7225
rect 7111 7183 7161 7225
rect 7329 7183 7379 7225
rect 27457 7605 27507 7647
rect 27675 7605 27725 7647
rect 27883 7605 27933 7647
rect 28816 7615 28866 7657
rect 29024 7615 29074 7657
rect 29242 7615 29292 7657
rect 9987 7183 10037 7225
rect 10205 7183 10255 7225
rect 10413 7183 10463 7225
rect 11280 7195 11330 7237
rect 11488 7195 11538 7237
rect 11706 7195 11756 7237
rect 17819 7354 17869 7396
rect 18037 7354 18087 7396
rect 18245 7354 18295 7396
rect 20873 7406 20923 7448
rect 21081 7406 21131 7448
rect 21299 7406 21349 7448
rect 31821 7618 31871 7660
rect 32039 7618 32089 7660
rect 32247 7618 32297 7660
rect 33180 7628 33230 7670
rect 33388 7628 33438 7670
rect 33606 7628 33656 7670
rect 22183 7367 22233 7409
rect 22401 7367 22451 7409
rect 22609 7367 22659 7409
rect 25237 7419 25287 7461
rect 25445 7419 25495 7461
rect 25663 7419 25713 7461
rect 449 6930 499 6972
rect 667 6930 717 6972
rect 875 6930 925 6972
rect 14351 7196 14401 7238
rect 14569 7196 14619 7238
rect 14777 7196 14827 7238
rect 15644 7208 15694 7250
rect 15852 7208 15902 7250
rect 16070 7208 16120 7250
rect 26560 7379 26610 7421
rect 26778 7379 26828 7421
rect 26986 7379 27036 7421
rect 29614 7431 29664 7473
rect 29822 7431 29872 7473
rect 30040 7431 30090 7473
rect 4813 6943 4863 6985
rect 5031 6943 5081 6985
rect 5239 6943 5289 6985
rect 18617 7170 18667 7212
rect 18835 7170 18885 7212
rect 19043 7170 19093 7212
rect 19910 7182 19960 7224
rect 20118 7182 20168 7224
rect 20336 7182 20386 7224
rect 30924 7392 30974 7434
rect 31142 7392 31192 7434
rect 31350 7392 31400 7434
rect 33978 7444 34028 7486
rect 34186 7444 34236 7486
rect 34404 7444 34454 7486
rect 9190 6955 9240 6997
rect 9408 6955 9458 6997
rect 9616 6955 9666 6997
rect 22981 7183 23031 7225
rect 23199 7183 23249 7225
rect 23407 7183 23457 7225
rect 24274 7195 24324 7237
rect 24482 7195 24532 7237
rect 24700 7195 24750 7237
rect 13554 6968 13604 7010
rect 13772 6968 13822 7010
rect 13980 6968 14030 7010
rect 27358 7195 27408 7237
rect 27576 7195 27626 7237
rect 27784 7195 27834 7237
rect 28651 7207 28701 7249
rect 28859 7207 28909 7249
rect 29077 7207 29127 7249
rect 17820 6942 17870 6984
rect 18038 6942 18088 6984
rect 18246 6942 18296 6984
rect 31722 7208 31772 7250
rect 31940 7208 31990 7250
rect 32148 7208 32198 7250
rect 33015 7220 33065 7262
rect 33223 7220 33273 7262
rect 33441 7220 33491 7262
rect 22184 6955 22234 6997
rect 22402 6955 22452 6997
rect 22610 6955 22660 6997
rect 26561 6967 26611 7009
rect 26779 6967 26829 7009
rect 26987 6967 27037 7009
rect 30925 6980 30975 7022
rect 31143 6980 31193 7022
rect 31351 6980 31401 7022
rect 3481 6788 3531 6830
rect 3689 6788 3739 6830
rect 3907 6788 3957 6830
rect 7845 6801 7895 6843
rect 8053 6801 8103 6843
rect 8271 6801 8321 6843
rect 12222 6813 12272 6855
rect 12430 6813 12480 6855
rect 12648 6813 12698 6855
rect 1391 6548 1441 6590
rect 1609 6548 1659 6590
rect 1817 6548 1867 6590
rect 2684 6560 2734 6602
rect 2892 6560 2942 6602
rect 3110 6560 3160 6602
rect 16586 6826 16636 6868
rect 16794 6826 16844 6868
rect 17012 6826 17062 6868
rect 5755 6561 5805 6603
rect 5973 6561 6023 6603
rect 6181 6561 6231 6603
rect 7048 6573 7098 6615
rect 7256 6573 7306 6615
rect 7474 6573 7524 6615
rect 20852 6800 20902 6842
rect 21060 6800 21110 6842
rect 21278 6800 21328 6842
rect 10132 6573 10182 6615
rect 10350 6573 10400 6615
rect 10558 6573 10608 6615
rect 11425 6585 11475 6627
rect 11633 6585 11683 6627
rect 11851 6585 11901 6627
rect 25216 6813 25266 6855
rect 25424 6813 25474 6855
rect 25642 6813 25692 6855
rect 428 6324 478 6366
rect 646 6324 696 6366
rect 854 6324 904 6366
rect 3482 6376 3532 6418
rect 3690 6376 3740 6418
rect 3908 6376 3958 6418
rect 14496 6586 14546 6628
rect 14714 6586 14764 6628
rect 14922 6586 14972 6628
rect 15789 6598 15839 6640
rect 15997 6598 16047 6640
rect 16215 6598 16265 6640
rect 29593 6825 29643 6867
rect 29801 6825 29851 6867
rect 30019 6825 30069 6867
rect 4792 6337 4842 6379
rect 5010 6337 5060 6379
rect 5218 6337 5268 6379
rect 7846 6389 7896 6431
rect 8054 6389 8104 6431
rect 8272 6389 8322 6431
rect 18762 6560 18812 6602
rect 18980 6560 19030 6602
rect 19188 6560 19238 6602
rect 20055 6572 20105 6614
rect 20263 6572 20313 6614
rect 20481 6572 20531 6614
rect 33957 6838 34007 6880
rect 34165 6838 34215 6880
rect 34383 6838 34433 6880
rect 9169 6349 9219 6391
rect 9387 6349 9437 6391
rect 9595 6349 9645 6391
rect 12223 6401 12273 6443
rect 12431 6401 12481 6443
rect 12649 6401 12699 6443
rect 1226 6140 1276 6182
rect 1444 6140 1494 6182
rect 1652 6140 1702 6182
rect 2585 6150 2635 6192
rect 2793 6150 2843 6192
rect 3011 6150 3061 6192
rect 13533 6362 13583 6404
rect 13751 6362 13801 6404
rect 13959 6362 14009 6404
rect 16587 6414 16637 6456
rect 16795 6414 16845 6456
rect 17013 6414 17063 6456
rect 23126 6573 23176 6615
rect 23344 6573 23394 6615
rect 23552 6573 23602 6615
rect 24419 6585 24469 6627
rect 24627 6585 24677 6627
rect 24845 6585 24895 6627
rect 5590 6153 5640 6195
rect 5808 6153 5858 6195
rect 6016 6153 6066 6195
rect 6949 6163 6999 6205
rect 7157 6163 7207 6205
rect 7375 6163 7425 6205
rect 27503 6585 27553 6627
rect 27721 6585 27771 6627
rect 27929 6585 27979 6627
rect 28796 6597 28846 6639
rect 29004 6597 29054 6639
rect 29222 6597 29272 6639
rect 9967 6165 10017 6207
rect 10185 6165 10235 6207
rect 10393 6165 10443 6207
rect 11326 6175 11376 6217
rect 11534 6175 11584 6217
rect 11752 6175 11802 6217
rect 17799 6336 17849 6378
rect 18017 6336 18067 6378
rect 18225 6336 18275 6378
rect 20853 6388 20903 6430
rect 21061 6388 21111 6430
rect 21279 6388 21329 6430
rect 31867 6598 31917 6640
rect 32085 6598 32135 6640
rect 32293 6598 32343 6640
rect 33160 6610 33210 6652
rect 33368 6610 33418 6652
rect 33586 6610 33636 6652
rect 22163 6349 22213 6391
rect 22381 6349 22431 6391
rect 22589 6349 22639 6391
rect 25217 6401 25267 6443
rect 25425 6401 25475 6443
rect 25643 6401 25693 6443
rect 429 5912 479 5954
rect 647 5912 697 5954
rect 855 5912 905 5954
rect 14331 6178 14381 6220
rect 14549 6178 14599 6220
rect 14757 6178 14807 6220
rect 15690 6188 15740 6230
rect 15898 6188 15948 6230
rect 16116 6188 16166 6230
rect 26540 6361 26590 6403
rect 26758 6361 26808 6403
rect 26966 6361 27016 6403
rect 29594 6413 29644 6455
rect 29802 6413 29852 6455
rect 30020 6413 30070 6455
rect 4793 5925 4843 5967
rect 5011 5925 5061 5967
rect 5219 5925 5269 5967
rect 18597 6152 18647 6194
rect 18815 6152 18865 6194
rect 19023 6152 19073 6194
rect 19956 6162 20006 6204
rect 20164 6162 20214 6204
rect 20382 6162 20432 6204
rect 30904 6374 30954 6416
rect 31122 6374 31172 6416
rect 31330 6374 31380 6416
rect 33958 6426 34008 6468
rect 34166 6426 34216 6468
rect 34384 6426 34434 6468
rect 9170 5937 9220 5979
rect 9388 5937 9438 5979
rect 9596 5937 9646 5979
rect 22961 6165 23011 6207
rect 23179 6165 23229 6207
rect 23387 6165 23437 6207
rect 24320 6175 24370 6217
rect 24528 6175 24578 6217
rect 24746 6175 24796 6217
rect 13534 5950 13584 5992
rect 13752 5950 13802 5992
rect 13960 5950 14010 5992
rect 27338 6177 27388 6219
rect 27556 6177 27606 6219
rect 27764 6177 27814 6219
rect 28697 6187 28747 6229
rect 28905 6187 28955 6229
rect 29123 6187 29173 6229
rect 17800 5924 17850 5966
rect 18018 5924 18068 5966
rect 18226 5924 18276 5966
rect 31702 6190 31752 6232
rect 31920 6190 31970 6232
rect 32128 6190 32178 6232
rect 33061 6200 33111 6242
rect 33269 6200 33319 6242
rect 33487 6200 33537 6242
rect 22164 5937 22214 5979
rect 22382 5937 22432 5979
rect 22590 5937 22640 5979
rect 26541 5949 26591 5991
rect 26759 5949 26809 5991
rect 26967 5949 27017 5991
rect 30905 5962 30955 6004
rect 31123 5962 31173 6004
rect 31331 5962 31381 6004
rect 3464 5770 3514 5812
rect 3672 5770 3722 5812
rect 3890 5770 3940 5812
rect 7828 5783 7878 5825
rect 8036 5783 8086 5825
rect 8254 5783 8304 5825
rect 12205 5795 12255 5837
rect 12413 5795 12463 5837
rect 12631 5795 12681 5837
rect 1308 5532 1358 5574
rect 1526 5532 1576 5574
rect 1734 5532 1784 5574
rect 2667 5542 2717 5584
rect 2875 5542 2925 5584
rect 3093 5542 3143 5584
rect 16569 5808 16619 5850
rect 16777 5808 16827 5850
rect 16995 5808 17045 5850
rect 5672 5545 5722 5587
rect 5890 5545 5940 5587
rect 6098 5545 6148 5587
rect 7031 5555 7081 5597
rect 7239 5555 7289 5597
rect 7457 5555 7507 5597
rect 20835 5782 20885 5824
rect 21043 5782 21093 5824
rect 21261 5782 21311 5824
rect 10049 5557 10099 5599
rect 10267 5557 10317 5599
rect 10475 5557 10525 5599
rect 11408 5567 11458 5609
rect 11616 5567 11666 5609
rect 11834 5567 11884 5609
rect 25199 5795 25249 5837
rect 25407 5795 25457 5837
rect 25625 5795 25675 5837
rect 411 5306 461 5348
rect 629 5306 679 5348
rect 837 5306 887 5348
rect 3465 5358 3515 5400
rect 3673 5358 3723 5400
rect 3891 5358 3941 5400
rect 14413 5570 14463 5612
rect 14631 5570 14681 5612
rect 14839 5570 14889 5612
rect 15772 5580 15822 5622
rect 15980 5580 16030 5622
rect 16198 5580 16248 5622
rect 29576 5807 29626 5849
rect 29784 5807 29834 5849
rect 30002 5807 30052 5849
rect 4775 5319 4825 5361
rect 4993 5319 5043 5361
rect 5201 5319 5251 5361
rect 7829 5371 7879 5413
rect 8037 5371 8087 5413
rect 8255 5371 8305 5413
rect 18679 5544 18729 5586
rect 18897 5544 18947 5586
rect 19105 5544 19155 5586
rect 20038 5554 20088 5596
rect 20246 5554 20296 5596
rect 20464 5554 20514 5596
rect 33940 5820 33990 5862
rect 34148 5820 34198 5862
rect 34366 5820 34416 5862
rect 9152 5331 9202 5373
rect 9370 5331 9420 5373
rect 9578 5331 9628 5373
rect 12206 5383 12256 5425
rect 12414 5383 12464 5425
rect 12632 5383 12682 5425
rect 1209 5122 1259 5164
rect 1427 5122 1477 5164
rect 1635 5122 1685 5164
rect 2363 5136 2413 5178
rect 2571 5136 2621 5178
rect 2789 5136 2839 5178
rect 13516 5344 13566 5386
rect 13734 5344 13784 5386
rect 13942 5344 13992 5386
rect 16570 5396 16620 5438
rect 16778 5396 16828 5438
rect 16996 5396 17046 5438
rect 23043 5557 23093 5599
rect 23261 5557 23311 5599
rect 23469 5557 23519 5599
rect 24402 5567 24452 5609
rect 24610 5567 24660 5609
rect 24828 5567 24878 5609
rect 5573 5135 5623 5177
rect 5791 5135 5841 5177
rect 5999 5135 6049 5177
rect 6727 5149 6777 5191
rect 6935 5149 6985 5191
rect 7153 5149 7203 5191
rect 27420 5569 27470 5611
rect 27638 5569 27688 5611
rect 27846 5569 27896 5611
rect 28779 5579 28829 5621
rect 28987 5579 29037 5621
rect 29205 5579 29255 5621
rect 9950 5147 10000 5189
rect 10168 5147 10218 5189
rect 10376 5147 10426 5189
rect 11104 5161 11154 5203
rect 11312 5161 11362 5203
rect 11530 5161 11580 5203
rect 17782 5318 17832 5360
rect 18000 5318 18050 5360
rect 18208 5318 18258 5360
rect 20836 5370 20886 5412
rect 21044 5370 21094 5412
rect 21262 5370 21312 5412
rect 31784 5582 31834 5624
rect 32002 5582 32052 5624
rect 32210 5582 32260 5624
rect 33143 5592 33193 5634
rect 33351 5592 33401 5634
rect 33569 5592 33619 5634
rect 22146 5331 22196 5373
rect 22364 5331 22414 5373
rect 22572 5331 22622 5373
rect 25200 5383 25250 5425
rect 25408 5383 25458 5425
rect 25626 5383 25676 5425
rect 412 4894 462 4936
rect 630 4894 680 4936
rect 838 4894 888 4936
rect 14314 5160 14364 5202
rect 14532 5160 14582 5202
rect 14740 5160 14790 5202
rect 15468 5174 15518 5216
rect 15676 5174 15726 5216
rect 15894 5174 15944 5216
rect 4776 4907 4826 4949
rect 4994 4907 5044 4949
rect 5202 4907 5252 4949
rect 26523 5343 26573 5385
rect 26741 5343 26791 5385
rect 26949 5343 26999 5385
rect 29577 5395 29627 5437
rect 29785 5395 29835 5437
rect 30003 5395 30053 5437
rect 18580 5134 18630 5176
rect 18798 5134 18848 5176
rect 19006 5134 19056 5176
rect 19734 5148 19784 5190
rect 19942 5148 19992 5190
rect 20160 5148 20210 5190
rect 30887 5356 30937 5398
rect 31105 5356 31155 5398
rect 31313 5356 31363 5398
rect 33941 5408 33991 5450
rect 34149 5408 34199 5450
rect 34367 5408 34417 5450
rect 9153 4919 9203 4961
rect 9371 4919 9421 4961
rect 9579 4919 9629 4961
rect 22944 5147 22994 5189
rect 23162 5147 23212 5189
rect 23370 5147 23420 5189
rect 24098 5161 24148 5203
rect 24306 5161 24356 5203
rect 24524 5161 24574 5203
rect 13517 4932 13567 4974
rect 13735 4932 13785 4974
rect 13943 4932 13993 4974
rect 27321 5159 27371 5201
rect 27539 5159 27589 5201
rect 27747 5159 27797 5201
rect 28475 5173 28525 5215
rect 28683 5173 28733 5215
rect 28901 5173 28951 5215
rect 17783 4906 17833 4948
rect 18001 4906 18051 4948
rect 18209 4906 18259 4948
rect 31685 5172 31735 5214
rect 31903 5172 31953 5214
rect 32111 5172 32161 5214
rect 32839 5186 32889 5228
rect 33047 5186 33097 5228
rect 33265 5186 33315 5228
rect 22147 4919 22197 4961
rect 22365 4919 22415 4961
rect 22573 4919 22623 4961
rect 26524 4931 26574 4973
rect 26742 4931 26792 4973
rect 26950 4931 27000 4973
rect 30888 4944 30938 4986
rect 31106 4944 31156 4986
rect 31314 4944 31364 4986
rect 3445 4752 3495 4794
rect 3653 4752 3703 4794
rect 3871 4752 3921 4794
rect 7809 4765 7859 4807
rect 8017 4765 8067 4807
rect 8235 4765 8285 4807
rect 12186 4777 12236 4819
rect 12394 4777 12444 4819
rect 12612 4777 12662 4819
rect 1494 4510 1544 4552
rect 1712 4510 1762 4552
rect 1920 4510 1970 4552
rect 2648 4524 2698 4566
rect 2856 4524 2906 4566
rect 3074 4524 3124 4566
rect 16550 4790 16600 4832
rect 16758 4790 16808 4832
rect 16976 4790 17026 4832
rect 5858 4523 5908 4565
rect 6076 4523 6126 4565
rect 6284 4523 6334 4565
rect 7012 4537 7062 4579
rect 7220 4537 7270 4579
rect 7438 4537 7488 4579
rect 20816 4764 20866 4806
rect 21024 4764 21074 4806
rect 21242 4764 21292 4806
rect 10235 4535 10285 4577
rect 10453 4535 10503 4577
rect 10661 4535 10711 4577
rect 11389 4549 11439 4591
rect 11597 4549 11647 4591
rect 11815 4549 11865 4591
rect 25180 4777 25230 4819
rect 25388 4777 25438 4819
rect 25606 4777 25656 4819
rect 392 4288 442 4330
rect 610 4288 660 4330
rect 818 4288 868 4330
rect 3446 4340 3496 4382
rect 3654 4340 3704 4382
rect 3872 4340 3922 4382
rect 14599 4548 14649 4590
rect 14817 4548 14867 4590
rect 15025 4548 15075 4590
rect 15753 4562 15803 4604
rect 15961 4562 16011 4604
rect 16179 4562 16229 4604
rect 4756 4301 4806 4343
rect 4974 4301 5024 4343
rect 5182 4301 5232 4343
rect 7810 4353 7860 4395
rect 8018 4353 8068 4395
rect 8236 4353 8286 4395
rect 29557 4789 29607 4831
rect 29765 4789 29815 4831
rect 29983 4789 30033 4831
rect 18865 4522 18915 4564
rect 19083 4522 19133 4564
rect 19291 4522 19341 4564
rect 20019 4536 20069 4578
rect 20227 4536 20277 4578
rect 20445 4536 20495 4578
rect 33921 4802 33971 4844
rect 34129 4802 34179 4844
rect 34347 4802 34397 4844
rect 9133 4313 9183 4355
rect 9351 4313 9401 4355
rect 9559 4313 9609 4355
rect 12187 4365 12237 4407
rect 12395 4365 12445 4407
rect 12613 4365 12663 4407
rect 1190 4104 1240 4146
rect 1408 4104 1458 4146
rect 1616 4104 1666 4146
rect 2549 4114 2599 4156
rect 2757 4114 2807 4156
rect 2975 4114 3025 4156
rect 13497 4326 13547 4368
rect 13715 4326 13765 4368
rect 13923 4326 13973 4368
rect 16551 4378 16601 4420
rect 16759 4378 16809 4420
rect 16977 4378 17027 4420
rect 23229 4535 23279 4577
rect 23447 4535 23497 4577
rect 23655 4535 23705 4577
rect 24383 4549 24433 4591
rect 24591 4549 24641 4591
rect 24809 4549 24859 4591
rect 5554 4117 5604 4159
rect 5772 4117 5822 4159
rect 5980 4117 6030 4159
rect 6913 4127 6963 4169
rect 7121 4127 7171 4169
rect 7339 4127 7389 4169
rect 27606 4547 27656 4589
rect 27824 4547 27874 4589
rect 28032 4547 28082 4589
rect 28760 4561 28810 4603
rect 28968 4561 29018 4603
rect 29186 4561 29236 4603
rect 9931 4129 9981 4171
rect 10149 4129 10199 4171
rect 10357 4129 10407 4171
rect 11290 4139 11340 4181
rect 11498 4139 11548 4181
rect 11716 4139 11766 4181
rect 17763 4300 17813 4342
rect 17981 4300 18031 4342
rect 18189 4300 18239 4342
rect 20817 4352 20867 4394
rect 21025 4352 21075 4394
rect 21243 4352 21293 4394
rect 31970 4560 32020 4602
rect 32188 4560 32238 4602
rect 32396 4560 32446 4602
rect 33124 4574 33174 4616
rect 33332 4574 33382 4616
rect 33550 4574 33600 4616
rect 22127 4313 22177 4355
rect 22345 4313 22395 4355
rect 22553 4313 22603 4355
rect 25181 4365 25231 4407
rect 25389 4365 25439 4407
rect 25607 4365 25657 4407
rect 393 3876 443 3918
rect 611 3876 661 3918
rect 819 3876 869 3918
rect 14295 4142 14345 4184
rect 14513 4142 14563 4184
rect 14721 4142 14771 4184
rect 15654 4152 15704 4194
rect 15862 4152 15912 4194
rect 16080 4152 16130 4194
rect 26504 4325 26554 4367
rect 26722 4325 26772 4367
rect 26930 4325 26980 4367
rect 29558 4377 29608 4419
rect 29766 4377 29816 4419
rect 29984 4377 30034 4419
rect 4757 3889 4807 3931
rect 4975 3889 5025 3931
rect 5183 3889 5233 3931
rect 18561 4116 18611 4158
rect 18779 4116 18829 4158
rect 18987 4116 19037 4158
rect 19920 4126 19970 4168
rect 20128 4126 20178 4168
rect 20346 4126 20396 4168
rect 30868 4338 30918 4380
rect 31086 4338 31136 4380
rect 31294 4338 31344 4380
rect 33922 4390 33972 4432
rect 34130 4390 34180 4432
rect 34348 4390 34398 4432
rect 9134 3901 9184 3943
rect 9352 3901 9402 3943
rect 9560 3901 9610 3943
rect 22925 4129 22975 4171
rect 23143 4129 23193 4171
rect 23351 4129 23401 4171
rect 24284 4139 24334 4181
rect 24492 4139 24542 4181
rect 24710 4139 24760 4181
rect 13498 3914 13548 3956
rect 13716 3914 13766 3956
rect 13924 3914 13974 3956
rect 27302 4141 27352 4183
rect 27520 4141 27570 4183
rect 27728 4141 27778 4183
rect 28661 4151 28711 4193
rect 28869 4151 28919 4193
rect 29087 4151 29137 4193
rect 17764 3888 17814 3930
rect 17982 3888 18032 3930
rect 18190 3888 18240 3930
rect 31666 4154 31716 4196
rect 31884 4154 31934 4196
rect 32092 4154 32142 4196
rect 33025 4164 33075 4206
rect 33233 4164 33283 4206
rect 33451 4164 33501 4206
rect 22128 3901 22178 3943
rect 22346 3901 22396 3943
rect 22554 3901 22604 3943
rect 26505 3913 26555 3955
rect 26723 3913 26773 3955
rect 26931 3913 26981 3955
rect 30869 3926 30919 3968
rect 31087 3926 31137 3968
rect 31295 3926 31345 3968
rect 3428 3734 3478 3776
rect 3636 3734 3686 3776
rect 3854 3734 3904 3776
rect 7792 3747 7842 3789
rect 8000 3747 8050 3789
rect 8218 3747 8268 3789
rect 12169 3759 12219 3801
rect 12377 3759 12427 3801
rect 12595 3759 12645 3801
rect 1272 3496 1322 3538
rect 1490 3496 1540 3538
rect 1698 3496 1748 3538
rect 2631 3506 2681 3548
rect 2839 3506 2889 3548
rect 3057 3506 3107 3548
rect 16533 3772 16583 3814
rect 16741 3772 16791 3814
rect 16959 3772 17009 3814
rect 5636 3509 5686 3551
rect 5854 3509 5904 3551
rect 6062 3509 6112 3551
rect 6995 3519 7045 3561
rect 7203 3519 7253 3561
rect 7421 3519 7471 3561
rect 20799 3746 20849 3788
rect 21007 3746 21057 3788
rect 21225 3746 21275 3788
rect 10013 3521 10063 3563
rect 10231 3521 10281 3563
rect 10439 3521 10489 3563
rect 11372 3531 11422 3573
rect 11580 3531 11630 3573
rect 11798 3531 11848 3573
rect 25163 3759 25213 3801
rect 25371 3759 25421 3801
rect 25589 3759 25639 3801
rect 375 3270 425 3312
rect 593 3270 643 3312
rect 801 3270 851 3312
rect 3429 3322 3479 3364
rect 3637 3322 3687 3364
rect 3855 3322 3905 3364
rect 14377 3534 14427 3576
rect 14595 3534 14645 3576
rect 14803 3534 14853 3576
rect 15736 3544 15786 3586
rect 15944 3544 15994 3586
rect 16162 3544 16212 3586
rect 29540 3771 29590 3813
rect 29748 3771 29798 3813
rect 29966 3771 30016 3813
rect 4739 3283 4789 3325
rect 4957 3283 5007 3325
rect 5165 3283 5215 3325
rect 7793 3335 7843 3377
rect 8001 3335 8051 3377
rect 8219 3335 8269 3377
rect 18643 3508 18693 3550
rect 18861 3508 18911 3550
rect 19069 3508 19119 3550
rect 20002 3518 20052 3560
rect 20210 3518 20260 3560
rect 20428 3518 20478 3560
rect 33904 3784 33954 3826
rect 34112 3784 34162 3826
rect 34330 3784 34380 3826
rect 9116 3295 9166 3337
rect 9334 3295 9384 3337
rect 9542 3295 9592 3337
rect 12170 3347 12220 3389
rect 12378 3347 12428 3389
rect 12596 3347 12646 3389
rect 1173 3086 1223 3128
rect 1391 3086 1441 3128
rect 1599 3086 1649 3128
rect 2466 3098 2516 3140
rect 2674 3098 2724 3140
rect 2892 3098 2942 3140
rect 13480 3308 13530 3350
rect 13698 3308 13748 3350
rect 13906 3308 13956 3350
rect 16534 3360 16584 3402
rect 16742 3360 16792 3402
rect 16960 3360 17010 3402
rect 23007 3521 23057 3563
rect 23225 3521 23275 3563
rect 23433 3521 23483 3563
rect 24366 3531 24416 3573
rect 24574 3531 24624 3573
rect 24792 3531 24842 3573
rect 5537 3099 5587 3141
rect 5755 3099 5805 3141
rect 5963 3099 6013 3141
rect 6830 3111 6880 3153
rect 7038 3111 7088 3153
rect 7256 3111 7306 3153
rect 27384 3533 27434 3575
rect 27602 3533 27652 3575
rect 27810 3533 27860 3575
rect 28743 3543 28793 3585
rect 28951 3543 29001 3585
rect 29169 3543 29219 3585
rect 9914 3111 9964 3153
rect 10132 3111 10182 3153
rect 10340 3111 10390 3153
rect 11207 3123 11257 3165
rect 11415 3123 11465 3165
rect 11633 3123 11683 3165
rect 17746 3282 17796 3324
rect 17964 3282 18014 3324
rect 18172 3282 18222 3324
rect 20800 3334 20850 3376
rect 21008 3334 21058 3376
rect 21226 3334 21276 3376
rect 31748 3546 31798 3588
rect 31966 3546 32016 3588
rect 32174 3546 32224 3588
rect 33107 3556 33157 3598
rect 33315 3556 33365 3598
rect 33533 3556 33583 3598
rect 22110 3295 22160 3337
rect 22328 3295 22378 3337
rect 22536 3295 22586 3337
rect 25164 3347 25214 3389
rect 25372 3347 25422 3389
rect 25590 3347 25640 3389
rect 376 2858 426 2900
rect 594 2858 644 2900
rect 802 2858 852 2900
rect 14278 3124 14328 3166
rect 14496 3124 14546 3166
rect 14704 3124 14754 3166
rect 15571 3136 15621 3178
rect 15779 3136 15829 3178
rect 15997 3136 16047 3178
rect 26487 3307 26537 3349
rect 26705 3307 26755 3349
rect 26913 3307 26963 3349
rect 29541 3359 29591 3401
rect 29749 3359 29799 3401
rect 29967 3359 30017 3401
rect 4740 2871 4790 2913
rect 4958 2871 5008 2913
rect 5166 2871 5216 2913
rect 18544 3098 18594 3140
rect 18762 3098 18812 3140
rect 18970 3098 19020 3140
rect 19837 3110 19887 3152
rect 20045 3110 20095 3152
rect 20263 3110 20313 3152
rect 30851 3320 30901 3362
rect 31069 3320 31119 3362
rect 31277 3320 31327 3362
rect 33905 3372 33955 3414
rect 34113 3372 34163 3414
rect 34331 3372 34381 3414
rect 9117 2883 9167 2925
rect 9335 2883 9385 2925
rect 9543 2883 9593 2925
rect 22908 3111 22958 3153
rect 23126 3111 23176 3153
rect 23334 3111 23384 3153
rect 24201 3123 24251 3165
rect 24409 3123 24459 3165
rect 24627 3123 24677 3165
rect 13481 2896 13531 2938
rect 13699 2896 13749 2938
rect 13907 2896 13957 2938
rect 27285 3123 27335 3165
rect 27503 3123 27553 3165
rect 27711 3123 27761 3165
rect 28578 3135 28628 3177
rect 28786 3135 28836 3177
rect 29004 3135 29054 3177
rect 17747 2870 17797 2912
rect 17965 2870 18015 2912
rect 18173 2870 18223 2912
rect 31649 3136 31699 3178
rect 31867 3136 31917 3178
rect 32075 3136 32125 3178
rect 32942 3148 32992 3190
rect 33150 3148 33200 3190
rect 33368 3148 33418 3190
rect 22111 2883 22161 2925
rect 22329 2883 22379 2925
rect 22537 2883 22587 2925
rect 26488 2895 26538 2937
rect 26706 2895 26756 2937
rect 26914 2895 26964 2937
rect 30852 2908 30902 2950
rect 31070 2908 31120 2950
rect 31278 2908 31328 2950
rect 3408 2716 3458 2758
rect 3616 2716 3666 2758
rect 3834 2716 3884 2758
rect 7772 2729 7822 2771
rect 7980 2729 8030 2771
rect 8198 2729 8248 2771
rect 12149 2741 12199 2783
rect 12357 2741 12407 2783
rect 12575 2741 12625 2783
rect 1318 2476 1368 2518
rect 1536 2476 1586 2518
rect 1744 2476 1794 2518
rect 2611 2488 2661 2530
rect 2819 2488 2869 2530
rect 3037 2488 3087 2530
rect 16513 2754 16563 2796
rect 16721 2754 16771 2796
rect 16939 2754 16989 2796
rect 5682 2489 5732 2531
rect 5900 2489 5950 2531
rect 6108 2489 6158 2531
rect 6975 2501 7025 2543
rect 7183 2501 7233 2543
rect 7401 2501 7451 2543
rect 20779 2728 20829 2770
rect 20987 2728 21037 2770
rect 21205 2728 21255 2770
rect 10059 2501 10109 2543
rect 10277 2501 10327 2543
rect 10485 2501 10535 2543
rect 11352 2513 11402 2555
rect 11560 2513 11610 2555
rect 11778 2513 11828 2555
rect 25143 2741 25193 2783
rect 25351 2741 25401 2783
rect 25569 2741 25619 2783
rect 355 2252 405 2294
rect 573 2252 623 2294
rect 781 2252 831 2294
rect 3409 2304 3459 2346
rect 3617 2304 3667 2346
rect 3835 2304 3885 2346
rect 14423 2514 14473 2556
rect 14641 2514 14691 2556
rect 14849 2514 14899 2556
rect 15716 2526 15766 2568
rect 15924 2526 15974 2568
rect 16142 2526 16192 2568
rect 29520 2753 29570 2795
rect 29728 2753 29778 2795
rect 29946 2753 29996 2795
rect 4719 2265 4769 2307
rect 4937 2265 4987 2307
rect 5145 2265 5195 2307
rect 7773 2317 7823 2359
rect 7981 2317 8031 2359
rect 8199 2317 8249 2359
rect 18689 2488 18739 2530
rect 18907 2488 18957 2530
rect 19115 2488 19165 2530
rect 19982 2500 20032 2542
rect 20190 2500 20240 2542
rect 20408 2500 20458 2542
rect 33884 2766 33934 2808
rect 34092 2766 34142 2808
rect 34310 2766 34360 2808
rect 9096 2277 9146 2319
rect 9314 2277 9364 2319
rect 9522 2277 9572 2319
rect 12150 2329 12200 2371
rect 12358 2329 12408 2371
rect 12576 2329 12626 2371
rect 1153 2068 1203 2110
rect 1371 2068 1421 2110
rect 1579 2068 1629 2110
rect 2512 2078 2562 2120
rect 2720 2078 2770 2120
rect 2938 2078 2988 2120
rect 13460 2290 13510 2332
rect 13678 2290 13728 2332
rect 13886 2290 13936 2332
rect 16514 2342 16564 2384
rect 16722 2342 16772 2384
rect 16940 2342 16990 2384
rect 23053 2501 23103 2543
rect 23271 2501 23321 2543
rect 23479 2501 23529 2543
rect 24346 2513 24396 2555
rect 24554 2513 24604 2555
rect 24772 2513 24822 2555
rect 5517 2081 5567 2123
rect 5735 2081 5785 2123
rect 5943 2081 5993 2123
rect 6876 2091 6926 2133
rect 7084 2091 7134 2133
rect 7302 2091 7352 2133
rect 27430 2513 27480 2555
rect 27648 2513 27698 2555
rect 27856 2513 27906 2555
rect 28723 2525 28773 2567
rect 28931 2525 28981 2567
rect 29149 2525 29199 2567
rect 9894 2093 9944 2135
rect 10112 2093 10162 2135
rect 10320 2093 10370 2135
rect 11253 2103 11303 2145
rect 11461 2103 11511 2145
rect 11679 2103 11729 2145
rect 17726 2264 17776 2306
rect 17944 2264 17994 2306
rect 18152 2264 18202 2306
rect 20780 2316 20830 2358
rect 20988 2316 21038 2358
rect 21206 2316 21256 2358
rect 31794 2526 31844 2568
rect 32012 2526 32062 2568
rect 32220 2526 32270 2568
rect 33087 2538 33137 2580
rect 33295 2538 33345 2580
rect 33513 2538 33563 2580
rect 22090 2277 22140 2319
rect 22308 2277 22358 2319
rect 22516 2277 22566 2319
rect 25144 2329 25194 2371
rect 25352 2329 25402 2371
rect 25570 2329 25620 2371
rect 356 1840 406 1882
rect 574 1840 624 1882
rect 782 1840 832 1882
rect 14258 2106 14308 2148
rect 14476 2106 14526 2148
rect 14684 2106 14734 2148
rect 15617 2116 15667 2158
rect 15825 2116 15875 2158
rect 16043 2116 16093 2158
rect 26467 2289 26517 2331
rect 26685 2289 26735 2331
rect 26893 2289 26943 2331
rect 29521 2341 29571 2383
rect 29729 2341 29779 2383
rect 29947 2341 29997 2383
rect 4720 1853 4770 1895
rect 4938 1853 4988 1895
rect 5146 1853 5196 1895
rect 18524 2080 18574 2122
rect 18742 2080 18792 2122
rect 18950 2080 19000 2122
rect 19883 2090 19933 2132
rect 20091 2090 20141 2132
rect 20309 2090 20359 2132
rect 30831 2302 30881 2344
rect 31049 2302 31099 2344
rect 31257 2302 31307 2344
rect 33885 2354 33935 2396
rect 34093 2354 34143 2396
rect 34311 2354 34361 2396
rect 9097 1865 9147 1907
rect 9315 1865 9365 1907
rect 9523 1865 9573 1907
rect 22888 2093 22938 2135
rect 23106 2093 23156 2135
rect 23314 2093 23364 2135
rect 24247 2103 24297 2145
rect 24455 2103 24505 2145
rect 24673 2103 24723 2145
rect 13461 1878 13511 1920
rect 13679 1878 13729 1920
rect 13887 1878 13937 1920
rect 27265 2105 27315 2147
rect 27483 2105 27533 2147
rect 27691 2105 27741 2147
rect 28624 2115 28674 2157
rect 28832 2115 28882 2157
rect 29050 2115 29100 2157
rect 17727 1852 17777 1894
rect 17945 1852 17995 1894
rect 18153 1852 18203 1894
rect 31629 2118 31679 2160
rect 31847 2118 31897 2160
rect 32055 2118 32105 2160
rect 32988 2128 33038 2170
rect 33196 2128 33246 2170
rect 33414 2128 33464 2170
rect 22091 1865 22141 1907
rect 22309 1865 22359 1907
rect 22517 1865 22567 1907
rect 26468 1877 26518 1919
rect 26686 1877 26736 1919
rect 26894 1877 26944 1919
rect 30832 1890 30882 1932
rect 31050 1890 31100 1932
rect 31258 1890 31308 1932
rect 3391 1698 3441 1740
rect 3599 1698 3649 1740
rect 3817 1698 3867 1740
rect 7755 1711 7805 1753
rect 7963 1711 8013 1753
rect 8181 1711 8231 1753
rect 12132 1723 12182 1765
rect 12340 1723 12390 1765
rect 12558 1723 12608 1765
rect 1235 1460 1285 1502
rect 1453 1460 1503 1502
rect 1661 1460 1711 1502
rect 2594 1470 2644 1512
rect 2802 1470 2852 1512
rect 3020 1470 3070 1512
rect 16496 1736 16546 1778
rect 16704 1736 16754 1778
rect 16922 1736 16972 1778
rect 5599 1473 5649 1515
rect 5817 1473 5867 1515
rect 6025 1473 6075 1515
rect 6958 1483 7008 1525
rect 7166 1483 7216 1525
rect 7384 1483 7434 1525
rect 20762 1710 20812 1752
rect 20970 1710 21020 1752
rect 21188 1710 21238 1752
rect 9976 1485 10026 1527
rect 10194 1485 10244 1527
rect 10402 1485 10452 1527
rect 11335 1495 11385 1537
rect 11543 1495 11593 1537
rect 11761 1495 11811 1537
rect 25126 1723 25176 1765
rect 25334 1723 25384 1765
rect 25552 1723 25602 1765
rect 338 1234 388 1276
rect 556 1234 606 1276
rect 764 1234 814 1276
rect 3392 1286 3442 1328
rect 3600 1286 3650 1328
rect 3818 1286 3868 1328
rect 14340 1498 14390 1540
rect 14558 1498 14608 1540
rect 14766 1498 14816 1540
rect 15699 1508 15749 1550
rect 15907 1508 15957 1550
rect 16125 1508 16175 1550
rect 29503 1735 29553 1777
rect 29711 1735 29761 1777
rect 29929 1735 29979 1777
rect 4702 1247 4752 1289
rect 4920 1247 4970 1289
rect 5128 1247 5178 1289
rect 7756 1299 7806 1341
rect 7964 1299 8014 1341
rect 8182 1299 8232 1341
rect 18606 1472 18656 1514
rect 18824 1472 18874 1514
rect 19032 1472 19082 1514
rect 19965 1482 20015 1524
rect 20173 1482 20223 1524
rect 20391 1482 20441 1524
rect 33867 1748 33917 1790
rect 34075 1748 34125 1790
rect 34293 1748 34343 1790
rect 9079 1259 9129 1301
rect 9297 1259 9347 1301
rect 9505 1259 9555 1301
rect 12133 1311 12183 1353
rect 12341 1311 12391 1353
rect 12559 1311 12609 1353
rect 13443 1272 13493 1314
rect 13661 1272 13711 1314
rect 13869 1272 13919 1314
rect 16497 1324 16547 1366
rect 16705 1324 16755 1366
rect 16923 1324 16973 1366
rect 22970 1485 23020 1527
rect 23188 1485 23238 1527
rect 23396 1485 23446 1527
rect 24329 1495 24379 1537
rect 24537 1495 24587 1537
rect 24755 1495 24805 1537
rect 27347 1497 27397 1539
rect 27565 1497 27615 1539
rect 27773 1497 27823 1539
rect 28706 1507 28756 1549
rect 28914 1507 28964 1549
rect 29132 1507 29182 1549
rect 17709 1246 17759 1288
rect 17927 1246 17977 1288
rect 18135 1246 18185 1288
rect 20763 1298 20813 1340
rect 20971 1298 21021 1340
rect 21189 1298 21239 1340
rect 31711 1510 31761 1552
rect 31929 1510 31979 1552
rect 32137 1510 32187 1552
rect 33070 1520 33120 1562
rect 33278 1520 33328 1562
rect 33496 1520 33546 1562
rect 22073 1259 22123 1301
rect 22291 1259 22341 1301
rect 22499 1259 22549 1301
rect 25127 1311 25177 1353
rect 25335 1311 25385 1353
rect 25553 1311 25603 1353
rect 1136 1050 1186 1092
rect 1354 1050 1404 1092
rect 1562 1050 1612 1092
rect 5500 1063 5550 1105
rect 5718 1063 5768 1105
rect 5926 1063 5976 1105
rect 9877 1075 9927 1117
rect 10095 1075 10145 1117
rect 10303 1075 10353 1117
rect 339 822 389 864
rect 557 822 607 864
rect 765 822 815 864
rect 14241 1088 14291 1130
rect 14459 1088 14509 1130
rect 14667 1088 14717 1130
rect 26450 1271 26500 1313
rect 26668 1271 26718 1313
rect 26876 1271 26926 1313
rect 29504 1323 29554 1365
rect 29712 1323 29762 1365
rect 29930 1323 29980 1365
rect 30814 1284 30864 1326
rect 31032 1284 31082 1326
rect 31240 1284 31290 1326
rect 33868 1336 33918 1378
rect 34076 1336 34126 1378
rect 34294 1336 34344 1378
rect 4703 835 4753 877
rect 4921 835 4971 877
rect 5129 835 5179 877
rect 18507 1062 18557 1104
rect 18725 1062 18775 1104
rect 18933 1062 18983 1104
rect 9080 847 9130 889
rect 9298 847 9348 889
rect 9506 847 9556 889
rect 22871 1075 22921 1117
rect 23089 1075 23139 1117
rect 23297 1075 23347 1117
rect 13444 860 13494 902
rect 13662 860 13712 902
rect 13870 860 13920 902
rect 27248 1087 27298 1129
rect 27466 1087 27516 1129
rect 27674 1087 27724 1129
rect 17710 834 17760 876
rect 17928 834 17978 876
rect 18136 834 18186 876
rect 31612 1100 31662 1142
rect 31830 1100 31880 1142
rect 32038 1100 32088 1142
rect 22074 847 22124 889
rect 22292 847 22342 889
rect 22500 847 22550 889
rect 26451 859 26501 901
rect 26669 859 26719 901
rect 26877 859 26927 901
rect 30815 872 30865 914
rect 31033 872 31083 914
rect 31241 872 31291 914
rect 1552 246 1602 288
rect 1770 246 1820 288
rect 1978 246 2028 288
rect 5916 259 5966 301
rect 6134 259 6184 301
rect 6342 259 6392 301
rect 10293 271 10343 313
rect 10511 271 10561 313
rect 10719 271 10769 313
rect 14657 284 14707 326
rect 14875 284 14925 326
rect 15083 284 15133 326
rect 18923 258 18973 300
rect 19141 258 19191 300
rect 19349 258 19399 300
rect 4041 172 4091 214
rect 4259 172 4309 214
rect 4467 172 4517 214
rect 8489 196 8539 238
rect 8707 196 8757 238
rect 8915 196 8965 238
rect 12782 197 12832 239
rect 13000 197 13050 239
rect 13208 197 13258 239
rect 23287 271 23337 313
rect 23505 271 23555 313
rect 23713 271 23763 313
rect 27664 283 27714 325
rect 27882 283 27932 325
rect 28090 283 28140 325
rect 32028 296 32078 338
rect 32246 296 32296 338
rect 32454 296 32504 338
rect 21412 184 21462 226
rect 21630 184 21680 226
rect 21838 184 21888 226
rect 25860 208 25910 250
rect 26078 208 26128 250
rect 26286 208 26336 250
rect 30153 209 30203 251
rect 30371 209 30421 251
rect 30579 209 30629 251
rect 16979 133 17029 175
rect 17197 133 17247 175
rect 17405 133 17455 175
<< pmos >>
rect 3518 8647 3568 8747
rect 3726 8647 3776 8747
rect 3944 8647 3994 8747
rect 7882 8660 7932 8760
rect 8090 8660 8140 8760
rect 8308 8660 8358 8760
rect 12259 8672 12309 8772
rect 12467 8672 12517 8772
rect 12685 8672 12735 8772
rect 16623 8685 16673 8785
rect 16831 8685 16881 8785
rect 17049 8685 17099 8785
rect 20889 8659 20939 8759
rect 21097 8659 21147 8759
rect 21315 8659 21365 8759
rect 465 8479 515 8579
rect 683 8479 733 8579
rect 891 8479 941 8579
rect 2721 8419 2771 8519
rect 2929 8419 2979 8519
rect 3147 8419 3197 8519
rect 4829 8492 4879 8592
rect 5047 8492 5097 8592
rect 5255 8492 5305 8592
rect 1263 8295 1313 8395
rect 1481 8295 1531 8395
rect 1689 8295 1739 8395
rect 7085 8432 7135 8532
rect 7293 8432 7343 8532
rect 7511 8432 7561 8532
rect 9206 8504 9256 8604
rect 9424 8504 9474 8604
rect 9632 8504 9682 8604
rect 3519 8235 3569 8335
rect 3727 8235 3777 8335
rect 3945 8235 3995 8335
rect 5627 8308 5677 8408
rect 5845 8308 5895 8408
rect 6053 8308 6103 8408
rect 11462 8444 11512 8544
rect 11670 8444 11720 8544
rect 11888 8444 11938 8544
rect 13570 8517 13620 8617
rect 13788 8517 13838 8617
rect 13996 8517 14046 8617
rect 25253 8672 25303 8772
rect 25461 8672 25511 8772
rect 25679 8672 25729 8772
rect 29630 8684 29680 8784
rect 29838 8684 29888 8784
rect 30056 8684 30106 8784
rect 33994 8697 34044 8797
rect 34202 8697 34252 8797
rect 34420 8697 34470 8797
rect 7883 8248 7933 8348
rect 8091 8248 8141 8348
rect 8309 8248 8359 8348
rect 10004 8320 10054 8420
rect 10222 8320 10272 8420
rect 10430 8320 10480 8420
rect 15826 8457 15876 8557
rect 16034 8457 16084 8557
rect 16252 8457 16302 8557
rect 17836 8491 17886 8591
rect 18054 8491 18104 8591
rect 18262 8491 18312 8591
rect 466 8067 516 8167
rect 684 8067 734 8167
rect 892 8067 942 8167
rect 12260 8260 12310 8360
rect 12468 8260 12518 8360
rect 12686 8260 12736 8360
rect 14368 8333 14418 8433
rect 14586 8333 14636 8433
rect 14794 8333 14844 8433
rect 20092 8431 20142 8531
rect 20300 8431 20350 8531
rect 20518 8431 20568 8531
rect 22200 8504 22250 8604
rect 22418 8504 22468 8604
rect 22626 8504 22676 8604
rect 2622 8009 2672 8109
rect 2830 8009 2880 8109
rect 3048 8009 3098 8109
rect 4830 8080 4880 8180
rect 5048 8080 5098 8180
rect 5256 8080 5306 8180
rect 16624 8273 16674 8373
rect 16832 8273 16882 8373
rect 17050 8273 17100 8373
rect 18634 8307 18684 8407
rect 18852 8307 18902 8407
rect 19060 8307 19110 8407
rect 24456 8444 24506 8544
rect 24664 8444 24714 8544
rect 24882 8444 24932 8544
rect 26577 8516 26627 8616
rect 26795 8516 26845 8616
rect 27003 8516 27053 8616
rect 6986 8022 7036 8122
rect 7194 8022 7244 8122
rect 7412 8022 7462 8122
rect 9207 8092 9257 8192
rect 9425 8092 9475 8192
rect 9633 8092 9683 8192
rect 20890 8247 20940 8347
rect 21098 8247 21148 8347
rect 21316 8247 21366 8347
rect 22998 8320 23048 8420
rect 23216 8320 23266 8420
rect 23424 8320 23474 8420
rect 28833 8456 28883 8556
rect 29041 8456 29091 8556
rect 29259 8456 29309 8556
rect 30941 8529 30991 8629
rect 31159 8529 31209 8629
rect 31367 8529 31417 8629
rect 11363 8034 11413 8134
rect 11571 8034 11621 8134
rect 11789 8034 11839 8134
rect 13571 8105 13621 8205
rect 13789 8105 13839 8205
rect 13997 8105 14047 8205
rect 25254 8260 25304 8360
rect 25462 8260 25512 8360
rect 25680 8260 25730 8360
rect 27375 8332 27425 8432
rect 27593 8332 27643 8432
rect 27801 8332 27851 8432
rect 33197 8469 33247 8569
rect 33405 8469 33455 8569
rect 33623 8469 33673 8569
rect 15727 8047 15777 8147
rect 15935 8047 15985 8147
rect 16153 8047 16203 8147
rect 17837 8079 17887 8179
rect 18055 8079 18105 8179
rect 18263 8079 18313 8179
rect 29631 8272 29681 8372
rect 29839 8272 29889 8372
rect 30057 8272 30107 8372
rect 31739 8345 31789 8445
rect 31957 8345 32007 8445
rect 32165 8345 32215 8445
rect 19993 8021 20043 8121
rect 20201 8021 20251 8121
rect 20419 8021 20469 8121
rect 22201 8092 22251 8192
rect 22419 8092 22469 8192
rect 22627 8092 22677 8192
rect 33995 8285 34045 8385
rect 34203 8285 34253 8385
rect 34421 8285 34471 8385
rect 24357 8034 24407 8134
rect 24565 8034 24615 8134
rect 24783 8034 24833 8134
rect 26578 8104 26628 8204
rect 26796 8104 26846 8204
rect 27004 8104 27054 8204
rect 28734 8046 28784 8146
rect 28942 8046 28992 8146
rect 29160 8046 29210 8146
rect 30942 8117 30992 8217
rect 31160 8117 31210 8217
rect 31368 8117 31418 8217
rect 33098 8059 33148 8159
rect 33306 8059 33356 8159
rect 33524 8059 33574 8159
rect 1345 7687 1395 7787
rect 1563 7687 1613 7787
rect 1771 7687 1821 7787
rect 3501 7629 3551 7729
rect 3709 7629 3759 7729
rect 3927 7629 3977 7729
rect 5709 7700 5759 7800
rect 5927 7700 5977 7800
rect 6135 7700 6185 7800
rect 7865 7642 7915 7742
rect 8073 7642 8123 7742
rect 8291 7642 8341 7742
rect 10086 7712 10136 7812
rect 10304 7712 10354 7812
rect 10512 7712 10562 7812
rect 448 7461 498 7561
rect 666 7461 716 7561
rect 874 7461 924 7561
rect 12242 7654 12292 7754
rect 12450 7654 12500 7754
rect 12668 7654 12718 7754
rect 14450 7725 14500 7825
rect 14668 7725 14718 7825
rect 14876 7725 14926 7825
rect 2704 7401 2754 7501
rect 2912 7401 2962 7501
rect 3130 7401 3180 7501
rect 4812 7474 4862 7574
rect 5030 7474 5080 7574
rect 5238 7474 5288 7574
rect 16606 7667 16656 7767
rect 16814 7667 16864 7767
rect 17032 7667 17082 7767
rect 18716 7699 18766 7799
rect 18934 7699 18984 7799
rect 19142 7699 19192 7799
rect 1246 7277 1296 7377
rect 1464 7277 1514 7377
rect 1672 7277 1722 7377
rect 7068 7414 7118 7514
rect 7276 7414 7326 7514
rect 7494 7414 7544 7514
rect 9189 7486 9239 7586
rect 9407 7486 9457 7586
rect 9615 7486 9665 7586
rect 20872 7641 20922 7741
rect 21080 7641 21130 7741
rect 21298 7641 21348 7741
rect 23080 7712 23130 7812
rect 23298 7712 23348 7812
rect 23506 7712 23556 7812
rect 3502 7217 3552 7317
rect 3710 7217 3760 7317
rect 3928 7217 3978 7317
rect 5610 7290 5660 7390
rect 5828 7290 5878 7390
rect 6036 7290 6086 7390
rect 11445 7426 11495 7526
rect 11653 7426 11703 7526
rect 11871 7426 11921 7526
rect 13553 7499 13603 7599
rect 13771 7499 13821 7599
rect 13979 7499 14029 7599
rect 25236 7654 25286 7754
rect 25444 7654 25494 7754
rect 25662 7654 25712 7754
rect 27457 7724 27507 7824
rect 27675 7724 27725 7824
rect 27883 7724 27933 7824
rect 7866 7230 7916 7330
rect 8074 7230 8124 7330
rect 8292 7230 8342 7330
rect 9987 7302 10037 7402
rect 10205 7302 10255 7402
rect 10413 7302 10463 7402
rect 15809 7439 15859 7539
rect 16017 7439 16067 7539
rect 16235 7439 16285 7539
rect 17819 7473 17869 7573
rect 18037 7473 18087 7573
rect 18245 7473 18295 7573
rect 29613 7666 29663 7766
rect 29821 7666 29871 7766
rect 30039 7666 30089 7766
rect 31821 7737 31871 7837
rect 32039 7737 32089 7837
rect 32247 7737 32297 7837
rect 449 7049 499 7149
rect 667 7049 717 7149
rect 875 7049 925 7149
rect 12243 7242 12293 7342
rect 12451 7242 12501 7342
rect 12669 7242 12719 7342
rect 14351 7315 14401 7415
rect 14569 7315 14619 7415
rect 14777 7315 14827 7415
rect 20075 7413 20125 7513
rect 20283 7413 20333 7513
rect 20501 7413 20551 7513
rect 22183 7486 22233 7586
rect 22401 7486 22451 7586
rect 22609 7486 22659 7586
rect 33977 7679 34027 7779
rect 34185 7679 34235 7779
rect 34403 7679 34453 7779
rect 2539 6993 2589 7093
rect 2747 6993 2797 7093
rect 2965 6993 3015 7093
rect 4813 7062 4863 7162
rect 5031 7062 5081 7162
rect 5239 7062 5289 7162
rect 16607 7255 16657 7355
rect 16815 7255 16865 7355
rect 17033 7255 17083 7355
rect 18617 7289 18667 7389
rect 18835 7289 18885 7389
rect 19043 7289 19093 7389
rect 24439 7426 24489 7526
rect 24647 7426 24697 7526
rect 24865 7426 24915 7526
rect 26560 7498 26610 7598
rect 26778 7498 26828 7598
rect 26986 7498 27036 7598
rect 6903 7006 6953 7106
rect 7111 7006 7161 7106
rect 7329 7006 7379 7106
rect 9190 7074 9240 7174
rect 9408 7074 9458 7174
rect 9616 7074 9666 7174
rect 20873 7229 20923 7329
rect 21081 7229 21131 7329
rect 21299 7229 21349 7329
rect 22981 7302 23031 7402
rect 23199 7302 23249 7402
rect 23407 7302 23457 7402
rect 28816 7438 28866 7538
rect 29024 7438 29074 7538
rect 29242 7438 29292 7538
rect 30924 7511 30974 7611
rect 31142 7511 31192 7611
rect 31350 7511 31400 7611
rect 11280 7018 11330 7118
rect 11488 7018 11538 7118
rect 11706 7018 11756 7118
rect 13554 7087 13604 7187
rect 13772 7087 13822 7187
rect 13980 7087 14030 7187
rect 25237 7242 25287 7342
rect 25445 7242 25495 7342
rect 25663 7242 25713 7342
rect 27358 7314 27408 7414
rect 27576 7314 27626 7414
rect 27784 7314 27834 7414
rect 33180 7451 33230 7551
rect 33388 7451 33438 7551
rect 33606 7451 33656 7551
rect 15644 7031 15694 7131
rect 15852 7031 15902 7131
rect 16070 7031 16120 7131
rect 17820 7061 17870 7161
rect 18038 7061 18088 7161
rect 18246 7061 18296 7161
rect 29614 7254 29664 7354
rect 29822 7254 29872 7354
rect 30040 7254 30090 7354
rect 31722 7327 31772 7427
rect 31940 7327 31990 7427
rect 32148 7327 32198 7427
rect 19910 7005 19960 7105
rect 20118 7005 20168 7105
rect 20336 7005 20386 7105
rect 22184 7074 22234 7174
rect 22402 7074 22452 7174
rect 22610 7074 22660 7174
rect 33978 7267 34028 7367
rect 34186 7267 34236 7367
rect 34404 7267 34454 7367
rect 24274 7018 24324 7118
rect 24482 7018 24532 7118
rect 24700 7018 24750 7118
rect 26561 7086 26611 7186
rect 26779 7086 26829 7186
rect 26987 7086 27037 7186
rect 28651 7030 28701 7130
rect 28859 7030 28909 7130
rect 29077 7030 29127 7130
rect 30925 7099 30975 7199
rect 31143 7099 31193 7199
rect 31351 7099 31401 7199
rect 33015 7043 33065 7143
rect 33223 7043 33273 7143
rect 33441 7043 33491 7143
rect 1391 6667 1441 6767
rect 1609 6667 1659 6767
rect 1817 6667 1867 6767
rect 3481 6611 3531 6711
rect 3689 6611 3739 6711
rect 3907 6611 3957 6711
rect 5755 6680 5805 6780
rect 5973 6680 6023 6780
rect 6181 6680 6231 6780
rect 7845 6624 7895 6724
rect 8053 6624 8103 6724
rect 8271 6624 8321 6724
rect 10132 6692 10182 6792
rect 10350 6692 10400 6792
rect 10558 6692 10608 6792
rect 428 6443 478 6543
rect 646 6443 696 6543
rect 854 6443 904 6543
rect 12222 6636 12272 6736
rect 12430 6636 12480 6736
rect 12648 6636 12698 6736
rect 14496 6705 14546 6805
rect 14714 6705 14764 6805
rect 14922 6705 14972 6805
rect 2684 6383 2734 6483
rect 2892 6383 2942 6483
rect 3110 6383 3160 6483
rect 4792 6456 4842 6556
rect 5010 6456 5060 6556
rect 5218 6456 5268 6556
rect 16586 6649 16636 6749
rect 16794 6649 16844 6749
rect 17012 6649 17062 6749
rect 18762 6679 18812 6779
rect 18980 6679 19030 6779
rect 19188 6679 19238 6779
rect 1226 6259 1276 6359
rect 1444 6259 1494 6359
rect 1652 6259 1702 6359
rect 7048 6396 7098 6496
rect 7256 6396 7306 6496
rect 7474 6396 7524 6496
rect 9169 6468 9219 6568
rect 9387 6468 9437 6568
rect 9595 6468 9645 6568
rect 20852 6623 20902 6723
rect 21060 6623 21110 6723
rect 21278 6623 21328 6723
rect 23126 6692 23176 6792
rect 23344 6692 23394 6792
rect 23552 6692 23602 6792
rect 3482 6199 3532 6299
rect 3690 6199 3740 6299
rect 3908 6199 3958 6299
rect 5590 6272 5640 6372
rect 5808 6272 5858 6372
rect 6016 6272 6066 6372
rect 11425 6408 11475 6508
rect 11633 6408 11683 6508
rect 11851 6408 11901 6508
rect 13533 6481 13583 6581
rect 13751 6481 13801 6581
rect 13959 6481 14009 6581
rect 25216 6636 25266 6736
rect 25424 6636 25474 6736
rect 25642 6636 25692 6736
rect 27503 6704 27553 6804
rect 27721 6704 27771 6804
rect 27929 6704 27979 6804
rect 7846 6212 7896 6312
rect 8054 6212 8104 6312
rect 8272 6212 8322 6312
rect 9967 6284 10017 6384
rect 10185 6284 10235 6384
rect 10393 6284 10443 6384
rect 15789 6421 15839 6521
rect 15997 6421 16047 6521
rect 16215 6421 16265 6521
rect 17799 6455 17849 6555
rect 18017 6455 18067 6555
rect 18225 6455 18275 6555
rect 29593 6648 29643 6748
rect 29801 6648 29851 6748
rect 30019 6648 30069 6748
rect 31867 6717 31917 6817
rect 32085 6717 32135 6817
rect 32293 6717 32343 6817
rect 429 6031 479 6131
rect 647 6031 697 6131
rect 855 6031 905 6131
rect 12223 6224 12273 6324
rect 12431 6224 12481 6324
rect 12649 6224 12699 6324
rect 14331 6297 14381 6397
rect 14549 6297 14599 6397
rect 14757 6297 14807 6397
rect 20055 6395 20105 6495
rect 20263 6395 20313 6495
rect 20481 6395 20531 6495
rect 22163 6468 22213 6568
rect 22381 6468 22431 6568
rect 22589 6468 22639 6568
rect 33957 6661 34007 6761
rect 34165 6661 34215 6761
rect 34383 6661 34433 6761
rect 2585 5973 2635 6073
rect 2793 5973 2843 6073
rect 3011 5973 3061 6073
rect 4793 6044 4843 6144
rect 5011 6044 5061 6144
rect 5219 6044 5269 6144
rect 16587 6237 16637 6337
rect 16795 6237 16845 6337
rect 17013 6237 17063 6337
rect 18597 6271 18647 6371
rect 18815 6271 18865 6371
rect 19023 6271 19073 6371
rect 24419 6408 24469 6508
rect 24627 6408 24677 6508
rect 24845 6408 24895 6508
rect 26540 6480 26590 6580
rect 26758 6480 26808 6580
rect 26966 6480 27016 6580
rect 6949 5986 6999 6086
rect 7157 5986 7207 6086
rect 7375 5986 7425 6086
rect 9170 6056 9220 6156
rect 9388 6056 9438 6156
rect 9596 6056 9646 6156
rect 20853 6211 20903 6311
rect 21061 6211 21111 6311
rect 21279 6211 21329 6311
rect 22961 6284 23011 6384
rect 23179 6284 23229 6384
rect 23387 6284 23437 6384
rect 28796 6420 28846 6520
rect 29004 6420 29054 6520
rect 29222 6420 29272 6520
rect 30904 6493 30954 6593
rect 31122 6493 31172 6593
rect 31330 6493 31380 6593
rect 11326 5998 11376 6098
rect 11534 5998 11584 6098
rect 11752 5998 11802 6098
rect 13534 6069 13584 6169
rect 13752 6069 13802 6169
rect 13960 6069 14010 6169
rect 25217 6224 25267 6324
rect 25425 6224 25475 6324
rect 25643 6224 25693 6324
rect 27338 6296 27388 6396
rect 27556 6296 27606 6396
rect 27764 6296 27814 6396
rect 33160 6433 33210 6533
rect 33368 6433 33418 6533
rect 33586 6433 33636 6533
rect 15690 6011 15740 6111
rect 15898 6011 15948 6111
rect 16116 6011 16166 6111
rect 17800 6043 17850 6143
rect 18018 6043 18068 6143
rect 18226 6043 18276 6143
rect 29594 6236 29644 6336
rect 29802 6236 29852 6336
rect 30020 6236 30070 6336
rect 31702 6309 31752 6409
rect 31920 6309 31970 6409
rect 32128 6309 32178 6409
rect 19956 5985 20006 6085
rect 20164 5985 20214 6085
rect 20382 5985 20432 6085
rect 22164 6056 22214 6156
rect 22382 6056 22432 6156
rect 22590 6056 22640 6156
rect 33958 6249 34008 6349
rect 34166 6249 34216 6349
rect 34384 6249 34434 6349
rect 24320 5998 24370 6098
rect 24528 5998 24578 6098
rect 24746 5998 24796 6098
rect 26541 6068 26591 6168
rect 26759 6068 26809 6168
rect 26967 6068 27017 6168
rect 28697 6010 28747 6110
rect 28905 6010 28955 6110
rect 29123 6010 29173 6110
rect 30905 6081 30955 6181
rect 31123 6081 31173 6181
rect 31331 6081 31381 6181
rect 33061 6023 33111 6123
rect 33269 6023 33319 6123
rect 33487 6023 33537 6123
rect 1308 5651 1358 5751
rect 1526 5651 1576 5751
rect 1734 5651 1784 5751
rect 3464 5593 3514 5693
rect 3672 5593 3722 5693
rect 3890 5593 3940 5693
rect 5672 5664 5722 5764
rect 5890 5664 5940 5764
rect 6098 5664 6148 5764
rect 7828 5606 7878 5706
rect 8036 5606 8086 5706
rect 8254 5606 8304 5706
rect 10049 5676 10099 5776
rect 10267 5676 10317 5776
rect 10475 5676 10525 5776
rect 411 5425 461 5525
rect 629 5425 679 5525
rect 837 5425 887 5525
rect 12205 5618 12255 5718
rect 12413 5618 12463 5718
rect 12631 5618 12681 5718
rect 14413 5689 14463 5789
rect 14631 5689 14681 5789
rect 14839 5689 14889 5789
rect 2667 5365 2717 5465
rect 2875 5365 2925 5465
rect 3093 5365 3143 5465
rect 4775 5438 4825 5538
rect 4993 5438 5043 5538
rect 5201 5438 5251 5538
rect 16569 5631 16619 5731
rect 16777 5631 16827 5731
rect 16995 5631 17045 5731
rect 18679 5663 18729 5763
rect 18897 5663 18947 5763
rect 19105 5663 19155 5763
rect 1209 5241 1259 5341
rect 1427 5241 1477 5341
rect 1635 5241 1685 5341
rect 7031 5378 7081 5478
rect 7239 5378 7289 5478
rect 7457 5378 7507 5478
rect 9152 5450 9202 5550
rect 9370 5450 9420 5550
rect 9578 5450 9628 5550
rect 20835 5605 20885 5705
rect 21043 5605 21093 5705
rect 21261 5605 21311 5705
rect 23043 5676 23093 5776
rect 23261 5676 23311 5776
rect 23469 5676 23519 5776
rect 3465 5181 3515 5281
rect 3673 5181 3723 5281
rect 3891 5181 3941 5281
rect 5573 5254 5623 5354
rect 5791 5254 5841 5354
rect 5999 5254 6049 5354
rect 11408 5390 11458 5490
rect 11616 5390 11666 5490
rect 11834 5390 11884 5490
rect 13516 5463 13566 5563
rect 13734 5463 13784 5563
rect 13942 5463 13992 5563
rect 25199 5618 25249 5718
rect 25407 5618 25457 5718
rect 25625 5618 25675 5718
rect 27420 5688 27470 5788
rect 27638 5688 27688 5788
rect 27846 5688 27896 5788
rect 7829 5194 7879 5294
rect 8037 5194 8087 5294
rect 8255 5194 8305 5294
rect 9950 5266 10000 5366
rect 10168 5266 10218 5366
rect 10376 5266 10426 5366
rect 15772 5403 15822 5503
rect 15980 5403 16030 5503
rect 16198 5403 16248 5503
rect 17782 5437 17832 5537
rect 18000 5437 18050 5537
rect 18208 5437 18258 5537
rect 29576 5630 29626 5730
rect 29784 5630 29834 5730
rect 30002 5630 30052 5730
rect 31784 5701 31834 5801
rect 32002 5701 32052 5801
rect 32210 5701 32260 5801
rect 412 5013 462 5113
rect 630 5013 680 5113
rect 838 5013 888 5113
rect 12206 5206 12256 5306
rect 12414 5206 12464 5306
rect 12632 5206 12682 5306
rect 14314 5279 14364 5379
rect 14532 5279 14582 5379
rect 14740 5279 14790 5379
rect 20038 5377 20088 5477
rect 20246 5377 20296 5477
rect 20464 5377 20514 5477
rect 22146 5450 22196 5550
rect 22364 5450 22414 5550
rect 22572 5450 22622 5550
rect 33940 5643 33990 5743
rect 34148 5643 34198 5743
rect 34366 5643 34416 5743
rect 2363 4959 2413 5059
rect 2571 4959 2621 5059
rect 2789 4959 2839 5059
rect 4776 5026 4826 5126
rect 4994 5026 5044 5126
rect 5202 5026 5252 5126
rect 16570 5219 16620 5319
rect 16778 5219 16828 5319
rect 16996 5219 17046 5319
rect 18580 5253 18630 5353
rect 18798 5253 18848 5353
rect 19006 5253 19056 5353
rect 24402 5390 24452 5490
rect 24610 5390 24660 5490
rect 24828 5390 24878 5490
rect 26523 5462 26573 5562
rect 26741 5462 26791 5562
rect 26949 5462 26999 5562
rect 6727 4972 6777 5072
rect 6935 4972 6985 5072
rect 7153 4972 7203 5072
rect 9153 5038 9203 5138
rect 9371 5038 9421 5138
rect 9579 5038 9629 5138
rect 11104 4984 11154 5084
rect 11312 4984 11362 5084
rect 11530 4984 11580 5084
rect 13517 5051 13567 5151
rect 13735 5051 13785 5151
rect 13943 5051 13993 5151
rect 20836 5193 20886 5293
rect 21044 5193 21094 5293
rect 21262 5193 21312 5293
rect 22944 5266 22994 5366
rect 23162 5266 23212 5366
rect 23370 5266 23420 5366
rect 28779 5402 28829 5502
rect 28987 5402 29037 5502
rect 29205 5402 29255 5502
rect 30887 5475 30937 5575
rect 31105 5475 31155 5575
rect 31313 5475 31363 5575
rect 25200 5206 25250 5306
rect 25408 5206 25458 5306
rect 25626 5206 25676 5306
rect 27321 5278 27371 5378
rect 27539 5278 27589 5378
rect 27747 5278 27797 5378
rect 33143 5415 33193 5515
rect 33351 5415 33401 5515
rect 33569 5415 33619 5515
rect 15468 4997 15518 5097
rect 15676 4997 15726 5097
rect 15894 4997 15944 5097
rect 17783 5025 17833 5125
rect 18001 5025 18051 5125
rect 18209 5025 18259 5125
rect 29577 5218 29627 5318
rect 29785 5218 29835 5318
rect 30003 5218 30053 5318
rect 31685 5291 31735 5391
rect 31903 5291 31953 5391
rect 32111 5291 32161 5391
rect 19734 4971 19784 5071
rect 19942 4971 19992 5071
rect 20160 4971 20210 5071
rect 22147 5038 22197 5138
rect 22365 5038 22415 5138
rect 22573 5038 22623 5138
rect 33941 5231 33991 5331
rect 34149 5231 34199 5331
rect 34367 5231 34417 5331
rect 24098 4984 24148 5084
rect 24306 4984 24356 5084
rect 24524 4984 24574 5084
rect 26524 5050 26574 5150
rect 26742 5050 26792 5150
rect 26950 5050 27000 5150
rect 28475 4996 28525 5096
rect 28683 4996 28733 5096
rect 28901 4996 28951 5096
rect 30888 5063 30938 5163
rect 31106 5063 31156 5163
rect 31314 5063 31364 5163
rect 32839 5009 32889 5109
rect 33047 5009 33097 5109
rect 33265 5009 33315 5109
rect 1494 4629 1544 4729
rect 1712 4629 1762 4729
rect 1920 4629 1970 4729
rect 3445 4575 3495 4675
rect 3653 4575 3703 4675
rect 3871 4575 3921 4675
rect 5858 4642 5908 4742
rect 6076 4642 6126 4742
rect 6284 4642 6334 4742
rect 7809 4588 7859 4688
rect 8017 4588 8067 4688
rect 8235 4588 8285 4688
rect 10235 4654 10285 4754
rect 10453 4654 10503 4754
rect 10661 4654 10711 4754
rect 392 4407 442 4507
rect 610 4407 660 4507
rect 818 4407 868 4507
rect 12186 4600 12236 4700
rect 12394 4600 12444 4700
rect 12612 4600 12662 4700
rect 14599 4667 14649 4767
rect 14817 4667 14867 4767
rect 15025 4667 15075 4767
rect 2648 4347 2698 4447
rect 2856 4347 2906 4447
rect 3074 4347 3124 4447
rect 4756 4420 4806 4520
rect 4974 4420 5024 4520
rect 5182 4420 5232 4520
rect 16550 4613 16600 4713
rect 16758 4613 16808 4713
rect 16976 4613 17026 4713
rect 18865 4641 18915 4741
rect 19083 4641 19133 4741
rect 19291 4641 19341 4741
rect 1190 4223 1240 4323
rect 1408 4223 1458 4323
rect 1616 4223 1666 4323
rect 7012 4360 7062 4460
rect 7220 4360 7270 4460
rect 7438 4360 7488 4460
rect 9133 4432 9183 4532
rect 9351 4432 9401 4532
rect 9559 4432 9609 4532
rect 3446 4163 3496 4263
rect 3654 4163 3704 4263
rect 3872 4163 3922 4263
rect 5554 4236 5604 4336
rect 5772 4236 5822 4336
rect 5980 4236 6030 4336
rect 11389 4372 11439 4472
rect 11597 4372 11647 4472
rect 11815 4372 11865 4472
rect 13497 4445 13547 4545
rect 13715 4445 13765 4545
rect 13923 4445 13973 4545
rect 20816 4587 20866 4687
rect 21024 4587 21074 4687
rect 21242 4587 21292 4687
rect 23229 4654 23279 4754
rect 23447 4654 23497 4754
rect 23655 4654 23705 4754
rect 25180 4600 25230 4700
rect 25388 4600 25438 4700
rect 25606 4600 25656 4700
rect 27606 4666 27656 4766
rect 27824 4666 27874 4766
rect 28032 4666 28082 4766
rect 7810 4176 7860 4276
rect 8018 4176 8068 4276
rect 8236 4176 8286 4276
rect 9931 4248 9981 4348
rect 10149 4248 10199 4348
rect 10357 4248 10407 4348
rect 15753 4385 15803 4485
rect 15961 4385 16011 4485
rect 16179 4385 16229 4485
rect 17763 4419 17813 4519
rect 17981 4419 18031 4519
rect 18189 4419 18239 4519
rect 29557 4612 29607 4712
rect 29765 4612 29815 4712
rect 29983 4612 30033 4712
rect 31970 4679 32020 4779
rect 32188 4679 32238 4779
rect 32396 4679 32446 4779
rect 393 3995 443 4095
rect 611 3995 661 4095
rect 819 3995 869 4095
rect 12187 4188 12237 4288
rect 12395 4188 12445 4288
rect 12613 4188 12663 4288
rect 14295 4261 14345 4361
rect 14513 4261 14563 4361
rect 14721 4261 14771 4361
rect 20019 4359 20069 4459
rect 20227 4359 20277 4459
rect 20445 4359 20495 4459
rect 22127 4432 22177 4532
rect 22345 4432 22395 4532
rect 22553 4432 22603 4532
rect 33921 4625 33971 4725
rect 34129 4625 34179 4725
rect 34347 4625 34397 4725
rect 2549 3937 2599 4037
rect 2757 3937 2807 4037
rect 2975 3937 3025 4037
rect 4757 4008 4807 4108
rect 4975 4008 5025 4108
rect 5183 4008 5233 4108
rect 16551 4201 16601 4301
rect 16759 4201 16809 4301
rect 16977 4201 17027 4301
rect 18561 4235 18611 4335
rect 18779 4235 18829 4335
rect 18987 4235 19037 4335
rect 24383 4372 24433 4472
rect 24591 4372 24641 4472
rect 24809 4372 24859 4472
rect 26504 4444 26554 4544
rect 26722 4444 26772 4544
rect 26930 4444 26980 4544
rect 6913 3950 6963 4050
rect 7121 3950 7171 4050
rect 7339 3950 7389 4050
rect 9134 4020 9184 4120
rect 9352 4020 9402 4120
rect 9560 4020 9610 4120
rect 20817 4175 20867 4275
rect 21025 4175 21075 4275
rect 21243 4175 21293 4275
rect 22925 4248 22975 4348
rect 23143 4248 23193 4348
rect 23351 4248 23401 4348
rect 28760 4384 28810 4484
rect 28968 4384 29018 4484
rect 29186 4384 29236 4484
rect 30868 4457 30918 4557
rect 31086 4457 31136 4557
rect 31294 4457 31344 4557
rect 11290 3962 11340 4062
rect 11498 3962 11548 4062
rect 11716 3962 11766 4062
rect 13498 4033 13548 4133
rect 13716 4033 13766 4133
rect 13924 4033 13974 4133
rect 25181 4188 25231 4288
rect 25389 4188 25439 4288
rect 25607 4188 25657 4288
rect 27302 4260 27352 4360
rect 27520 4260 27570 4360
rect 27728 4260 27778 4360
rect 33124 4397 33174 4497
rect 33332 4397 33382 4497
rect 33550 4397 33600 4497
rect 15654 3975 15704 4075
rect 15862 3975 15912 4075
rect 16080 3975 16130 4075
rect 17764 4007 17814 4107
rect 17982 4007 18032 4107
rect 18190 4007 18240 4107
rect 29558 4200 29608 4300
rect 29766 4200 29816 4300
rect 29984 4200 30034 4300
rect 31666 4273 31716 4373
rect 31884 4273 31934 4373
rect 32092 4273 32142 4373
rect 19920 3949 19970 4049
rect 20128 3949 20178 4049
rect 20346 3949 20396 4049
rect 22128 4020 22178 4120
rect 22346 4020 22396 4120
rect 22554 4020 22604 4120
rect 33922 4213 33972 4313
rect 34130 4213 34180 4313
rect 34348 4213 34398 4313
rect 24284 3962 24334 4062
rect 24492 3962 24542 4062
rect 24710 3962 24760 4062
rect 26505 4032 26555 4132
rect 26723 4032 26773 4132
rect 26931 4032 26981 4132
rect 28661 3974 28711 4074
rect 28869 3974 28919 4074
rect 29087 3974 29137 4074
rect 30869 4045 30919 4145
rect 31087 4045 31137 4145
rect 31295 4045 31345 4145
rect 33025 3987 33075 4087
rect 33233 3987 33283 4087
rect 33451 3987 33501 4087
rect 1272 3615 1322 3715
rect 1490 3615 1540 3715
rect 1698 3615 1748 3715
rect 3428 3557 3478 3657
rect 3636 3557 3686 3657
rect 3854 3557 3904 3657
rect 5636 3628 5686 3728
rect 5854 3628 5904 3728
rect 6062 3628 6112 3728
rect 7792 3570 7842 3670
rect 8000 3570 8050 3670
rect 8218 3570 8268 3670
rect 10013 3640 10063 3740
rect 10231 3640 10281 3740
rect 10439 3640 10489 3740
rect 375 3389 425 3489
rect 593 3389 643 3489
rect 801 3389 851 3489
rect 12169 3582 12219 3682
rect 12377 3582 12427 3682
rect 12595 3582 12645 3682
rect 14377 3653 14427 3753
rect 14595 3653 14645 3753
rect 14803 3653 14853 3753
rect 2631 3329 2681 3429
rect 2839 3329 2889 3429
rect 3057 3329 3107 3429
rect 4739 3402 4789 3502
rect 4957 3402 5007 3502
rect 5165 3402 5215 3502
rect 16533 3595 16583 3695
rect 16741 3595 16791 3695
rect 16959 3595 17009 3695
rect 18643 3627 18693 3727
rect 18861 3627 18911 3727
rect 19069 3627 19119 3727
rect 1173 3205 1223 3305
rect 1391 3205 1441 3305
rect 1599 3205 1649 3305
rect 6995 3342 7045 3442
rect 7203 3342 7253 3442
rect 7421 3342 7471 3442
rect 9116 3414 9166 3514
rect 9334 3414 9384 3514
rect 9542 3414 9592 3514
rect 20799 3569 20849 3669
rect 21007 3569 21057 3669
rect 21225 3569 21275 3669
rect 23007 3640 23057 3740
rect 23225 3640 23275 3740
rect 23433 3640 23483 3740
rect 3429 3145 3479 3245
rect 3637 3145 3687 3245
rect 3855 3145 3905 3245
rect 5537 3218 5587 3318
rect 5755 3218 5805 3318
rect 5963 3218 6013 3318
rect 11372 3354 11422 3454
rect 11580 3354 11630 3454
rect 11798 3354 11848 3454
rect 13480 3427 13530 3527
rect 13698 3427 13748 3527
rect 13906 3427 13956 3527
rect 25163 3582 25213 3682
rect 25371 3582 25421 3682
rect 25589 3582 25639 3682
rect 27384 3652 27434 3752
rect 27602 3652 27652 3752
rect 27810 3652 27860 3752
rect 7793 3158 7843 3258
rect 8001 3158 8051 3258
rect 8219 3158 8269 3258
rect 9914 3230 9964 3330
rect 10132 3230 10182 3330
rect 10340 3230 10390 3330
rect 15736 3367 15786 3467
rect 15944 3367 15994 3467
rect 16162 3367 16212 3467
rect 17746 3401 17796 3501
rect 17964 3401 18014 3501
rect 18172 3401 18222 3501
rect 29540 3594 29590 3694
rect 29748 3594 29798 3694
rect 29966 3594 30016 3694
rect 31748 3665 31798 3765
rect 31966 3665 32016 3765
rect 32174 3665 32224 3765
rect 376 2977 426 3077
rect 594 2977 644 3077
rect 802 2977 852 3077
rect 12170 3170 12220 3270
rect 12378 3170 12428 3270
rect 12596 3170 12646 3270
rect 14278 3243 14328 3343
rect 14496 3243 14546 3343
rect 14704 3243 14754 3343
rect 20002 3341 20052 3441
rect 20210 3341 20260 3441
rect 20428 3341 20478 3441
rect 22110 3414 22160 3514
rect 22328 3414 22378 3514
rect 22536 3414 22586 3514
rect 33904 3607 33954 3707
rect 34112 3607 34162 3707
rect 34330 3607 34380 3707
rect 2466 2921 2516 3021
rect 2674 2921 2724 3021
rect 2892 2921 2942 3021
rect 4740 2990 4790 3090
rect 4958 2990 5008 3090
rect 5166 2990 5216 3090
rect 16534 3183 16584 3283
rect 16742 3183 16792 3283
rect 16960 3183 17010 3283
rect 18544 3217 18594 3317
rect 18762 3217 18812 3317
rect 18970 3217 19020 3317
rect 24366 3354 24416 3454
rect 24574 3354 24624 3454
rect 24792 3354 24842 3454
rect 26487 3426 26537 3526
rect 26705 3426 26755 3526
rect 26913 3426 26963 3526
rect 6830 2934 6880 3034
rect 7038 2934 7088 3034
rect 7256 2934 7306 3034
rect 9117 3002 9167 3102
rect 9335 3002 9385 3102
rect 9543 3002 9593 3102
rect 20800 3157 20850 3257
rect 21008 3157 21058 3257
rect 21226 3157 21276 3257
rect 22908 3230 22958 3330
rect 23126 3230 23176 3330
rect 23334 3230 23384 3330
rect 28743 3366 28793 3466
rect 28951 3366 29001 3466
rect 29169 3366 29219 3466
rect 30851 3439 30901 3539
rect 31069 3439 31119 3539
rect 31277 3439 31327 3539
rect 11207 2946 11257 3046
rect 11415 2946 11465 3046
rect 11633 2946 11683 3046
rect 13481 3015 13531 3115
rect 13699 3015 13749 3115
rect 13907 3015 13957 3115
rect 25164 3170 25214 3270
rect 25372 3170 25422 3270
rect 25590 3170 25640 3270
rect 27285 3242 27335 3342
rect 27503 3242 27553 3342
rect 27711 3242 27761 3342
rect 33107 3379 33157 3479
rect 33315 3379 33365 3479
rect 33533 3379 33583 3479
rect 15571 2959 15621 3059
rect 15779 2959 15829 3059
rect 15997 2959 16047 3059
rect 17747 2989 17797 3089
rect 17965 2989 18015 3089
rect 18173 2989 18223 3089
rect 29541 3182 29591 3282
rect 29749 3182 29799 3282
rect 29967 3182 30017 3282
rect 31649 3255 31699 3355
rect 31867 3255 31917 3355
rect 32075 3255 32125 3355
rect 19837 2933 19887 3033
rect 20045 2933 20095 3033
rect 20263 2933 20313 3033
rect 22111 3002 22161 3102
rect 22329 3002 22379 3102
rect 22537 3002 22587 3102
rect 33905 3195 33955 3295
rect 34113 3195 34163 3295
rect 34331 3195 34381 3295
rect 24201 2946 24251 3046
rect 24409 2946 24459 3046
rect 24627 2946 24677 3046
rect 26488 3014 26538 3114
rect 26706 3014 26756 3114
rect 26914 3014 26964 3114
rect 28578 2958 28628 3058
rect 28786 2958 28836 3058
rect 29004 2958 29054 3058
rect 30852 3027 30902 3127
rect 31070 3027 31120 3127
rect 31278 3027 31328 3127
rect 32942 2971 32992 3071
rect 33150 2971 33200 3071
rect 33368 2971 33418 3071
rect 1318 2595 1368 2695
rect 1536 2595 1586 2695
rect 1744 2595 1794 2695
rect 3408 2539 3458 2639
rect 3616 2539 3666 2639
rect 3834 2539 3884 2639
rect 5682 2608 5732 2708
rect 5900 2608 5950 2708
rect 6108 2608 6158 2708
rect 7772 2552 7822 2652
rect 7980 2552 8030 2652
rect 8198 2552 8248 2652
rect 10059 2620 10109 2720
rect 10277 2620 10327 2720
rect 10485 2620 10535 2720
rect 355 2371 405 2471
rect 573 2371 623 2471
rect 781 2371 831 2471
rect 12149 2564 12199 2664
rect 12357 2564 12407 2664
rect 12575 2564 12625 2664
rect 14423 2633 14473 2733
rect 14641 2633 14691 2733
rect 14849 2633 14899 2733
rect 2611 2311 2661 2411
rect 2819 2311 2869 2411
rect 3037 2311 3087 2411
rect 4719 2384 4769 2484
rect 4937 2384 4987 2484
rect 5145 2384 5195 2484
rect 16513 2577 16563 2677
rect 16721 2577 16771 2677
rect 16939 2577 16989 2677
rect 18689 2607 18739 2707
rect 18907 2607 18957 2707
rect 19115 2607 19165 2707
rect 1153 2187 1203 2287
rect 1371 2187 1421 2287
rect 1579 2187 1629 2287
rect 6975 2324 7025 2424
rect 7183 2324 7233 2424
rect 7401 2324 7451 2424
rect 9096 2396 9146 2496
rect 9314 2396 9364 2496
rect 9522 2396 9572 2496
rect 20779 2551 20829 2651
rect 20987 2551 21037 2651
rect 21205 2551 21255 2651
rect 23053 2620 23103 2720
rect 23271 2620 23321 2720
rect 23479 2620 23529 2720
rect 3409 2127 3459 2227
rect 3617 2127 3667 2227
rect 3835 2127 3885 2227
rect 5517 2200 5567 2300
rect 5735 2200 5785 2300
rect 5943 2200 5993 2300
rect 11352 2336 11402 2436
rect 11560 2336 11610 2436
rect 11778 2336 11828 2436
rect 13460 2409 13510 2509
rect 13678 2409 13728 2509
rect 13886 2409 13936 2509
rect 25143 2564 25193 2664
rect 25351 2564 25401 2664
rect 25569 2564 25619 2664
rect 27430 2632 27480 2732
rect 27648 2632 27698 2732
rect 27856 2632 27906 2732
rect 7773 2140 7823 2240
rect 7981 2140 8031 2240
rect 8199 2140 8249 2240
rect 9894 2212 9944 2312
rect 10112 2212 10162 2312
rect 10320 2212 10370 2312
rect 15716 2349 15766 2449
rect 15924 2349 15974 2449
rect 16142 2349 16192 2449
rect 17726 2383 17776 2483
rect 17944 2383 17994 2483
rect 18152 2383 18202 2483
rect 29520 2576 29570 2676
rect 29728 2576 29778 2676
rect 29946 2576 29996 2676
rect 31794 2645 31844 2745
rect 32012 2645 32062 2745
rect 32220 2645 32270 2745
rect 356 1959 406 2059
rect 574 1959 624 2059
rect 782 1959 832 2059
rect 12150 2152 12200 2252
rect 12358 2152 12408 2252
rect 12576 2152 12626 2252
rect 14258 2225 14308 2325
rect 14476 2225 14526 2325
rect 14684 2225 14734 2325
rect 19982 2323 20032 2423
rect 20190 2323 20240 2423
rect 20408 2323 20458 2423
rect 22090 2396 22140 2496
rect 22308 2396 22358 2496
rect 22516 2396 22566 2496
rect 33884 2589 33934 2689
rect 34092 2589 34142 2689
rect 34310 2589 34360 2689
rect 2512 1901 2562 2001
rect 2720 1901 2770 2001
rect 2938 1901 2988 2001
rect 4720 1972 4770 2072
rect 4938 1972 4988 2072
rect 5146 1972 5196 2072
rect 16514 2165 16564 2265
rect 16722 2165 16772 2265
rect 16940 2165 16990 2265
rect 18524 2199 18574 2299
rect 18742 2199 18792 2299
rect 18950 2199 19000 2299
rect 24346 2336 24396 2436
rect 24554 2336 24604 2436
rect 24772 2336 24822 2436
rect 26467 2408 26517 2508
rect 26685 2408 26735 2508
rect 26893 2408 26943 2508
rect 6876 1914 6926 2014
rect 7084 1914 7134 2014
rect 7302 1914 7352 2014
rect 9097 1984 9147 2084
rect 9315 1984 9365 2084
rect 9523 1984 9573 2084
rect 20780 2139 20830 2239
rect 20988 2139 21038 2239
rect 21206 2139 21256 2239
rect 22888 2212 22938 2312
rect 23106 2212 23156 2312
rect 23314 2212 23364 2312
rect 28723 2348 28773 2448
rect 28931 2348 28981 2448
rect 29149 2348 29199 2448
rect 30831 2421 30881 2521
rect 31049 2421 31099 2521
rect 31257 2421 31307 2521
rect 11253 1926 11303 2026
rect 11461 1926 11511 2026
rect 11679 1926 11729 2026
rect 13461 1997 13511 2097
rect 13679 1997 13729 2097
rect 13887 1997 13937 2097
rect 25144 2152 25194 2252
rect 25352 2152 25402 2252
rect 25570 2152 25620 2252
rect 27265 2224 27315 2324
rect 27483 2224 27533 2324
rect 27691 2224 27741 2324
rect 33087 2361 33137 2461
rect 33295 2361 33345 2461
rect 33513 2361 33563 2461
rect 15617 1939 15667 2039
rect 15825 1939 15875 2039
rect 16043 1939 16093 2039
rect 17727 1971 17777 2071
rect 17945 1971 17995 2071
rect 18153 1971 18203 2071
rect 29521 2164 29571 2264
rect 29729 2164 29779 2264
rect 29947 2164 29997 2264
rect 31629 2237 31679 2337
rect 31847 2237 31897 2337
rect 32055 2237 32105 2337
rect 19883 1913 19933 2013
rect 20091 1913 20141 2013
rect 20309 1913 20359 2013
rect 22091 1984 22141 2084
rect 22309 1984 22359 2084
rect 22517 1984 22567 2084
rect 33885 2177 33935 2277
rect 34093 2177 34143 2277
rect 34311 2177 34361 2277
rect 24247 1926 24297 2026
rect 24455 1926 24505 2026
rect 24673 1926 24723 2026
rect 26468 1996 26518 2096
rect 26686 1996 26736 2096
rect 26894 1996 26944 2096
rect 28624 1938 28674 2038
rect 28832 1938 28882 2038
rect 29050 1938 29100 2038
rect 30832 2009 30882 2109
rect 31050 2009 31100 2109
rect 31258 2009 31308 2109
rect 32988 1951 33038 2051
rect 33196 1951 33246 2051
rect 33414 1951 33464 2051
rect 1235 1579 1285 1679
rect 1453 1579 1503 1679
rect 1661 1579 1711 1679
rect 3391 1521 3441 1621
rect 3599 1521 3649 1621
rect 3817 1521 3867 1621
rect 5599 1592 5649 1692
rect 5817 1592 5867 1692
rect 6025 1592 6075 1692
rect 7755 1534 7805 1634
rect 7963 1534 8013 1634
rect 8181 1534 8231 1634
rect 9976 1604 10026 1704
rect 10194 1604 10244 1704
rect 10402 1604 10452 1704
rect 338 1353 388 1453
rect 556 1353 606 1453
rect 764 1353 814 1453
rect 12132 1546 12182 1646
rect 12340 1546 12390 1646
rect 12558 1546 12608 1646
rect 14340 1617 14390 1717
rect 14558 1617 14608 1717
rect 14766 1617 14816 1717
rect 2594 1293 2644 1393
rect 2802 1293 2852 1393
rect 3020 1293 3070 1393
rect 4702 1366 4752 1466
rect 4920 1366 4970 1466
rect 5128 1366 5178 1466
rect 16496 1559 16546 1659
rect 16704 1559 16754 1659
rect 16922 1559 16972 1659
rect 18606 1591 18656 1691
rect 18824 1591 18874 1691
rect 19032 1591 19082 1691
rect 1136 1169 1186 1269
rect 1354 1169 1404 1269
rect 1562 1169 1612 1269
rect 6958 1306 7008 1406
rect 7166 1306 7216 1406
rect 7384 1306 7434 1406
rect 9079 1378 9129 1478
rect 9297 1378 9347 1478
rect 9505 1378 9555 1478
rect 20762 1533 20812 1633
rect 20970 1533 21020 1633
rect 21188 1533 21238 1633
rect 22970 1604 23020 1704
rect 23188 1604 23238 1704
rect 23396 1604 23446 1704
rect 3392 1109 3442 1209
rect 3600 1109 3650 1209
rect 3818 1109 3868 1209
rect 5500 1182 5550 1282
rect 5718 1182 5768 1282
rect 5926 1182 5976 1282
rect 11335 1318 11385 1418
rect 11543 1318 11593 1418
rect 11761 1318 11811 1418
rect 13443 1391 13493 1491
rect 13661 1391 13711 1491
rect 13869 1391 13919 1491
rect 25126 1546 25176 1646
rect 25334 1546 25384 1646
rect 25552 1546 25602 1646
rect 27347 1616 27397 1716
rect 27565 1616 27615 1716
rect 27773 1616 27823 1716
rect 7756 1122 7806 1222
rect 7964 1122 8014 1222
rect 8182 1122 8232 1222
rect 9877 1194 9927 1294
rect 10095 1194 10145 1294
rect 10303 1194 10353 1294
rect 15699 1331 15749 1431
rect 15907 1331 15957 1431
rect 16125 1331 16175 1431
rect 17709 1365 17759 1465
rect 17927 1365 17977 1465
rect 18135 1365 18185 1465
rect 29503 1558 29553 1658
rect 29711 1558 29761 1658
rect 29929 1558 29979 1658
rect 31711 1629 31761 1729
rect 31929 1629 31979 1729
rect 32137 1629 32187 1729
rect 12133 1134 12183 1234
rect 12341 1134 12391 1234
rect 12559 1134 12609 1234
rect 14241 1207 14291 1307
rect 14459 1207 14509 1307
rect 14667 1207 14717 1307
rect 19965 1305 20015 1405
rect 20173 1305 20223 1405
rect 20391 1305 20441 1405
rect 22073 1378 22123 1478
rect 22291 1378 22341 1478
rect 22499 1378 22549 1478
rect 33867 1571 33917 1671
rect 34075 1571 34125 1671
rect 34293 1571 34343 1671
rect 16497 1147 16547 1247
rect 16705 1147 16755 1247
rect 16923 1147 16973 1247
rect 18507 1181 18557 1281
rect 18725 1181 18775 1281
rect 18933 1181 18983 1281
rect 24329 1318 24379 1418
rect 24537 1318 24587 1418
rect 24755 1318 24805 1418
rect 26450 1390 26500 1490
rect 26668 1390 26718 1490
rect 26876 1390 26926 1490
rect 339 941 389 1041
rect 557 941 607 1041
rect 765 941 815 1041
rect 4703 954 4753 1054
rect 4921 954 4971 1054
rect 5129 954 5179 1054
rect 9080 966 9130 1066
rect 9298 966 9348 1066
rect 9506 966 9556 1066
rect 20763 1121 20813 1221
rect 20971 1121 21021 1221
rect 21189 1121 21239 1221
rect 22871 1194 22921 1294
rect 23089 1194 23139 1294
rect 23297 1194 23347 1294
rect 28706 1330 28756 1430
rect 28914 1330 28964 1430
rect 29132 1330 29182 1430
rect 30814 1403 30864 1503
rect 31032 1403 31082 1503
rect 31240 1403 31290 1503
rect 25127 1134 25177 1234
rect 25335 1134 25385 1234
rect 25553 1134 25603 1234
rect 27248 1206 27298 1306
rect 27466 1206 27516 1306
rect 27674 1206 27724 1306
rect 33070 1343 33120 1443
rect 33278 1343 33328 1443
rect 33496 1343 33546 1443
rect 29504 1146 29554 1246
rect 29712 1146 29762 1246
rect 29930 1146 29980 1246
rect 31612 1219 31662 1319
rect 31830 1219 31880 1319
rect 32038 1219 32088 1319
rect 33868 1159 33918 1259
rect 34076 1159 34126 1259
rect 34294 1159 34344 1259
rect 13444 979 13494 1079
rect 13662 979 13712 1079
rect 13870 979 13920 1079
rect 17710 953 17760 1053
rect 17928 953 17978 1053
rect 18136 953 18186 1053
rect 22074 966 22124 1066
rect 22292 966 22342 1066
rect 22500 966 22550 1066
rect 26451 978 26501 1078
rect 26669 978 26719 1078
rect 26877 978 26927 1078
rect 30815 991 30865 1091
rect 31033 991 31083 1091
rect 31241 991 31291 1091
rect 1552 365 1602 465
rect 1770 365 1820 465
rect 1978 365 2028 465
rect 4041 291 4091 391
rect 4259 291 4309 391
rect 4467 291 4517 391
rect 5916 378 5966 478
rect 6134 378 6184 478
rect 6342 378 6392 478
rect 8489 315 8539 415
rect 8707 315 8757 415
rect 8915 315 8965 415
rect 10293 390 10343 490
rect 10511 390 10561 490
rect 10719 390 10769 490
rect 12782 316 12832 416
rect 13000 316 13050 416
rect 13208 316 13258 416
rect 14657 403 14707 503
rect 14875 403 14925 503
rect 15083 403 15133 503
rect 18923 377 18973 477
rect 19141 377 19191 477
rect 19349 377 19399 477
rect 16979 252 17029 352
rect 17197 252 17247 352
rect 17405 252 17455 352
rect 21412 303 21462 403
rect 21630 303 21680 403
rect 21838 303 21888 403
rect 23287 390 23337 490
rect 23505 390 23555 490
rect 23713 390 23763 490
rect 25860 327 25910 427
rect 26078 327 26128 427
rect 26286 327 26336 427
rect 27664 402 27714 502
rect 27882 402 27932 502
rect 28090 402 28140 502
rect 30153 328 30203 428
rect 30371 328 30421 428
rect 30579 328 30629 428
rect 32028 415 32078 515
rect 32246 415 32296 515
rect 32454 415 32504 515
<< ndiff >>
rect 3469 8854 3518 8866
rect 3469 8834 3480 8854
rect 3500 8834 3518 8854
rect 3469 8824 3518 8834
rect 3568 8850 3612 8866
rect 3568 8830 3583 8850
rect 3603 8830 3612 8850
rect 3568 8824 3612 8830
rect 3682 8850 3726 8866
rect 3682 8830 3691 8850
rect 3711 8830 3726 8850
rect 3682 8824 3726 8830
rect 3776 8854 3825 8866
rect 3776 8834 3794 8854
rect 3814 8834 3825 8854
rect 3776 8824 3825 8834
rect 3900 8850 3944 8866
rect 3900 8830 3909 8850
rect 3929 8830 3944 8850
rect 3900 8824 3944 8830
rect 3994 8854 4043 8866
rect 3994 8834 4012 8854
rect 4032 8834 4043 8854
rect 3994 8824 4043 8834
rect 7833 8867 7882 8879
rect 7833 8847 7844 8867
rect 7864 8847 7882 8867
rect 7833 8837 7882 8847
rect 7932 8863 7976 8879
rect 7932 8843 7947 8863
rect 7967 8843 7976 8863
rect 7932 8837 7976 8843
rect 8046 8863 8090 8879
rect 8046 8843 8055 8863
rect 8075 8843 8090 8863
rect 8046 8837 8090 8843
rect 8140 8867 8189 8879
rect 8140 8847 8158 8867
rect 8178 8847 8189 8867
rect 8140 8837 8189 8847
rect 8264 8863 8308 8879
rect 8264 8843 8273 8863
rect 8293 8843 8308 8863
rect 8264 8837 8308 8843
rect 8358 8867 8407 8879
rect 8358 8847 8376 8867
rect 8396 8847 8407 8867
rect 8358 8837 8407 8847
rect 12210 8879 12259 8891
rect 12210 8859 12221 8879
rect 12241 8859 12259 8879
rect 12210 8849 12259 8859
rect 12309 8875 12353 8891
rect 12309 8855 12324 8875
rect 12344 8855 12353 8875
rect 12309 8849 12353 8855
rect 12423 8875 12467 8891
rect 12423 8855 12432 8875
rect 12452 8855 12467 8875
rect 12423 8849 12467 8855
rect 12517 8879 12566 8891
rect 12517 8859 12535 8879
rect 12555 8859 12566 8879
rect 12517 8849 12566 8859
rect 12641 8875 12685 8891
rect 12641 8855 12650 8875
rect 12670 8855 12685 8875
rect 12641 8849 12685 8855
rect 12735 8879 12784 8891
rect 12735 8859 12753 8879
rect 12773 8859 12784 8879
rect 12735 8849 12784 8859
rect 16574 8892 16623 8904
rect 2672 8626 2721 8638
rect 2672 8606 2683 8626
rect 2703 8606 2721 8626
rect 2672 8596 2721 8606
rect 2771 8622 2815 8638
rect 2771 8602 2786 8622
rect 2806 8602 2815 8622
rect 2771 8596 2815 8602
rect 2885 8622 2929 8638
rect 2885 8602 2894 8622
rect 2914 8602 2929 8622
rect 2885 8596 2929 8602
rect 2979 8626 3028 8638
rect 2979 8606 2997 8626
rect 3017 8606 3028 8626
rect 2979 8596 3028 8606
rect 3103 8622 3147 8638
rect 3103 8602 3112 8622
rect 3132 8602 3147 8622
rect 3103 8596 3147 8602
rect 3197 8626 3246 8638
rect 16574 8872 16585 8892
rect 16605 8872 16623 8892
rect 16574 8862 16623 8872
rect 16673 8888 16717 8904
rect 16673 8868 16688 8888
rect 16708 8868 16717 8888
rect 16673 8862 16717 8868
rect 16787 8888 16831 8904
rect 16787 8868 16796 8888
rect 16816 8868 16831 8888
rect 16787 8862 16831 8868
rect 16881 8892 16930 8904
rect 16881 8872 16899 8892
rect 16919 8872 16930 8892
rect 16881 8862 16930 8872
rect 17005 8888 17049 8904
rect 17005 8868 17014 8888
rect 17034 8868 17049 8888
rect 17005 8862 17049 8868
rect 17099 8892 17148 8904
rect 17099 8872 17117 8892
rect 17137 8872 17148 8892
rect 17099 8862 17148 8872
rect 3197 8606 3215 8626
rect 3235 8606 3246 8626
rect 3197 8596 3246 8606
rect 7036 8639 7085 8651
rect 7036 8619 7047 8639
rect 7067 8619 7085 8639
rect 7036 8609 7085 8619
rect 7135 8635 7179 8651
rect 7135 8615 7150 8635
rect 7170 8615 7179 8635
rect 7135 8609 7179 8615
rect 7249 8635 7293 8651
rect 7249 8615 7258 8635
rect 7278 8615 7293 8635
rect 7249 8609 7293 8615
rect 7343 8639 7392 8651
rect 7343 8619 7361 8639
rect 7381 8619 7392 8639
rect 7343 8609 7392 8619
rect 7467 8635 7511 8651
rect 7467 8615 7476 8635
rect 7496 8615 7511 8635
rect 7467 8609 7511 8615
rect 7561 8639 7610 8651
rect 20840 8866 20889 8878
rect 20840 8846 20851 8866
rect 20871 8846 20889 8866
rect 20840 8836 20889 8846
rect 20939 8862 20983 8878
rect 20939 8842 20954 8862
rect 20974 8842 20983 8862
rect 20939 8836 20983 8842
rect 21053 8862 21097 8878
rect 21053 8842 21062 8862
rect 21082 8842 21097 8862
rect 21053 8836 21097 8842
rect 21147 8866 21196 8878
rect 21147 8846 21165 8866
rect 21185 8846 21196 8866
rect 21147 8836 21196 8846
rect 21271 8862 21315 8878
rect 21271 8842 21280 8862
rect 21300 8842 21315 8862
rect 21271 8836 21315 8842
rect 21365 8866 21414 8878
rect 21365 8846 21383 8866
rect 21403 8846 21414 8866
rect 21365 8836 21414 8846
rect 25204 8879 25253 8891
rect 7561 8619 7579 8639
rect 7599 8619 7610 8639
rect 7561 8609 7610 8619
rect 11413 8651 11462 8663
rect 11413 8631 11424 8651
rect 11444 8631 11462 8651
rect 11413 8621 11462 8631
rect 11512 8647 11556 8663
rect 11512 8627 11527 8647
rect 11547 8627 11556 8647
rect 11512 8621 11556 8627
rect 11626 8647 11670 8663
rect 11626 8627 11635 8647
rect 11655 8627 11670 8647
rect 11626 8621 11670 8627
rect 11720 8651 11769 8663
rect 11720 8631 11738 8651
rect 11758 8631 11769 8651
rect 11720 8621 11769 8631
rect 11844 8647 11888 8663
rect 11844 8627 11853 8647
rect 11873 8627 11888 8647
rect 11844 8621 11888 8627
rect 11938 8651 11987 8663
rect 25204 8859 25215 8879
rect 25235 8859 25253 8879
rect 25204 8849 25253 8859
rect 25303 8875 25347 8891
rect 25303 8855 25318 8875
rect 25338 8855 25347 8875
rect 25303 8849 25347 8855
rect 25417 8875 25461 8891
rect 25417 8855 25426 8875
rect 25446 8855 25461 8875
rect 25417 8849 25461 8855
rect 25511 8879 25560 8891
rect 25511 8859 25529 8879
rect 25549 8859 25560 8879
rect 25511 8849 25560 8859
rect 25635 8875 25679 8891
rect 25635 8855 25644 8875
rect 25664 8855 25679 8875
rect 25635 8849 25679 8855
rect 25729 8879 25778 8891
rect 25729 8859 25747 8879
rect 25767 8859 25778 8879
rect 25729 8849 25778 8859
rect 29581 8891 29630 8903
rect 11938 8631 11956 8651
rect 11976 8631 11987 8651
rect 11938 8621 11987 8631
rect 15777 8664 15826 8676
rect 15777 8644 15788 8664
rect 15808 8644 15826 8664
rect 15777 8634 15826 8644
rect 15876 8660 15920 8676
rect 15876 8640 15891 8660
rect 15911 8640 15920 8660
rect 15876 8634 15920 8640
rect 15990 8660 16034 8676
rect 15990 8640 15999 8660
rect 16019 8640 16034 8660
rect 15990 8634 16034 8640
rect 16084 8664 16133 8676
rect 16084 8644 16102 8664
rect 16122 8644 16133 8664
rect 16084 8634 16133 8644
rect 16208 8660 16252 8676
rect 16208 8640 16217 8660
rect 16237 8640 16252 8660
rect 16208 8634 16252 8640
rect 16302 8664 16351 8676
rect 16302 8644 16320 8664
rect 16340 8644 16351 8664
rect 16302 8634 16351 8644
rect 29581 8871 29592 8891
rect 29612 8871 29630 8891
rect 29581 8861 29630 8871
rect 29680 8887 29724 8903
rect 29680 8867 29695 8887
rect 29715 8867 29724 8887
rect 29680 8861 29724 8867
rect 29794 8887 29838 8903
rect 29794 8867 29803 8887
rect 29823 8867 29838 8887
rect 29794 8861 29838 8867
rect 29888 8891 29937 8903
rect 29888 8871 29906 8891
rect 29926 8871 29937 8891
rect 29888 8861 29937 8871
rect 30012 8887 30056 8903
rect 30012 8867 30021 8887
rect 30041 8867 30056 8887
rect 30012 8861 30056 8867
rect 30106 8891 30155 8903
rect 30106 8871 30124 8891
rect 30144 8871 30155 8891
rect 30106 8861 30155 8871
rect 33945 8904 33994 8916
rect 3470 8442 3519 8454
rect 3470 8422 3481 8442
rect 3501 8422 3519 8442
rect 416 8392 465 8402
rect 416 8372 427 8392
rect 447 8372 465 8392
rect 416 8360 465 8372
rect 515 8396 559 8402
rect 515 8376 530 8396
rect 550 8376 559 8396
rect 515 8360 559 8376
rect 634 8392 683 8402
rect 634 8372 645 8392
rect 665 8372 683 8392
rect 634 8360 683 8372
rect 733 8396 777 8402
rect 733 8376 748 8396
rect 768 8376 777 8396
rect 733 8360 777 8376
rect 847 8396 891 8402
rect 847 8376 856 8396
rect 876 8376 891 8396
rect 847 8360 891 8376
rect 941 8392 990 8402
rect 3470 8412 3519 8422
rect 3569 8438 3613 8454
rect 3569 8418 3584 8438
rect 3604 8418 3613 8438
rect 3569 8412 3613 8418
rect 3683 8438 3727 8454
rect 3683 8418 3692 8438
rect 3712 8418 3727 8438
rect 3683 8412 3727 8418
rect 3777 8442 3826 8454
rect 3777 8422 3795 8442
rect 3815 8422 3826 8442
rect 3777 8412 3826 8422
rect 3901 8438 3945 8454
rect 3901 8418 3910 8438
rect 3930 8418 3945 8438
rect 3901 8412 3945 8418
rect 3995 8442 4044 8454
rect 3995 8422 4013 8442
rect 4033 8422 4044 8442
rect 3995 8412 4044 8422
rect 941 8372 959 8392
rect 979 8372 990 8392
rect 941 8360 990 8372
rect 7834 8455 7883 8467
rect 7834 8435 7845 8455
rect 7865 8435 7883 8455
rect 4780 8405 4829 8415
rect 4780 8385 4791 8405
rect 4811 8385 4829 8405
rect 4780 8373 4829 8385
rect 4879 8409 4923 8415
rect 4879 8389 4894 8409
rect 4914 8389 4923 8409
rect 4879 8373 4923 8389
rect 4998 8405 5047 8415
rect 4998 8385 5009 8405
rect 5029 8385 5047 8405
rect 4998 8373 5047 8385
rect 5097 8409 5141 8415
rect 5097 8389 5112 8409
rect 5132 8389 5141 8409
rect 5097 8373 5141 8389
rect 5211 8409 5255 8415
rect 5211 8389 5220 8409
rect 5240 8389 5255 8409
rect 5211 8373 5255 8389
rect 5305 8405 5354 8415
rect 7834 8425 7883 8435
rect 7933 8451 7977 8467
rect 7933 8431 7948 8451
rect 7968 8431 7977 8451
rect 7933 8425 7977 8431
rect 8047 8451 8091 8467
rect 8047 8431 8056 8451
rect 8076 8431 8091 8451
rect 8047 8425 8091 8431
rect 8141 8455 8190 8467
rect 8141 8435 8159 8455
rect 8179 8435 8190 8455
rect 8141 8425 8190 8435
rect 8265 8451 8309 8467
rect 8265 8431 8274 8451
rect 8294 8431 8309 8451
rect 8265 8425 8309 8431
rect 8359 8455 8408 8467
rect 8359 8435 8377 8455
rect 8397 8435 8408 8455
rect 8359 8425 8408 8435
rect 5305 8385 5323 8405
rect 5343 8385 5354 8405
rect 5305 8373 5354 8385
rect 20043 8638 20092 8650
rect 20043 8618 20054 8638
rect 20074 8618 20092 8638
rect 20043 8608 20092 8618
rect 20142 8634 20186 8650
rect 20142 8614 20157 8634
rect 20177 8614 20186 8634
rect 20142 8608 20186 8614
rect 20256 8634 20300 8650
rect 20256 8614 20265 8634
rect 20285 8614 20300 8634
rect 20256 8608 20300 8614
rect 20350 8638 20399 8650
rect 20350 8618 20368 8638
rect 20388 8618 20399 8638
rect 20350 8608 20399 8618
rect 20474 8634 20518 8650
rect 20474 8614 20483 8634
rect 20503 8614 20518 8634
rect 20474 8608 20518 8614
rect 20568 8638 20617 8650
rect 33945 8884 33956 8904
rect 33976 8884 33994 8904
rect 33945 8874 33994 8884
rect 34044 8900 34088 8916
rect 34044 8880 34059 8900
rect 34079 8880 34088 8900
rect 34044 8874 34088 8880
rect 34158 8900 34202 8916
rect 34158 8880 34167 8900
rect 34187 8880 34202 8900
rect 34158 8874 34202 8880
rect 34252 8904 34301 8916
rect 34252 8884 34270 8904
rect 34290 8884 34301 8904
rect 34252 8874 34301 8884
rect 34376 8900 34420 8916
rect 34376 8880 34385 8900
rect 34405 8880 34420 8900
rect 34376 8874 34420 8880
rect 34470 8904 34519 8916
rect 34470 8884 34488 8904
rect 34508 8884 34519 8904
rect 34470 8874 34519 8884
rect 20568 8618 20586 8638
rect 20606 8618 20617 8638
rect 20568 8608 20617 8618
rect 24407 8651 24456 8663
rect 24407 8631 24418 8651
rect 24438 8631 24456 8651
rect 24407 8621 24456 8631
rect 24506 8647 24550 8663
rect 24506 8627 24521 8647
rect 24541 8627 24550 8647
rect 24506 8621 24550 8627
rect 24620 8647 24664 8663
rect 24620 8627 24629 8647
rect 24649 8627 24664 8647
rect 24620 8621 24664 8627
rect 24714 8651 24763 8663
rect 24714 8631 24732 8651
rect 24752 8631 24763 8651
rect 24714 8621 24763 8631
rect 24838 8647 24882 8663
rect 24838 8627 24847 8647
rect 24867 8627 24882 8647
rect 24838 8621 24882 8627
rect 24932 8651 24981 8663
rect 24932 8631 24950 8651
rect 24970 8631 24981 8651
rect 24932 8621 24981 8631
rect 28784 8663 28833 8675
rect 28784 8643 28795 8663
rect 28815 8643 28833 8663
rect 28784 8633 28833 8643
rect 28883 8659 28927 8675
rect 28883 8639 28898 8659
rect 28918 8639 28927 8659
rect 28883 8633 28927 8639
rect 28997 8659 29041 8675
rect 28997 8639 29006 8659
rect 29026 8639 29041 8659
rect 28997 8633 29041 8639
rect 29091 8663 29140 8675
rect 29091 8643 29109 8663
rect 29129 8643 29140 8663
rect 29091 8633 29140 8643
rect 29215 8659 29259 8675
rect 29215 8639 29224 8659
rect 29244 8639 29259 8659
rect 29215 8633 29259 8639
rect 29309 8663 29358 8675
rect 29309 8643 29327 8663
rect 29347 8643 29358 8663
rect 29309 8633 29358 8643
rect 33148 8676 33197 8688
rect 33148 8656 33159 8676
rect 33179 8656 33197 8676
rect 33148 8646 33197 8656
rect 33247 8672 33291 8688
rect 33247 8652 33262 8672
rect 33282 8652 33291 8672
rect 33247 8646 33291 8652
rect 33361 8672 33405 8688
rect 33361 8652 33370 8672
rect 33390 8652 33405 8672
rect 33361 8646 33405 8652
rect 33455 8676 33504 8688
rect 33455 8656 33473 8676
rect 33493 8656 33504 8676
rect 33455 8646 33504 8656
rect 33579 8672 33623 8688
rect 33579 8652 33588 8672
rect 33608 8652 33623 8672
rect 33579 8646 33623 8652
rect 33673 8676 33722 8688
rect 33673 8656 33691 8676
rect 33711 8656 33722 8676
rect 33673 8646 33722 8656
rect 12211 8467 12260 8479
rect 12211 8447 12222 8467
rect 12242 8447 12260 8467
rect 9157 8417 9206 8427
rect 9157 8397 9168 8417
rect 9188 8397 9206 8417
rect 9157 8385 9206 8397
rect 9256 8421 9300 8427
rect 9256 8401 9271 8421
rect 9291 8401 9300 8421
rect 9256 8385 9300 8401
rect 9375 8417 9424 8427
rect 9375 8397 9386 8417
rect 9406 8397 9424 8417
rect 9375 8385 9424 8397
rect 9474 8421 9518 8427
rect 9474 8401 9489 8421
rect 9509 8401 9518 8421
rect 9474 8385 9518 8401
rect 9588 8421 9632 8427
rect 9588 8401 9597 8421
rect 9617 8401 9632 8421
rect 9588 8385 9632 8401
rect 9682 8417 9731 8427
rect 12211 8437 12260 8447
rect 12310 8463 12354 8479
rect 12310 8443 12325 8463
rect 12345 8443 12354 8463
rect 12310 8437 12354 8443
rect 12424 8463 12468 8479
rect 12424 8443 12433 8463
rect 12453 8443 12468 8463
rect 12424 8437 12468 8443
rect 12518 8467 12567 8479
rect 12518 8447 12536 8467
rect 12556 8447 12567 8467
rect 12518 8437 12567 8447
rect 12642 8463 12686 8479
rect 12642 8443 12651 8463
rect 12671 8443 12686 8463
rect 12642 8437 12686 8443
rect 12736 8467 12785 8479
rect 12736 8447 12754 8467
rect 12774 8447 12785 8467
rect 12736 8437 12785 8447
rect 9682 8397 9700 8417
rect 9720 8397 9731 8417
rect 9682 8385 9731 8397
rect 1214 8208 1263 8218
rect 1214 8188 1225 8208
rect 1245 8188 1263 8208
rect 1214 8176 1263 8188
rect 1313 8212 1357 8218
rect 1313 8192 1328 8212
rect 1348 8192 1357 8212
rect 1313 8176 1357 8192
rect 1432 8208 1481 8218
rect 1432 8188 1443 8208
rect 1463 8188 1481 8208
rect 1432 8176 1481 8188
rect 1531 8212 1575 8218
rect 1531 8192 1546 8212
rect 1566 8192 1575 8212
rect 1531 8176 1575 8192
rect 1645 8212 1689 8218
rect 1645 8192 1654 8212
rect 1674 8192 1689 8212
rect 1645 8176 1689 8192
rect 1739 8208 1788 8218
rect 1739 8188 1757 8208
rect 1777 8188 1788 8208
rect 1739 8176 1788 8188
rect 2573 8216 2622 8228
rect 2573 8196 2584 8216
rect 2604 8196 2622 8216
rect 2573 8186 2622 8196
rect 2672 8212 2716 8228
rect 2672 8192 2687 8212
rect 2707 8192 2716 8212
rect 2672 8186 2716 8192
rect 2786 8212 2830 8228
rect 2786 8192 2795 8212
rect 2815 8192 2830 8212
rect 2786 8186 2830 8192
rect 2880 8216 2929 8228
rect 2880 8196 2898 8216
rect 2918 8196 2929 8216
rect 2880 8186 2929 8196
rect 3004 8212 3048 8228
rect 3004 8192 3013 8212
rect 3033 8192 3048 8212
rect 3004 8186 3048 8192
rect 3098 8216 3147 8228
rect 16575 8480 16624 8492
rect 16575 8460 16586 8480
rect 16606 8460 16624 8480
rect 13521 8430 13570 8440
rect 13521 8410 13532 8430
rect 13552 8410 13570 8430
rect 13521 8398 13570 8410
rect 13620 8434 13664 8440
rect 13620 8414 13635 8434
rect 13655 8414 13664 8434
rect 13620 8398 13664 8414
rect 13739 8430 13788 8440
rect 13739 8410 13750 8430
rect 13770 8410 13788 8430
rect 13739 8398 13788 8410
rect 13838 8434 13882 8440
rect 13838 8414 13853 8434
rect 13873 8414 13882 8434
rect 13838 8398 13882 8414
rect 13952 8434 13996 8440
rect 13952 8414 13961 8434
rect 13981 8414 13996 8434
rect 13952 8398 13996 8414
rect 14046 8430 14095 8440
rect 16575 8450 16624 8460
rect 16674 8476 16718 8492
rect 16674 8456 16689 8476
rect 16709 8456 16718 8476
rect 16674 8450 16718 8456
rect 16788 8476 16832 8492
rect 16788 8456 16797 8476
rect 16817 8456 16832 8476
rect 16788 8450 16832 8456
rect 16882 8480 16931 8492
rect 16882 8460 16900 8480
rect 16920 8460 16931 8480
rect 16882 8450 16931 8460
rect 17006 8476 17050 8492
rect 17006 8456 17015 8476
rect 17035 8456 17050 8476
rect 17006 8450 17050 8456
rect 17100 8480 17149 8492
rect 17100 8460 17118 8480
rect 17138 8460 17149 8480
rect 17100 8450 17149 8460
rect 14046 8410 14064 8430
rect 14084 8410 14095 8430
rect 14046 8398 14095 8410
rect 3098 8196 3116 8216
rect 3136 8196 3147 8216
rect 3098 8186 3147 8196
rect 5578 8221 5627 8231
rect 5578 8201 5589 8221
rect 5609 8201 5627 8221
rect 5578 8189 5627 8201
rect 5677 8225 5721 8231
rect 5677 8205 5692 8225
rect 5712 8205 5721 8225
rect 5677 8189 5721 8205
rect 5796 8221 5845 8231
rect 5796 8201 5807 8221
rect 5827 8201 5845 8221
rect 5796 8189 5845 8201
rect 5895 8225 5939 8231
rect 5895 8205 5910 8225
rect 5930 8205 5939 8225
rect 5895 8189 5939 8205
rect 6009 8225 6053 8231
rect 6009 8205 6018 8225
rect 6038 8205 6053 8225
rect 6009 8189 6053 8205
rect 6103 8221 6152 8231
rect 6103 8201 6121 8221
rect 6141 8201 6152 8221
rect 6103 8189 6152 8201
rect 6937 8229 6986 8241
rect 6937 8209 6948 8229
rect 6968 8209 6986 8229
rect 6937 8199 6986 8209
rect 7036 8225 7080 8241
rect 7036 8205 7051 8225
rect 7071 8205 7080 8225
rect 7036 8199 7080 8205
rect 7150 8225 7194 8241
rect 7150 8205 7159 8225
rect 7179 8205 7194 8225
rect 7150 8199 7194 8205
rect 7244 8229 7293 8241
rect 7244 8209 7262 8229
rect 7282 8209 7293 8229
rect 7244 8199 7293 8209
rect 7368 8225 7412 8241
rect 7368 8205 7377 8225
rect 7397 8205 7412 8225
rect 7368 8199 7412 8205
rect 7462 8229 7511 8241
rect 20841 8454 20890 8466
rect 20841 8434 20852 8454
rect 20872 8434 20890 8454
rect 7462 8209 7480 8229
rect 7500 8209 7511 8229
rect 7462 8199 7511 8209
rect 9955 8233 10004 8243
rect 9955 8213 9966 8233
rect 9986 8213 10004 8233
rect 9955 8201 10004 8213
rect 10054 8237 10098 8243
rect 10054 8217 10069 8237
rect 10089 8217 10098 8237
rect 10054 8201 10098 8217
rect 10173 8233 10222 8243
rect 10173 8213 10184 8233
rect 10204 8213 10222 8233
rect 10173 8201 10222 8213
rect 10272 8237 10316 8243
rect 10272 8217 10287 8237
rect 10307 8217 10316 8237
rect 10272 8201 10316 8217
rect 10386 8237 10430 8243
rect 10386 8217 10395 8237
rect 10415 8217 10430 8237
rect 10386 8201 10430 8217
rect 10480 8233 10529 8243
rect 10480 8213 10498 8233
rect 10518 8213 10529 8233
rect 10480 8201 10529 8213
rect 11314 8241 11363 8253
rect 11314 8221 11325 8241
rect 11345 8221 11363 8241
rect 11314 8211 11363 8221
rect 11413 8237 11457 8253
rect 11413 8217 11428 8237
rect 11448 8217 11457 8237
rect 11413 8211 11457 8217
rect 11527 8237 11571 8253
rect 11527 8217 11536 8237
rect 11556 8217 11571 8237
rect 11527 8211 11571 8217
rect 11621 8241 11670 8253
rect 11621 8221 11639 8241
rect 11659 8221 11670 8241
rect 11621 8211 11670 8221
rect 11745 8237 11789 8253
rect 11745 8217 11754 8237
rect 11774 8217 11789 8237
rect 11745 8211 11789 8217
rect 11839 8241 11888 8253
rect 17787 8404 17836 8414
rect 17787 8384 17798 8404
rect 17818 8384 17836 8404
rect 17787 8372 17836 8384
rect 17886 8408 17930 8414
rect 17886 8388 17901 8408
rect 17921 8388 17930 8408
rect 17886 8372 17930 8388
rect 18005 8404 18054 8414
rect 18005 8384 18016 8404
rect 18036 8384 18054 8404
rect 18005 8372 18054 8384
rect 18104 8408 18148 8414
rect 18104 8388 18119 8408
rect 18139 8388 18148 8408
rect 18104 8372 18148 8388
rect 18218 8408 18262 8414
rect 18218 8388 18227 8408
rect 18247 8388 18262 8408
rect 18218 8372 18262 8388
rect 18312 8404 18361 8414
rect 20841 8424 20890 8434
rect 20940 8450 20984 8466
rect 20940 8430 20955 8450
rect 20975 8430 20984 8450
rect 20940 8424 20984 8430
rect 21054 8450 21098 8466
rect 21054 8430 21063 8450
rect 21083 8430 21098 8450
rect 21054 8424 21098 8430
rect 21148 8454 21197 8466
rect 21148 8434 21166 8454
rect 21186 8434 21197 8454
rect 21148 8424 21197 8434
rect 21272 8450 21316 8466
rect 21272 8430 21281 8450
rect 21301 8430 21316 8450
rect 21272 8424 21316 8430
rect 21366 8454 21415 8466
rect 21366 8434 21384 8454
rect 21404 8434 21415 8454
rect 21366 8424 21415 8434
rect 18312 8384 18330 8404
rect 18350 8384 18361 8404
rect 18312 8372 18361 8384
rect 25205 8467 25254 8479
rect 25205 8447 25216 8467
rect 25236 8447 25254 8467
rect 22151 8417 22200 8427
rect 22151 8397 22162 8417
rect 22182 8397 22200 8417
rect 22151 8385 22200 8397
rect 22250 8421 22294 8427
rect 22250 8401 22265 8421
rect 22285 8401 22294 8421
rect 22250 8385 22294 8401
rect 22369 8417 22418 8427
rect 22369 8397 22380 8417
rect 22400 8397 22418 8417
rect 22369 8385 22418 8397
rect 22468 8421 22512 8427
rect 22468 8401 22483 8421
rect 22503 8401 22512 8421
rect 22468 8385 22512 8401
rect 22582 8421 22626 8427
rect 22582 8401 22591 8421
rect 22611 8401 22626 8421
rect 22582 8385 22626 8401
rect 22676 8417 22725 8427
rect 25205 8437 25254 8447
rect 25304 8463 25348 8479
rect 25304 8443 25319 8463
rect 25339 8443 25348 8463
rect 25304 8437 25348 8443
rect 25418 8463 25462 8479
rect 25418 8443 25427 8463
rect 25447 8443 25462 8463
rect 25418 8437 25462 8443
rect 25512 8467 25561 8479
rect 25512 8447 25530 8467
rect 25550 8447 25561 8467
rect 25512 8437 25561 8447
rect 25636 8463 25680 8479
rect 25636 8443 25645 8463
rect 25665 8443 25680 8463
rect 25636 8437 25680 8443
rect 25730 8467 25779 8479
rect 25730 8447 25748 8467
rect 25768 8447 25779 8467
rect 25730 8437 25779 8447
rect 22676 8397 22694 8417
rect 22714 8397 22725 8417
rect 22676 8385 22725 8397
rect 11839 8221 11857 8241
rect 11877 8221 11888 8241
rect 11839 8211 11888 8221
rect 14319 8246 14368 8256
rect 14319 8226 14330 8246
rect 14350 8226 14368 8246
rect 417 7980 466 7990
rect 417 7960 428 7980
rect 448 7960 466 7980
rect 417 7948 466 7960
rect 516 7984 560 7990
rect 516 7964 531 7984
rect 551 7964 560 7984
rect 516 7948 560 7964
rect 635 7980 684 7990
rect 635 7960 646 7980
rect 666 7960 684 7980
rect 635 7948 684 7960
rect 734 7984 778 7990
rect 734 7964 749 7984
rect 769 7964 778 7984
rect 734 7948 778 7964
rect 848 7984 892 7990
rect 848 7964 857 7984
rect 877 7964 892 7984
rect 848 7948 892 7964
rect 942 7980 991 7990
rect 942 7960 960 7980
rect 980 7960 991 7980
rect 14319 8214 14368 8226
rect 14418 8250 14462 8256
rect 14418 8230 14433 8250
rect 14453 8230 14462 8250
rect 14418 8214 14462 8230
rect 14537 8246 14586 8256
rect 14537 8226 14548 8246
rect 14568 8226 14586 8246
rect 14537 8214 14586 8226
rect 14636 8250 14680 8256
rect 14636 8230 14651 8250
rect 14671 8230 14680 8250
rect 14636 8214 14680 8230
rect 14750 8250 14794 8256
rect 14750 8230 14759 8250
rect 14779 8230 14794 8250
rect 14750 8214 14794 8230
rect 14844 8246 14893 8256
rect 14844 8226 14862 8246
rect 14882 8226 14893 8246
rect 14844 8214 14893 8226
rect 15678 8254 15727 8266
rect 15678 8234 15689 8254
rect 15709 8234 15727 8254
rect 15678 8224 15727 8234
rect 15777 8250 15821 8266
rect 15777 8230 15792 8250
rect 15812 8230 15821 8250
rect 15777 8224 15821 8230
rect 15891 8250 15935 8266
rect 15891 8230 15900 8250
rect 15920 8230 15935 8250
rect 15891 8224 15935 8230
rect 15985 8254 16034 8266
rect 15985 8234 16003 8254
rect 16023 8234 16034 8254
rect 15985 8224 16034 8234
rect 16109 8250 16153 8266
rect 16109 8230 16118 8250
rect 16138 8230 16153 8250
rect 16109 8224 16153 8230
rect 16203 8254 16252 8266
rect 16203 8234 16221 8254
rect 16241 8234 16252 8254
rect 16203 8224 16252 8234
rect 29582 8479 29631 8491
rect 29582 8459 29593 8479
rect 29613 8459 29631 8479
rect 26528 8429 26577 8439
rect 26528 8409 26539 8429
rect 26559 8409 26577 8429
rect 26528 8397 26577 8409
rect 26627 8433 26671 8439
rect 26627 8413 26642 8433
rect 26662 8413 26671 8433
rect 26627 8397 26671 8413
rect 26746 8429 26795 8439
rect 26746 8409 26757 8429
rect 26777 8409 26795 8429
rect 26746 8397 26795 8409
rect 26845 8433 26889 8439
rect 26845 8413 26860 8433
rect 26880 8413 26889 8433
rect 26845 8397 26889 8413
rect 26959 8433 27003 8439
rect 26959 8413 26968 8433
rect 26988 8413 27003 8433
rect 26959 8397 27003 8413
rect 27053 8429 27102 8439
rect 29582 8449 29631 8459
rect 29681 8475 29725 8491
rect 29681 8455 29696 8475
rect 29716 8455 29725 8475
rect 29681 8449 29725 8455
rect 29795 8475 29839 8491
rect 29795 8455 29804 8475
rect 29824 8455 29839 8475
rect 29795 8449 29839 8455
rect 29889 8479 29938 8491
rect 29889 8459 29907 8479
rect 29927 8459 29938 8479
rect 29889 8449 29938 8459
rect 30013 8475 30057 8491
rect 30013 8455 30022 8475
rect 30042 8455 30057 8475
rect 30013 8449 30057 8455
rect 30107 8479 30156 8491
rect 30107 8459 30125 8479
rect 30145 8459 30156 8479
rect 30107 8449 30156 8459
rect 27053 8409 27071 8429
rect 27091 8409 27102 8429
rect 27053 8397 27102 8409
rect 942 7948 991 7960
rect 4781 7993 4830 8003
rect 4781 7973 4792 7993
rect 4812 7973 4830 7993
rect 4781 7961 4830 7973
rect 4880 7997 4924 8003
rect 4880 7977 4895 7997
rect 4915 7977 4924 7997
rect 4880 7961 4924 7977
rect 4999 7993 5048 8003
rect 4999 7973 5010 7993
rect 5030 7973 5048 7993
rect 4999 7961 5048 7973
rect 5098 7997 5142 8003
rect 5098 7977 5113 7997
rect 5133 7977 5142 7997
rect 5098 7961 5142 7977
rect 5212 7997 5256 8003
rect 5212 7977 5221 7997
rect 5241 7977 5256 7997
rect 5212 7961 5256 7977
rect 5306 7993 5355 8003
rect 5306 7973 5324 7993
rect 5344 7973 5355 7993
rect 18585 8220 18634 8230
rect 18585 8200 18596 8220
rect 18616 8200 18634 8220
rect 18585 8188 18634 8200
rect 18684 8224 18728 8230
rect 18684 8204 18699 8224
rect 18719 8204 18728 8224
rect 18684 8188 18728 8204
rect 18803 8220 18852 8230
rect 18803 8200 18814 8220
rect 18834 8200 18852 8220
rect 18803 8188 18852 8200
rect 18902 8224 18946 8230
rect 18902 8204 18917 8224
rect 18937 8204 18946 8224
rect 18902 8188 18946 8204
rect 19016 8224 19060 8230
rect 19016 8204 19025 8224
rect 19045 8204 19060 8224
rect 19016 8188 19060 8204
rect 19110 8220 19159 8230
rect 19110 8200 19128 8220
rect 19148 8200 19159 8220
rect 19110 8188 19159 8200
rect 19944 8228 19993 8240
rect 19944 8208 19955 8228
rect 19975 8208 19993 8228
rect 19944 8198 19993 8208
rect 20043 8224 20087 8240
rect 20043 8204 20058 8224
rect 20078 8204 20087 8224
rect 20043 8198 20087 8204
rect 20157 8224 20201 8240
rect 20157 8204 20166 8224
rect 20186 8204 20201 8224
rect 20157 8198 20201 8204
rect 20251 8228 20300 8240
rect 20251 8208 20269 8228
rect 20289 8208 20300 8228
rect 20251 8198 20300 8208
rect 20375 8224 20419 8240
rect 20375 8204 20384 8224
rect 20404 8204 20419 8224
rect 20375 8198 20419 8204
rect 20469 8228 20518 8240
rect 33946 8492 33995 8504
rect 33946 8472 33957 8492
rect 33977 8472 33995 8492
rect 30892 8442 30941 8452
rect 30892 8422 30903 8442
rect 30923 8422 30941 8442
rect 30892 8410 30941 8422
rect 30991 8446 31035 8452
rect 30991 8426 31006 8446
rect 31026 8426 31035 8446
rect 30991 8410 31035 8426
rect 31110 8442 31159 8452
rect 31110 8422 31121 8442
rect 31141 8422 31159 8442
rect 31110 8410 31159 8422
rect 31209 8446 31253 8452
rect 31209 8426 31224 8446
rect 31244 8426 31253 8446
rect 31209 8410 31253 8426
rect 31323 8446 31367 8452
rect 31323 8426 31332 8446
rect 31352 8426 31367 8446
rect 31323 8410 31367 8426
rect 31417 8442 31466 8452
rect 33946 8462 33995 8472
rect 34045 8488 34089 8504
rect 34045 8468 34060 8488
rect 34080 8468 34089 8488
rect 34045 8462 34089 8468
rect 34159 8488 34203 8504
rect 34159 8468 34168 8488
rect 34188 8468 34203 8488
rect 34159 8462 34203 8468
rect 34253 8492 34302 8504
rect 34253 8472 34271 8492
rect 34291 8472 34302 8492
rect 34253 8462 34302 8472
rect 34377 8488 34421 8504
rect 34377 8468 34386 8488
rect 34406 8468 34421 8488
rect 34377 8462 34421 8468
rect 34471 8492 34520 8504
rect 34471 8472 34489 8492
rect 34509 8472 34520 8492
rect 34471 8462 34520 8472
rect 31417 8422 31435 8442
rect 31455 8422 31466 8442
rect 31417 8410 31466 8422
rect 20469 8208 20487 8228
rect 20507 8208 20518 8228
rect 20469 8198 20518 8208
rect 22949 8233 22998 8243
rect 22949 8213 22960 8233
rect 22980 8213 22998 8233
rect 5306 7961 5355 7973
rect 9158 8005 9207 8015
rect 9158 7985 9169 8005
rect 9189 7985 9207 8005
rect 9158 7973 9207 7985
rect 9257 8009 9301 8015
rect 9257 7989 9272 8009
rect 9292 7989 9301 8009
rect 9257 7973 9301 7989
rect 9376 8005 9425 8015
rect 9376 7985 9387 8005
rect 9407 7985 9425 8005
rect 9376 7973 9425 7985
rect 9475 8009 9519 8015
rect 9475 7989 9490 8009
rect 9510 7989 9519 8009
rect 9475 7973 9519 7989
rect 9589 8009 9633 8015
rect 9589 7989 9598 8009
rect 9618 7989 9633 8009
rect 9589 7973 9633 7989
rect 9683 8005 9732 8015
rect 9683 7985 9701 8005
rect 9721 7985 9732 8005
rect 22949 8201 22998 8213
rect 23048 8237 23092 8243
rect 23048 8217 23063 8237
rect 23083 8217 23092 8237
rect 23048 8201 23092 8217
rect 23167 8233 23216 8243
rect 23167 8213 23178 8233
rect 23198 8213 23216 8233
rect 23167 8201 23216 8213
rect 23266 8237 23310 8243
rect 23266 8217 23281 8237
rect 23301 8217 23310 8237
rect 23266 8201 23310 8217
rect 23380 8237 23424 8243
rect 23380 8217 23389 8237
rect 23409 8217 23424 8237
rect 23380 8201 23424 8217
rect 23474 8233 23523 8243
rect 23474 8213 23492 8233
rect 23512 8213 23523 8233
rect 23474 8201 23523 8213
rect 24308 8241 24357 8253
rect 24308 8221 24319 8241
rect 24339 8221 24357 8241
rect 24308 8211 24357 8221
rect 24407 8237 24451 8253
rect 24407 8217 24422 8237
rect 24442 8217 24451 8237
rect 24407 8211 24451 8217
rect 24521 8237 24565 8253
rect 24521 8217 24530 8237
rect 24550 8217 24565 8237
rect 24521 8211 24565 8217
rect 24615 8241 24664 8253
rect 24615 8221 24633 8241
rect 24653 8221 24664 8241
rect 24615 8211 24664 8221
rect 24739 8237 24783 8253
rect 24739 8217 24748 8237
rect 24768 8217 24783 8237
rect 24739 8211 24783 8217
rect 24833 8241 24882 8253
rect 24833 8221 24851 8241
rect 24871 8221 24882 8241
rect 24833 8211 24882 8221
rect 9683 7973 9732 7985
rect 13522 8018 13571 8028
rect 13522 7998 13533 8018
rect 13553 7998 13571 8018
rect 13522 7986 13571 7998
rect 13621 8022 13665 8028
rect 13621 8002 13636 8022
rect 13656 8002 13665 8022
rect 13621 7986 13665 8002
rect 13740 8018 13789 8028
rect 13740 7998 13751 8018
rect 13771 7998 13789 8018
rect 13740 7986 13789 7998
rect 13839 8022 13883 8028
rect 13839 8002 13854 8022
rect 13874 8002 13883 8022
rect 13839 7986 13883 8002
rect 13953 8022 13997 8028
rect 13953 8002 13962 8022
rect 13982 8002 13997 8022
rect 13953 7986 13997 8002
rect 14047 8018 14096 8028
rect 14047 7998 14065 8018
rect 14085 7998 14096 8018
rect 14047 7986 14096 7998
rect 27326 8245 27375 8255
rect 27326 8225 27337 8245
rect 27357 8225 27375 8245
rect 27326 8213 27375 8225
rect 27425 8249 27469 8255
rect 27425 8229 27440 8249
rect 27460 8229 27469 8249
rect 27425 8213 27469 8229
rect 27544 8245 27593 8255
rect 27544 8225 27555 8245
rect 27575 8225 27593 8245
rect 27544 8213 27593 8225
rect 27643 8249 27687 8255
rect 27643 8229 27658 8249
rect 27678 8229 27687 8249
rect 27643 8213 27687 8229
rect 27757 8249 27801 8255
rect 27757 8229 27766 8249
rect 27786 8229 27801 8249
rect 27757 8213 27801 8229
rect 27851 8245 27900 8255
rect 27851 8225 27869 8245
rect 27889 8225 27900 8245
rect 27851 8213 27900 8225
rect 28685 8253 28734 8265
rect 28685 8233 28696 8253
rect 28716 8233 28734 8253
rect 28685 8223 28734 8233
rect 28784 8249 28828 8265
rect 28784 8229 28799 8249
rect 28819 8229 28828 8249
rect 28784 8223 28828 8229
rect 28898 8249 28942 8265
rect 28898 8229 28907 8249
rect 28927 8229 28942 8249
rect 28898 8223 28942 8229
rect 28992 8253 29041 8265
rect 28992 8233 29010 8253
rect 29030 8233 29041 8253
rect 28992 8223 29041 8233
rect 29116 8249 29160 8265
rect 29116 8229 29125 8249
rect 29145 8229 29160 8249
rect 29116 8223 29160 8229
rect 29210 8253 29259 8265
rect 29210 8233 29228 8253
rect 29248 8233 29259 8253
rect 29210 8223 29259 8233
rect 31690 8258 31739 8268
rect 31690 8238 31701 8258
rect 31721 8238 31739 8258
rect 17788 7992 17837 8002
rect 17788 7972 17799 7992
rect 17819 7972 17837 7992
rect 17788 7960 17837 7972
rect 17887 7996 17931 8002
rect 17887 7976 17902 7996
rect 17922 7976 17931 7996
rect 17887 7960 17931 7976
rect 18006 7992 18055 8002
rect 18006 7972 18017 7992
rect 18037 7972 18055 7992
rect 18006 7960 18055 7972
rect 18105 7996 18149 8002
rect 18105 7976 18120 7996
rect 18140 7976 18149 7996
rect 18105 7960 18149 7976
rect 18219 7996 18263 8002
rect 18219 7976 18228 7996
rect 18248 7976 18263 7996
rect 18219 7960 18263 7976
rect 18313 7992 18362 8002
rect 18313 7972 18331 7992
rect 18351 7972 18362 7992
rect 31690 8226 31739 8238
rect 31789 8262 31833 8268
rect 31789 8242 31804 8262
rect 31824 8242 31833 8262
rect 31789 8226 31833 8242
rect 31908 8258 31957 8268
rect 31908 8238 31919 8258
rect 31939 8238 31957 8258
rect 31908 8226 31957 8238
rect 32007 8262 32051 8268
rect 32007 8242 32022 8262
rect 32042 8242 32051 8262
rect 32007 8226 32051 8242
rect 32121 8262 32165 8268
rect 32121 8242 32130 8262
rect 32150 8242 32165 8262
rect 32121 8226 32165 8242
rect 32215 8258 32264 8268
rect 32215 8238 32233 8258
rect 32253 8238 32264 8258
rect 32215 8226 32264 8238
rect 33049 8266 33098 8278
rect 33049 8246 33060 8266
rect 33080 8246 33098 8266
rect 33049 8236 33098 8246
rect 33148 8262 33192 8278
rect 33148 8242 33163 8262
rect 33183 8242 33192 8262
rect 33148 8236 33192 8242
rect 33262 8262 33306 8278
rect 33262 8242 33271 8262
rect 33291 8242 33306 8262
rect 33262 8236 33306 8242
rect 33356 8266 33405 8278
rect 33356 8246 33374 8266
rect 33394 8246 33405 8266
rect 33356 8236 33405 8246
rect 33480 8262 33524 8278
rect 33480 8242 33489 8262
rect 33509 8242 33524 8262
rect 33480 8236 33524 8242
rect 33574 8266 33623 8278
rect 33574 8246 33592 8266
rect 33612 8246 33623 8266
rect 33574 8236 33623 8246
rect 18313 7960 18362 7972
rect 22152 8005 22201 8015
rect 22152 7985 22163 8005
rect 22183 7985 22201 8005
rect 22152 7973 22201 7985
rect 22251 8009 22295 8015
rect 22251 7989 22266 8009
rect 22286 7989 22295 8009
rect 22251 7973 22295 7989
rect 22370 8005 22419 8015
rect 22370 7985 22381 8005
rect 22401 7985 22419 8005
rect 22370 7973 22419 7985
rect 22469 8009 22513 8015
rect 22469 7989 22484 8009
rect 22504 7989 22513 8009
rect 22469 7973 22513 7989
rect 22583 8009 22627 8015
rect 22583 7989 22592 8009
rect 22612 7989 22627 8009
rect 22583 7973 22627 7989
rect 22677 8005 22726 8015
rect 22677 7985 22695 8005
rect 22715 7985 22726 8005
rect 22677 7973 22726 7985
rect 26529 8017 26578 8027
rect 26529 7997 26540 8017
rect 26560 7997 26578 8017
rect 26529 7985 26578 7997
rect 26628 8021 26672 8027
rect 26628 8001 26643 8021
rect 26663 8001 26672 8021
rect 26628 7985 26672 8001
rect 26747 8017 26796 8027
rect 26747 7997 26758 8017
rect 26778 7997 26796 8017
rect 26747 7985 26796 7997
rect 26846 8021 26890 8027
rect 26846 8001 26861 8021
rect 26881 8001 26890 8021
rect 26846 7985 26890 8001
rect 26960 8021 27004 8027
rect 26960 8001 26969 8021
rect 26989 8001 27004 8021
rect 26960 7985 27004 8001
rect 27054 8017 27103 8027
rect 27054 7997 27072 8017
rect 27092 7997 27103 8017
rect 27054 7985 27103 7997
rect 30893 8030 30942 8040
rect 30893 8010 30904 8030
rect 30924 8010 30942 8030
rect 30893 7998 30942 8010
rect 30992 8034 31036 8040
rect 30992 8014 31007 8034
rect 31027 8014 31036 8034
rect 30992 7998 31036 8014
rect 31111 8030 31160 8040
rect 31111 8010 31122 8030
rect 31142 8010 31160 8030
rect 31111 7998 31160 8010
rect 31210 8034 31254 8040
rect 31210 8014 31225 8034
rect 31245 8014 31254 8034
rect 31210 7998 31254 8014
rect 31324 8034 31368 8040
rect 31324 8014 31333 8034
rect 31353 8014 31368 8034
rect 31324 7998 31368 8014
rect 31418 8030 31467 8040
rect 31418 8010 31436 8030
rect 31456 8010 31467 8030
rect 31418 7998 31467 8010
rect 3452 7836 3501 7848
rect 3452 7816 3463 7836
rect 3483 7816 3501 7836
rect 3452 7806 3501 7816
rect 3551 7832 3595 7848
rect 3551 7812 3566 7832
rect 3586 7812 3595 7832
rect 3551 7806 3595 7812
rect 3665 7832 3709 7848
rect 3665 7812 3674 7832
rect 3694 7812 3709 7832
rect 3665 7806 3709 7812
rect 3759 7836 3808 7848
rect 3759 7816 3777 7836
rect 3797 7816 3808 7836
rect 3759 7806 3808 7816
rect 3883 7832 3927 7848
rect 3883 7812 3892 7832
rect 3912 7812 3927 7832
rect 3883 7806 3927 7812
rect 3977 7836 4026 7848
rect 3977 7816 3995 7836
rect 4015 7816 4026 7836
rect 3977 7806 4026 7816
rect 7816 7849 7865 7861
rect 7816 7829 7827 7849
rect 7847 7829 7865 7849
rect 7816 7819 7865 7829
rect 7915 7845 7959 7861
rect 7915 7825 7930 7845
rect 7950 7825 7959 7845
rect 7915 7819 7959 7825
rect 8029 7845 8073 7861
rect 8029 7825 8038 7845
rect 8058 7825 8073 7845
rect 8029 7819 8073 7825
rect 8123 7849 8172 7861
rect 8123 7829 8141 7849
rect 8161 7829 8172 7849
rect 8123 7819 8172 7829
rect 8247 7845 8291 7861
rect 8247 7825 8256 7845
rect 8276 7825 8291 7845
rect 8247 7819 8291 7825
rect 8341 7849 8390 7861
rect 8341 7829 8359 7849
rect 8379 7829 8390 7849
rect 8341 7819 8390 7829
rect 12193 7861 12242 7873
rect 12193 7841 12204 7861
rect 12224 7841 12242 7861
rect 12193 7831 12242 7841
rect 12292 7857 12336 7873
rect 12292 7837 12307 7857
rect 12327 7837 12336 7857
rect 12292 7831 12336 7837
rect 12406 7857 12450 7873
rect 12406 7837 12415 7857
rect 12435 7837 12450 7857
rect 12406 7831 12450 7837
rect 12500 7861 12549 7873
rect 12500 7841 12518 7861
rect 12538 7841 12549 7861
rect 12500 7831 12549 7841
rect 12624 7857 12668 7873
rect 12624 7837 12633 7857
rect 12653 7837 12668 7857
rect 12624 7831 12668 7837
rect 12718 7861 12767 7873
rect 12718 7841 12736 7861
rect 12756 7841 12767 7861
rect 12718 7831 12767 7841
rect 16557 7874 16606 7886
rect 1296 7600 1345 7610
rect 1296 7580 1307 7600
rect 1327 7580 1345 7600
rect 1296 7568 1345 7580
rect 1395 7604 1439 7610
rect 1395 7584 1410 7604
rect 1430 7584 1439 7604
rect 1395 7568 1439 7584
rect 1514 7600 1563 7610
rect 1514 7580 1525 7600
rect 1545 7580 1563 7600
rect 1514 7568 1563 7580
rect 1613 7604 1657 7610
rect 1613 7584 1628 7604
rect 1648 7584 1657 7604
rect 1613 7568 1657 7584
rect 1727 7604 1771 7610
rect 1727 7584 1736 7604
rect 1756 7584 1771 7604
rect 1727 7568 1771 7584
rect 1821 7600 1870 7610
rect 1821 7580 1839 7600
rect 1859 7580 1870 7600
rect 1821 7568 1870 7580
rect 2655 7608 2704 7620
rect 2655 7588 2666 7608
rect 2686 7588 2704 7608
rect 2655 7578 2704 7588
rect 2754 7604 2798 7620
rect 2754 7584 2769 7604
rect 2789 7584 2798 7604
rect 2754 7578 2798 7584
rect 2868 7604 2912 7620
rect 2868 7584 2877 7604
rect 2897 7584 2912 7604
rect 2868 7578 2912 7584
rect 2962 7608 3011 7620
rect 2962 7588 2980 7608
rect 3000 7588 3011 7608
rect 2962 7578 3011 7588
rect 3086 7604 3130 7620
rect 3086 7584 3095 7604
rect 3115 7584 3130 7604
rect 3086 7578 3130 7584
rect 3180 7608 3229 7620
rect 16557 7854 16568 7874
rect 16588 7854 16606 7874
rect 16557 7844 16606 7854
rect 16656 7870 16700 7886
rect 16656 7850 16671 7870
rect 16691 7850 16700 7870
rect 16656 7844 16700 7850
rect 16770 7870 16814 7886
rect 16770 7850 16779 7870
rect 16799 7850 16814 7870
rect 16770 7844 16814 7850
rect 16864 7874 16913 7886
rect 16864 7854 16882 7874
rect 16902 7854 16913 7874
rect 16864 7844 16913 7854
rect 16988 7870 17032 7886
rect 16988 7850 16997 7870
rect 17017 7850 17032 7870
rect 16988 7844 17032 7850
rect 17082 7874 17131 7886
rect 17082 7854 17100 7874
rect 17120 7854 17131 7874
rect 17082 7844 17131 7854
rect 3180 7588 3198 7608
rect 3218 7588 3229 7608
rect 3180 7578 3229 7588
rect 5660 7613 5709 7623
rect 5660 7593 5671 7613
rect 5691 7593 5709 7613
rect 5660 7581 5709 7593
rect 5759 7617 5803 7623
rect 5759 7597 5774 7617
rect 5794 7597 5803 7617
rect 5759 7581 5803 7597
rect 5878 7613 5927 7623
rect 5878 7593 5889 7613
rect 5909 7593 5927 7613
rect 5878 7581 5927 7593
rect 5977 7617 6021 7623
rect 5977 7597 5992 7617
rect 6012 7597 6021 7617
rect 5977 7581 6021 7597
rect 6091 7617 6135 7623
rect 6091 7597 6100 7617
rect 6120 7597 6135 7617
rect 6091 7581 6135 7597
rect 6185 7613 6234 7623
rect 6185 7593 6203 7613
rect 6223 7593 6234 7613
rect 6185 7581 6234 7593
rect 7019 7621 7068 7633
rect 7019 7601 7030 7621
rect 7050 7601 7068 7621
rect 7019 7591 7068 7601
rect 7118 7617 7162 7633
rect 7118 7597 7133 7617
rect 7153 7597 7162 7617
rect 7118 7591 7162 7597
rect 7232 7617 7276 7633
rect 7232 7597 7241 7617
rect 7261 7597 7276 7617
rect 7232 7591 7276 7597
rect 7326 7621 7375 7633
rect 7326 7601 7344 7621
rect 7364 7601 7375 7621
rect 7326 7591 7375 7601
rect 7450 7617 7494 7633
rect 7450 7597 7459 7617
rect 7479 7597 7494 7617
rect 7450 7591 7494 7597
rect 7544 7621 7593 7633
rect 7544 7601 7562 7621
rect 7582 7601 7593 7621
rect 7544 7591 7593 7601
rect 20823 7848 20872 7860
rect 20823 7828 20834 7848
rect 20854 7828 20872 7848
rect 20823 7818 20872 7828
rect 20922 7844 20966 7860
rect 20922 7824 20937 7844
rect 20957 7824 20966 7844
rect 20922 7818 20966 7824
rect 21036 7844 21080 7860
rect 21036 7824 21045 7844
rect 21065 7824 21080 7844
rect 21036 7818 21080 7824
rect 21130 7848 21179 7860
rect 21130 7828 21148 7848
rect 21168 7828 21179 7848
rect 21130 7818 21179 7828
rect 21254 7844 21298 7860
rect 21254 7824 21263 7844
rect 21283 7824 21298 7844
rect 21254 7818 21298 7824
rect 21348 7848 21397 7860
rect 21348 7828 21366 7848
rect 21386 7828 21397 7848
rect 21348 7818 21397 7828
rect 25187 7861 25236 7873
rect 10037 7625 10086 7635
rect 10037 7605 10048 7625
rect 10068 7605 10086 7625
rect 10037 7593 10086 7605
rect 10136 7629 10180 7635
rect 10136 7609 10151 7629
rect 10171 7609 10180 7629
rect 10136 7593 10180 7609
rect 10255 7625 10304 7635
rect 10255 7605 10266 7625
rect 10286 7605 10304 7625
rect 10255 7593 10304 7605
rect 10354 7629 10398 7635
rect 10354 7609 10369 7629
rect 10389 7609 10398 7629
rect 10354 7593 10398 7609
rect 10468 7629 10512 7635
rect 10468 7609 10477 7629
rect 10497 7609 10512 7629
rect 10468 7593 10512 7609
rect 10562 7625 10611 7635
rect 10562 7605 10580 7625
rect 10600 7605 10611 7625
rect 10562 7593 10611 7605
rect 11396 7633 11445 7645
rect 11396 7613 11407 7633
rect 11427 7613 11445 7633
rect 11396 7603 11445 7613
rect 11495 7629 11539 7645
rect 11495 7609 11510 7629
rect 11530 7609 11539 7629
rect 11495 7603 11539 7609
rect 11609 7629 11653 7645
rect 11609 7609 11618 7629
rect 11638 7609 11653 7629
rect 11609 7603 11653 7609
rect 11703 7633 11752 7645
rect 11703 7613 11721 7633
rect 11741 7613 11752 7633
rect 11703 7603 11752 7613
rect 11827 7629 11871 7645
rect 11827 7609 11836 7629
rect 11856 7609 11871 7629
rect 11827 7603 11871 7609
rect 11921 7633 11970 7645
rect 25187 7841 25198 7861
rect 25218 7841 25236 7861
rect 25187 7831 25236 7841
rect 25286 7857 25330 7873
rect 25286 7837 25301 7857
rect 25321 7837 25330 7857
rect 25286 7831 25330 7837
rect 25400 7857 25444 7873
rect 25400 7837 25409 7857
rect 25429 7837 25444 7857
rect 25400 7831 25444 7837
rect 25494 7861 25543 7873
rect 25494 7841 25512 7861
rect 25532 7841 25543 7861
rect 25494 7831 25543 7841
rect 25618 7857 25662 7873
rect 25618 7837 25627 7857
rect 25647 7837 25662 7857
rect 25618 7831 25662 7837
rect 25712 7861 25761 7873
rect 25712 7841 25730 7861
rect 25750 7841 25761 7861
rect 25712 7831 25761 7841
rect 29564 7873 29613 7885
rect 11921 7613 11939 7633
rect 11959 7613 11970 7633
rect 11921 7603 11970 7613
rect 14401 7638 14450 7648
rect 14401 7618 14412 7638
rect 14432 7618 14450 7638
rect 3453 7424 3502 7436
rect 3453 7404 3464 7424
rect 3484 7404 3502 7424
rect 399 7374 448 7384
rect 399 7354 410 7374
rect 430 7354 448 7374
rect 399 7342 448 7354
rect 498 7378 542 7384
rect 498 7358 513 7378
rect 533 7358 542 7378
rect 498 7342 542 7358
rect 617 7374 666 7384
rect 617 7354 628 7374
rect 648 7354 666 7374
rect 617 7342 666 7354
rect 716 7378 760 7384
rect 716 7358 731 7378
rect 751 7358 760 7378
rect 716 7342 760 7358
rect 830 7378 874 7384
rect 830 7358 839 7378
rect 859 7358 874 7378
rect 830 7342 874 7358
rect 924 7374 973 7384
rect 3453 7394 3502 7404
rect 3552 7420 3596 7436
rect 3552 7400 3567 7420
rect 3587 7400 3596 7420
rect 3552 7394 3596 7400
rect 3666 7420 3710 7436
rect 3666 7400 3675 7420
rect 3695 7400 3710 7420
rect 3666 7394 3710 7400
rect 3760 7424 3809 7436
rect 3760 7404 3778 7424
rect 3798 7404 3809 7424
rect 3760 7394 3809 7404
rect 3884 7420 3928 7436
rect 3884 7400 3893 7420
rect 3913 7400 3928 7420
rect 3884 7394 3928 7400
rect 3978 7424 4027 7436
rect 3978 7404 3996 7424
rect 4016 7404 4027 7424
rect 3978 7394 4027 7404
rect 924 7354 942 7374
rect 962 7354 973 7374
rect 924 7342 973 7354
rect 14401 7606 14450 7618
rect 14500 7642 14544 7648
rect 14500 7622 14515 7642
rect 14535 7622 14544 7642
rect 14500 7606 14544 7622
rect 14619 7638 14668 7648
rect 14619 7618 14630 7638
rect 14650 7618 14668 7638
rect 14619 7606 14668 7618
rect 14718 7642 14762 7648
rect 14718 7622 14733 7642
rect 14753 7622 14762 7642
rect 14718 7606 14762 7622
rect 14832 7642 14876 7648
rect 14832 7622 14841 7642
rect 14861 7622 14876 7642
rect 14832 7606 14876 7622
rect 14926 7638 14975 7648
rect 14926 7618 14944 7638
rect 14964 7618 14975 7638
rect 14926 7606 14975 7618
rect 15760 7646 15809 7658
rect 15760 7626 15771 7646
rect 15791 7626 15809 7646
rect 15760 7616 15809 7626
rect 15859 7642 15903 7658
rect 15859 7622 15874 7642
rect 15894 7622 15903 7642
rect 15859 7616 15903 7622
rect 15973 7642 16017 7658
rect 15973 7622 15982 7642
rect 16002 7622 16017 7642
rect 15973 7616 16017 7622
rect 16067 7646 16116 7658
rect 16067 7626 16085 7646
rect 16105 7626 16116 7646
rect 16067 7616 16116 7626
rect 16191 7642 16235 7658
rect 16191 7622 16200 7642
rect 16220 7622 16235 7642
rect 16191 7616 16235 7622
rect 16285 7646 16334 7658
rect 16285 7626 16303 7646
rect 16323 7626 16334 7646
rect 16285 7616 16334 7626
rect 29564 7853 29575 7873
rect 29595 7853 29613 7873
rect 29564 7843 29613 7853
rect 29663 7869 29707 7885
rect 29663 7849 29678 7869
rect 29698 7849 29707 7869
rect 29663 7843 29707 7849
rect 29777 7869 29821 7885
rect 29777 7849 29786 7869
rect 29806 7849 29821 7869
rect 29777 7843 29821 7849
rect 29871 7873 29920 7885
rect 29871 7853 29889 7873
rect 29909 7853 29920 7873
rect 29871 7843 29920 7853
rect 29995 7869 30039 7885
rect 29995 7849 30004 7869
rect 30024 7849 30039 7869
rect 29995 7843 30039 7849
rect 30089 7873 30138 7885
rect 30089 7853 30107 7873
rect 30127 7853 30138 7873
rect 30089 7843 30138 7853
rect 33928 7886 33977 7898
rect 7817 7437 7866 7449
rect 7817 7417 7828 7437
rect 7848 7417 7866 7437
rect 4763 7387 4812 7397
rect 4763 7367 4774 7387
rect 4794 7367 4812 7387
rect 4763 7355 4812 7367
rect 4862 7391 4906 7397
rect 4862 7371 4877 7391
rect 4897 7371 4906 7391
rect 4862 7355 4906 7371
rect 4981 7387 5030 7397
rect 4981 7367 4992 7387
rect 5012 7367 5030 7387
rect 4981 7355 5030 7367
rect 5080 7391 5124 7397
rect 5080 7371 5095 7391
rect 5115 7371 5124 7391
rect 5080 7355 5124 7371
rect 5194 7391 5238 7397
rect 5194 7371 5203 7391
rect 5223 7371 5238 7391
rect 5194 7355 5238 7371
rect 5288 7387 5337 7397
rect 7817 7407 7866 7417
rect 7916 7433 7960 7449
rect 7916 7413 7931 7433
rect 7951 7413 7960 7433
rect 7916 7407 7960 7413
rect 8030 7433 8074 7449
rect 8030 7413 8039 7433
rect 8059 7413 8074 7433
rect 8030 7407 8074 7413
rect 8124 7437 8173 7449
rect 8124 7417 8142 7437
rect 8162 7417 8173 7437
rect 8124 7407 8173 7417
rect 8248 7433 8292 7449
rect 8248 7413 8257 7433
rect 8277 7413 8292 7433
rect 8248 7407 8292 7413
rect 8342 7437 8391 7449
rect 8342 7417 8360 7437
rect 8380 7417 8391 7437
rect 8342 7407 8391 7417
rect 5288 7367 5306 7387
rect 5326 7367 5337 7387
rect 5288 7355 5337 7367
rect 18667 7612 18716 7622
rect 18667 7592 18678 7612
rect 18698 7592 18716 7612
rect 18667 7580 18716 7592
rect 18766 7616 18810 7622
rect 18766 7596 18781 7616
rect 18801 7596 18810 7616
rect 18766 7580 18810 7596
rect 18885 7612 18934 7622
rect 18885 7592 18896 7612
rect 18916 7592 18934 7612
rect 18885 7580 18934 7592
rect 18984 7616 19028 7622
rect 18984 7596 18999 7616
rect 19019 7596 19028 7616
rect 18984 7580 19028 7596
rect 19098 7616 19142 7622
rect 19098 7596 19107 7616
rect 19127 7596 19142 7616
rect 19098 7580 19142 7596
rect 19192 7612 19241 7622
rect 19192 7592 19210 7612
rect 19230 7592 19241 7612
rect 19192 7580 19241 7592
rect 20026 7620 20075 7632
rect 20026 7600 20037 7620
rect 20057 7600 20075 7620
rect 20026 7590 20075 7600
rect 20125 7616 20169 7632
rect 20125 7596 20140 7616
rect 20160 7596 20169 7616
rect 20125 7590 20169 7596
rect 20239 7616 20283 7632
rect 20239 7596 20248 7616
rect 20268 7596 20283 7616
rect 20239 7590 20283 7596
rect 20333 7620 20382 7632
rect 20333 7600 20351 7620
rect 20371 7600 20382 7620
rect 20333 7590 20382 7600
rect 20457 7616 20501 7632
rect 20457 7596 20466 7616
rect 20486 7596 20501 7616
rect 20457 7590 20501 7596
rect 20551 7620 20600 7632
rect 33928 7866 33939 7886
rect 33959 7866 33977 7886
rect 33928 7856 33977 7866
rect 34027 7882 34071 7898
rect 34027 7862 34042 7882
rect 34062 7862 34071 7882
rect 34027 7856 34071 7862
rect 34141 7882 34185 7898
rect 34141 7862 34150 7882
rect 34170 7862 34185 7882
rect 34141 7856 34185 7862
rect 34235 7886 34284 7898
rect 34235 7866 34253 7886
rect 34273 7866 34284 7886
rect 34235 7856 34284 7866
rect 34359 7882 34403 7898
rect 34359 7862 34368 7882
rect 34388 7862 34403 7882
rect 34359 7856 34403 7862
rect 34453 7886 34502 7898
rect 34453 7866 34471 7886
rect 34491 7866 34502 7886
rect 34453 7856 34502 7866
rect 20551 7600 20569 7620
rect 20589 7600 20600 7620
rect 20551 7590 20600 7600
rect 23031 7625 23080 7635
rect 23031 7605 23042 7625
rect 23062 7605 23080 7625
rect 12194 7449 12243 7461
rect 12194 7429 12205 7449
rect 12225 7429 12243 7449
rect 9140 7399 9189 7409
rect 9140 7379 9151 7399
rect 9171 7379 9189 7399
rect 9140 7367 9189 7379
rect 9239 7403 9283 7409
rect 9239 7383 9254 7403
rect 9274 7383 9283 7403
rect 9239 7367 9283 7383
rect 9358 7399 9407 7409
rect 9358 7379 9369 7399
rect 9389 7379 9407 7399
rect 9358 7367 9407 7379
rect 9457 7403 9501 7409
rect 9457 7383 9472 7403
rect 9492 7383 9501 7403
rect 9457 7367 9501 7383
rect 9571 7403 9615 7409
rect 9571 7383 9580 7403
rect 9600 7383 9615 7403
rect 9571 7367 9615 7383
rect 9665 7399 9714 7409
rect 12194 7419 12243 7429
rect 12293 7445 12337 7461
rect 12293 7425 12308 7445
rect 12328 7425 12337 7445
rect 12293 7419 12337 7425
rect 12407 7445 12451 7461
rect 12407 7425 12416 7445
rect 12436 7425 12451 7445
rect 12407 7419 12451 7425
rect 12501 7449 12550 7461
rect 12501 7429 12519 7449
rect 12539 7429 12550 7449
rect 12501 7419 12550 7429
rect 12625 7445 12669 7461
rect 12625 7425 12634 7445
rect 12654 7425 12669 7445
rect 12625 7419 12669 7425
rect 12719 7449 12768 7461
rect 12719 7429 12737 7449
rect 12757 7429 12768 7449
rect 12719 7419 12768 7429
rect 9665 7379 9683 7399
rect 9703 7379 9714 7399
rect 9665 7367 9714 7379
rect 2490 7200 2539 7212
rect 1197 7190 1246 7200
rect 1197 7170 1208 7190
rect 1228 7170 1246 7190
rect 1197 7158 1246 7170
rect 1296 7194 1340 7200
rect 1296 7174 1311 7194
rect 1331 7174 1340 7194
rect 1296 7158 1340 7174
rect 1415 7190 1464 7200
rect 1415 7170 1426 7190
rect 1446 7170 1464 7190
rect 1415 7158 1464 7170
rect 1514 7194 1558 7200
rect 1514 7174 1529 7194
rect 1549 7174 1558 7194
rect 1514 7158 1558 7174
rect 1628 7194 1672 7200
rect 1628 7174 1637 7194
rect 1657 7174 1672 7194
rect 1628 7158 1672 7174
rect 1722 7190 1771 7200
rect 1722 7170 1740 7190
rect 1760 7170 1771 7190
rect 2490 7180 2501 7200
rect 2521 7180 2539 7200
rect 2490 7170 2539 7180
rect 2589 7196 2633 7212
rect 2589 7176 2604 7196
rect 2624 7176 2633 7196
rect 2589 7170 2633 7176
rect 2703 7196 2747 7212
rect 2703 7176 2712 7196
rect 2732 7176 2747 7196
rect 2703 7170 2747 7176
rect 2797 7200 2846 7212
rect 2797 7180 2815 7200
rect 2835 7180 2846 7200
rect 2797 7170 2846 7180
rect 2921 7196 2965 7212
rect 2921 7176 2930 7196
rect 2950 7176 2965 7196
rect 2921 7170 2965 7176
rect 3015 7200 3064 7212
rect 16558 7462 16607 7474
rect 16558 7442 16569 7462
rect 16589 7442 16607 7462
rect 13504 7412 13553 7422
rect 13504 7392 13515 7412
rect 13535 7392 13553 7412
rect 13504 7380 13553 7392
rect 13603 7416 13647 7422
rect 13603 7396 13618 7416
rect 13638 7396 13647 7416
rect 13603 7380 13647 7396
rect 13722 7412 13771 7422
rect 13722 7392 13733 7412
rect 13753 7392 13771 7412
rect 13722 7380 13771 7392
rect 13821 7416 13865 7422
rect 13821 7396 13836 7416
rect 13856 7396 13865 7416
rect 13821 7380 13865 7396
rect 13935 7416 13979 7422
rect 13935 7396 13944 7416
rect 13964 7396 13979 7416
rect 13935 7380 13979 7396
rect 14029 7412 14078 7422
rect 16558 7432 16607 7442
rect 16657 7458 16701 7474
rect 16657 7438 16672 7458
rect 16692 7438 16701 7458
rect 16657 7432 16701 7438
rect 16771 7458 16815 7474
rect 16771 7438 16780 7458
rect 16800 7438 16815 7458
rect 16771 7432 16815 7438
rect 16865 7462 16914 7474
rect 16865 7442 16883 7462
rect 16903 7442 16914 7462
rect 16865 7432 16914 7442
rect 16989 7458 17033 7474
rect 16989 7438 16998 7458
rect 17018 7438 17033 7458
rect 16989 7432 17033 7438
rect 17083 7462 17132 7474
rect 17083 7442 17101 7462
rect 17121 7442 17132 7462
rect 17083 7432 17132 7442
rect 23031 7593 23080 7605
rect 23130 7629 23174 7635
rect 23130 7609 23145 7629
rect 23165 7609 23174 7629
rect 23130 7593 23174 7609
rect 23249 7625 23298 7635
rect 23249 7605 23260 7625
rect 23280 7605 23298 7625
rect 23249 7593 23298 7605
rect 23348 7629 23392 7635
rect 23348 7609 23363 7629
rect 23383 7609 23392 7629
rect 23348 7593 23392 7609
rect 23462 7629 23506 7635
rect 23462 7609 23471 7629
rect 23491 7609 23506 7629
rect 23462 7593 23506 7609
rect 23556 7625 23605 7635
rect 23556 7605 23574 7625
rect 23594 7605 23605 7625
rect 23556 7593 23605 7605
rect 24390 7633 24439 7645
rect 24390 7613 24401 7633
rect 24421 7613 24439 7633
rect 24390 7603 24439 7613
rect 24489 7629 24533 7645
rect 24489 7609 24504 7629
rect 24524 7609 24533 7629
rect 24489 7603 24533 7609
rect 24603 7629 24647 7645
rect 24603 7609 24612 7629
rect 24632 7609 24647 7629
rect 24603 7603 24647 7609
rect 24697 7633 24746 7645
rect 24697 7613 24715 7633
rect 24735 7613 24746 7633
rect 24697 7603 24746 7613
rect 24821 7629 24865 7645
rect 24821 7609 24830 7629
rect 24850 7609 24865 7629
rect 24821 7603 24865 7609
rect 24915 7633 24964 7645
rect 24915 7613 24933 7633
rect 24953 7613 24964 7633
rect 24915 7603 24964 7613
rect 27408 7637 27457 7647
rect 27408 7617 27419 7637
rect 27439 7617 27457 7637
rect 14029 7392 14047 7412
rect 14067 7392 14078 7412
rect 14029 7380 14078 7392
rect 6854 7213 6903 7225
rect 3015 7180 3033 7200
rect 3053 7180 3064 7200
rect 3015 7170 3064 7180
rect 1722 7158 1771 7170
rect 5561 7203 5610 7213
rect 5561 7183 5572 7203
rect 5592 7183 5610 7203
rect 5561 7171 5610 7183
rect 5660 7207 5704 7213
rect 5660 7187 5675 7207
rect 5695 7187 5704 7207
rect 5660 7171 5704 7187
rect 5779 7203 5828 7213
rect 5779 7183 5790 7203
rect 5810 7183 5828 7203
rect 5779 7171 5828 7183
rect 5878 7207 5922 7213
rect 5878 7187 5893 7207
rect 5913 7187 5922 7207
rect 5878 7171 5922 7187
rect 5992 7207 6036 7213
rect 5992 7187 6001 7207
rect 6021 7187 6036 7207
rect 5992 7171 6036 7187
rect 6086 7203 6135 7213
rect 6086 7183 6104 7203
rect 6124 7183 6135 7203
rect 6854 7193 6865 7213
rect 6885 7193 6903 7213
rect 6854 7183 6903 7193
rect 6953 7209 6997 7225
rect 6953 7189 6968 7209
rect 6988 7189 6997 7209
rect 6953 7183 6997 7189
rect 7067 7209 7111 7225
rect 7067 7189 7076 7209
rect 7096 7189 7111 7209
rect 7067 7183 7111 7189
rect 7161 7213 7210 7225
rect 7161 7193 7179 7213
rect 7199 7193 7210 7213
rect 7161 7183 7210 7193
rect 7285 7209 7329 7225
rect 7285 7189 7294 7209
rect 7314 7189 7329 7209
rect 7285 7183 7329 7189
rect 7379 7213 7428 7225
rect 27408 7605 27457 7617
rect 27507 7641 27551 7647
rect 27507 7621 27522 7641
rect 27542 7621 27551 7641
rect 27507 7605 27551 7621
rect 27626 7637 27675 7647
rect 27626 7617 27637 7637
rect 27657 7617 27675 7637
rect 27626 7605 27675 7617
rect 27725 7641 27769 7647
rect 27725 7621 27740 7641
rect 27760 7621 27769 7641
rect 27725 7605 27769 7621
rect 27839 7641 27883 7647
rect 27839 7621 27848 7641
rect 27868 7621 27883 7641
rect 27839 7605 27883 7621
rect 27933 7637 27982 7647
rect 27933 7617 27951 7637
rect 27971 7617 27982 7637
rect 27933 7605 27982 7617
rect 28767 7645 28816 7657
rect 28767 7625 28778 7645
rect 28798 7625 28816 7645
rect 28767 7615 28816 7625
rect 28866 7641 28910 7657
rect 28866 7621 28881 7641
rect 28901 7621 28910 7641
rect 28866 7615 28910 7621
rect 28980 7641 29024 7657
rect 28980 7621 28989 7641
rect 29009 7621 29024 7641
rect 28980 7615 29024 7621
rect 29074 7645 29123 7657
rect 29074 7625 29092 7645
rect 29112 7625 29123 7645
rect 29074 7615 29123 7625
rect 29198 7641 29242 7657
rect 29198 7621 29207 7641
rect 29227 7621 29242 7641
rect 29198 7615 29242 7621
rect 29292 7645 29341 7657
rect 29292 7625 29310 7645
rect 29330 7625 29341 7645
rect 29292 7615 29341 7625
rect 31772 7650 31821 7660
rect 31772 7630 31783 7650
rect 31803 7630 31821 7650
rect 20824 7436 20873 7448
rect 20824 7416 20835 7436
rect 20855 7416 20873 7436
rect 11231 7225 11280 7237
rect 7379 7193 7397 7213
rect 7417 7193 7428 7213
rect 7379 7183 7428 7193
rect 6086 7171 6135 7183
rect 9938 7215 9987 7225
rect 9938 7195 9949 7215
rect 9969 7195 9987 7215
rect 9938 7183 9987 7195
rect 10037 7219 10081 7225
rect 10037 7199 10052 7219
rect 10072 7199 10081 7219
rect 10037 7183 10081 7199
rect 10156 7215 10205 7225
rect 10156 7195 10167 7215
rect 10187 7195 10205 7215
rect 10156 7183 10205 7195
rect 10255 7219 10299 7225
rect 10255 7199 10270 7219
rect 10290 7199 10299 7219
rect 10255 7183 10299 7199
rect 10369 7219 10413 7225
rect 10369 7199 10378 7219
rect 10398 7199 10413 7219
rect 10369 7183 10413 7199
rect 10463 7215 10512 7225
rect 10463 7195 10481 7215
rect 10501 7195 10512 7215
rect 11231 7205 11242 7225
rect 11262 7205 11280 7225
rect 11231 7195 11280 7205
rect 11330 7221 11374 7237
rect 11330 7201 11345 7221
rect 11365 7201 11374 7221
rect 11330 7195 11374 7201
rect 11444 7221 11488 7237
rect 11444 7201 11453 7221
rect 11473 7201 11488 7221
rect 11444 7195 11488 7201
rect 11538 7225 11587 7237
rect 11538 7205 11556 7225
rect 11576 7205 11587 7225
rect 11538 7195 11587 7205
rect 11662 7221 11706 7237
rect 11662 7201 11671 7221
rect 11691 7201 11706 7221
rect 11662 7195 11706 7201
rect 11756 7225 11805 7237
rect 17770 7386 17819 7396
rect 17770 7366 17781 7386
rect 17801 7366 17819 7386
rect 17770 7354 17819 7366
rect 17869 7390 17913 7396
rect 17869 7370 17884 7390
rect 17904 7370 17913 7390
rect 17869 7354 17913 7370
rect 17988 7386 18037 7396
rect 17988 7366 17999 7386
rect 18019 7366 18037 7386
rect 17988 7354 18037 7366
rect 18087 7390 18131 7396
rect 18087 7370 18102 7390
rect 18122 7370 18131 7390
rect 18087 7354 18131 7370
rect 18201 7390 18245 7396
rect 18201 7370 18210 7390
rect 18230 7370 18245 7390
rect 18201 7354 18245 7370
rect 18295 7386 18344 7396
rect 20824 7406 20873 7416
rect 20923 7432 20967 7448
rect 20923 7412 20938 7432
rect 20958 7412 20967 7432
rect 20923 7406 20967 7412
rect 21037 7432 21081 7448
rect 21037 7412 21046 7432
rect 21066 7412 21081 7432
rect 21037 7406 21081 7412
rect 21131 7436 21180 7448
rect 21131 7416 21149 7436
rect 21169 7416 21180 7436
rect 21131 7406 21180 7416
rect 21255 7432 21299 7448
rect 21255 7412 21264 7432
rect 21284 7412 21299 7432
rect 21255 7406 21299 7412
rect 21349 7436 21398 7448
rect 21349 7416 21367 7436
rect 21387 7416 21398 7436
rect 21349 7406 21398 7416
rect 18295 7366 18313 7386
rect 18333 7366 18344 7386
rect 18295 7354 18344 7366
rect 31772 7618 31821 7630
rect 31871 7654 31915 7660
rect 31871 7634 31886 7654
rect 31906 7634 31915 7654
rect 31871 7618 31915 7634
rect 31990 7650 32039 7660
rect 31990 7630 32001 7650
rect 32021 7630 32039 7650
rect 31990 7618 32039 7630
rect 32089 7654 32133 7660
rect 32089 7634 32104 7654
rect 32124 7634 32133 7654
rect 32089 7618 32133 7634
rect 32203 7654 32247 7660
rect 32203 7634 32212 7654
rect 32232 7634 32247 7654
rect 32203 7618 32247 7634
rect 32297 7650 32346 7660
rect 32297 7630 32315 7650
rect 32335 7630 32346 7650
rect 32297 7618 32346 7630
rect 33131 7658 33180 7670
rect 33131 7638 33142 7658
rect 33162 7638 33180 7658
rect 33131 7628 33180 7638
rect 33230 7654 33274 7670
rect 33230 7634 33245 7654
rect 33265 7634 33274 7654
rect 33230 7628 33274 7634
rect 33344 7654 33388 7670
rect 33344 7634 33353 7654
rect 33373 7634 33388 7654
rect 33344 7628 33388 7634
rect 33438 7658 33487 7670
rect 33438 7638 33456 7658
rect 33476 7638 33487 7658
rect 33438 7628 33487 7638
rect 33562 7654 33606 7670
rect 33562 7634 33571 7654
rect 33591 7634 33606 7654
rect 33562 7628 33606 7634
rect 33656 7658 33705 7670
rect 33656 7638 33674 7658
rect 33694 7638 33705 7658
rect 33656 7628 33705 7638
rect 25188 7449 25237 7461
rect 25188 7429 25199 7449
rect 25219 7429 25237 7449
rect 22134 7399 22183 7409
rect 22134 7379 22145 7399
rect 22165 7379 22183 7399
rect 22134 7367 22183 7379
rect 22233 7403 22277 7409
rect 22233 7383 22248 7403
rect 22268 7383 22277 7403
rect 22233 7367 22277 7383
rect 22352 7399 22401 7409
rect 22352 7379 22363 7399
rect 22383 7379 22401 7399
rect 22352 7367 22401 7379
rect 22451 7403 22495 7409
rect 22451 7383 22466 7403
rect 22486 7383 22495 7403
rect 22451 7367 22495 7383
rect 22565 7403 22609 7409
rect 22565 7383 22574 7403
rect 22594 7383 22609 7403
rect 22565 7367 22609 7383
rect 22659 7399 22708 7409
rect 25188 7419 25237 7429
rect 25287 7445 25331 7461
rect 25287 7425 25302 7445
rect 25322 7425 25331 7445
rect 25287 7419 25331 7425
rect 25401 7445 25445 7461
rect 25401 7425 25410 7445
rect 25430 7425 25445 7445
rect 25401 7419 25445 7425
rect 25495 7449 25544 7461
rect 25495 7429 25513 7449
rect 25533 7429 25544 7449
rect 25495 7419 25544 7429
rect 25619 7445 25663 7461
rect 25619 7425 25628 7445
rect 25648 7425 25663 7445
rect 25619 7419 25663 7425
rect 25713 7449 25762 7461
rect 25713 7429 25731 7449
rect 25751 7429 25762 7449
rect 25713 7419 25762 7429
rect 22659 7379 22677 7399
rect 22697 7379 22708 7399
rect 22659 7367 22708 7379
rect 15595 7238 15644 7250
rect 11756 7205 11774 7225
rect 11794 7205 11805 7225
rect 11756 7195 11805 7205
rect 10463 7183 10512 7195
rect 400 6962 449 6972
rect 400 6942 411 6962
rect 431 6942 449 6962
rect 400 6930 449 6942
rect 499 6966 543 6972
rect 499 6946 514 6966
rect 534 6946 543 6966
rect 499 6930 543 6946
rect 618 6962 667 6972
rect 618 6942 629 6962
rect 649 6942 667 6962
rect 618 6930 667 6942
rect 717 6966 761 6972
rect 717 6946 732 6966
rect 752 6946 761 6966
rect 717 6930 761 6946
rect 831 6966 875 6972
rect 831 6946 840 6966
rect 860 6946 875 6966
rect 831 6930 875 6946
rect 925 6962 974 6972
rect 925 6942 943 6962
rect 963 6942 974 6962
rect 14302 7228 14351 7238
rect 14302 7208 14313 7228
rect 14333 7208 14351 7228
rect 14302 7196 14351 7208
rect 14401 7232 14445 7238
rect 14401 7212 14416 7232
rect 14436 7212 14445 7232
rect 14401 7196 14445 7212
rect 14520 7228 14569 7238
rect 14520 7208 14531 7228
rect 14551 7208 14569 7228
rect 14520 7196 14569 7208
rect 14619 7232 14663 7238
rect 14619 7212 14634 7232
rect 14654 7212 14663 7232
rect 14619 7196 14663 7212
rect 14733 7232 14777 7238
rect 14733 7212 14742 7232
rect 14762 7212 14777 7232
rect 14733 7196 14777 7212
rect 14827 7228 14876 7238
rect 14827 7208 14845 7228
rect 14865 7208 14876 7228
rect 15595 7218 15606 7238
rect 15626 7218 15644 7238
rect 15595 7208 15644 7218
rect 15694 7234 15738 7250
rect 15694 7214 15709 7234
rect 15729 7214 15738 7234
rect 15694 7208 15738 7214
rect 15808 7234 15852 7250
rect 15808 7214 15817 7234
rect 15837 7214 15852 7234
rect 15808 7208 15852 7214
rect 15902 7238 15951 7250
rect 15902 7218 15920 7238
rect 15940 7218 15951 7238
rect 15902 7208 15951 7218
rect 16026 7234 16070 7250
rect 16026 7214 16035 7234
rect 16055 7214 16070 7234
rect 16026 7208 16070 7214
rect 16120 7238 16169 7250
rect 16120 7218 16138 7238
rect 16158 7218 16169 7238
rect 16120 7208 16169 7218
rect 29565 7461 29614 7473
rect 29565 7441 29576 7461
rect 29596 7441 29614 7461
rect 26511 7411 26560 7421
rect 26511 7391 26522 7411
rect 26542 7391 26560 7411
rect 26511 7379 26560 7391
rect 26610 7415 26654 7421
rect 26610 7395 26625 7415
rect 26645 7395 26654 7415
rect 26610 7379 26654 7395
rect 26729 7411 26778 7421
rect 26729 7391 26740 7411
rect 26760 7391 26778 7411
rect 26729 7379 26778 7391
rect 26828 7415 26872 7421
rect 26828 7395 26843 7415
rect 26863 7395 26872 7415
rect 26828 7379 26872 7395
rect 26942 7415 26986 7421
rect 26942 7395 26951 7415
rect 26971 7395 26986 7415
rect 26942 7379 26986 7395
rect 27036 7411 27085 7421
rect 29565 7431 29614 7441
rect 29664 7457 29708 7473
rect 29664 7437 29679 7457
rect 29699 7437 29708 7457
rect 29664 7431 29708 7437
rect 29778 7457 29822 7473
rect 29778 7437 29787 7457
rect 29807 7437 29822 7457
rect 29778 7431 29822 7437
rect 29872 7461 29921 7473
rect 29872 7441 29890 7461
rect 29910 7441 29921 7461
rect 29872 7431 29921 7441
rect 29996 7457 30040 7473
rect 29996 7437 30005 7457
rect 30025 7437 30040 7457
rect 29996 7431 30040 7437
rect 30090 7461 30139 7473
rect 30090 7441 30108 7461
rect 30128 7441 30139 7461
rect 30090 7431 30139 7441
rect 27036 7391 27054 7411
rect 27074 7391 27085 7411
rect 27036 7379 27085 7391
rect 19861 7212 19910 7224
rect 14827 7196 14876 7208
rect 925 6930 974 6942
rect 4764 6975 4813 6985
rect 4764 6955 4775 6975
rect 4795 6955 4813 6975
rect 4764 6943 4813 6955
rect 4863 6979 4907 6985
rect 4863 6959 4878 6979
rect 4898 6959 4907 6979
rect 4863 6943 4907 6959
rect 4982 6975 5031 6985
rect 4982 6955 4993 6975
rect 5013 6955 5031 6975
rect 4982 6943 5031 6955
rect 5081 6979 5125 6985
rect 5081 6959 5096 6979
rect 5116 6959 5125 6979
rect 5081 6943 5125 6959
rect 5195 6979 5239 6985
rect 5195 6959 5204 6979
rect 5224 6959 5239 6979
rect 5195 6943 5239 6959
rect 5289 6975 5338 6985
rect 5289 6955 5307 6975
rect 5327 6955 5338 6975
rect 18568 7202 18617 7212
rect 18568 7182 18579 7202
rect 18599 7182 18617 7202
rect 18568 7170 18617 7182
rect 18667 7206 18711 7212
rect 18667 7186 18682 7206
rect 18702 7186 18711 7206
rect 18667 7170 18711 7186
rect 18786 7202 18835 7212
rect 18786 7182 18797 7202
rect 18817 7182 18835 7202
rect 18786 7170 18835 7182
rect 18885 7206 18929 7212
rect 18885 7186 18900 7206
rect 18920 7186 18929 7206
rect 18885 7170 18929 7186
rect 18999 7206 19043 7212
rect 18999 7186 19008 7206
rect 19028 7186 19043 7206
rect 18999 7170 19043 7186
rect 19093 7202 19142 7212
rect 19093 7182 19111 7202
rect 19131 7182 19142 7202
rect 19861 7192 19872 7212
rect 19892 7192 19910 7212
rect 19861 7182 19910 7192
rect 19960 7208 20004 7224
rect 19960 7188 19975 7208
rect 19995 7188 20004 7208
rect 19960 7182 20004 7188
rect 20074 7208 20118 7224
rect 20074 7188 20083 7208
rect 20103 7188 20118 7208
rect 20074 7182 20118 7188
rect 20168 7212 20217 7224
rect 20168 7192 20186 7212
rect 20206 7192 20217 7212
rect 20168 7182 20217 7192
rect 20292 7208 20336 7224
rect 20292 7188 20301 7208
rect 20321 7188 20336 7208
rect 20292 7182 20336 7188
rect 20386 7212 20435 7224
rect 33929 7474 33978 7486
rect 33929 7454 33940 7474
rect 33960 7454 33978 7474
rect 30875 7424 30924 7434
rect 30875 7404 30886 7424
rect 30906 7404 30924 7424
rect 30875 7392 30924 7404
rect 30974 7428 31018 7434
rect 30974 7408 30989 7428
rect 31009 7408 31018 7428
rect 30974 7392 31018 7408
rect 31093 7424 31142 7434
rect 31093 7404 31104 7424
rect 31124 7404 31142 7424
rect 31093 7392 31142 7404
rect 31192 7428 31236 7434
rect 31192 7408 31207 7428
rect 31227 7408 31236 7428
rect 31192 7392 31236 7408
rect 31306 7428 31350 7434
rect 31306 7408 31315 7428
rect 31335 7408 31350 7428
rect 31306 7392 31350 7408
rect 31400 7424 31449 7434
rect 33929 7444 33978 7454
rect 34028 7470 34072 7486
rect 34028 7450 34043 7470
rect 34063 7450 34072 7470
rect 34028 7444 34072 7450
rect 34142 7470 34186 7486
rect 34142 7450 34151 7470
rect 34171 7450 34186 7470
rect 34142 7444 34186 7450
rect 34236 7474 34285 7486
rect 34236 7454 34254 7474
rect 34274 7454 34285 7474
rect 34236 7444 34285 7454
rect 34360 7470 34404 7486
rect 34360 7450 34369 7470
rect 34389 7450 34404 7470
rect 34360 7444 34404 7450
rect 34454 7474 34503 7486
rect 34454 7454 34472 7474
rect 34492 7454 34503 7474
rect 34454 7444 34503 7454
rect 31400 7404 31418 7424
rect 31438 7404 31449 7424
rect 31400 7392 31449 7404
rect 24225 7225 24274 7237
rect 20386 7192 20404 7212
rect 20424 7192 20435 7212
rect 20386 7182 20435 7192
rect 19093 7170 19142 7182
rect 5289 6943 5338 6955
rect 9141 6987 9190 6997
rect 9141 6967 9152 6987
rect 9172 6967 9190 6987
rect 9141 6955 9190 6967
rect 9240 6991 9284 6997
rect 9240 6971 9255 6991
rect 9275 6971 9284 6991
rect 9240 6955 9284 6971
rect 9359 6987 9408 6997
rect 9359 6967 9370 6987
rect 9390 6967 9408 6987
rect 9359 6955 9408 6967
rect 9458 6991 9502 6997
rect 9458 6971 9473 6991
rect 9493 6971 9502 6991
rect 9458 6955 9502 6971
rect 9572 6991 9616 6997
rect 9572 6971 9581 6991
rect 9601 6971 9616 6991
rect 9572 6955 9616 6971
rect 9666 6987 9715 6997
rect 9666 6967 9684 6987
rect 9704 6967 9715 6987
rect 22932 7215 22981 7225
rect 22932 7195 22943 7215
rect 22963 7195 22981 7215
rect 22932 7183 22981 7195
rect 23031 7219 23075 7225
rect 23031 7199 23046 7219
rect 23066 7199 23075 7219
rect 23031 7183 23075 7199
rect 23150 7215 23199 7225
rect 23150 7195 23161 7215
rect 23181 7195 23199 7215
rect 23150 7183 23199 7195
rect 23249 7219 23293 7225
rect 23249 7199 23264 7219
rect 23284 7199 23293 7219
rect 23249 7183 23293 7199
rect 23363 7219 23407 7225
rect 23363 7199 23372 7219
rect 23392 7199 23407 7219
rect 23363 7183 23407 7199
rect 23457 7215 23506 7225
rect 23457 7195 23475 7215
rect 23495 7195 23506 7215
rect 24225 7205 24236 7225
rect 24256 7205 24274 7225
rect 24225 7195 24274 7205
rect 24324 7221 24368 7237
rect 24324 7201 24339 7221
rect 24359 7201 24368 7221
rect 24324 7195 24368 7201
rect 24438 7221 24482 7237
rect 24438 7201 24447 7221
rect 24467 7201 24482 7221
rect 24438 7195 24482 7201
rect 24532 7225 24581 7237
rect 24532 7205 24550 7225
rect 24570 7205 24581 7225
rect 24532 7195 24581 7205
rect 24656 7221 24700 7237
rect 24656 7201 24665 7221
rect 24685 7201 24700 7221
rect 24656 7195 24700 7201
rect 24750 7225 24799 7237
rect 28602 7237 28651 7249
rect 24750 7205 24768 7225
rect 24788 7205 24799 7225
rect 24750 7195 24799 7205
rect 23457 7183 23506 7195
rect 9666 6955 9715 6967
rect 13505 7000 13554 7010
rect 13505 6980 13516 7000
rect 13536 6980 13554 7000
rect 13505 6968 13554 6980
rect 13604 7004 13648 7010
rect 13604 6984 13619 7004
rect 13639 6984 13648 7004
rect 13604 6968 13648 6984
rect 13723 7000 13772 7010
rect 13723 6980 13734 7000
rect 13754 6980 13772 7000
rect 13723 6968 13772 6980
rect 13822 7004 13866 7010
rect 13822 6984 13837 7004
rect 13857 6984 13866 7004
rect 13822 6968 13866 6984
rect 13936 7004 13980 7010
rect 13936 6984 13945 7004
rect 13965 6984 13980 7004
rect 13936 6968 13980 6984
rect 14030 7000 14079 7010
rect 14030 6980 14048 7000
rect 14068 6980 14079 7000
rect 14030 6968 14079 6980
rect 27309 7227 27358 7237
rect 27309 7207 27320 7227
rect 27340 7207 27358 7227
rect 27309 7195 27358 7207
rect 27408 7231 27452 7237
rect 27408 7211 27423 7231
rect 27443 7211 27452 7231
rect 27408 7195 27452 7211
rect 27527 7227 27576 7237
rect 27527 7207 27538 7227
rect 27558 7207 27576 7227
rect 27527 7195 27576 7207
rect 27626 7231 27670 7237
rect 27626 7211 27641 7231
rect 27661 7211 27670 7231
rect 27626 7195 27670 7211
rect 27740 7231 27784 7237
rect 27740 7211 27749 7231
rect 27769 7211 27784 7231
rect 27740 7195 27784 7211
rect 27834 7227 27883 7237
rect 27834 7207 27852 7227
rect 27872 7207 27883 7227
rect 28602 7217 28613 7237
rect 28633 7217 28651 7237
rect 28602 7207 28651 7217
rect 28701 7233 28745 7249
rect 28701 7213 28716 7233
rect 28736 7213 28745 7233
rect 28701 7207 28745 7213
rect 28815 7233 28859 7249
rect 28815 7213 28824 7233
rect 28844 7213 28859 7233
rect 28815 7207 28859 7213
rect 28909 7237 28958 7249
rect 28909 7217 28927 7237
rect 28947 7217 28958 7237
rect 28909 7207 28958 7217
rect 29033 7233 29077 7249
rect 29033 7213 29042 7233
rect 29062 7213 29077 7233
rect 29033 7207 29077 7213
rect 29127 7237 29176 7249
rect 32966 7250 33015 7262
rect 29127 7217 29145 7237
rect 29165 7217 29176 7237
rect 29127 7207 29176 7217
rect 27834 7195 27883 7207
rect 17771 6974 17820 6984
rect 17771 6954 17782 6974
rect 17802 6954 17820 6974
rect 17771 6942 17820 6954
rect 17870 6978 17914 6984
rect 17870 6958 17885 6978
rect 17905 6958 17914 6978
rect 17870 6942 17914 6958
rect 17989 6974 18038 6984
rect 17989 6954 18000 6974
rect 18020 6954 18038 6974
rect 17989 6942 18038 6954
rect 18088 6978 18132 6984
rect 18088 6958 18103 6978
rect 18123 6958 18132 6978
rect 18088 6942 18132 6958
rect 18202 6978 18246 6984
rect 18202 6958 18211 6978
rect 18231 6958 18246 6978
rect 18202 6942 18246 6958
rect 18296 6974 18345 6984
rect 18296 6954 18314 6974
rect 18334 6954 18345 6974
rect 31673 7240 31722 7250
rect 31673 7220 31684 7240
rect 31704 7220 31722 7240
rect 31673 7208 31722 7220
rect 31772 7244 31816 7250
rect 31772 7224 31787 7244
rect 31807 7224 31816 7244
rect 31772 7208 31816 7224
rect 31891 7240 31940 7250
rect 31891 7220 31902 7240
rect 31922 7220 31940 7240
rect 31891 7208 31940 7220
rect 31990 7244 32034 7250
rect 31990 7224 32005 7244
rect 32025 7224 32034 7244
rect 31990 7208 32034 7224
rect 32104 7244 32148 7250
rect 32104 7224 32113 7244
rect 32133 7224 32148 7244
rect 32104 7208 32148 7224
rect 32198 7240 32247 7250
rect 32198 7220 32216 7240
rect 32236 7220 32247 7240
rect 32966 7230 32977 7250
rect 32997 7230 33015 7250
rect 32966 7220 33015 7230
rect 33065 7246 33109 7262
rect 33065 7226 33080 7246
rect 33100 7226 33109 7246
rect 33065 7220 33109 7226
rect 33179 7246 33223 7262
rect 33179 7226 33188 7246
rect 33208 7226 33223 7246
rect 33179 7220 33223 7226
rect 33273 7250 33322 7262
rect 33273 7230 33291 7250
rect 33311 7230 33322 7250
rect 33273 7220 33322 7230
rect 33397 7246 33441 7262
rect 33397 7226 33406 7246
rect 33426 7226 33441 7246
rect 33397 7220 33441 7226
rect 33491 7250 33540 7262
rect 33491 7230 33509 7250
rect 33529 7230 33540 7250
rect 33491 7220 33540 7230
rect 32198 7208 32247 7220
rect 18296 6942 18345 6954
rect 22135 6987 22184 6997
rect 22135 6967 22146 6987
rect 22166 6967 22184 6987
rect 22135 6955 22184 6967
rect 22234 6991 22278 6997
rect 22234 6971 22249 6991
rect 22269 6971 22278 6991
rect 22234 6955 22278 6971
rect 22353 6987 22402 6997
rect 22353 6967 22364 6987
rect 22384 6967 22402 6987
rect 22353 6955 22402 6967
rect 22452 6991 22496 6997
rect 22452 6971 22467 6991
rect 22487 6971 22496 6991
rect 22452 6955 22496 6971
rect 22566 6991 22610 6997
rect 22566 6971 22575 6991
rect 22595 6971 22610 6991
rect 22566 6955 22610 6971
rect 22660 6987 22709 6997
rect 22660 6967 22678 6987
rect 22698 6967 22709 6987
rect 22660 6955 22709 6967
rect 26512 6999 26561 7009
rect 26512 6979 26523 6999
rect 26543 6979 26561 6999
rect 26512 6967 26561 6979
rect 26611 7003 26655 7009
rect 26611 6983 26626 7003
rect 26646 6983 26655 7003
rect 26611 6967 26655 6983
rect 26730 6999 26779 7009
rect 26730 6979 26741 6999
rect 26761 6979 26779 6999
rect 26730 6967 26779 6979
rect 26829 7003 26873 7009
rect 26829 6983 26844 7003
rect 26864 6983 26873 7003
rect 26829 6967 26873 6983
rect 26943 7003 26987 7009
rect 26943 6983 26952 7003
rect 26972 6983 26987 7003
rect 26943 6967 26987 6983
rect 27037 6999 27086 7009
rect 27037 6979 27055 6999
rect 27075 6979 27086 6999
rect 27037 6967 27086 6979
rect 30876 7012 30925 7022
rect 30876 6992 30887 7012
rect 30907 6992 30925 7012
rect 30876 6980 30925 6992
rect 30975 7016 31019 7022
rect 30975 6996 30990 7016
rect 31010 6996 31019 7016
rect 30975 6980 31019 6996
rect 31094 7012 31143 7022
rect 31094 6992 31105 7012
rect 31125 6992 31143 7012
rect 31094 6980 31143 6992
rect 31193 7016 31237 7022
rect 31193 6996 31208 7016
rect 31228 6996 31237 7016
rect 31193 6980 31237 6996
rect 31307 7016 31351 7022
rect 31307 6996 31316 7016
rect 31336 6996 31351 7016
rect 31307 6980 31351 6996
rect 31401 7012 31450 7022
rect 31401 6992 31419 7012
rect 31439 6992 31450 7012
rect 31401 6980 31450 6992
rect 3432 6818 3481 6830
rect 3432 6798 3443 6818
rect 3463 6798 3481 6818
rect 3432 6788 3481 6798
rect 3531 6814 3575 6830
rect 3531 6794 3546 6814
rect 3566 6794 3575 6814
rect 3531 6788 3575 6794
rect 3645 6814 3689 6830
rect 3645 6794 3654 6814
rect 3674 6794 3689 6814
rect 3645 6788 3689 6794
rect 3739 6818 3788 6830
rect 3739 6798 3757 6818
rect 3777 6798 3788 6818
rect 3739 6788 3788 6798
rect 3863 6814 3907 6830
rect 3863 6794 3872 6814
rect 3892 6794 3907 6814
rect 3863 6788 3907 6794
rect 3957 6818 4006 6830
rect 3957 6798 3975 6818
rect 3995 6798 4006 6818
rect 3957 6788 4006 6798
rect 7796 6831 7845 6843
rect 7796 6811 7807 6831
rect 7827 6811 7845 6831
rect 7796 6801 7845 6811
rect 7895 6827 7939 6843
rect 7895 6807 7910 6827
rect 7930 6807 7939 6827
rect 7895 6801 7939 6807
rect 8009 6827 8053 6843
rect 8009 6807 8018 6827
rect 8038 6807 8053 6827
rect 8009 6801 8053 6807
rect 8103 6831 8152 6843
rect 8103 6811 8121 6831
rect 8141 6811 8152 6831
rect 8103 6801 8152 6811
rect 8227 6827 8271 6843
rect 8227 6807 8236 6827
rect 8256 6807 8271 6827
rect 8227 6801 8271 6807
rect 8321 6831 8370 6843
rect 8321 6811 8339 6831
rect 8359 6811 8370 6831
rect 8321 6801 8370 6811
rect 12173 6843 12222 6855
rect 12173 6823 12184 6843
rect 12204 6823 12222 6843
rect 12173 6813 12222 6823
rect 12272 6839 12316 6855
rect 12272 6819 12287 6839
rect 12307 6819 12316 6839
rect 12272 6813 12316 6819
rect 12386 6839 12430 6855
rect 12386 6819 12395 6839
rect 12415 6819 12430 6839
rect 12386 6813 12430 6819
rect 12480 6843 12529 6855
rect 12480 6823 12498 6843
rect 12518 6823 12529 6843
rect 12480 6813 12529 6823
rect 12604 6839 12648 6855
rect 12604 6819 12613 6839
rect 12633 6819 12648 6839
rect 12604 6813 12648 6819
rect 12698 6843 12747 6855
rect 12698 6823 12716 6843
rect 12736 6823 12747 6843
rect 12698 6813 12747 6823
rect 16537 6856 16586 6868
rect 2635 6590 2684 6602
rect 1342 6580 1391 6590
rect 1342 6560 1353 6580
rect 1373 6560 1391 6580
rect 1342 6548 1391 6560
rect 1441 6584 1485 6590
rect 1441 6564 1456 6584
rect 1476 6564 1485 6584
rect 1441 6548 1485 6564
rect 1560 6580 1609 6590
rect 1560 6560 1571 6580
rect 1591 6560 1609 6580
rect 1560 6548 1609 6560
rect 1659 6584 1703 6590
rect 1659 6564 1674 6584
rect 1694 6564 1703 6584
rect 1659 6548 1703 6564
rect 1773 6584 1817 6590
rect 1773 6564 1782 6584
rect 1802 6564 1817 6584
rect 1773 6548 1817 6564
rect 1867 6580 1916 6590
rect 1867 6560 1885 6580
rect 1905 6560 1916 6580
rect 2635 6570 2646 6590
rect 2666 6570 2684 6590
rect 2635 6560 2684 6570
rect 2734 6586 2778 6602
rect 2734 6566 2749 6586
rect 2769 6566 2778 6586
rect 2734 6560 2778 6566
rect 2848 6586 2892 6602
rect 2848 6566 2857 6586
rect 2877 6566 2892 6586
rect 2848 6560 2892 6566
rect 2942 6590 2991 6602
rect 2942 6570 2960 6590
rect 2980 6570 2991 6590
rect 2942 6560 2991 6570
rect 3066 6586 3110 6602
rect 3066 6566 3075 6586
rect 3095 6566 3110 6586
rect 3066 6560 3110 6566
rect 3160 6590 3209 6602
rect 3160 6570 3178 6590
rect 3198 6570 3209 6590
rect 3160 6560 3209 6570
rect 16537 6836 16548 6856
rect 16568 6836 16586 6856
rect 16537 6826 16586 6836
rect 16636 6852 16680 6868
rect 16636 6832 16651 6852
rect 16671 6832 16680 6852
rect 16636 6826 16680 6832
rect 16750 6852 16794 6868
rect 16750 6832 16759 6852
rect 16779 6832 16794 6852
rect 16750 6826 16794 6832
rect 16844 6856 16893 6868
rect 16844 6836 16862 6856
rect 16882 6836 16893 6856
rect 16844 6826 16893 6836
rect 16968 6852 17012 6868
rect 16968 6832 16977 6852
rect 16997 6832 17012 6852
rect 16968 6826 17012 6832
rect 17062 6856 17111 6868
rect 17062 6836 17080 6856
rect 17100 6836 17111 6856
rect 17062 6826 17111 6836
rect 6999 6603 7048 6615
rect 5706 6593 5755 6603
rect 5706 6573 5717 6593
rect 5737 6573 5755 6593
rect 1867 6548 1916 6560
rect 5706 6561 5755 6573
rect 5805 6597 5849 6603
rect 5805 6577 5820 6597
rect 5840 6577 5849 6597
rect 5805 6561 5849 6577
rect 5924 6593 5973 6603
rect 5924 6573 5935 6593
rect 5955 6573 5973 6593
rect 5924 6561 5973 6573
rect 6023 6597 6067 6603
rect 6023 6577 6038 6597
rect 6058 6577 6067 6597
rect 6023 6561 6067 6577
rect 6137 6597 6181 6603
rect 6137 6577 6146 6597
rect 6166 6577 6181 6597
rect 6137 6561 6181 6577
rect 6231 6593 6280 6603
rect 6231 6573 6249 6593
rect 6269 6573 6280 6593
rect 6999 6583 7010 6603
rect 7030 6583 7048 6603
rect 6999 6573 7048 6583
rect 7098 6599 7142 6615
rect 7098 6579 7113 6599
rect 7133 6579 7142 6599
rect 7098 6573 7142 6579
rect 7212 6599 7256 6615
rect 7212 6579 7221 6599
rect 7241 6579 7256 6599
rect 7212 6573 7256 6579
rect 7306 6603 7355 6615
rect 7306 6583 7324 6603
rect 7344 6583 7355 6603
rect 7306 6573 7355 6583
rect 7430 6599 7474 6615
rect 7430 6579 7439 6599
rect 7459 6579 7474 6599
rect 7430 6573 7474 6579
rect 7524 6603 7573 6615
rect 7524 6583 7542 6603
rect 7562 6583 7573 6603
rect 7524 6573 7573 6583
rect 20803 6830 20852 6842
rect 20803 6810 20814 6830
rect 20834 6810 20852 6830
rect 20803 6800 20852 6810
rect 20902 6826 20946 6842
rect 20902 6806 20917 6826
rect 20937 6806 20946 6826
rect 20902 6800 20946 6806
rect 21016 6826 21060 6842
rect 21016 6806 21025 6826
rect 21045 6806 21060 6826
rect 21016 6800 21060 6806
rect 21110 6830 21159 6842
rect 21110 6810 21128 6830
rect 21148 6810 21159 6830
rect 21110 6800 21159 6810
rect 21234 6826 21278 6842
rect 21234 6806 21243 6826
rect 21263 6806 21278 6826
rect 21234 6800 21278 6806
rect 21328 6830 21377 6842
rect 21328 6810 21346 6830
rect 21366 6810 21377 6830
rect 21328 6800 21377 6810
rect 25167 6843 25216 6855
rect 11376 6615 11425 6627
rect 10083 6605 10132 6615
rect 10083 6585 10094 6605
rect 10114 6585 10132 6605
rect 6231 6561 6280 6573
rect 10083 6573 10132 6585
rect 10182 6609 10226 6615
rect 10182 6589 10197 6609
rect 10217 6589 10226 6609
rect 10182 6573 10226 6589
rect 10301 6605 10350 6615
rect 10301 6585 10312 6605
rect 10332 6585 10350 6605
rect 10301 6573 10350 6585
rect 10400 6609 10444 6615
rect 10400 6589 10415 6609
rect 10435 6589 10444 6609
rect 10400 6573 10444 6589
rect 10514 6609 10558 6615
rect 10514 6589 10523 6609
rect 10543 6589 10558 6609
rect 10514 6573 10558 6589
rect 10608 6605 10657 6615
rect 10608 6585 10626 6605
rect 10646 6585 10657 6605
rect 11376 6595 11387 6615
rect 11407 6595 11425 6615
rect 11376 6585 11425 6595
rect 11475 6611 11519 6627
rect 11475 6591 11490 6611
rect 11510 6591 11519 6611
rect 11475 6585 11519 6591
rect 11589 6611 11633 6627
rect 11589 6591 11598 6611
rect 11618 6591 11633 6611
rect 11589 6585 11633 6591
rect 11683 6615 11732 6627
rect 11683 6595 11701 6615
rect 11721 6595 11732 6615
rect 11683 6585 11732 6595
rect 11807 6611 11851 6627
rect 11807 6591 11816 6611
rect 11836 6591 11851 6611
rect 11807 6585 11851 6591
rect 11901 6615 11950 6627
rect 11901 6595 11919 6615
rect 11939 6595 11950 6615
rect 11901 6585 11950 6595
rect 25167 6823 25178 6843
rect 25198 6823 25216 6843
rect 25167 6813 25216 6823
rect 25266 6839 25310 6855
rect 25266 6819 25281 6839
rect 25301 6819 25310 6839
rect 25266 6813 25310 6819
rect 25380 6839 25424 6855
rect 25380 6819 25389 6839
rect 25409 6819 25424 6839
rect 25380 6813 25424 6819
rect 25474 6843 25523 6855
rect 25474 6823 25492 6843
rect 25512 6823 25523 6843
rect 25474 6813 25523 6823
rect 25598 6839 25642 6855
rect 25598 6819 25607 6839
rect 25627 6819 25642 6839
rect 25598 6813 25642 6819
rect 25692 6843 25741 6855
rect 25692 6823 25710 6843
rect 25730 6823 25741 6843
rect 25692 6813 25741 6823
rect 29544 6855 29593 6867
rect 15740 6628 15789 6640
rect 14447 6618 14496 6628
rect 14447 6598 14458 6618
rect 14478 6598 14496 6618
rect 10608 6573 10657 6585
rect 3433 6406 3482 6418
rect 3433 6386 3444 6406
rect 3464 6386 3482 6406
rect 379 6356 428 6366
rect 379 6336 390 6356
rect 410 6336 428 6356
rect 379 6324 428 6336
rect 478 6360 522 6366
rect 478 6340 493 6360
rect 513 6340 522 6360
rect 478 6324 522 6340
rect 597 6356 646 6366
rect 597 6336 608 6356
rect 628 6336 646 6356
rect 597 6324 646 6336
rect 696 6360 740 6366
rect 696 6340 711 6360
rect 731 6340 740 6360
rect 696 6324 740 6340
rect 810 6360 854 6366
rect 810 6340 819 6360
rect 839 6340 854 6360
rect 810 6324 854 6340
rect 904 6356 953 6366
rect 3433 6376 3482 6386
rect 3532 6402 3576 6418
rect 3532 6382 3547 6402
rect 3567 6382 3576 6402
rect 3532 6376 3576 6382
rect 3646 6402 3690 6418
rect 3646 6382 3655 6402
rect 3675 6382 3690 6402
rect 3646 6376 3690 6382
rect 3740 6406 3789 6418
rect 3740 6386 3758 6406
rect 3778 6386 3789 6406
rect 3740 6376 3789 6386
rect 3864 6402 3908 6418
rect 3864 6382 3873 6402
rect 3893 6382 3908 6402
rect 3864 6376 3908 6382
rect 3958 6406 4007 6418
rect 3958 6386 3976 6406
rect 3996 6386 4007 6406
rect 3958 6376 4007 6386
rect 904 6336 922 6356
rect 942 6336 953 6356
rect 904 6324 953 6336
rect 14447 6586 14496 6598
rect 14546 6622 14590 6628
rect 14546 6602 14561 6622
rect 14581 6602 14590 6622
rect 14546 6586 14590 6602
rect 14665 6618 14714 6628
rect 14665 6598 14676 6618
rect 14696 6598 14714 6618
rect 14665 6586 14714 6598
rect 14764 6622 14808 6628
rect 14764 6602 14779 6622
rect 14799 6602 14808 6622
rect 14764 6586 14808 6602
rect 14878 6622 14922 6628
rect 14878 6602 14887 6622
rect 14907 6602 14922 6622
rect 14878 6586 14922 6602
rect 14972 6618 15021 6628
rect 14972 6598 14990 6618
rect 15010 6598 15021 6618
rect 15740 6608 15751 6628
rect 15771 6608 15789 6628
rect 15740 6598 15789 6608
rect 15839 6624 15883 6640
rect 15839 6604 15854 6624
rect 15874 6604 15883 6624
rect 15839 6598 15883 6604
rect 15953 6624 15997 6640
rect 15953 6604 15962 6624
rect 15982 6604 15997 6624
rect 15953 6598 15997 6604
rect 16047 6628 16096 6640
rect 16047 6608 16065 6628
rect 16085 6608 16096 6628
rect 16047 6598 16096 6608
rect 16171 6624 16215 6640
rect 16171 6604 16180 6624
rect 16200 6604 16215 6624
rect 16171 6598 16215 6604
rect 16265 6628 16314 6640
rect 16265 6608 16283 6628
rect 16303 6608 16314 6628
rect 16265 6598 16314 6608
rect 29544 6835 29555 6855
rect 29575 6835 29593 6855
rect 29544 6825 29593 6835
rect 29643 6851 29687 6867
rect 29643 6831 29658 6851
rect 29678 6831 29687 6851
rect 29643 6825 29687 6831
rect 29757 6851 29801 6867
rect 29757 6831 29766 6851
rect 29786 6831 29801 6851
rect 29757 6825 29801 6831
rect 29851 6855 29900 6867
rect 29851 6835 29869 6855
rect 29889 6835 29900 6855
rect 29851 6825 29900 6835
rect 29975 6851 30019 6867
rect 29975 6831 29984 6851
rect 30004 6831 30019 6851
rect 29975 6825 30019 6831
rect 30069 6855 30118 6867
rect 30069 6835 30087 6855
rect 30107 6835 30118 6855
rect 30069 6825 30118 6835
rect 33908 6868 33957 6880
rect 20006 6602 20055 6614
rect 14972 6586 15021 6598
rect 7797 6419 7846 6431
rect 7797 6399 7808 6419
rect 7828 6399 7846 6419
rect 4743 6369 4792 6379
rect 4743 6349 4754 6369
rect 4774 6349 4792 6369
rect 4743 6337 4792 6349
rect 4842 6373 4886 6379
rect 4842 6353 4857 6373
rect 4877 6353 4886 6373
rect 4842 6337 4886 6353
rect 4961 6369 5010 6379
rect 4961 6349 4972 6369
rect 4992 6349 5010 6369
rect 4961 6337 5010 6349
rect 5060 6373 5104 6379
rect 5060 6353 5075 6373
rect 5095 6353 5104 6373
rect 5060 6337 5104 6353
rect 5174 6373 5218 6379
rect 5174 6353 5183 6373
rect 5203 6353 5218 6373
rect 5174 6337 5218 6353
rect 5268 6369 5317 6379
rect 7797 6389 7846 6399
rect 7896 6415 7940 6431
rect 7896 6395 7911 6415
rect 7931 6395 7940 6415
rect 7896 6389 7940 6395
rect 8010 6415 8054 6431
rect 8010 6395 8019 6415
rect 8039 6395 8054 6415
rect 8010 6389 8054 6395
rect 8104 6419 8153 6431
rect 8104 6399 8122 6419
rect 8142 6399 8153 6419
rect 8104 6389 8153 6399
rect 8228 6415 8272 6431
rect 8228 6395 8237 6415
rect 8257 6395 8272 6415
rect 8228 6389 8272 6395
rect 8322 6419 8371 6431
rect 8322 6399 8340 6419
rect 8360 6399 8371 6419
rect 8322 6389 8371 6399
rect 5268 6349 5286 6369
rect 5306 6349 5317 6369
rect 5268 6337 5317 6349
rect 18713 6592 18762 6602
rect 18713 6572 18724 6592
rect 18744 6572 18762 6592
rect 18713 6560 18762 6572
rect 18812 6596 18856 6602
rect 18812 6576 18827 6596
rect 18847 6576 18856 6596
rect 18812 6560 18856 6576
rect 18931 6592 18980 6602
rect 18931 6572 18942 6592
rect 18962 6572 18980 6592
rect 18931 6560 18980 6572
rect 19030 6596 19074 6602
rect 19030 6576 19045 6596
rect 19065 6576 19074 6596
rect 19030 6560 19074 6576
rect 19144 6596 19188 6602
rect 19144 6576 19153 6596
rect 19173 6576 19188 6596
rect 19144 6560 19188 6576
rect 19238 6592 19287 6602
rect 19238 6572 19256 6592
rect 19276 6572 19287 6592
rect 20006 6582 20017 6602
rect 20037 6582 20055 6602
rect 20006 6572 20055 6582
rect 20105 6598 20149 6614
rect 20105 6578 20120 6598
rect 20140 6578 20149 6598
rect 20105 6572 20149 6578
rect 20219 6598 20263 6614
rect 20219 6578 20228 6598
rect 20248 6578 20263 6598
rect 20219 6572 20263 6578
rect 20313 6602 20362 6614
rect 20313 6582 20331 6602
rect 20351 6582 20362 6602
rect 20313 6572 20362 6582
rect 20437 6598 20481 6614
rect 20437 6578 20446 6598
rect 20466 6578 20481 6598
rect 20437 6572 20481 6578
rect 20531 6602 20580 6614
rect 20531 6582 20549 6602
rect 20569 6582 20580 6602
rect 20531 6572 20580 6582
rect 33908 6848 33919 6868
rect 33939 6848 33957 6868
rect 33908 6838 33957 6848
rect 34007 6864 34051 6880
rect 34007 6844 34022 6864
rect 34042 6844 34051 6864
rect 34007 6838 34051 6844
rect 34121 6864 34165 6880
rect 34121 6844 34130 6864
rect 34150 6844 34165 6864
rect 34121 6838 34165 6844
rect 34215 6868 34264 6880
rect 34215 6848 34233 6868
rect 34253 6848 34264 6868
rect 34215 6838 34264 6848
rect 34339 6864 34383 6880
rect 34339 6844 34348 6864
rect 34368 6844 34383 6864
rect 34339 6838 34383 6844
rect 34433 6868 34482 6880
rect 34433 6848 34451 6868
rect 34471 6848 34482 6868
rect 34433 6838 34482 6848
rect 24370 6615 24419 6627
rect 23077 6605 23126 6615
rect 23077 6585 23088 6605
rect 23108 6585 23126 6605
rect 19238 6560 19287 6572
rect 12174 6431 12223 6443
rect 12174 6411 12185 6431
rect 12205 6411 12223 6431
rect 9120 6381 9169 6391
rect 9120 6361 9131 6381
rect 9151 6361 9169 6381
rect 9120 6349 9169 6361
rect 9219 6385 9263 6391
rect 9219 6365 9234 6385
rect 9254 6365 9263 6385
rect 9219 6349 9263 6365
rect 9338 6381 9387 6391
rect 9338 6361 9349 6381
rect 9369 6361 9387 6381
rect 9338 6349 9387 6361
rect 9437 6385 9481 6391
rect 9437 6365 9452 6385
rect 9472 6365 9481 6385
rect 9437 6349 9481 6365
rect 9551 6385 9595 6391
rect 9551 6365 9560 6385
rect 9580 6365 9595 6385
rect 9551 6349 9595 6365
rect 9645 6381 9694 6391
rect 12174 6401 12223 6411
rect 12273 6427 12317 6443
rect 12273 6407 12288 6427
rect 12308 6407 12317 6427
rect 12273 6401 12317 6407
rect 12387 6427 12431 6443
rect 12387 6407 12396 6427
rect 12416 6407 12431 6427
rect 12387 6401 12431 6407
rect 12481 6431 12530 6443
rect 12481 6411 12499 6431
rect 12519 6411 12530 6431
rect 12481 6401 12530 6411
rect 12605 6427 12649 6443
rect 12605 6407 12614 6427
rect 12634 6407 12649 6427
rect 12605 6401 12649 6407
rect 12699 6431 12748 6443
rect 12699 6411 12717 6431
rect 12737 6411 12748 6431
rect 12699 6401 12748 6411
rect 9645 6361 9663 6381
rect 9683 6361 9694 6381
rect 9645 6349 9694 6361
rect 1177 6172 1226 6182
rect 1177 6152 1188 6172
rect 1208 6152 1226 6172
rect 1177 6140 1226 6152
rect 1276 6176 1320 6182
rect 1276 6156 1291 6176
rect 1311 6156 1320 6176
rect 1276 6140 1320 6156
rect 1395 6172 1444 6182
rect 1395 6152 1406 6172
rect 1426 6152 1444 6172
rect 1395 6140 1444 6152
rect 1494 6176 1538 6182
rect 1494 6156 1509 6176
rect 1529 6156 1538 6176
rect 1494 6140 1538 6156
rect 1608 6176 1652 6182
rect 1608 6156 1617 6176
rect 1637 6156 1652 6176
rect 1608 6140 1652 6156
rect 1702 6172 1751 6182
rect 1702 6152 1720 6172
rect 1740 6152 1751 6172
rect 1702 6140 1751 6152
rect 2536 6180 2585 6192
rect 2536 6160 2547 6180
rect 2567 6160 2585 6180
rect 2536 6150 2585 6160
rect 2635 6176 2679 6192
rect 2635 6156 2650 6176
rect 2670 6156 2679 6176
rect 2635 6150 2679 6156
rect 2749 6176 2793 6192
rect 2749 6156 2758 6176
rect 2778 6156 2793 6176
rect 2749 6150 2793 6156
rect 2843 6180 2892 6192
rect 2843 6160 2861 6180
rect 2881 6160 2892 6180
rect 2843 6150 2892 6160
rect 2967 6176 3011 6192
rect 2967 6156 2976 6176
rect 2996 6156 3011 6176
rect 2967 6150 3011 6156
rect 3061 6180 3110 6192
rect 16538 6444 16587 6456
rect 16538 6424 16549 6444
rect 16569 6424 16587 6444
rect 13484 6394 13533 6404
rect 13484 6374 13495 6394
rect 13515 6374 13533 6394
rect 13484 6362 13533 6374
rect 13583 6398 13627 6404
rect 13583 6378 13598 6398
rect 13618 6378 13627 6398
rect 13583 6362 13627 6378
rect 13702 6394 13751 6404
rect 13702 6374 13713 6394
rect 13733 6374 13751 6394
rect 13702 6362 13751 6374
rect 13801 6398 13845 6404
rect 13801 6378 13816 6398
rect 13836 6378 13845 6398
rect 13801 6362 13845 6378
rect 13915 6398 13959 6404
rect 13915 6378 13924 6398
rect 13944 6378 13959 6398
rect 13915 6362 13959 6378
rect 14009 6394 14058 6404
rect 16538 6414 16587 6424
rect 16637 6440 16681 6456
rect 16637 6420 16652 6440
rect 16672 6420 16681 6440
rect 16637 6414 16681 6420
rect 16751 6440 16795 6456
rect 16751 6420 16760 6440
rect 16780 6420 16795 6440
rect 16751 6414 16795 6420
rect 16845 6444 16894 6456
rect 16845 6424 16863 6444
rect 16883 6424 16894 6444
rect 16845 6414 16894 6424
rect 16969 6440 17013 6456
rect 16969 6420 16978 6440
rect 16998 6420 17013 6440
rect 16969 6414 17013 6420
rect 17063 6444 17112 6456
rect 17063 6424 17081 6444
rect 17101 6424 17112 6444
rect 17063 6414 17112 6424
rect 23077 6573 23126 6585
rect 23176 6609 23220 6615
rect 23176 6589 23191 6609
rect 23211 6589 23220 6609
rect 23176 6573 23220 6589
rect 23295 6605 23344 6615
rect 23295 6585 23306 6605
rect 23326 6585 23344 6605
rect 23295 6573 23344 6585
rect 23394 6609 23438 6615
rect 23394 6589 23409 6609
rect 23429 6589 23438 6609
rect 23394 6573 23438 6589
rect 23508 6609 23552 6615
rect 23508 6589 23517 6609
rect 23537 6589 23552 6609
rect 23508 6573 23552 6589
rect 23602 6605 23651 6615
rect 23602 6585 23620 6605
rect 23640 6585 23651 6605
rect 24370 6595 24381 6615
rect 24401 6595 24419 6615
rect 24370 6585 24419 6595
rect 24469 6611 24513 6627
rect 24469 6591 24484 6611
rect 24504 6591 24513 6611
rect 24469 6585 24513 6591
rect 24583 6611 24627 6627
rect 24583 6591 24592 6611
rect 24612 6591 24627 6611
rect 24583 6585 24627 6591
rect 24677 6615 24726 6627
rect 24677 6595 24695 6615
rect 24715 6595 24726 6615
rect 24677 6585 24726 6595
rect 24801 6611 24845 6627
rect 24801 6591 24810 6611
rect 24830 6591 24845 6611
rect 24801 6585 24845 6591
rect 24895 6615 24944 6627
rect 24895 6595 24913 6615
rect 24933 6595 24944 6615
rect 24895 6585 24944 6595
rect 28747 6627 28796 6639
rect 27454 6617 27503 6627
rect 27454 6597 27465 6617
rect 27485 6597 27503 6617
rect 23602 6573 23651 6585
rect 14009 6374 14027 6394
rect 14047 6374 14058 6394
rect 14009 6362 14058 6374
rect 3061 6160 3079 6180
rect 3099 6160 3110 6180
rect 3061 6150 3110 6160
rect 5541 6185 5590 6195
rect 5541 6165 5552 6185
rect 5572 6165 5590 6185
rect 5541 6153 5590 6165
rect 5640 6189 5684 6195
rect 5640 6169 5655 6189
rect 5675 6169 5684 6189
rect 5640 6153 5684 6169
rect 5759 6185 5808 6195
rect 5759 6165 5770 6185
rect 5790 6165 5808 6185
rect 5759 6153 5808 6165
rect 5858 6189 5902 6195
rect 5858 6169 5873 6189
rect 5893 6169 5902 6189
rect 5858 6153 5902 6169
rect 5972 6189 6016 6195
rect 5972 6169 5981 6189
rect 6001 6169 6016 6189
rect 5972 6153 6016 6169
rect 6066 6185 6115 6195
rect 6066 6165 6084 6185
rect 6104 6165 6115 6185
rect 6066 6153 6115 6165
rect 6900 6193 6949 6205
rect 6900 6173 6911 6193
rect 6931 6173 6949 6193
rect 6900 6163 6949 6173
rect 6999 6189 7043 6205
rect 6999 6169 7014 6189
rect 7034 6169 7043 6189
rect 6999 6163 7043 6169
rect 7113 6189 7157 6205
rect 7113 6169 7122 6189
rect 7142 6169 7157 6189
rect 7113 6163 7157 6169
rect 7207 6193 7256 6205
rect 7207 6173 7225 6193
rect 7245 6173 7256 6193
rect 7207 6163 7256 6173
rect 7331 6189 7375 6205
rect 7331 6169 7340 6189
rect 7360 6169 7375 6189
rect 7331 6163 7375 6169
rect 7425 6193 7474 6205
rect 27454 6585 27503 6597
rect 27553 6621 27597 6627
rect 27553 6601 27568 6621
rect 27588 6601 27597 6621
rect 27553 6585 27597 6601
rect 27672 6617 27721 6627
rect 27672 6597 27683 6617
rect 27703 6597 27721 6617
rect 27672 6585 27721 6597
rect 27771 6621 27815 6627
rect 27771 6601 27786 6621
rect 27806 6601 27815 6621
rect 27771 6585 27815 6601
rect 27885 6621 27929 6627
rect 27885 6601 27894 6621
rect 27914 6601 27929 6621
rect 27885 6585 27929 6601
rect 27979 6617 28028 6627
rect 27979 6597 27997 6617
rect 28017 6597 28028 6617
rect 28747 6607 28758 6627
rect 28778 6607 28796 6627
rect 28747 6597 28796 6607
rect 28846 6623 28890 6639
rect 28846 6603 28861 6623
rect 28881 6603 28890 6623
rect 28846 6597 28890 6603
rect 28960 6623 29004 6639
rect 28960 6603 28969 6623
rect 28989 6603 29004 6623
rect 28960 6597 29004 6603
rect 29054 6627 29103 6639
rect 29054 6607 29072 6627
rect 29092 6607 29103 6627
rect 29054 6597 29103 6607
rect 29178 6623 29222 6639
rect 29178 6603 29187 6623
rect 29207 6603 29222 6623
rect 29178 6597 29222 6603
rect 29272 6627 29321 6639
rect 29272 6607 29290 6627
rect 29310 6607 29321 6627
rect 29272 6597 29321 6607
rect 33111 6640 33160 6652
rect 31818 6630 31867 6640
rect 31818 6610 31829 6630
rect 31849 6610 31867 6630
rect 27979 6585 28028 6597
rect 20804 6418 20853 6430
rect 20804 6398 20815 6418
rect 20835 6398 20853 6418
rect 7425 6173 7443 6193
rect 7463 6173 7474 6193
rect 7425 6163 7474 6173
rect 9918 6197 9967 6207
rect 9918 6177 9929 6197
rect 9949 6177 9967 6197
rect 9918 6165 9967 6177
rect 10017 6201 10061 6207
rect 10017 6181 10032 6201
rect 10052 6181 10061 6201
rect 10017 6165 10061 6181
rect 10136 6197 10185 6207
rect 10136 6177 10147 6197
rect 10167 6177 10185 6197
rect 10136 6165 10185 6177
rect 10235 6201 10279 6207
rect 10235 6181 10250 6201
rect 10270 6181 10279 6201
rect 10235 6165 10279 6181
rect 10349 6201 10393 6207
rect 10349 6181 10358 6201
rect 10378 6181 10393 6201
rect 10349 6165 10393 6181
rect 10443 6197 10492 6207
rect 10443 6177 10461 6197
rect 10481 6177 10492 6197
rect 10443 6165 10492 6177
rect 11277 6205 11326 6217
rect 11277 6185 11288 6205
rect 11308 6185 11326 6205
rect 11277 6175 11326 6185
rect 11376 6201 11420 6217
rect 11376 6181 11391 6201
rect 11411 6181 11420 6201
rect 11376 6175 11420 6181
rect 11490 6201 11534 6217
rect 11490 6181 11499 6201
rect 11519 6181 11534 6201
rect 11490 6175 11534 6181
rect 11584 6205 11633 6217
rect 11584 6185 11602 6205
rect 11622 6185 11633 6205
rect 11584 6175 11633 6185
rect 11708 6201 11752 6217
rect 11708 6181 11717 6201
rect 11737 6181 11752 6201
rect 11708 6175 11752 6181
rect 11802 6205 11851 6217
rect 17750 6368 17799 6378
rect 17750 6348 17761 6368
rect 17781 6348 17799 6368
rect 17750 6336 17799 6348
rect 17849 6372 17893 6378
rect 17849 6352 17864 6372
rect 17884 6352 17893 6372
rect 17849 6336 17893 6352
rect 17968 6368 18017 6378
rect 17968 6348 17979 6368
rect 17999 6348 18017 6368
rect 17968 6336 18017 6348
rect 18067 6372 18111 6378
rect 18067 6352 18082 6372
rect 18102 6352 18111 6372
rect 18067 6336 18111 6352
rect 18181 6372 18225 6378
rect 18181 6352 18190 6372
rect 18210 6352 18225 6372
rect 18181 6336 18225 6352
rect 18275 6368 18324 6378
rect 20804 6388 20853 6398
rect 20903 6414 20947 6430
rect 20903 6394 20918 6414
rect 20938 6394 20947 6414
rect 20903 6388 20947 6394
rect 21017 6414 21061 6430
rect 21017 6394 21026 6414
rect 21046 6394 21061 6414
rect 21017 6388 21061 6394
rect 21111 6418 21160 6430
rect 21111 6398 21129 6418
rect 21149 6398 21160 6418
rect 21111 6388 21160 6398
rect 21235 6414 21279 6430
rect 21235 6394 21244 6414
rect 21264 6394 21279 6414
rect 21235 6388 21279 6394
rect 21329 6418 21378 6430
rect 21329 6398 21347 6418
rect 21367 6398 21378 6418
rect 21329 6388 21378 6398
rect 18275 6348 18293 6368
rect 18313 6348 18324 6368
rect 18275 6336 18324 6348
rect 31818 6598 31867 6610
rect 31917 6634 31961 6640
rect 31917 6614 31932 6634
rect 31952 6614 31961 6634
rect 31917 6598 31961 6614
rect 32036 6630 32085 6640
rect 32036 6610 32047 6630
rect 32067 6610 32085 6630
rect 32036 6598 32085 6610
rect 32135 6634 32179 6640
rect 32135 6614 32150 6634
rect 32170 6614 32179 6634
rect 32135 6598 32179 6614
rect 32249 6634 32293 6640
rect 32249 6614 32258 6634
rect 32278 6614 32293 6634
rect 32249 6598 32293 6614
rect 32343 6630 32392 6640
rect 32343 6610 32361 6630
rect 32381 6610 32392 6630
rect 33111 6620 33122 6640
rect 33142 6620 33160 6640
rect 33111 6610 33160 6620
rect 33210 6636 33254 6652
rect 33210 6616 33225 6636
rect 33245 6616 33254 6636
rect 33210 6610 33254 6616
rect 33324 6636 33368 6652
rect 33324 6616 33333 6636
rect 33353 6616 33368 6636
rect 33324 6610 33368 6616
rect 33418 6640 33467 6652
rect 33418 6620 33436 6640
rect 33456 6620 33467 6640
rect 33418 6610 33467 6620
rect 33542 6636 33586 6652
rect 33542 6616 33551 6636
rect 33571 6616 33586 6636
rect 33542 6610 33586 6616
rect 33636 6640 33685 6652
rect 33636 6620 33654 6640
rect 33674 6620 33685 6640
rect 33636 6610 33685 6620
rect 32343 6598 32392 6610
rect 25168 6431 25217 6443
rect 25168 6411 25179 6431
rect 25199 6411 25217 6431
rect 22114 6381 22163 6391
rect 22114 6361 22125 6381
rect 22145 6361 22163 6381
rect 22114 6349 22163 6361
rect 22213 6385 22257 6391
rect 22213 6365 22228 6385
rect 22248 6365 22257 6385
rect 22213 6349 22257 6365
rect 22332 6381 22381 6391
rect 22332 6361 22343 6381
rect 22363 6361 22381 6381
rect 22332 6349 22381 6361
rect 22431 6385 22475 6391
rect 22431 6365 22446 6385
rect 22466 6365 22475 6385
rect 22431 6349 22475 6365
rect 22545 6385 22589 6391
rect 22545 6365 22554 6385
rect 22574 6365 22589 6385
rect 22545 6349 22589 6365
rect 22639 6381 22688 6391
rect 25168 6401 25217 6411
rect 25267 6427 25311 6443
rect 25267 6407 25282 6427
rect 25302 6407 25311 6427
rect 25267 6401 25311 6407
rect 25381 6427 25425 6443
rect 25381 6407 25390 6427
rect 25410 6407 25425 6427
rect 25381 6401 25425 6407
rect 25475 6431 25524 6443
rect 25475 6411 25493 6431
rect 25513 6411 25524 6431
rect 25475 6401 25524 6411
rect 25599 6427 25643 6443
rect 25599 6407 25608 6427
rect 25628 6407 25643 6427
rect 25599 6401 25643 6407
rect 25693 6431 25742 6443
rect 25693 6411 25711 6431
rect 25731 6411 25742 6431
rect 25693 6401 25742 6411
rect 22639 6361 22657 6381
rect 22677 6361 22688 6381
rect 22639 6349 22688 6361
rect 11802 6185 11820 6205
rect 11840 6185 11851 6205
rect 11802 6175 11851 6185
rect 14282 6210 14331 6220
rect 14282 6190 14293 6210
rect 14313 6190 14331 6210
rect 380 5944 429 5954
rect 380 5924 391 5944
rect 411 5924 429 5944
rect 380 5912 429 5924
rect 479 5948 523 5954
rect 479 5928 494 5948
rect 514 5928 523 5948
rect 479 5912 523 5928
rect 598 5944 647 5954
rect 598 5924 609 5944
rect 629 5924 647 5944
rect 598 5912 647 5924
rect 697 5948 741 5954
rect 697 5928 712 5948
rect 732 5928 741 5948
rect 697 5912 741 5928
rect 811 5948 855 5954
rect 811 5928 820 5948
rect 840 5928 855 5948
rect 811 5912 855 5928
rect 905 5944 954 5954
rect 905 5924 923 5944
rect 943 5924 954 5944
rect 14282 6178 14331 6190
rect 14381 6214 14425 6220
rect 14381 6194 14396 6214
rect 14416 6194 14425 6214
rect 14381 6178 14425 6194
rect 14500 6210 14549 6220
rect 14500 6190 14511 6210
rect 14531 6190 14549 6210
rect 14500 6178 14549 6190
rect 14599 6214 14643 6220
rect 14599 6194 14614 6214
rect 14634 6194 14643 6214
rect 14599 6178 14643 6194
rect 14713 6214 14757 6220
rect 14713 6194 14722 6214
rect 14742 6194 14757 6214
rect 14713 6178 14757 6194
rect 14807 6210 14856 6220
rect 14807 6190 14825 6210
rect 14845 6190 14856 6210
rect 14807 6178 14856 6190
rect 15641 6218 15690 6230
rect 15641 6198 15652 6218
rect 15672 6198 15690 6218
rect 15641 6188 15690 6198
rect 15740 6214 15784 6230
rect 15740 6194 15755 6214
rect 15775 6194 15784 6214
rect 15740 6188 15784 6194
rect 15854 6214 15898 6230
rect 15854 6194 15863 6214
rect 15883 6194 15898 6214
rect 15854 6188 15898 6194
rect 15948 6218 15997 6230
rect 15948 6198 15966 6218
rect 15986 6198 15997 6218
rect 15948 6188 15997 6198
rect 16072 6214 16116 6230
rect 16072 6194 16081 6214
rect 16101 6194 16116 6214
rect 16072 6188 16116 6194
rect 16166 6218 16215 6230
rect 16166 6198 16184 6218
rect 16204 6198 16215 6218
rect 16166 6188 16215 6198
rect 29545 6443 29594 6455
rect 29545 6423 29556 6443
rect 29576 6423 29594 6443
rect 26491 6393 26540 6403
rect 26491 6373 26502 6393
rect 26522 6373 26540 6393
rect 26491 6361 26540 6373
rect 26590 6397 26634 6403
rect 26590 6377 26605 6397
rect 26625 6377 26634 6397
rect 26590 6361 26634 6377
rect 26709 6393 26758 6403
rect 26709 6373 26720 6393
rect 26740 6373 26758 6393
rect 26709 6361 26758 6373
rect 26808 6397 26852 6403
rect 26808 6377 26823 6397
rect 26843 6377 26852 6397
rect 26808 6361 26852 6377
rect 26922 6397 26966 6403
rect 26922 6377 26931 6397
rect 26951 6377 26966 6397
rect 26922 6361 26966 6377
rect 27016 6393 27065 6403
rect 29545 6413 29594 6423
rect 29644 6439 29688 6455
rect 29644 6419 29659 6439
rect 29679 6419 29688 6439
rect 29644 6413 29688 6419
rect 29758 6439 29802 6455
rect 29758 6419 29767 6439
rect 29787 6419 29802 6439
rect 29758 6413 29802 6419
rect 29852 6443 29901 6455
rect 29852 6423 29870 6443
rect 29890 6423 29901 6443
rect 29852 6413 29901 6423
rect 29976 6439 30020 6455
rect 29976 6419 29985 6439
rect 30005 6419 30020 6439
rect 29976 6413 30020 6419
rect 30070 6443 30119 6455
rect 30070 6423 30088 6443
rect 30108 6423 30119 6443
rect 30070 6413 30119 6423
rect 27016 6373 27034 6393
rect 27054 6373 27065 6393
rect 27016 6361 27065 6373
rect 905 5912 954 5924
rect 4744 5957 4793 5967
rect 4744 5937 4755 5957
rect 4775 5937 4793 5957
rect 4744 5925 4793 5937
rect 4843 5961 4887 5967
rect 4843 5941 4858 5961
rect 4878 5941 4887 5961
rect 4843 5925 4887 5941
rect 4962 5957 5011 5967
rect 4962 5937 4973 5957
rect 4993 5937 5011 5957
rect 4962 5925 5011 5937
rect 5061 5961 5105 5967
rect 5061 5941 5076 5961
rect 5096 5941 5105 5961
rect 5061 5925 5105 5941
rect 5175 5961 5219 5967
rect 5175 5941 5184 5961
rect 5204 5941 5219 5961
rect 5175 5925 5219 5941
rect 5269 5957 5318 5967
rect 5269 5937 5287 5957
rect 5307 5937 5318 5957
rect 18548 6184 18597 6194
rect 18548 6164 18559 6184
rect 18579 6164 18597 6184
rect 18548 6152 18597 6164
rect 18647 6188 18691 6194
rect 18647 6168 18662 6188
rect 18682 6168 18691 6188
rect 18647 6152 18691 6168
rect 18766 6184 18815 6194
rect 18766 6164 18777 6184
rect 18797 6164 18815 6184
rect 18766 6152 18815 6164
rect 18865 6188 18909 6194
rect 18865 6168 18880 6188
rect 18900 6168 18909 6188
rect 18865 6152 18909 6168
rect 18979 6188 19023 6194
rect 18979 6168 18988 6188
rect 19008 6168 19023 6188
rect 18979 6152 19023 6168
rect 19073 6184 19122 6194
rect 19073 6164 19091 6184
rect 19111 6164 19122 6184
rect 19073 6152 19122 6164
rect 19907 6192 19956 6204
rect 19907 6172 19918 6192
rect 19938 6172 19956 6192
rect 19907 6162 19956 6172
rect 20006 6188 20050 6204
rect 20006 6168 20021 6188
rect 20041 6168 20050 6188
rect 20006 6162 20050 6168
rect 20120 6188 20164 6204
rect 20120 6168 20129 6188
rect 20149 6168 20164 6188
rect 20120 6162 20164 6168
rect 20214 6192 20263 6204
rect 20214 6172 20232 6192
rect 20252 6172 20263 6192
rect 20214 6162 20263 6172
rect 20338 6188 20382 6204
rect 20338 6168 20347 6188
rect 20367 6168 20382 6188
rect 20338 6162 20382 6168
rect 20432 6192 20481 6204
rect 33909 6456 33958 6468
rect 33909 6436 33920 6456
rect 33940 6436 33958 6456
rect 30855 6406 30904 6416
rect 30855 6386 30866 6406
rect 30886 6386 30904 6406
rect 30855 6374 30904 6386
rect 30954 6410 30998 6416
rect 30954 6390 30969 6410
rect 30989 6390 30998 6410
rect 30954 6374 30998 6390
rect 31073 6406 31122 6416
rect 31073 6386 31084 6406
rect 31104 6386 31122 6406
rect 31073 6374 31122 6386
rect 31172 6410 31216 6416
rect 31172 6390 31187 6410
rect 31207 6390 31216 6410
rect 31172 6374 31216 6390
rect 31286 6410 31330 6416
rect 31286 6390 31295 6410
rect 31315 6390 31330 6410
rect 31286 6374 31330 6390
rect 31380 6406 31429 6416
rect 33909 6426 33958 6436
rect 34008 6452 34052 6468
rect 34008 6432 34023 6452
rect 34043 6432 34052 6452
rect 34008 6426 34052 6432
rect 34122 6452 34166 6468
rect 34122 6432 34131 6452
rect 34151 6432 34166 6452
rect 34122 6426 34166 6432
rect 34216 6456 34265 6468
rect 34216 6436 34234 6456
rect 34254 6436 34265 6456
rect 34216 6426 34265 6436
rect 34340 6452 34384 6468
rect 34340 6432 34349 6452
rect 34369 6432 34384 6452
rect 34340 6426 34384 6432
rect 34434 6456 34483 6468
rect 34434 6436 34452 6456
rect 34472 6436 34483 6456
rect 34434 6426 34483 6436
rect 31380 6386 31398 6406
rect 31418 6386 31429 6406
rect 31380 6374 31429 6386
rect 20432 6172 20450 6192
rect 20470 6172 20481 6192
rect 20432 6162 20481 6172
rect 22912 6197 22961 6207
rect 22912 6177 22923 6197
rect 22943 6177 22961 6197
rect 5269 5925 5318 5937
rect 9121 5969 9170 5979
rect 9121 5949 9132 5969
rect 9152 5949 9170 5969
rect 9121 5937 9170 5949
rect 9220 5973 9264 5979
rect 9220 5953 9235 5973
rect 9255 5953 9264 5973
rect 9220 5937 9264 5953
rect 9339 5969 9388 5979
rect 9339 5949 9350 5969
rect 9370 5949 9388 5969
rect 9339 5937 9388 5949
rect 9438 5973 9482 5979
rect 9438 5953 9453 5973
rect 9473 5953 9482 5973
rect 9438 5937 9482 5953
rect 9552 5973 9596 5979
rect 9552 5953 9561 5973
rect 9581 5953 9596 5973
rect 9552 5937 9596 5953
rect 9646 5969 9695 5979
rect 9646 5949 9664 5969
rect 9684 5949 9695 5969
rect 22912 6165 22961 6177
rect 23011 6201 23055 6207
rect 23011 6181 23026 6201
rect 23046 6181 23055 6201
rect 23011 6165 23055 6181
rect 23130 6197 23179 6207
rect 23130 6177 23141 6197
rect 23161 6177 23179 6197
rect 23130 6165 23179 6177
rect 23229 6201 23273 6207
rect 23229 6181 23244 6201
rect 23264 6181 23273 6201
rect 23229 6165 23273 6181
rect 23343 6201 23387 6207
rect 23343 6181 23352 6201
rect 23372 6181 23387 6201
rect 23343 6165 23387 6181
rect 23437 6197 23486 6207
rect 23437 6177 23455 6197
rect 23475 6177 23486 6197
rect 23437 6165 23486 6177
rect 24271 6205 24320 6217
rect 24271 6185 24282 6205
rect 24302 6185 24320 6205
rect 24271 6175 24320 6185
rect 24370 6201 24414 6217
rect 24370 6181 24385 6201
rect 24405 6181 24414 6201
rect 24370 6175 24414 6181
rect 24484 6201 24528 6217
rect 24484 6181 24493 6201
rect 24513 6181 24528 6201
rect 24484 6175 24528 6181
rect 24578 6205 24627 6217
rect 24578 6185 24596 6205
rect 24616 6185 24627 6205
rect 24578 6175 24627 6185
rect 24702 6201 24746 6217
rect 24702 6181 24711 6201
rect 24731 6181 24746 6201
rect 24702 6175 24746 6181
rect 24796 6205 24845 6217
rect 24796 6185 24814 6205
rect 24834 6185 24845 6205
rect 24796 6175 24845 6185
rect 9646 5937 9695 5949
rect 13485 5982 13534 5992
rect 13485 5962 13496 5982
rect 13516 5962 13534 5982
rect 13485 5950 13534 5962
rect 13584 5986 13628 5992
rect 13584 5966 13599 5986
rect 13619 5966 13628 5986
rect 13584 5950 13628 5966
rect 13703 5982 13752 5992
rect 13703 5962 13714 5982
rect 13734 5962 13752 5982
rect 13703 5950 13752 5962
rect 13802 5986 13846 5992
rect 13802 5966 13817 5986
rect 13837 5966 13846 5986
rect 13802 5950 13846 5966
rect 13916 5986 13960 5992
rect 13916 5966 13925 5986
rect 13945 5966 13960 5986
rect 13916 5950 13960 5966
rect 14010 5982 14059 5992
rect 14010 5962 14028 5982
rect 14048 5962 14059 5982
rect 14010 5950 14059 5962
rect 27289 6209 27338 6219
rect 27289 6189 27300 6209
rect 27320 6189 27338 6209
rect 27289 6177 27338 6189
rect 27388 6213 27432 6219
rect 27388 6193 27403 6213
rect 27423 6193 27432 6213
rect 27388 6177 27432 6193
rect 27507 6209 27556 6219
rect 27507 6189 27518 6209
rect 27538 6189 27556 6209
rect 27507 6177 27556 6189
rect 27606 6213 27650 6219
rect 27606 6193 27621 6213
rect 27641 6193 27650 6213
rect 27606 6177 27650 6193
rect 27720 6213 27764 6219
rect 27720 6193 27729 6213
rect 27749 6193 27764 6213
rect 27720 6177 27764 6193
rect 27814 6209 27863 6219
rect 27814 6189 27832 6209
rect 27852 6189 27863 6209
rect 27814 6177 27863 6189
rect 28648 6217 28697 6229
rect 28648 6197 28659 6217
rect 28679 6197 28697 6217
rect 28648 6187 28697 6197
rect 28747 6213 28791 6229
rect 28747 6193 28762 6213
rect 28782 6193 28791 6213
rect 28747 6187 28791 6193
rect 28861 6213 28905 6229
rect 28861 6193 28870 6213
rect 28890 6193 28905 6213
rect 28861 6187 28905 6193
rect 28955 6217 29004 6229
rect 28955 6197 28973 6217
rect 28993 6197 29004 6217
rect 28955 6187 29004 6197
rect 29079 6213 29123 6229
rect 29079 6193 29088 6213
rect 29108 6193 29123 6213
rect 29079 6187 29123 6193
rect 29173 6217 29222 6229
rect 29173 6197 29191 6217
rect 29211 6197 29222 6217
rect 29173 6187 29222 6197
rect 31653 6222 31702 6232
rect 31653 6202 31664 6222
rect 31684 6202 31702 6222
rect 17751 5956 17800 5966
rect 17751 5936 17762 5956
rect 17782 5936 17800 5956
rect 17751 5924 17800 5936
rect 17850 5960 17894 5966
rect 17850 5940 17865 5960
rect 17885 5940 17894 5960
rect 17850 5924 17894 5940
rect 17969 5956 18018 5966
rect 17969 5936 17980 5956
rect 18000 5936 18018 5956
rect 17969 5924 18018 5936
rect 18068 5960 18112 5966
rect 18068 5940 18083 5960
rect 18103 5940 18112 5960
rect 18068 5924 18112 5940
rect 18182 5960 18226 5966
rect 18182 5940 18191 5960
rect 18211 5940 18226 5960
rect 18182 5924 18226 5940
rect 18276 5956 18325 5966
rect 18276 5936 18294 5956
rect 18314 5936 18325 5956
rect 31653 6190 31702 6202
rect 31752 6226 31796 6232
rect 31752 6206 31767 6226
rect 31787 6206 31796 6226
rect 31752 6190 31796 6206
rect 31871 6222 31920 6232
rect 31871 6202 31882 6222
rect 31902 6202 31920 6222
rect 31871 6190 31920 6202
rect 31970 6226 32014 6232
rect 31970 6206 31985 6226
rect 32005 6206 32014 6226
rect 31970 6190 32014 6206
rect 32084 6226 32128 6232
rect 32084 6206 32093 6226
rect 32113 6206 32128 6226
rect 32084 6190 32128 6206
rect 32178 6222 32227 6232
rect 32178 6202 32196 6222
rect 32216 6202 32227 6222
rect 32178 6190 32227 6202
rect 33012 6230 33061 6242
rect 33012 6210 33023 6230
rect 33043 6210 33061 6230
rect 33012 6200 33061 6210
rect 33111 6226 33155 6242
rect 33111 6206 33126 6226
rect 33146 6206 33155 6226
rect 33111 6200 33155 6206
rect 33225 6226 33269 6242
rect 33225 6206 33234 6226
rect 33254 6206 33269 6226
rect 33225 6200 33269 6206
rect 33319 6230 33368 6242
rect 33319 6210 33337 6230
rect 33357 6210 33368 6230
rect 33319 6200 33368 6210
rect 33443 6226 33487 6242
rect 33443 6206 33452 6226
rect 33472 6206 33487 6226
rect 33443 6200 33487 6206
rect 33537 6230 33586 6242
rect 33537 6210 33555 6230
rect 33575 6210 33586 6230
rect 33537 6200 33586 6210
rect 18276 5924 18325 5936
rect 22115 5969 22164 5979
rect 22115 5949 22126 5969
rect 22146 5949 22164 5969
rect 22115 5937 22164 5949
rect 22214 5973 22258 5979
rect 22214 5953 22229 5973
rect 22249 5953 22258 5973
rect 22214 5937 22258 5953
rect 22333 5969 22382 5979
rect 22333 5949 22344 5969
rect 22364 5949 22382 5969
rect 22333 5937 22382 5949
rect 22432 5973 22476 5979
rect 22432 5953 22447 5973
rect 22467 5953 22476 5973
rect 22432 5937 22476 5953
rect 22546 5973 22590 5979
rect 22546 5953 22555 5973
rect 22575 5953 22590 5973
rect 22546 5937 22590 5953
rect 22640 5969 22689 5979
rect 22640 5949 22658 5969
rect 22678 5949 22689 5969
rect 22640 5937 22689 5949
rect 26492 5981 26541 5991
rect 26492 5961 26503 5981
rect 26523 5961 26541 5981
rect 26492 5949 26541 5961
rect 26591 5985 26635 5991
rect 26591 5965 26606 5985
rect 26626 5965 26635 5985
rect 26591 5949 26635 5965
rect 26710 5981 26759 5991
rect 26710 5961 26721 5981
rect 26741 5961 26759 5981
rect 26710 5949 26759 5961
rect 26809 5985 26853 5991
rect 26809 5965 26824 5985
rect 26844 5965 26853 5985
rect 26809 5949 26853 5965
rect 26923 5985 26967 5991
rect 26923 5965 26932 5985
rect 26952 5965 26967 5985
rect 26923 5949 26967 5965
rect 27017 5981 27066 5991
rect 27017 5961 27035 5981
rect 27055 5961 27066 5981
rect 27017 5949 27066 5961
rect 30856 5994 30905 6004
rect 30856 5974 30867 5994
rect 30887 5974 30905 5994
rect 30856 5962 30905 5974
rect 30955 5998 30999 6004
rect 30955 5978 30970 5998
rect 30990 5978 30999 5998
rect 30955 5962 30999 5978
rect 31074 5994 31123 6004
rect 31074 5974 31085 5994
rect 31105 5974 31123 5994
rect 31074 5962 31123 5974
rect 31173 5998 31217 6004
rect 31173 5978 31188 5998
rect 31208 5978 31217 5998
rect 31173 5962 31217 5978
rect 31287 5998 31331 6004
rect 31287 5978 31296 5998
rect 31316 5978 31331 5998
rect 31287 5962 31331 5978
rect 31381 5994 31430 6004
rect 31381 5974 31399 5994
rect 31419 5974 31430 5994
rect 31381 5962 31430 5974
rect 3415 5800 3464 5812
rect 3415 5780 3426 5800
rect 3446 5780 3464 5800
rect 3415 5770 3464 5780
rect 3514 5796 3558 5812
rect 3514 5776 3529 5796
rect 3549 5776 3558 5796
rect 3514 5770 3558 5776
rect 3628 5796 3672 5812
rect 3628 5776 3637 5796
rect 3657 5776 3672 5796
rect 3628 5770 3672 5776
rect 3722 5800 3771 5812
rect 3722 5780 3740 5800
rect 3760 5780 3771 5800
rect 3722 5770 3771 5780
rect 3846 5796 3890 5812
rect 3846 5776 3855 5796
rect 3875 5776 3890 5796
rect 3846 5770 3890 5776
rect 3940 5800 3989 5812
rect 3940 5780 3958 5800
rect 3978 5780 3989 5800
rect 3940 5770 3989 5780
rect 7779 5813 7828 5825
rect 7779 5793 7790 5813
rect 7810 5793 7828 5813
rect 7779 5783 7828 5793
rect 7878 5809 7922 5825
rect 7878 5789 7893 5809
rect 7913 5789 7922 5809
rect 7878 5783 7922 5789
rect 7992 5809 8036 5825
rect 7992 5789 8001 5809
rect 8021 5789 8036 5809
rect 7992 5783 8036 5789
rect 8086 5813 8135 5825
rect 8086 5793 8104 5813
rect 8124 5793 8135 5813
rect 8086 5783 8135 5793
rect 8210 5809 8254 5825
rect 8210 5789 8219 5809
rect 8239 5789 8254 5809
rect 8210 5783 8254 5789
rect 8304 5813 8353 5825
rect 8304 5793 8322 5813
rect 8342 5793 8353 5813
rect 8304 5783 8353 5793
rect 12156 5825 12205 5837
rect 12156 5805 12167 5825
rect 12187 5805 12205 5825
rect 12156 5795 12205 5805
rect 12255 5821 12299 5837
rect 12255 5801 12270 5821
rect 12290 5801 12299 5821
rect 12255 5795 12299 5801
rect 12369 5821 12413 5837
rect 12369 5801 12378 5821
rect 12398 5801 12413 5821
rect 12369 5795 12413 5801
rect 12463 5825 12512 5837
rect 12463 5805 12481 5825
rect 12501 5805 12512 5825
rect 12463 5795 12512 5805
rect 12587 5821 12631 5837
rect 12587 5801 12596 5821
rect 12616 5801 12631 5821
rect 12587 5795 12631 5801
rect 12681 5825 12730 5837
rect 12681 5805 12699 5825
rect 12719 5805 12730 5825
rect 12681 5795 12730 5805
rect 16520 5838 16569 5850
rect 1259 5564 1308 5574
rect 1259 5544 1270 5564
rect 1290 5544 1308 5564
rect 1259 5532 1308 5544
rect 1358 5568 1402 5574
rect 1358 5548 1373 5568
rect 1393 5548 1402 5568
rect 1358 5532 1402 5548
rect 1477 5564 1526 5574
rect 1477 5544 1488 5564
rect 1508 5544 1526 5564
rect 1477 5532 1526 5544
rect 1576 5568 1620 5574
rect 1576 5548 1591 5568
rect 1611 5548 1620 5568
rect 1576 5532 1620 5548
rect 1690 5568 1734 5574
rect 1690 5548 1699 5568
rect 1719 5548 1734 5568
rect 1690 5532 1734 5548
rect 1784 5564 1833 5574
rect 1784 5544 1802 5564
rect 1822 5544 1833 5564
rect 1784 5532 1833 5544
rect 2618 5572 2667 5584
rect 2618 5552 2629 5572
rect 2649 5552 2667 5572
rect 2618 5542 2667 5552
rect 2717 5568 2761 5584
rect 2717 5548 2732 5568
rect 2752 5548 2761 5568
rect 2717 5542 2761 5548
rect 2831 5568 2875 5584
rect 2831 5548 2840 5568
rect 2860 5548 2875 5568
rect 2831 5542 2875 5548
rect 2925 5572 2974 5584
rect 2925 5552 2943 5572
rect 2963 5552 2974 5572
rect 2925 5542 2974 5552
rect 3049 5568 3093 5584
rect 3049 5548 3058 5568
rect 3078 5548 3093 5568
rect 3049 5542 3093 5548
rect 3143 5572 3192 5584
rect 16520 5818 16531 5838
rect 16551 5818 16569 5838
rect 16520 5808 16569 5818
rect 16619 5834 16663 5850
rect 16619 5814 16634 5834
rect 16654 5814 16663 5834
rect 16619 5808 16663 5814
rect 16733 5834 16777 5850
rect 16733 5814 16742 5834
rect 16762 5814 16777 5834
rect 16733 5808 16777 5814
rect 16827 5838 16876 5850
rect 16827 5818 16845 5838
rect 16865 5818 16876 5838
rect 16827 5808 16876 5818
rect 16951 5834 16995 5850
rect 16951 5814 16960 5834
rect 16980 5814 16995 5834
rect 16951 5808 16995 5814
rect 17045 5838 17094 5850
rect 17045 5818 17063 5838
rect 17083 5818 17094 5838
rect 17045 5808 17094 5818
rect 3143 5552 3161 5572
rect 3181 5552 3192 5572
rect 3143 5542 3192 5552
rect 5623 5577 5672 5587
rect 5623 5557 5634 5577
rect 5654 5557 5672 5577
rect 5623 5545 5672 5557
rect 5722 5581 5766 5587
rect 5722 5561 5737 5581
rect 5757 5561 5766 5581
rect 5722 5545 5766 5561
rect 5841 5577 5890 5587
rect 5841 5557 5852 5577
rect 5872 5557 5890 5577
rect 5841 5545 5890 5557
rect 5940 5581 5984 5587
rect 5940 5561 5955 5581
rect 5975 5561 5984 5581
rect 5940 5545 5984 5561
rect 6054 5581 6098 5587
rect 6054 5561 6063 5581
rect 6083 5561 6098 5581
rect 6054 5545 6098 5561
rect 6148 5577 6197 5587
rect 6148 5557 6166 5577
rect 6186 5557 6197 5577
rect 6148 5545 6197 5557
rect 6982 5585 7031 5597
rect 6982 5565 6993 5585
rect 7013 5565 7031 5585
rect 6982 5555 7031 5565
rect 7081 5581 7125 5597
rect 7081 5561 7096 5581
rect 7116 5561 7125 5581
rect 7081 5555 7125 5561
rect 7195 5581 7239 5597
rect 7195 5561 7204 5581
rect 7224 5561 7239 5581
rect 7195 5555 7239 5561
rect 7289 5585 7338 5597
rect 7289 5565 7307 5585
rect 7327 5565 7338 5585
rect 7289 5555 7338 5565
rect 7413 5581 7457 5597
rect 7413 5561 7422 5581
rect 7442 5561 7457 5581
rect 7413 5555 7457 5561
rect 7507 5585 7556 5597
rect 7507 5565 7525 5585
rect 7545 5565 7556 5585
rect 7507 5555 7556 5565
rect 20786 5812 20835 5824
rect 20786 5792 20797 5812
rect 20817 5792 20835 5812
rect 20786 5782 20835 5792
rect 20885 5808 20929 5824
rect 20885 5788 20900 5808
rect 20920 5788 20929 5808
rect 20885 5782 20929 5788
rect 20999 5808 21043 5824
rect 20999 5788 21008 5808
rect 21028 5788 21043 5808
rect 20999 5782 21043 5788
rect 21093 5812 21142 5824
rect 21093 5792 21111 5812
rect 21131 5792 21142 5812
rect 21093 5782 21142 5792
rect 21217 5808 21261 5824
rect 21217 5788 21226 5808
rect 21246 5788 21261 5808
rect 21217 5782 21261 5788
rect 21311 5812 21360 5824
rect 21311 5792 21329 5812
rect 21349 5792 21360 5812
rect 21311 5782 21360 5792
rect 25150 5825 25199 5837
rect 10000 5589 10049 5599
rect 10000 5569 10011 5589
rect 10031 5569 10049 5589
rect 10000 5557 10049 5569
rect 10099 5593 10143 5599
rect 10099 5573 10114 5593
rect 10134 5573 10143 5593
rect 10099 5557 10143 5573
rect 10218 5589 10267 5599
rect 10218 5569 10229 5589
rect 10249 5569 10267 5589
rect 10218 5557 10267 5569
rect 10317 5593 10361 5599
rect 10317 5573 10332 5593
rect 10352 5573 10361 5593
rect 10317 5557 10361 5573
rect 10431 5593 10475 5599
rect 10431 5573 10440 5593
rect 10460 5573 10475 5593
rect 10431 5557 10475 5573
rect 10525 5589 10574 5599
rect 10525 5569 10543 5589
rect 10563 5569 10574 5589
rect 10525 5557 10574 5569
rect 11359 5597 11408 5609
rect 11359 5577 11370 5597
rect 11390 5577 11408 5597
rect 11359 5567 11408 5577
rect 11458 5593 11502 5609
rect 11458 5573 11473 5593
rect 11493 5573 11502 5593
rect 11458 5567 11502 5573
rect 11572 5593 11616 5609
rect 11572 5573 11581 5593
rect 11601 5573 11616 5593
rect 11572 5567 11616 5573
rect 11666 5597 11715 5609
rect 11666 5577 11684 5597
rect 11704 5577 11715 5597
rect 11666 5567 11715 5577
rect 11790 5593 11834 5609
rect 11790 5573 11799 5593
rect 11819 5573 11834 5593
rect 11790 5567 11834 5573
rect 11884 5597 11933 5609
rect 25150 5805 25161 5825
rect 25181 5805 25199 5825
rect 25150 5795 25199 5805
rect 25249 5821 25293 5837
rect 25249 5801 25264 5821
rect 25284 5801 25293 5821
rect 25249 5795 25293 5801
rect 25363 5821 25407 5837
rect 25363 5801 25372 5821
rect 25392 5801 25407 5821
rect 25363 5795 25407 5801
rect 25457 5825 25506 5837
rect 25457 5805 25475 5825
rect 25495 5805 25506 5825
rect 25457 5795 25506 5805
rect 25581 5821 25625 5837
rect 25581 5801 25590 5821
rect 25610 5801 25625 5821
rect 25581 5795 25625 5801
rect 25675 5825 25724 5837
rect 25675 5805 25693 5825
rect 25713 5805 25724 5825
rect 25675 5795 25724 5805
rect 29527 5837 29576 5849
rect 11884 5577 11902 5597
rect 11922 5577 11933 5597
rect 11884 5567 11933 5577
rect 14364 5602 14413 5612
rect 14364 5582 14375 5602
rect 14395 5582 14413 5602
rect 3416 5388 3465 5400
rect 3416 5368 3427 5388
rect 3447 5368 3465 5388
rect 362 5338 411 5348
rect 362 5318 373 5338
rect 393 5318 411 5338
rect 362 5306 411 5318
rect 461 5342 505 5348
rect 461 5322 476 5342
rect 496 5322 505 5342
rect 461 5306 505 5322
rect 580 5338 629 5348
rect 580 5318 591 5338
rect 611 5318 629 5338
rect 580 5306 629 5318
rect 679 5342 723 5348
rect 679 5322 694 5342
rect 714 5322 723 5342
rect 679 5306 723 5322
rect 793 5342 837 5348
rect 793 5322 802 5342
rect 822 5322 837 5342
rect 793 5306 837 5322
rect 887 5338 936 5348
rect 3416 5358 3465 5368
rect 3515 5384 3559 5400
rect 3515 5364 3530 5384
rect 3550 5364 3559 5384
rect 3515 5358 3559 5364
rect 3629 5384 3673 5400
rect 3629 5364 3638 5384
rect 3658 5364 3673 5384
rect 3629 5358 3673 5364
rect 3723 5388 3772 5400
rect 3723 5368 3741 5388
rect 3761 5368 3772 5388
rect 3723 5358 3772 5368
rect 3847 5384 3891 5400
rect 3847 5364 3856 5384
rect 3876 5364 3891 5384
rect 3847 5358 3891 5364
rect 3941 5388 3990 5400
rect 3941 5368 3959 5388
rect 3979 5368 3990 5388
rect 3941 5358 3990 5368
rect 887 5318 905 5338
rect 925 5318 936 5338
rect 887 5306 936 5318
rect 14364 5570 14413 5582
rect 14463 5606 14507 5612
rect 14463 5586 14478 5606
rect 14498 5586 14507 5606
rect 14463 5570 14507 5586
rect 14582 5602 14631 5612
rect 14582 5582 14593 5602
rect 14613 5582 14631 5602
rect 14582 5570 14631 5582
rect 14681 5606 14725 5612
rect 14681 5586 14696 5606
rect 14716 5586 14725 5606
rect 14681 5570 14725 5586
rect 14795 5606 14839 5612
rect 14795 5586 14804 5606
rect 14824 5586 14839 5606
rect 14795 5570 14839 5586
rect 14889 5602 14938 5612
rect 14889 5582 14907 5602
rect 14927 5582 14938 5602
rect 14889 5570 14938 5582
rect 15723 5610 15772 5622
rect 15723 5590 15734 5610
rect 15754 5590 15772 5610
rect 15723 5580 15772 5590
rect 15822 5606 15866 5622
rect 15822 5586 15837 5606
rect 15857 5586 15866 5606
rect 15822 5580 15866 5586
rect 15936 5606 15980 5622
rect 15936 5586 15945 5606
rect 15965 5586 15980 5606
rect 15936 5580 15980 5586
rect 16030 5610 16079 5622
rect 16030 5590 16048 5610
rect 16068 5590 16079 5610
rect 16030 5580 16079 5590
rect 16154 5606 16198 5622
rect 16154 5586 16163 5606
rect 16183 5586 16198 5606
rect 16154 5580 16198 5586
rect 16248 5610 16297 5622
rect 16248 5590 16266 5610
rect 16286 5590 16297 5610
rect 16248 5580 16297 5590
rect 29527 5817 29538 5837
rect 29558 5817 29576 5837
rect 29527 5807 29576 5817
rect 29626 5833 29670 5849
rect 29626 5813 29641 5833
rect 29661 5813 29670 5833
rect 29626 5807 29670 5813
rect 29740 5833 29784 5849
rect 29740 5813 29749 5833
rect 29769 5813 29784 5833
rect 29740 5807 29784 5813
rect 29834 5837 29883 5849
rect 29834 5817 29852 5837
rect 29872 5817 29883 5837
rect 29834 5807 29883 5817
rect 29958 5833 30002 5849
rect 29958 5813 29967 5833
rect 29987 5813 30002 5833
rect 29958 5807 30002 5813
rect 30052 5837 30101 5849
rect 30052 5817 30070 5837
rect 30090 5817 30101 5837
rect 30052 5807 30101 5817
rect 33891 5850 33940 5862
rect 7780 5401 7829 5413
rect 7780 5381 7791 5401
rect 7811 5381 7829 5401
rect 4726 5351 4775 5361
rect 4726 5331 4737 5351
rect 4757 5331 4775 5351
rect 4726 5319 4775 5331
rect 4825 5355 4869 5361
rect 4825 5335 4840 5355
rect 4860 5335 4869 5355
rect 4825 5319 4869 5335
rect 4944 5351 4993 5361
rect 4944 5331 4955 5351
rect 4975 5331 4993 5351
rect 4944 5319 4993 5331
rect 5043 5355 5087 5361
rect 5043 5335 5058 5355
rect 5078 5335 5087 5355
rect 5043 5319 5087 5335
rect 5157 5355 5201 5361
rect 5157 5335 5166 5355
rect 5186 5335 5201 5355
rect 5157 5319 5201 5335
rect 5251 5351 5300 5361
rect 7780 5371 7829 5381
rect 7879 5397 7923 5413
rect 7879 5377 7894 5397
rect 7914 5377 7923 5397
rect 7879 5371 7923 5377
rect 7993 5397 8037 5413
rect 7993 5377 8002 5397
rect 8022 5377 8037 5397
rect 7993 5371 8037 5377
rect 8087 5401 8136 5413
rect 8087 5381 8105 5401
rect 8125 5381 8136 5401
rect 8087 5371 8136 5381
rect 8211 5397 8255 5413
rect 8211 5377 8220 5397
rect 8240 5377 8255 5397
rect 8211 5371 8255 5377
rect 8305 5401 8354 5413
rect 8305 5381 8323 5401
rect 8343 5381 8354 5401
rect 8305 5371 8354 5381
rect 5251 5331 5269 5351
rect 5289 5331 5300 5351
rect 5251 5319 5300 5331
rect 18630 5576 18679 5586
rect 18630 5556 18641 5576
rect 18661 5556 18679 5576
rect 18630 5544 18679 5556
rect 18729 5580 18773 5586
rect 18729 5560 18744 5580
rect 18764 5560 18773 5580
rect 18729 5544 18773 5560
rect 18848 5576 18897 5586
rect 18848 5556 18859 5576
rect 18879 5556 18897 5576
rect 18848 5544 18897 5556
rect 18947 5580 18991 5586
rect 18947 5560 18962 5580
rect 18982 5560 18991 5580
rect 18947 5544 18991 5560
rect 19061 5580 19105 5586
rect 19061 5560 19070 5580
rect 19090 5560 19105 5580
rect 19061 5544 19105 5560
rect 19155 5576 19204 5586
rect 19155 5556 19173 5576
rect 19193 5556 19204 5576
rect 19155 5544 19204 5556
rect 19989 5584 20038 5596
rect 19989 5564 20000 5584
rect 20020 5564 20038 5584
rect 19989 5554 20038 5564
rect 20088 5580 20132 5596
rect 20088 5560 20103 5580
rect 20123 5560 20132 5580
rect 20088 5554 20132 5560
rect 20202 5580 20246 5596
rect 20202 5560 20211 5580
rect 20231 5560 20246 5580
rect 20202 5554 20246 5560
rect 20296 5584 20345 5596
rect 20296 5564 20314 5584
rect 20334 5564 20345 5584
rect 20296 5554 20345 5564
rect 20420 5580 20464 5596
rect 20420 5560 20429 5580
rect 20449 5560 20464 5580
rect 20420 5554 20464 5560
rect 20514 5584 20563 5596
rect 33891 5830 33902 5850
rect 33922 5830 33940 5850
rect 33891 5820 33940 5830
rect 33990 5846 34034 5862
rect 33990 5826 34005 5846
rect 34025 5826 34034 5846
rect 33990 5820 34034 5826
rect 34104 5846 34148 5862
rect 34104 5826 34113 5846
rect 34133 5826 34148 5846
rect 34104 5820 34148 5826
rect 34198 5850 34247 5862
rect 34198 5830 34216 5850
rect 34236 5830 34247 5850
rect 34198 5820 34247 5830
rect 34322 5846 34366 5862
rect 34322 5826 34331 5846
rect 34351 5826 34366 5846
rect 34322 5820 34366 5826
rect 34416 5850 34465 5862
rect 34416 5830 34434 5850
rect 34454 5830 34465 5850
rect 34416 5820 34465 5830
rect 20514 5564 20532 5584
rect 20552 5564 20563 5584
rect 20514 5554 20563 5564
rect 22994 5589 23043 5599
rect 22994 5569 23005 5589
rect 23025 5569 23043 5589
rect 12157 5413 12206 5425
rect 12157 5393 12168 5413
rect 12188 5393 12206 5413
rect 9103 5363 9152 5373
rect 9103 5343 9114 5363
rect 9134 5343 9152 5363
rect 9103 5331 9152 5343
rect 9202 5367 9246 5373
rect 9202 5347 9217 5367
rect 9237 5347 9246 5367
rect 9202 5331 9246 5347
rect 9321 5363 9370 5373
rect 9321 5343 9332 5363
rect 9352 5343 9370 5363
rect 9321 5331 9370 5343
rect 9420 5367 9464 5373
rect 9420 5347 9435 5367
rect 9455 5347 9464 5367
rect 9420 5331 9464 5347
rect 9534 5367 9578 5373
rect 9534 5347 9543 5367
rect 9563 5347 9578 5367
rect 9534 5331 9578 5347
rect 9628 5363 9677 5373
rect 12157 5383 12206 5393
rect 12256 5409 12300 5425
rect 12256 5389 12271 5409
rect 12291 5389 12300 5409
rect 12256 5383 12300 5389
rect 12370 5409 12414 5425
rect 12370 5389 12379 5409
rect 12399 5389 12414 5409
rect 12370 5383 12414 5389
rect 12464 5413 12513 5425
rect 12464 5393 12482 5413
rect 12502 5393 12513 5413
rect 12464 5383 12513 5393
rect 12588 5409 12632 5425
rect 12588 5389 12597 5409
rect 12617 5389 12632 5409
rect 12588 5383 12632 5389
rect 12682 5413 12731 5425
rect 12682 5393 12700 5413
rect 12720 5393 12731 5413
rect 12682 5383 12731 5393
rect 9628 5343 9646 5363
rect 9666 5343 9677 5363
rect 9628 5331 9677 5343
rect 2314 5166 2363 5178
rect 1160 5154 1209 5164
rect 1160 5134 1171 5154
rect 1191 5134 1209 5154
rect 1160 5122 1209 5134
rect 1259 5158 1303 5164
rect 1259 5138 1274 5158
rect 1294 5138 1303 5158
rect 1259 5122 1303 5138
rect 1378 5154 1427 5164
rect 1378 5134 1389 5154
rect 1409 5134 1427 5154
rect 1378 5122 1427 5134
rect 1477 5158 1521 5164
rect 1477 5138 1492 5158
rect 1512 5138 1521 5158
rect 1477 5122 1521 5138
rect 1591 5158 1635 5164
rect 1591 5138 1600 5158
rect 1620 5138 1635 5158
rect 1591 5122 1635 5138
rect 1685 5154 1734 5164
rect 1685 5134 1703 5154
rect 1723 5134 1734 5154
rect 2314 5146 2325 5166
rect 2345 5146 2363 5166
rect 2314 5136 2363 5146
rect 2413 5162 2457 5178
rect 2413 5142 2428 5162
rect 2448 5142 2457 5162
rect 2413 5136 2457 5142
rect 2527 5162 2571 5178
rect 2527 5142 2536 5162
rect 2556 5142 2571 5162
rect 2527 5136 2571 5142
rect 2621 5166 2670 5178
rect 2621 5146 2639 5166
rect 2659 5146 2670 5166
rect 2621 5136 2670 5146
rect 2745 5162 2789 5178
rect 2745 5142 2754 5162
rect 2774 5142 2789 5162
rect 2745 5136 2789 5142
rect 2839 5166 2888 5178
rect 16521 5426 16570 5438
rect 16521 5406 16532 5426
rect 16552 5406 16570 5426
rect 13467 5376 13516 5386
rect 13467 5356 13478 5376
rect 13498 5356 13516 5376
rect 13467 5344 13516 5356
rect 13566 5380 13610 5386
rect 13566 5360 13581 5380
rect 13601 5360 13610 5380
rect 13566 5344 13610 5360
rect 13685 5376 13734 5386
rect 13685 5356 13696 5376
rect 13716 5356 13734 5376
rect 13685 5344 13734 5356
rect 13784 5380 13828 5386
rect 13784 5360 13799 5380
rect 13819 5360 13828 5380
rect 13784 5344 13828 5360
rect 13898 5380 13942 5386
rect 13898 5360 13907 5380
rect 13927 5360 13942 5380
rect 13898 5344 13942 5360
rect 13992 5376 14041 5386
rect 16521 5396 16570 5406
rect 16620 5422 16664 5438
rect 16620 5402 16635 5422
rect 16655 5402 16664 5422
rect 16620 5396 16664 5402
rect 16734 5422 16778 5438
rect 16734 5402 16743 5422
rect 16763 5402 16778 5422
rect 16734 5396 16778 5402
rect 16828 5426 16877 5438
rect 16828 5406 16846 5426
rect 16866 5406 16877 5426
rect 16828 5396 16877 5406
rect 16952 5422 16996 5438
rect 16952 5402 16961 5422
rect 16981 5402 16996 5422
rect 16952 5396 16996 5402
rect 17046 5426 17095 5438
rect 17046 5406 17064 5426
rect 17084 5406 17095 5426
rect 17046 5396 17095 5406
rect 22994 5557 23043 5569
rect 23093 5593 23137 5599
rect 23093 5573 23108 5593
rect 23128 5573 23137 5593
rect 23093 5557 23137 5573
rect 23212 5589 23261 5599
rect 23212 5569 23223 5589
rect 23243 5569 23261 5589
rect 23212 5557 23261 5569
rect 23311 5593 23355 5599
rect 23311 5573 23326 5593
rect 23346 5573 23355 5593
rect 23311 5557 23355 5573
rect 23425 5593 23469 5599
rect 23425 5573 23434 5593
rect 23454 5573 23469 5593
rect 23425 5557 23469 5573
rect 23519 5589 23568 5599
rect 23519 5569 23537 5589
rect 23557 5569 23568 5589
rect 23519 5557 23568 5569
rect 24353 5597 24402 5609
rect 24353 5577 24364 5597
rect 24384 5577 24402 5597
rect 24353 5567 24402 5577
rect 24452 5593 24496 5609
rect 24452 5573 24467 5593
rect 24487 5573 24496 5593
rect 24452 5567 24496 5573
rect 24566 5593 24610 5609
rect 24566 5573 24575 5593
rect 24595 5573 24610 5593
rect 24566 5567 24610 5573
rect 24660 5597 24709 5609
rect 24660 5577 24678 5597
rect 24698 5577 24709 5597
rect 24660 5567 24709 5577
rect 24784 5593 24828 5609
rect 24784 5573 24793 5593
rect 24813 5573 24828 5593
rect 24784 5567 24828 5573
rect 24878 5597 24927 5609
rect 24878 5577 24896 5597
rect 24916 5577 24927 5597
rect 24878 5567 24927 5577
rect 27371 5601 27420 5611
rect 27371 5581 27382 5601
rect 27402 5581 27420 5601
rect 13992 5356 14010 5376
rect 14030 5356 14041 5376
rect 13992 5344 14041 5356
rect 6678 5179 6727 5191
rect 2839 5146 2857 5166
rect 2877 5146 2888 5166
rect 2839 5136 2888 5146
rect 1685 5122 1734 5134
rect 5524 5167 5573 5177
rect 5524 5147 5535 5167
rect 5555 5147 5573 5167
rect 5524 5135 5573 5147
rect 5623 5171 5667 5177
rect 5623 5151 5638 5171
rect 5658 5151 5667 5171
rect 5623 5135 5667 5151
rect 5742 5167 5791 5177
rect 5742 5147 5753 5167
rect 5773 5147 5791 5167
rect 5742 5135 5791 5147
rect 5841 5171 5885 5177
rect 5841 5151 5856 5171
rect 5876 5151 5885 5171
rect 5841 5135 5885 5151
rect 5955 5171 5999 5177
rect 5955 5151 5964 5171
rect 5984 5151 5999 5171
rect 5955 5135 5999 5151
rect 6049 5167 6098 5177
rect 6049 5147 6067 5167
rect 6087 5147 6098 5167
rect 6678 5159 6689 5179
rect 6709 5159 6727 5179
rect 6678 5149 6727 5159
rect 6777 5175 6821 5191
rect 6777 5155 6792 5175
rect 6812 5155 6821 5175
rect 6777 5149 6821 5155
rect 6891 5175 6935 5191
rect 6891 5155 6900 5175
rect 6920 5155 6935 5175
rect 6891 5149 6935 5155
rect 6985 5179 7034 5191
rect 6985 5159 7003 5179
rect 7023 5159 7034 5179
rect 6985 5149 7034 5159
rect 7109 5175 7153 5191
rect 7109 5155 7118 5175
rect 7138 5155 7153 5175
rect 7109 5149 7153 5155
rect 7203 5179 7252 5191
rect 27371 5569 27420 5581
rect 27470 5605 27514 5611
rect 27470 5585 27485 5605
rect 27505 5585 27514 5605
rect 27470 5569 27514 5585
rect 27589 5601 27638 5611
rect 27589 5581 27600 5601
rect 27620 5581 27638 5601
rect 27589 5569 27638 5581
rect 27688 5605 27732 5611
rect 27688 5585 27703 5605
rect 27723 5585 27732 5605
rect 27688 5569 27732 5585
rect 27802 5605 27846 5611
rect 27802 5585 27811 5605
rect 27831 5585 27846 5605
rect 27802 5569 27846 5585
rect 27896 5601 27945 5611
rect 27896 5581 27914 5601
rect 27934 5581 27945 5601
rect 27896 5569 27945 5581
rect 28730 5609 28779 5621
rect 28730 5589 28741 5609
rect 28761 5589 28779 5609
rect 28730 5579 28779 5589
rect 28829 5605 28873 5621
rect 28829 5585 28844 5605
rect 28864 5585 28873 5605
rect 28829 5579 28873 5585
rect 28943 5605 28987 5621
rect 28943 5585 28952 5605
rect 28972 5585 28987 5605
rect 28943 5579 28987 5585
rect 29037 5609 29086 5621
rect 29037 5589 29055 5609
rect 29075 5589 29086 5609
rect 29037 5579 29086 5589
rect 29161 5605 29205 5621
rect 29161 5585 29170 5605
rect 29190 5585 29205 5605
rect 29161 5579 29205 5585
rect 29255 5609 29304 5621
rect 29255 5589 29273 5609
rect 29293 5589 29304 5609
rect 29255 5579 29304 5589
rect 31735 5614 31784 5624
rect 31735 5594 31746 5614
rect 31766 5594 31784 5614
rect 20787 5400 20836 5412
rect 20787 5380 20798 5400
rect 20818 5380 20836 5400
rect 11055 5191 11104 5203
rect 7203 5159 7221 5179
rect 7241 5159 7252 5179
rect 7203 5149 7252 5159
rect 6049 5135 6098 5147
rect 9901 5179 9950 5189
rect 9901 5159 9912 5179
rect 9932 5159 9950 5179
rect 9901 5147 9950 5159
rect 10000 5183 10044 5189
rect 10000 5163 10015 5183
rect 10035 5163 10044 5183
rect 10000 5147 10044 5163
rect 10119 5179 10168 5189
rect 10119 5159 10130 5179
rect 10150 5159 10168 5179
rect 10119 5147 10168 5159
rect 10218 5183 10262 5189
rect 10218 5163 10233 5183
rect 10253 5163 10262 5183
rect 10218 5147 10262 5163
rect 10332 5183 10376 5189
rect 10332 5163 10341 5183
rect 10361 5163 10376 5183
rect 10332 5147 10376 5163
rect 10426 5179 10475 5189
rect 10426 5159 10444 5179
rect 10464 5159 10475 5179
rect 11055 5171 11066 5191
rect 11086 5171 11104 5191
rect 11055 5161 11104 5171
rect 11154 5187 11198 5203
rect 11154 5167 11169 5187
rect 11189 5167 11198 5187
rect 11154 5161 11198 5167
rect 11268 5187 11312 5203
rect 11268 5167 11277 5187
rect 11297 5167 11312 5187
rect 11268 5161 11312 5167
rect 11362 5191 11411 5203
rect 11362 5171 11380 5191
rect 11400 5171 11411 5191
rect 11362 5161 11411 5171
rect 11486 5187 11530 5203
rect 11486 5167 11495 5187
rect 11515 5167 11530 5187
rect 11486 5161 11530 5167
rect 11580 5191 11629 5203
rect 17733 5350 17782 5360
rect 17733 5330 17744 5350
rect 17764 5330 17782 5350
rect 17733 5318 17782 5330
rect 17832 5354 17876 5360
rect 17832 5334 17847 5354
rect 17867 5334 17876 5354
rect 17832 5318 17876 5334
rect 17951 5350 18000 5360
rect 17951 5330 17962 5350
rect 17982 5330 18000 5350
rect 17951 5318 18000 5330
rect 18050 5354 18094 5360
rect 18050 5334 18065 5354
rect 18085 5334 18094 5354
rect 18050 5318 18094 5334
rect 18164 5354 18208 5360
rect 18164 5334 18173 5354
rect 18193 5334 18208 5354
rect 18164 5318 18208 5334
rect 18258 5350 18307 5360
rect 20787 5370 20836 5380
rect 20886 5396 20930 5412
rect 20886 5376 20901 5396
rect 20921 5376 20930 5396
rect 20886 5370 20930 5376
rect 21000 5396 21044 5412
rect 21000 5376 21009 5396
rect 21029 5376 21044 5396
rect 21000 5370 21044 5376
rect 21094 5400 21143 5412
rect 21094 5380 21112 5400
rect 21132 5380 21143 5400
rect 21094 5370 21143 5380
rect 21218 5396 21262 5412
rect 21218 5376 21227 5396
rect 21247 5376 21262 5396
rect 21218 5370 21262 5376
rect 21312 5400 21361 5412
rect 21312 5380 21330 5400
rect 21350 5380 21361 5400
rect 21312 5370 21361 5380
rect 18258 5330 18276 5350
rect 18296 5330 18307 5350
rect 18258 5318 18307 5330
rect 31735 5582 31784 5594
rect 31834 5618 31878 5624
rect 31834 5598 31849 5618
rect 31869 5598 31878 5618
rect 31834 5582 31878 5598
rect 31953 5614 32002 5624
rect 31953 5594 31964 5614
rect 31984 5594 32002 5614
rect 31953 5582 32002 5594
rect 32052 5618 32096 5624
rect 32052 5598 32067 5618
rect 32087 5598 32096 5618
rect 32052 5582 32096 5598
rect 32166 5618 32210 5624
rect 32166 5598 32175 5618
rect 32195 5598 32210 5618
rect 32166 5582 32210 5598
rect 32260 5614 32309 5624
rect 32260 5594 32278 5614
rect 32298 5594 32309 5614
rect 32260 5582 32309 5594
rect 33094 5622 33143 5634
rect 33094 5602 33105 5622
rect 33125 5602 33143 5622
rect 33094 5592 33143 5602
rect 33193 5618 33237 5634
rect 33193 5598 33208 5618
rect 33228 5598 33237 5618
rect 33193 5592 33237 5598
rect 33307 5618 33351 5634
rect 33307 5598 33316 5618
rect 33336 5598 33351 5618
rect 33307 5592 33351 5598
rect 33401 5622 33450 5634
rect 33401 5602 33419 5622
rect 33439 5602 33450 5622
rect 33401 5592 33450 5602
rect 33525 5618 33569 5634
rect 33525 5598 33534 5618
rect 33554 5598 33569 5618
rect 33525 5592 33569 5598
rect 33619 5622 33668 5634
rect 33619 5602 33637 5622
rect 33657 5602 33668 5622
rect 33619 5592 33668 5602
rect 25151 5413 25200 5425
rect 25151 5393 25162 5413
rect 25182 5393 25200 5413
rect 22097 5363 22146 5373
rect 22097 5343 22108 5363
rect 22128 5343 22146 5363
rect 22097 5331 22146 5343
rect 22196 5367 22240 5373
rect 22196 5347 22211 5367
rect 22231 5347 22240 5367
rect 22196 5331 22240 5347
rect 22315 5363 22364 5373
rect 22315 5343 22326 5363
rect 22346 5343 22364 5363
rect 22315 5331 22364 5343
rect 22414 5367 22458 5373
rect 22414 5347 22429 5367
rect 22449 5347 22458 5367
rect 22414 5331 22458 5347
rect 22528 5367 22572 5373
rect 22528 5347 22537 5367
rect 22557 5347 22572 5367
rect 22528 5331 22572 5347
rect 22622 5363 22671 5373
rect 25151 5383 25200 5393
rect 25250 5409 25294 5425
rect 25250 5389 25265 5409
rect 25285 5389 25294 5409
rect 25250 5383 25294 5389
rect 25364 5409 25408 5425
rect 25364 5389 25373 5409
rect 25393 5389 25408 5409
rect 25364 5383 25408 5389
rect 25458 5413 25507 5425
rect 25458 5393 25476 5413
rect 25496 5393 25507 5413
rect 25458 5383 25507 5393
rect 25582 5409 25626 5425
rect 25582 5389 25591 5409
rect 25611 5389 25626 5409
rect 25582 5383 25626 5389
rect 25676 5413 25725 5425
rect 25676 5393 25694 5413
rect 25714 5393 25725 5413
rect 25676 5383 25725 5393
rect 22622 5343 22640 5363
rect 22660 5343 22671 5363
rect 22622 5331 22671 5343
rect 15419 5204 15468 5216
rect 11580 5171 11598 5191
rect 11618 5171 11629 5191
rect 11580 5161 11629 5171
rect 10426 5147 10475 5159
rect 363 4926 412 4936
rect 363 4906 374 4926
rect 394 4906 412 4926
rect 363 4894 412 4906
rect 462 4930 506 4936
rect 462 4910 477 4930
rect 497 4910 506 4930
rect 462 4894 506 4910
rect 581 4926 630 4936
rect 581 4906 592 4926
rect 612 4906 630 4926
rect 581 4894 630 4906
rect 680 4930 724 4936
rect 680 4910 695 4930
rect 715 4910 724 4930
rect 680 4894 724 4910
rect 794 4930 838 4936
rect 794 4910 803 4930
rect 823 4910 838 4930
rect 794 4894 838 4910
rect 888 4926 937 4936
rect 888 4906 906 4926
rect 926 4906 937 4926
rect 14265 5192 14314 5202
rect 14265 5172 14276 5192
rect 14296 5172 14314 5192
rect 14265 5160 14314 5172
rect 14364 5196 14408 5202
rect 14364 5176 14379 5196
rect 14399 5176 14408 5196
rect 14364 5160 14408 5176
rect 14483 5192 14532 5202
rect 14483 5172 14494 5192
rect 14514 5172 14532 5192
rect 14483 5160 14532 5172
rect 14582 5196 14626 5202
rect 14582 5176 14597 5196
rect 14617 5176 14626 5196
rect 14582 5160 14626 5176
rect 14696 5196 14740 5202
rect 14696 5176 14705 5196
rect 14725 5176 14740 5196
rect 14696 5160 14740 5176
rect 14790 5192 14839 5202
rect 14790 5172 14808 5192
rect 14828 5172 14839 5192
rect 15419 5184 15430 5204
rect 15450 5184 15468 5204
rect 15419 5174 15468 5184
rect 15518 5200 15562 5216
rect 15518 5180 15533 5200
rect 15553 5180 15562 5200
rect 15518 5174 15562 5180
rect 15632 5200 15676 5216
rect 15632 5180 15641 5200
rect 15661 5180 15676 5200
rect 15632 5174 15676 5180
rect 15726 5204 15775 5216
rect 15726 5184 15744 5204
rect 15764 5184 15775 5204
rect 15726 5174 15775 5184
rect 15850 5200 15894 5216
rect 15850 5180 15859 5200
rect 15879 5180 15894 5200
rect 15850 5174 15894 5180
rect 15944 5204 15993 5216
rect 15944 5184 15962 5204
rect 15982 5184 15993 5204
rect 15944 5174 15993 5184
rect 14790 5160 14839 5172
rect 888 4894 937 4906
rect 4727 4939 4776 4949
rect 4727 4919 4738 4939
rect 4758 4919 4776 4939
rect 4727 4907 4776 4919
rect 4826 4943 4870 4949
rect 4826 4923 4841 4943
rect 4861 4923 4870 4943
rect 4826 4907 4870 4923
rect 4945 4939 4994 4949
rect 4945 4919 4956 4939
rect 4976 4919 4994 4939
rect 4945 4907 4994 4919
rect 5044 4943 5088 4949
rect 5044 4923 5059 4943
rect 5079 4923 5088 4943
rect 5044 4907 5088 4923
rect 5158 4943 5202 4949
rect 5158 4923 5167 4943
rect 5187 4923 5202 4943
rect 5158 4907 5202 4923
rect 5252 4939 5301 4949
rect 5252 4919 5270 4939
rect 5290 4919 5301 4939
rect 29528 5425 29577 5437
rect 29528 5405 29539 5425
rect 29559 5405 29577 5425
rect 26474 5375 26523 5385
rect 26474 5355 26485 5375
rect 26505 5355 26523 5375
rect 26474 5343 26523 5355
rect 26573 5379 26617 5385
rect 26573 5359 26588 5379
rect 26608 5359 26617 5379
rect 26573 5343 26617 5359
rect 26692 5375 26741 5385
rect 26692 5355 26703 5375
rect 26723 5355 26741 5375
rect 26692 5343 26741 5355
rect 26791 5379 26835 5385
rect 26791 5359 26806 5379
rect 26826 5359 26835 5379
rect 26791 5343 26835 5359
rect 26905 5379 26949 5385
rect 26905 5359 26914 5379
rect 26934 5359 26949 5379
rect 26905 5343 26949 5359
rect 26999 5375 27048 5385
rect 29528 5395 29577 5405
rect 29627 5421 29671 5437
rect 29627 5401 29642 5421
rect 29662 5401 29671 5421
rect 29627 5395 29671 5401
rect 29741 5421 29785 5437
rect 29741 5401 29750 5421
rect 29770 5401 29785 5421
rect 29741 5395 29785 5401
rect 29835 5425 29884 5437
rect 29835 5405 29853 5425
rect 29873 5405 29884 5425
rect 29835 5395 29884 5405
rect 29959 5421 30003 5437
rect 29959 5401 29968 5421
rect 29988 5401 30003 5421
rect 29959 5395 30003 5401
rect 30053 5425 30102 5437
rect 30053 5405 30071 5425
rect 30091 5405 30102 5425
rect 30053 5395 30102 5405
rect 26999 5355 27017 5375
rect 27037 5355 27048 5375
rect 26999 5343 27048 5355
rect 19685 5178 19734 5190
rect 18531 5166 18580 5176
rect 18531 5146 18542 5166
rect 18562 5146 18580 5166
rect 18531 5134 18580 5146
rect 18630 5170 18674 5176
rect 18630 5150 18645 5170
rect 18665 5150 18674 5170
rect 18630 5134 18674 5150
rect 18749 5166 18798 5176
rect 18749 5146 18760 5166
rect 18780 5146 18798 5166
rect 18749 5134 18798 5146
rect 18848 5170 18892 5176
rect 18848 5150 18863 5170
rect 18883 5150 18892 5170
rect 18848 5134 18892 5150
rect 18962 5170 19006 5176
rect 18962 5150 18971 5170
rect 18991 5150 19006 5170
rect 18962 5134 19006 5150
rect 19056 5166 19105 5176
rect 19056 5146 19074 5166
rect 19094 5146 19105 5166
rect 19685 5158 19696 5178
rect 19716 5158 19734 5178
rect 19685 5148 19734 5158
rect 19784 5174 19828 5190
rect 19784 5154 19799 5174
rect 19819 5154 19828 5174
rect 19784 5148 19828 5154
rect 19898 5174 19942 5190
rect 19898 5154 19907 5174
rect 19927 5154 19942 5174
rect 19898 5148 19942 5154
rect 19992 5178 20041 5190
rect 19992 5158 20010 5178
rect 20030 5158 20041 5178
rect 19992 5148 20041 5158
rect 20116 5174 20160 5190
rect 20116 5154 20125 5174
rect 20145 5154 20160 5174
rect 20116 5148 20160 5154
rect 20210 5178 20259 5190
rect 33892 5438 33941 5450
rect 33892 5418 33903 5438
rect 33923 5418 33941 5438
rect 30838 5388 30887 5398
rect 30838 5368 30849 5388
rect 30869 5368 30887 5388
rect 30838 5356 30887 5368
rect 30937 5392 30981 5398
rect 30937 5372 30952 5392
rect 30972 5372 30981 5392
rect 30937 5356 30981 5372
rect 31056 5388 31105 5398
rect 31056 5368 31067 5388
rect 31087 5368 31105 5388
rect 31056 5356 31105 5368
rect 31155 5392 31199 5398
rect 31155 5372 31170 5392
rect 31190 5372 31199 5392
rect 31155 5356 31199 5372
rect 31269 5392 31313 5398
rect 31269 5372 31278 5392
rect 31298 5372 31313 5392
rect 31269 5356 31313 5372
rect 31363 5388 31412 5398
rect 33892 5408 33941 5418
rect 33991 5434 34035 5450
rect 33991 5414 34006 5434
rect 34026 5414 34035 5434
rect 33991 5408 34035 5414
rect 34105 5434 34149 5450
rect 34105 5414 34114 5434
rect 34134 5414 34149 5434
rect 34105 5408 34149 5414
rect 34199 5438 34248 5450
rect 34199 5418 34217 5438
rect 34237 5418 34248 5438
rect 34199 5408 34248 5418
rect 34323 5434 34367 5450
rect 34323 5414 34332 5434
rect 34352 5414 34367 5434
rect 34323 5408 34367 5414
rect 34417 5438 34466 5450
rect 34417 5418 34435 5438
rect 34455 5418 34466 5438
rect 34417 5408 34466 5418
rect 31363 5368 31381 5388
rect 31401 5368 31412 5388
rect 31363 5356 31412 5368
rect 24049 5191 24098 5203
rect 20210 5158 20228 5178
rect 20248 5158 20259 5178
rect 20210 5148 20259 5158
rect 19056 5134 19105 5146
rect 5252 4907 5301 4919
rect 9104 4951 9153 4961
rect 9104 4931 9115 4951
rect 9135 4931 9153 4951
rect 9104 4919 9153 4931
rect 9203 4955 9247 4961
rect 9203 4935 9218 4955
rect 9238 4935 9247 4955
rect 9203 4919 9247 4935
rect 9322 4951 9371 4961
rect 9322 4931 9333 4951
rect 9353 4931 9371 4951
rect 9322 4919 9371 4931
rect 9421 4955 9465 4961
rect 9421 4935 9436 4955
rect 9456 4935 9465 4955
rect 9421 4919 9465 4935
rect 9535 4955 9579 4961
rect 9535 4935 9544 4955
rect 9564 4935 9579 4955
rect 9535 4919 9579 4935
rect 9629 4951 9678 4961
rect 9629 4931 9647 4951
rect 9667 4931 9678 4951
rect 22895 5179 22944 5189
rect 22895 5159 22906 5179
rect 22926 5159 22944 5179
rect 22895 5147 22944 5159
rect 22994 5183 23038 5189
rect 22994 5163 23009 5183
rect 23029 5163 23038 5183
rect 22994 5147 23038 5163
rect 23113 5179 23162 5189
rect 23113 5159 23124 5179
rect 23144 5159 23162 5179
rect 23113 5147 23162 5159
rect 23212 5183 23256 5189
rect 23212 5163 23227 5183
rect 23247 5163 23256 5183
rect 23212 5147 23256 5163
rect 23326 5183 23370 5189
rect 23326 5163 23335 5183
rect 23355 5163 23370 5183
rect 23326 5147 23370 5163
rect 23420 5179 23469 5189
rect 23420 5159 23438 5179
rect 23458 5159 23469 5179
rect 24049 5171 24060 5191
rect 24080 5171 24098 5191
rect 24049 5161 24098 5171
rect 24148 5187 24192 5203
rect 24148 5167 24163 5187
rect 24183 5167 24192 5187
rect 24148 5161 24192 5167
rect 24262 5187 24306 5203
rect 24262 5167 24271 5187
rect 24291 5167 24306 5187
rect 24262 5161 24306 5167
rect 24356 5191 24405 5203
rect 24356 5171 24374 5191
rect 24394 5171 24405 5191
rect 24356 5161 24405 5171
rect 24480 5187 24524 5203
rect 24480 5167 24489 5187
rect 24509 5167 24524 5187
rect 24480 5161 24524 5167
rect 24574 5191 24623 5203
rect 28426 5203 28475 5215
rect 24574 5171 24592 5191
rect 24612 5171 24623 5191
rect 24574 5161 24623 5171
rect 23420 5147 23469 5159
rect 9629 4919 9678 4931
rect 13468 4964 13517 4974
rect 13468 4944 13479 4964
rect 13499 4944 13517 4964
rect 13468 4932 13517 4944
rect 13567 4968 13611 4974
rect 13567 4948 13582 4968
rect 13602 4948 13611 4968
rect 13567 4932 13611 4948
rect 13686 4964 13735 4974
rect 13686 4944 13697 4964
rect 13717 4944 13735 4964
rect 13686 4932 13735 4944
rect 13785 4968 13829 4974
rect 13785 4948 13800 4968
rect 13820 4948 13829 4968
rect 13785 4932 13829 4948
rect 13899 4968 13943 4974
rect 13899 4948 13908 4968
rect 13928 4948 13943 4968
rect 13899 4932 13943 4948
rect 13993 4964 14042 4974
rect 13993 4944 14011 4964
rect 14031 4944 14042 4964
rect 13993 4932 14042 4944
rect 27272 5191 27321 5201
rect 27272 5171 27283 5191
rect 27303 5171 27321 5191
rect 27272 5159 27321 5171
rect 27371 5195 27415 5201
rect 27371 5175 27386 5195
rect 27406 5175 27415 5195
rect 27371 5159 27415 5175
rect 27490 5191 27539 5201
rect 27490 5171 27501 5191
rect 27521 5171 27539 5191
rect 27490 5159 27539 5171
rect 27589 5195 27633 5201
rect 27589 5175 27604 5195
rect 27624 5175 27633 5195
rect 27589 5159 27633 5175
rect 27703 5195 27747 5201
rect 27703 5175 27712 5195
rect 27732 5175 27747 5195
rect 27703 5159 27747 5175
rect 27797 5191 27846 5201
rect 27797 5171 27815 5191
rect 27835 5171 27846 5191
rect 28426 5183 28437 5203
rect 28457 5183 28475 5203
rect 28426 5173 28475 5183
rect 28525 5199 28569 5215
rect 28525 5179 28540 5199
rect 28560 5179 28569 5199
rect 28525 5173 28569 5179
rect 28639 5199 28683 5215
rect 28639 5179 28648 5199
rect 28668 5179 28683 5199
rect 28639 5173 28683 5179
rect 28733 5203 28782 5215
rect 28733 5183 28751 5203
rect 28771 5183 28782 5203
rect 28733 5173 28782 5183
rect 28857 5199 28901 5215
rect 28857 5179 28866 5199
rect 28886 5179 28901 5199
rect 28857 5173 28901 5179
rect 28951 5203 29000 5215
rect 32790 5216 32839 5228
rect 28951 5183 28969 5203
rect 28989 5183 29000 5203
rect 28951 5173 29000 5183
rect 27797 5159 27846 5171
rect 17734 4938 17783 4948
rect 17734 4918 17745 4938
rect 17765 4918 17783 4938
rect 17734 4906 17783 4918
rect 17833 4942 17877 4948
rect 17833 4922 17848 4942
rect 17868 4922 17877 4942
rect 17833 4906 17877 4922
rect 17952 4938 18001 4948
rect 17952 4918 17963 4938
rect 17983 4918 18001 4938
rect 17952 4906 18001 4918
rect 18051 4942 18095 4948
rect 18051 4922 18066 4942
rect 18086 4922 18095 4942
rect 18051 4906 18095 4922
rect 18165 4942 18209 4948
rect 18165 4922 18174 4942
rect 18194 4922 18209 4942
rect 18165 4906 18209 4922
rect 18259 4938 18308 4948
rect 18259 4918 18277 4938
rect 18297 4918 18308 4938
rect 31636 5204 31685 5214
rect 31636 5184 31647 5204
rect 31667 5184 31685 5204
rect 31636 5172 31685 5184
rect 31735 5208 31779 5214
rect 31735 5188 31750 5208
rect 31770 5188 31779 5208
rect 31735 5172 31779 5188
rect 31854 5204 31903 5214
rect 31854 5184 31865 5204
rect 31885 5184 31903 5204
rect 31854 5172 31903 5184
rect 31953 5208 31997 5214
rect 31953 5188 31968 5208
rect 31988 5188 31997 5208
rect 31953 5172 31997 5188
rect 32067 5208 32111 5214
rect 32067 5188 32076 5208
rect 32096 5188 32111 5208
rect 32067 5172 32111 5188
rect 32161 5204 32210 5214
rect 32161 5184 32179 5204
rect 32199 5184 32210 5204
rect 32790 5196 32801 5216
rect 32821 5196 32839 5216
rect 32790 5186 32839 5196
rect 32889 5212 32933 5228
rect 32889 5192 32904 5212
rect 32924 5192 32933 5212
rect 32889 5186 32933 5192
rect 33003 5212 33047 5228
rect 33003 5192 33012 5212
rect 33032 5192 33047 5212
rect 33003 5186 33047 5192
rect 33097 5216 33146 5228
rect 33097 5196 33115 5216
rect 33135 5196 33146 5216
rect 33097 5186 33146 5196
rect 33221 5212 33265 5228
rect 33221 5192 33230 5212
rect 33250 5192 33265 5212
rect 33221 5186 33265 5192
rect 33315 5216 33364 5228
rect 33315 5196 33333 5216
rect 33353 5196 33364 5216
rect 33315 5186 33364 5196
rect 32161 5172 32210 5184
rect 18259 4906 18308 4918
rect 22098 4951 22147 4961
rect 22098 4931 22109 4951
rect 22129 4931 22147 4951
rect 22098 4919 22147 4931
rect 22197 4955 22241 4961
rect 22197 4935 22212 4955
rect 22232 4935 22241 4955
rect 22197 4919 22241 4935
rect 22316 4951 22365 4961
rect 22316 4931 22327 4951
rect 22347 4931 22365 4951
rect 22316 4919 22365 4931
rect 22415 4955 22459 4961
rect 22415 4935 22430 4955
rect 22450 4935 22459 4955
rect 22415 4919 22459 4935
rect 22529 4955 22573 4961
rect 22529 4935 22538 4955
rect 22558 4935 22573 4955
rect 22529 4919 22573 4935
rect 22623 4951 22672 4961
rect 22623 4931 22641 4951
rect 22661 4931 22672 4951
rect 22623 4919 22672 4931
rect 26475 4963 26524 4973
rect 26475 4943 26486 4963
rect 26506 4943 26524 4963
rect 26475 4931 26524 4943
rect 26574 4967 26618 4973
rect 26574 4947 26589 4967
rect 26609 4947 26618 4967
rect 26574 4931 26618 4947
rect 26693 4963 26742 4973
rect 26693 4943 26704 4963
rect 26724 4943 26742 4963
rect 26693 4931 26742 4943
rect 26792 4967 26836 4973
rect 26792 4947 26807 4967
rect 26827 4947 26836 4967
rect 26792 4931 26836 4947
rect 26906 4967 26950 4973
rect 26906 4947 26915 4967
rect 26935 4947 26950 4967
rect 26906 4931 26950 4947
rect 27000 4963 27049 4973
rect 27000 4943 27018 4963
rect 27038 4943 27049 4963
rect 27000 4931 27049 4943
rect 30839 4976 30888 4986
rect 30839 4956 30850 4976
rect 30870 4956 30888 4976
rect 30839 4944 30888 4956
rect 30938 4980 30982 4986
rect 30938 4960 30953 4980
rect 30973 4960 30982 4980
rect 30938 4944 30982 4960
rect 31057 4976 31106 4986
rect 31057 4956 31068 4976
rect 31088 4956 31106 4976
rect 31057 4944 31106 4956
rect 31156 4980 31200 4986
rect 31156 4960 31171 4980
rect 31191 4960 31200 4980
rect 31156 4944 31200 4960
rect 31270 4980 31314 4986
rect 31270 4960 31279 4980
rect 31299 4960 31314 4980
rect 31270 4944 31314 4960
rect 31364 4976 31413 4986
rect 31364 4956 31382 4976
rect 31402 4956 31413 4976
rect 31364 4944 31413 4956
rect 3396 4782 3445 4794
rect 3396 4762 3407 4782
rect 3427 4762 3445 4782
rect 3396 4752 3445 4762
rect 3495 4778 3539 4794
rect 3495 4758 3510 4778
rect 3530 4758 3539 4778
rect 3495 4752 3539 4758
rect 3609 4778 3653 4794
rect 3609 4758 3618 4778
rect 3638 4758 3653 4778
rect 3609 4752 3653 4758
rect 3703 4782 3752 4794
rect 3703 4762 3721 4782
rect 3741 4762 3752 4782
rect 3703 4752 3752 4762
rect 3827 4778 3871 4794
rect 3827 4758 3836 4778
rect 3856 4758 3871 4778
rect 3827 4752 3871 4758
rect 3921 4782 3970 4794
rect 3921 4762 3939 4782
rect 3959 4762 3970 4782
rect 3921 4752 3970 4762
rect 7760 4795 7809 4807
rect 7760 4775 7771 4795
rect 7791 4775 7809 4795
rect 7760 4765 7809 4775
rect 7859 4791 7903 4807
rect 7859 4771 7874 4791
rect 7894 4771 7903 4791
rect 7859 4765 7903 4771
rect 7973 4791 8017 4807
rect 7973 4771 7982 4791
rect 8002 4771 8017 4791
rect 7973 4765 8017 4771
rect 8067 4795 8116 4807
rect 8067 4775 8085 4795
rect 8105 4775 8116 4795
rect 8067 4765 8116 4775
rect 8191 4791 8235 4807
rect 8191 4771 8200 4791
rect 8220 4771 8235 4791
rect 8191 4765 8235 4771
rect 8285 4795 8334 4807
rect 8285 4775 8303 4795
rect 8323 4775 8334 4795
rect 8285 4765 8334 4775
rect 12137 4807 12186 4819
rect 12137 4787 12148 4807
rect 12168 4787 12186 4807
rect 12137 4777 12186 4787
rect 12236 4803 12280 4819
rect 12236 4783 12251 4803
rect 12271 4783 12280 4803
rect 12236 4777 12280 4783
rect 12350 4803 12394 4819
rect 12350 4783 12359 4803
rect 12379 4783 12394 4803
rect 12350 4777 12394 4783
rect 12444 4807 12493 4819
rect 12444 4787 12462 4807
rect 12482 4787 12493 4807
rect 12444 4777 12493 4787
rect 12568 4803 12612 4819
rect 12568 4783 12577 4803
rect 12597 4783 12612 4803
rect 12568 4777 12612 4783
rect 12662 4807 12711 4819
rect 12662 4787 12680 4807
rect 12700 4787 12711 4807
rect 12662 4777 12711 4787
rect 16501 4820 16550 4832
rect 2599 4554 2648 4566
rect 1445 4542 1494 4552
rect 1445 4522 1456 4542
rect 1476 4522 1494 4542
rect 1445 4510 1494 4522
rect 1544 4546 1588 4552
rect 1544 4526 1559 4546
rect 1579 4526 1588 4546
rect 1544 4510 1588 4526
rect 1663 4542 1712 4552
rect 1663 4522 1674 4542
rect 1694 4522 1712 4542
rect 1663 4510 1712 4522
rect 1762 4546 1806 4552
rect 1762 4526 1777 4546
rect 1797 4526 1806 4546
rect 1762 4510 1806 4526
rect 1876 4546 1920 4552
rect 1876 4526 1885 4546
rect 1905 4526 1920 4546
rect 1876 4510 1920 4526
rect 1970 4542 2019 4552
rect 1970 4522 1988 4542
rect 2008 4522 2019 4542
rect 2599 4534 2610 4554
rect 2630 4534 2648 4554
rect 2599 4524 2648 4534
rect 2698 4550 2742 4566
rect 2698 4530 2713 4550
rect 2733 4530 2742 4550
rect 2698 4524 2742 4530
rect 2812 4550 2856 4566
rect 2812 4530 2821 4550
rect 2841 4530 2856 4550
rect 2812 4524 2856 4530
rect 2906 4554 2955 4566
rect 2906 4534 2924 4554
rect 2944 4534 2955 4554
rect 2906 4524 2955 4534
rect 3030 4550 3074 4566
rect 3030 4530 3039 4550
rect 3059 4530 3074 4550
rect 3030 4524 3074 4530
rect 3124 4554 3173 4566
rect 3124 4534 3142 4554
rect 3162 4534 3173 4554
rect 3124 4524 3173 4534
rect 16501 4800 16512 4820
rect 16532 4800 16550 4820
rect 16501 4790 16550 4800
rect 16600 4816 16644 4832
rect 16600 4796 16615 4816
rect 16635 4796 16644 4816
rect 16600 4790 16644 4796
rect 16714 4816 16758 4832
rect 16714 4796 16723 4816
rect 16743 4796 16758 4816
rect 16714 4790 16758 4796
rect 16808 4820 16857 4832
rect 16808 4800 16826 4820
rect 16846 4800 16857 4820
rect 16808 4790 16857 4800
rect 16932 4816 16976 4832
rect 16932 4796 16941 4816
rect 16961 4796 16976 4816
rect 16932 4790 16976 4796
rect 17026 4820 17075 4832
rect 17026 4800 17044 4820
rect 17064 4800 17075 4820
rect 17026 4790 17075 4800
rect 6963 4567 7012 4579
rect 5809 4555 5858 4565
rect 5809 4535 5820 4555
rect 5840 4535 5858 4555
rect 1970 4510 2019 4522
rect 5809 4523 5858 4535
rect 5908 4559 5952 4565
rect 5908 4539 5923 4559
rect 5943 4539 5952 4559
rect 5908 4523 5952 4539
rect 6027 4555 6076 4565
rect 6027 4535 6038 4555
rect 6058 4535 6076 4555
rect 6027 4523 6076 4535
rect 6126 4559 6170 4565
rect 6126 4539 6141 4559
rect 6161 4539 6170 4559
rect 6126 4523 6170 4539
rect 6240 4559 6284 4565
rect 6240 4539 6249 4559
rect 6269 4539 6284 4559
rect 6240 4523 6284 4539
rect 6334 4555 6383 4565
rect 6334 4535 6352 4555
rect 6372 4535 6383 4555
rect 6963 4547 6974 4567
rect 6994 4547 7012 4567
rect 6963 4537 7012 4547
rect 7062 4563 7106 4579
rect 7062 4543 7077 4563
rect 7097 4543 7106 4563
rect 7062 4537 7106 4543
rect 7176 4563 7220 4579
rect 7176 4543 7185 4563
rect 7205 4543 7220 4563
rect 7176 4537 7220 4543
rect 7270 4567 7319 4579
rect 7270 4547 7288 4567
rect 7308 4547 7319 4567
rect 7270 4537 7319 4547
rect 7394 4563 7438 4579
rect 7394 4543 7403 4563
rect 7423 4543 7438 4563
rect 7394 4537 7438 4543
rect 7488 4567 7537 4579
rect 7488 4547 7506 4567
rect 7526 4547 7537 4567
rect 7488 4537 7537 4547
rect 20767 4794 20816 4806
rect 20767 4774 20778 4794
rect 20798 4774 20816 4794
rect 20767 4764 20816 4774
rect 20866 4790 20910 4806
rect 20866 4770 20881 4790
rect 20901 4770 20910 4790
rect 20866 4764 20910 4770
rect 20980 4790 21024 4806
rect 20980 4770 20989 4790
rect 21009 4770 21024 4790
rect 20980 4764 21024 4770
rect 21074 4794 21123 4806
rect 21074 4774 21092 4794
rect 21112 4774 21123 4794
rect 21074 4764 21123 4774
rect 21198 4790 21242 4806
rect 21198 4770 21207 4790
rect 21227 4770 21242 4790
rect 21198 4764 21242 4770
rect 21292 4794 21341 4806
rect 21292 4774 21310 4794
rect 21330 4774 21341 4794
rect 21292 4764 21341 4774
rect 25131 4807 25180 4819
rect 11340 4579 11389 4591
rect 10186 4567 10235 4577
rect 10186 4547 10197 4567
rect 10217 4547 10235 4567
rect 6334 4523 6383 4535
rect 10186 4535 10235 4547
rect 10285 4571 10329 4577
rect 10285 4551 10300 4571
rect 10320 4551 10329 4571
rect 10285 4535 10329 4551
rect 10404 4567 10453 4577
rect 10404 4547 10415 4567
rect 10435 4547 10453 4567
rect 10404 4535 10453 4547
rect 10503 4571 10547 4577
rect 10503 4551 10518 4571
rect 10538 4551 10547 4571
rect 10503 4535 10547 4551
rect 10617 4571 10661 4577
rect 10617 4551 10626 4571
rect 10646 4551 10661 4571
rect 10617 4535 10661 4551
rect 10711 4567 10760 4577
rect 10711 4547 10729 4567
rect 10749 4547 10760 4567
rect 11340 4559 11351 4579
rect 11371 4559 11389 4579
rect 11340 4549 11389 4559
rect 11439 4575 11483 4591
rect 11439 4555 11454 4575
rect 11474 4555 11483 4575
rect 11439 4549 11483 4555
rect 11553 4575 11597 4591
rect 11553 4555 11562 4575
rect 11582 4555 11597 4575
rect 11553 4549 11597 4555
rect 11647 4579 11696 4591
rect 11647 4559 11665 4579
rect 11685 4559 11696 4579
rect 11647 4549 11696 4559
rect 11771 4575 11815 4591
rect 11771 4555 11780 4575
rect 11800 4555 11815 4575
rect 11771 4549 11815 4555
rect 11865 4579 11914 4591
rect 11865 4559 11883 4579
rect 11903 4559 11914 4579
rect 11865 4549 11914 4559
rect 25131 4787 25142 4807
rect 25162 4787 25180 4807
rect 25131 4777 25180 4787
rect 25230 4803 25274 4819
rect 25230 4783 25245 4803
rect 25265 4783 25274 4803
rect 25230 4777 25274 4783
rect 25344 4803 25388 4819
rect 25344 4783 25353 4803
rect 25373 4783 25388 4803
rect 25344 4777 25388 4783
rect 25438 4807 25487 4819
rect 25438 4787 25456 4807
rect 25476 4787 25487 4807
rect 25438 4777 25487 4787
rect 25562 4803 25606 4819
rect 25562 4783 25571 4803
rect 25591 4783 25606 4803
rect 25562 4777 25606 4783
rect 25656 4807 25705 4819
rect 25656 4787 25674 4807
rect 25694 4787 25705 4807
rect 25656 4777 25705 4787
rect 29508 4819 29557 4831
rect 15704 4592 15753 4604
rect 14550 4580 14599 4590
rect 14550 4560 14561 4580
rect 14581 4560 14599 4580
rect 10711 4535 10760 4547
rect 3397 4370 3446 4382
rect 3397 4350 3408 4370
rect 3428 4350 3446 4370
rect 343 4320 392 4330
rect 343 4300 354 4320
rect 374 4300 392 4320
rect 343 4288 392 4300
rect 442 4324 486 4330
rect 442 4304 457 4324
rect 477 4304 486 4324
rect 442 4288 486 4304
rect 561 4320 610 4330
rect 561 4300 572 4320
rect 592 4300 610 4320
rect 561 4288 610 4300
rect 660 4324 704 4330
rect 660 4304 675 4324
rect 695 4304 704 4324
rect 660 4288 704 4304
rect 774 4324 818 4330
rect 774 4304 783 4324
rect 803 4304 818 4324
rect 774 4288 818 4304
rect 868 4320 917 4330
rect 3397 4340 3446 4350
rect 3496 4366 3540 4382
rect 3496 4346 3511 4366
rect 3531 4346 3540 4366
rect 3496 4340 3540 4346
rect 3610 4366 3654 4382
rect 3610 4346 3619 4366
rect 3639 4346 3654 4366
rect 3610 4340 3654 4346
rect 3704 4370 3753 4382
rect 3704 4350 3722 4370
rect 3742 4350 3753 4370
rect 3704 4340 3753 4350
rect 3828 4366 3872 4382
rect 3828 4346 3837 4366
rect 3857 4346 3872 4366
rect 3828 4340 3872 4346
rect 3922 4370 3971 4382
rect 3922 4350 3940 4370
rect 3960 4350 3971 4370
rect 3922 4340 3971 4350
rect 868 4300 886 4320
rect 906 4300 917 4320
rect 868 4288 917 4300
rect 14550 4548 14599 4560
rect 14649 4584 14693 4590
rect 14649 4564 14664 4584
rect 14684 4564 14693 4584
rect 14649 4548 14693 4564
rect 14768 4580 14817 4590
rect 14768 4560 14779 4580
rect 14799 4560 14817 4580
rect 14768 4548 14817 4560
rect 14867 4584 14911 4590
rect 14867 4564 14882 4584
rect 14902 4564 14911 4584
rect 14867 4548 14911 4564
rect 14981 4584 15025 4590
rect 14981 4564 14990 4584
rect 15010 4564 15025 4584
rect 14981 4548 15025 4564
rect 15075 4580 15124 4590
rect 15075 4560 15093 4580
rect 15113 4560 15124 4580
rect 15704 4572 15715 4592
rect 15735 4572 15753 4592
rect 15704 4562 15753 4572
rect 15803 4588 15847 4604
rect 15803 4568 15818 4588
rect 15838 4568 15847 4588
rect 15803 4562 15847 4568
rect 15917 4588 15961 4604
rect 15917 4568 15926 4588
rect 15946 4568 15961 4588
rect 15917 4562 15961 4568
rect 16011 4592 16060 4604
rect 16011 4572 16029 4592
rect 16049 4572 16060 4592
rect 16011 4562 16060 4572
rect 16135 4588 16179 4604
rect 16135 4568 16144 4588
rect 16164 4568 16179 4588
rect 16135 4562 16179 4568
rect 16229 4592 16278 4604
rect 16229 4572 16247 4592
rect 16267 4572 16278 4592
rect 16229 4562 16278 4572
rect 15075 4548 15124 4560
rect 7761 4383 7810 4395
rect 7761 4363 7772 4383
rect 7792 4363 7810 4383
rect 4707 4333 4756 4343
rect 4707 4313 4718 4333
rect 4738 4313 4756 4333
rect 4707 4301 4756 4313
rect 4806 4337 4850 4343
rect 4806 4317 4821 4337
rect 4841 4317 4850 4337
rect 4806 4301 4850 4317
rect 4925 4333 4974 4343
rect 4925 4313 4936 4333
rect 4956 4313 4974 4333
rect 4925 4301 4974 4313
rect 5024 4337 5068 4343
rect 5024 4317 5039 4337
rect 5059 4317 5068 4337
rect 5024 4301 5068 4317
rect 5138 4337 5182 4343
rect 5138 4317 5147 4337
rect 5167 4317 5182 4337
rect 5138 4301 5182 4317
rect 5232 4333 5281 4343
rect 7761 4353 7810 4363
rect 7860 4379 7904 4395
rect 7860 4359 7875 4379
rect 7895 4359 7904 4379
rect 7860 4353 7904 4359
rect 7974 4379 8018 4395
rect 7974 4359 7983 4379
rect 8003 4359 8018 4379
rect 7974 4353 8018 4359
rect 8068 4383 8117 4395
rect 8068 4363 8086 4383
rect 8106 4363 8117 4383
rect 8068 4353 8117 4363
rect 8192 4379 8236 4395
rect 8192 4359 8201 4379
rect 8221 4359 8236 4379
rect 8192 4353 8236 4359
rect 8286 4383 8335 4395
rect 8286 4363 8304 4383
rect 8324 4363 8335 4383
rect 8286 4353 8335 4363
rect 5232 4313 5250 4333
rect 5270 4313 5281 4333
rect 5232 4301 5281 4313
rect 29508 4799 29519 4819
rect 29539 4799 29557 4819
rect 29508 4789 29557 4799
rect 29607 4815 29651 4831
rect 29607 4795 29622 4815
rect 29642 4795 29651 4815
rect 29607 4789 29651 4795
rect 29721 4815 29765 4831
rect 29721 4795 29730 4815
rect 29750 4795 29765 4815
rect 29721 4789 29765 4795
rect 29815 4819 29864 4831
rect 29815 4799 29833 4819
rect 29853 4799 29864 4819
rect 29815 4789 29864 4799
rect 29939 4815 29983 4831
rect 29939 4795 29948 4815
rect 29968 4795 29983 4815
rect 29939 4789 29983 4795
rect 30033 4819 30082 4831
rect 30033 4799 30051 4819
rect 30071 4799 30082 4819
rect 30033 4789 30082 4799
rect 33872 4832 33921 4844
rect 19970 4566 20019 4578
rect 18816 4554 18865 4564
rect 18816 4534 18827 4554
rect 18847 4534 18865 4554
rect 18816 4522 18865 4534
rect 18915 4558 18959 4564
rect 18915 4538 18930 4558
rect 18950 4538 18959 4558
rect 18915 4522 18959 4538
rect 19034 4554 19083 4564
rect 19034 4534 19045 4554
rect 19065 4534 19083 4554
rect 19034 4522 19083 4534
rect 19133 4558 19177 4564
rect 19133 4538 19148 4558
rect 19168 4538 19177 4558
rect 19133 4522 19177 4538
rect 19247 4558 19291 4564
rect 19247 4538 19256 4558
rect 19276 4538 19291 4558
rect 19247 4522 19291 4538
rect 19341 4554 19390 4564
rect 19341 4534 19359 4554
rect 19379 4534 19390 4554
rect 19970 4546 19981 4566
rect 20001 4546 20019 4566
rect 19970 4536 20019 4546
rect 20069 4562 20113 4578
rect 20069 4542 20084 4562
rect 20104 4542 20113 4562
rect 20069 4536 20113 4542
rect 20183 4562 20227 4578
rect 20183 4542 20192 4562
rect 20212 4542 20227 4562
rect 20183 4536 20227 4542
rect 20277 4566 20326 4578
rect 20277 4546 20295 4566
rect 20315 4546 20326 4566
rect 20277 4536 20326 4546
rect 20401 4562 20445 4578
rect 20401 4542 20410 4562
rect 20430 4542 20445 4562
rect 20401 4536 20445 4542
rect 20495 4566 20544 4578
rect 20495 4546 20513 4566
rect 20533 4546 20544 4566
rect 20495 4536 20544 4546
rect 33872 4812 33883 4832
rect 33903 4812 33921 4832
rect 33872 4802 33921 4812
rect 33971 4828 34015 4844
rect 33971 4808 33986 4828
rect 34006 4808 34015 4828
rect 33971 4802 34015 4808
rect 34085 4828 34129 4844
rect 34085 4808 34094 4828
rect 34114 4808 34129 4828
rect 34085 4802 34129 4808
rect 34179 4832 34228 4844
rect 34179 4812 34197 4832
rect 34217 4812 34228 4832
rect 34179 4802 34228 4812
rect 34303 4828 34347 4844
rect 34303 4808 34312 4828
rect 34332 4808 34347 4828
rect 34303 4802 34347 4808
rect 34397 4832 34446 4844
rect 34397 4812 34415 4832
rect 34435 4812 34446 4832
rect 34397 4802 34446 4812
rect 24334 4579 24383 4591
rect 23180 4567 23229 4577
rect 23180 4547 23191 4567
rect 23211 4547 23229 4567
rect 19341 4522 19390 4534
rect 12138 4395 12187 4407
rect 12138 4375 12149 4395
rect 12169 4375 12187 4395
rect 9084 4345 9133 4355
rect 9084 4325 9095 4345
rect 9115 4325 9133 4345
rect 9084 4313 9133 4325
rect 9183 4349 9227 4355
rect 9183 4329 9198 4349
rect 9218 4329 9227 4349
rect 9183 4313 9227 4329
rect 9302 4345 9351 4355
rect 9302 4325 9313 4345
rect 9333 4325 9351 4345
rect 9302 4313 9351 4325
rect 9401 4349 9445 4355
rect 9401 4329 9416 4349
rect 9436 4329 9445 4349
rect 9401 4313 9445 4329
rect 9515 4349 9559 4355
rect 9515 4329 9524 4349
rect 9544 4329 9559 4349
rect 9515 4313 9559 4329
rect 9609 4345 9658 4355
rect 12138 4365 12187 4375
rect 12237 4391 12281 4407
rect 12237 4371 12252 4391
rect 12272 4371 12281 4391
rect 12237 4365 12281 4371
rect 12351 4391 12395 4407
rect 12351 4371 12360 4391
rect 12380 4371 12395 4391
rect 12351 4365 12395 4371
rect 12445 4395 12494 4407
rect 12445 4375 12463 4395
rect 12483 4375 12494 4395
rect 12445 4365 12494 4375
rect 12569 4391 12613 4407
rect 12569 4371 12578 4391
rect 12598 4371 12613 4391
rect 12569 4365 12613 4371
rect 12663 4395 12712 4407
rect 12663 4375 12681 4395
rect 12701 4375 12712 4395
rect 12663 4365 12712 4375
rect 9609 4325 9627 4345
rect 9647 4325 9658 4345
rect 9609 4313 9658 4325
rect 1141 4136 1190 4146
rect 1141 4116 1152 4136
rect 1172 4116 1190 4136
rect 1141 4104 1190 4116
rect 1240 4140 1284 4146
rect 1240 4120 1255 4140
rect 1275 4120 1284 4140
rect 1240 4104 1284 4120
rect 1359 4136 1408 4146
rect 1359 4116 1370 4136
rect 1390 4116 1408 4136
rect 1359 4104 1408 4116
rect 1458 4140 1502 4146
rect 1458 4120 1473 4140
rect 1493 4120 1502 4140
rect 1458 4104 1502 4120
rect 1572 4140 1616 4146
rect 1572 4120 1581 4140
rect 1601 4120 1616 4140
rect 1572 4104 1616 4120
rect 1666 4136 1715 4146
rect 1666 4116 1684 4136
rect 1704 4116 1715 4136
rect 1666 4104 1715 4116
rect 2500 4144 2549 4156
rect 2500 4124 2511 4144
rect 2531 4124 2549 4144
rect 2500 4114 2549 4124
rect 2599 4140 2643 4156
rect 2599 4120 2614 4140
rect 2634 4120 2643 4140
rect 2599 4114 2643 4120
rect 2713 4140 2757 4156
rect 2713 4120 2722 4140
rect 2742 4120 2757 4140
rect 2713 4114 2757 4120
rect 2807 4144 2856 4156
rect 2807 4124 2825 4144
rect 2845 4124 2856 4144
rect 2807 4114 2856 4124
rect 2931 4140 2975 4156
rect 2931 4120 2940 4140
rect 2960 4120 2975 4140
rect 2931 4114 2975 4120
rect 3025 4144 3074 4156
rect 16502 4408 16551 4420
rect 16502 4388 16513 4408
rect 16533 4388 16551 4408
rect 13448 4358 13497 4368
rect 13448 4338 13459 4358
rect 13479 4338 13497 4358
rect 13448 4326 13497 4338
rect 13547 4362 13591 4368
rect 13547 4342 13562 4362
rect 13582 4342 13591 4362
rect 13547 4326 13591 4342
rect 13666 4358 13715 4368
rect 13666 4338 13677 4358
rect 13697 4338 13715 4358
rect 13666 4326 13715 4338
rect 13765 4362 13809 4368
rect 13765 4342 13780 4362
rect 13800 4342 13809 4362
rect 13765 4326 13809 4342
rect 13879 4362 13923 4368
rect 13879 4342 13888 4362
rect 13908 4342 13923 4362
rect 13879 4326 13923 4342
rect 13973 4358 14022 4368
rect 16502 4378 16551 4388
rect 16601 4404 16645 4420
rect 16601 4384 16616 4404
rect 16636 4384 16645 4404
rect 16601 4378 16645 4384
rect 16715 4404 16759 4420
rect 16715 4384 16724 4404
rect 16744 4384 16759 4404
rect 16715 4378 16759 4384
rect 16809 4408 16858 4420
rect 16809 4388 16827 4408
rect 16847 4388 16858 4408
rect 16809 4378 16858 4388
rect 16933 4404 16977 4420
rect 16933 4384 16942 4404
rect 16962 4384 16977 4404
rect 16933 4378 16977 4384
rect 17027 4408 17076 4420
rect 17027 4388 17045 4408
rect 17065 4388 17076 4408
rect 17027 4378 17076 4388
rect 23180 4535 23229 4547
rect 23279 4571 23323 4577
rect 23279 4551 23294 4571
rect 23314 4551 23323 4571
rect 23279 4535 23323 4551
rect 23398 4567 23447 4577
rect 23398 4547 23409 4567
rect 23429 4547 23447 4567
rect 23398 4535 23447 4547
rect 23497 4571 23541 4577
rect 23497 4551 23512 4571
rect 23532 4551 23541 4571
rect 23497 4535 23541 4551
rect 23611 4571 23655 4577
rect 23611 4551 23620 4571
rect 23640 4551 23655 4571
rect 23611 4535 23655 4551
rect 23705 4567 23754 4577
rect 23705 4547 23723 4567
rect 23743 4547 23754 4567
rect 24334 4559 24345 4579
rect 24365 4559 24383 4579
rect 24334 4549 24383 4559
rect 24433 4575 24477 4591
rect 24433 4555 24448 4575
rect 24468 4555 24477 4575
rect 24433 4549 24477 4555
rect 24547 4575 24591 4591
rect 24547 4555 24556 4575
rect 24576 4555 24591 4575
rect 24547 4549 24591 4555
rect 24641 4579 24690 4591
rect 24641 4559 24659 4579
rect 24679 4559 24690 4579
rect 24641 4549 24690 4559
rect 24765 4575 24809 4591
rect 24765 4555 24774 4575
rect 24794 4555 24809 4575
rect 24765 4549 24809 4555
rect 24859 4579 24908 4591
rect 24859 4559 24877 4579
rect 24897 4559 24908 4579
rect 24859 4549 24908 4559
rect 28711 4591 28760 4603
rect 27557 4579 27606 4589
rect 27557 4559 27568 4579
rect 27588 4559 27606 4579
rect 23705 4535 23754 4547
rect 13973 4338 13991 4358
rect 14011 4338 14022 4358
rect 13973 4326 14022 4338
rect 3025 4124 3043 4144
rect 3063 4124 3074 4144
rect 3025 4114 3074 4124
rect 5505 4149 5554 4159
rect 5505 4129 5516 4149
rect 5536 4129 5554 4149
rect 5505 4117 5554 4129
rect 5604 4153 5648 4159
rect 5604 4133 5619 4153
rect 5639 4133 5648 4153
rect 5604 4117 5648 4133
rect 5723 4149 5772 4159
rect 5723 4129 5734 4149
rect 5754 4129 5772 4149
rect 5723 4117 5772 4129
rect 5822 4153 5866 4159
rect 5822 4133 5837 4153
rect 5857 4133 5866 4153
rect 5822 4117 5866 4133
rect 5936 4153 5980 4159
rect 5936 4133 5945 4153
rect 5965 4133 5980 4153
rect 5936 4117 5980 4133
rect 6030 4149 6079 4159
rect 6030 4129 6048 4149
rect 6068 4129 6079 4149
rect 6030 4117 6079 4129
rect 6864 4157 6913 4169
rect 6864 4137 6875 4157
rect 6895 4137 6913 4157
rect 6864 4127 6913 4137
rect 6963 4153 7007 4169
rect 6963 4133 6978 4153
rect 6998 4133 7007 4153
rect 6963 4127 7007 4133
rect 7077 4153 7121 4169
rect 7077 4133 7086 4153
rect 7106 4133 7121 4153
rect 7077 4127 7121 4133
rect 7171 4157 7220 4169
rect 7171 4137 7189 4157
rect 7209 4137 7220 4157
rect 7171 4127 7220 4137
rect 7295 4153 7339 4169
rect 7295 4133 7304 4153
rect 7324 4133 7339 4153
rect 7295 4127 7339 4133
rect 7389 4157 7438 4169
rect 27557 4547 27606 4559
rect 27656 4583 27700 4589
rect 27656 4563 27671 4583
rect 27691 4563 27700 4583
rect 27656 4547 27700 4563
rect 27775 4579 27824 4589
rect 27775 4559 27786 4579
rect 27806 4559 27824 4579
rect 27775 4547 27824 4559
rect 27874 4583 27918 4589
rect 27874 4563 27889 4583
rect 27909 4563 27918 4583
rect 27874 4547 27918 4563
rect 27988 4583 28032 4589
rect 27988 4563 27997 4583
rect 28017 4563 28032 4583
rect 27988 4547 28032 4563
rect 28082 4579 28131 4589
rect 28082 4559 28100 4579
rect 28120 4559 28131 4579
rect 28711 4571 28722 4591
rect 28742 4571 28760 4591
rect 28711 4561 28760 4571
rect 28810 4587 28854 4603
rect 28810 4567 28825 4587
rect 28845 4567 28854 4587
rect 28810 4561 28854 4567
rect 28924 4587 28968 4603
rect 28924 4567 28933 4587
rect 28953 4567 28968 4587
rect 28924 4561 28968 4567
rect 29018 4591 29067 4603
rect 29018 4571 29036 4591
rect 29056 4571 29067 4591
rect 29018 4561 29067 4571
rect 29142 4587 29186 4603
rect 29142 4567 29151 4587
rect 29171 4567 29186 4587
rect 29142 4561 29186 4567
rect 29236 4591 29285 4603
rect 29236 4571 29254 4591
rect 29274 4571 29285 4591
rect 29236 4561 29285 4571
rect 33075 4604 33124 4616
rect 31921 4592 31970 4602
rect 31921 4572 31932 4592
rect 31952 4572 31970 4592
rect 28082 4547 28131 4559
rect 20768 4382 20817 4394
rect 20768 4362 20779 4382
rect 20799 4362 20817 4382
rect 7389 4137 7407 4157
rect 7427 4137 7438 4157
rect 7389 4127 7438 4137
rect 9882 4161 9931 4171
rect 9882 4141 9893 4161
rect 9913 4141 9931 4161
rect 9882 4129 9931 4141
rect 9981 4165 10025 4171
rect 9981 4145 9996 4165
rect 10016 4145 10025 4165
rect 9981 4129 10025 4145
rect 10100 4161 10149 4171
rect 10100 4141 10111 4161
rect 10131 4141 10149 4161
rect 10100 4129 10149 4141
rect 10199 4165 10243 4171
rect 10199 4145 10214 4165
rect 10234 4145 10243 4165
rect 10199 4129 10243 4145
rect 10313 4165 10357 4171
rect 10313 4145 10322 4165
rect 10342 4145 10357 4165
rect 10313 4129 10357 4145
rect 10407 4161 10456 4171
rect 10407 4141 10425 4161
rect 10445 4141 10456 4161
rect 10407 4129 10456 4141
rect 11241 4169 11290 4181
rect 11241 4149 11252 4169
rect 11272 4149 11290 4169
rect 11241 4139 11290 4149
rect 11340 4165 11384 4181
rect 11340 4145 11355 4165
rect 11375 4145 11384 4165
rect 11340 4139 11384 4145
rect 11454 4165 11498 4181
rect 11454 4145 11463 4165
rect 11483 4145 11498 4165
rect 11454 4139 11498 4145
rect 11548 4169 11597 4181
rect 11548 4149 11566 4169
rect 11586 4149 11597 4169
rect 11548 4139 11597 4149
rect 11672 4165 11716 4181
rect 11672 4145 11681 4165
rect 11701 4145 11716 4165
rect 11672 4139 11716 4145
rect 11766 4169 11815 4181
rect 17714 4332 17763 4342
rect 17714 4312 17725 4332
rect 17745 4312 17763 4332
rect 17714 4300 17763 4312
rect 17813 4336 17857 4342
rect 17813 4316 17828 4336
rect 17848 4316 17857 4336
rect 17813 4300 17857 4316
rect 17932 4332 17981 4342
rect 17932 4312 17943 4332
rect 17963 4312 17981 4332
rect 17932 4300 17981 4312
rect 18031 4336 18075 4342
rect 18031 4316 18046 4336
rect 18066 4316 18075 4336
rect 18031 4300 18075 4316
rect 18145 4336 18189 4342
rect 18145 4316 18154 4336
rect 18174 4316 18189 4336
rect 18145 4300 18189 4316
rect 18239 4332 18288 4342
rect 20768 4352 20817 4362
rect 20867 4378 20911 4394
rect 20867 4358 20882 4378
rect 20902 4358 20911 4378
rect 20867 4352 20911 4358
rect 20981 4378 21025 4394
rect 20981 4358 20990 4378
rect 21010 4358 21025 4378
rect 20981 4352 21025 4358
rect 21075 4382 21124 4394
rect 21075 4362 21093 4382
rect 21113 4362 21124 4382
rect 21075 4352 21124 4362
rect 21199 4378 21243 4394
rect 21199 4358 21208 4378
rect 21228 4358 21243 4378
rect 21199 4352 21243 4358
rect 21293 4382 21342 4394
rect 21293 4362 21311 4382
rect 21331 4362 21342 4382
rect 21293 4352 21342 4362
rect 18239 4312 18257 4332
rect 18277 4312 18288 4332
rect 18239 4300 18288 4312
rect 31921 4560 31970 4572
rect 32020 4596 32064 4602
rect 32020 4576 32035 4596
rect 32055 4576 32064 4596
rect 32020 4560 32064 4576
rect 32139 4592 32188 4602
rect 32139 4572 32150 4592
rect 32170 4572 32188 4592
rect 32139 4560 32188 4572
rect 32238 4596 32282 4602
rect 32238 4576 32253 4596
rect 32273 4576 32282 4596
rect 32238 4560 32282 4576
rect 32352 4596 32396 4602
rect 32352 4576 32361 4596
rect 32381 4576 32396 4596
rect 32352 4560 32396 4576
rect 32446 4592 32495 4602
rect 32446 4572 32464 4592
rect 32484 4572 32495 4592
rect 33075 4584 33086 4604
rect 33106 4584 33124 4604
rect 33075 4574 33124 4584
rect 33174 4600 33218 4616
rect 33174 4580 33189 4600
rect 33209 4580 33218 4600
rect 33174 4574 33218 4580
rect 33288 4600 33332 4616
rect 33288 4580 33297 4600
rect 33317 4580 33332 4600
rect 33288 4574 33332 4580
rect 33382 4604 33431 4616
rect 33382 4584 33400 4604
rect 33420 4584 33431 4604
rect 33382 4574 33431 4584
rect 33506 4600 33550 4616
rect 33506 4580 33515 4600
rect 33535 4580 33550 4600
rect 33506 4574 33550 4580
rect 33600 4604 33649 4616
rect 33600 4584 33618 4604
rect 33638 4584 33649 4604
rect 33600 4574 33649 4584
rect 32446 4560 32495 4572
rect 25132 4395 25181 4407
rect 25132 4375 25143 4395
rect 25163 4375 25181 4395
rect 22078 4345 22127 4355
rect 22078 4325 22089 4345
rect 22109 4325 22127 4345
rect 22078 4313 22127 4325
rect 22177 4349 22221 4355
rect 22177 4329 22192 4349
rect 22212 4329 22221 4349
rect 22177 4313 22221 4329
rect 22296 4345 22345 4355
rect 22296 4325 22307 4345
rect 22327 4325 22345 4345
rect 22296 4313 22345 4325
rect 22395 4349 22439 4355
rect 22395 4329 22410 4349
rect 22430 4329 22439 4349
rect 22395 4313 22439 4329
rect 22509 4349 22553 4355
rect 22509 4329 22518 4349
rect 22538 4329 22553 4349
rect 22509 4313 22553 4329
rect 22603 4345 22652 4355
rect 25132 4365 25181 4375
rect 25231 4391 25275 4407
rect 25231 4371 25246 4391
rect 25266 4371 25275 4391
rect 25231 4365 25275 4371
rect 25345 4391 25389 4407
rect 25345 4371 25354 4391
rect 25374 4371 25389 4391
rect 25345 4365 25389 4371
rect 25439 4395 25488 4407
rect 25439 4375 25457 4395
rect 25477 4375 25488 4395
rect 25439 4365 25488 4375
rect 25563 4391 25607 4407
rect 25563 4371 25572 4391
rect 25592 4371 25607 4391
rect 25563 4365 25607 4371
rect 25657 4395 25706 4407
rect 25657 4375 25675 4395
rect 25695 4375 25706 4395
rect 25657 4365 25706 4375
rect 22603 4325 22621 4345
rect 22641 4325 22652 4345
rect 22603 4313 22652 4325
rect 11766 4149 11784 4169
rect 11804 4149 11815 4169
rect 11766 4139 11815 4149
rect 14246 4174 14295 4184
rect 14246 4154 14257 4174
rect 14277 4154 14295 4174
rect 344 3908 393 3918
rect 344 3888 355 3908
rect 375 3888 393 3908
rect 344 3876 393 3888
rect 443 3912 487 3918
rect 443 3892 458 3912
rect 478 3892 487 3912
rect 443 3876 487 3892
rect 562 3908 611 3918
rect 562 3888 573 3908
rect 593 3888 611 3908
rect 562 3876 611 3888
rect 661 3912 705 3918
rect 661 3892 676 3912
rect 696 3892 705 3912
rect 661 3876 705 3892
rect 775 3912 819 3918
rect 775 3892 784 3912
rect 804 3892 819 3912
rect 775 3876 819 3892
rect 869 3908 918 3918
rect 869 3888 887 3908
rect 907 3888 918 3908
rect 14246 4142 14295 4154
rect 14345 4178 14389 4184
rect 14345 4158 14360 4178
rect 14380 4158 14389 4178
rect 14345 4142 14389 4158
rect 14464 4174 14513 4184
rect 14464 4154 14475 4174
rect 14495 4154 14513 4174
rect 14464 4142 14513 4154
rect 14563 4178 14607 4184
rect 14563 4158 14578 4178
rect 14598 4158 14607 4178
rect 14563 4142 14607 4158
rect 14677 4178 14721 4184
rect 14677 4158 14686 4178
rect 14706 4158 14721 4178
rect 14677 4142 14721 4158
rect 14771 4174 14820 4184
rect 14771 4154 14789 4174
rect 14809 4154 14820 4174
rect 14771 4142 14820 4154
rect 15605 4182 15654 4194
rect 15605 4162 15616 4182
rect 15636 4162 15654 4182
rect 15605 4152 15654 4162
rect 15704 4178 15748 4194
rect 15704 4158 15719 4178
rect 15739 4158 15748 4178
rect 15704 4152 15748 4158
rect 15818 4178 15862 4194
rect 15818 4158 15827 4178
rect 15847 4158 15862 4178
rect 15818 4152 15862 4158
rect 15912 4182 15961 4194
rect 15912 4162 15930 4182
rect 15950 4162 15961 4182
rect 15912 4152 15961 4162
rect 16036 4178 16080 4194
rect 16036 4158 16045 4178
rect 16065 4158 16080 4178
rect 16036 4152 16080 4158
rect 16130 4182 16179 4194
rect 16130 4162 16148 4182
rect 16168 4162 16179 4182
rect 16130 4152 16179 4162
rect 29509 4407 29558 4419
rect 29509 4387 29520 4407
rect 29540 4387 29558 4407
rect 26455 4357 26504 4367
rect 26455 4337 26466 4357
rect 26486 4337 26504 4357
rect 26455 4325 26504 4337
rect 26554 4361 26598 4367
rect 26554 4341 26569 4361
rect 26589 4341 26598 4361
rect 26554 4325 26598 4341
rect 26673 4357 26722 4367
rect 26673 4337 26684 4357
rect 26704 4337 26722 4357
rect 26673 4325 26722 4337
rect 26772 4361 26816 4367
rect 26772 4341 26787 4361
rect 26807 4341 26816 4361
rect 26772 4325 26816 4341
rect 26886 4361 26930 4367
rect 26886 4341 26895 4361
rect 26915 4341 26930 4361
rect 26886 4325 26930 4341
rect 26980 4357 27029 4367
rect 29509 4377 29558 4387
rect 29608 4403 29652 4419
rect 29608 4383 29623 4403
rect 29643 4383 29652 4403
rect 29608 4377 29652 4383
rect 29722 4403 29766 4419
rect 29722 4383 29731 4403
rect 29751 4383 29766 4403
rect 29722 4377 29766 4383
rect 29816 4407 29865 4419
rect 29816 4387 29834 4407
rect 29854 4387 29865 4407
rect 29816 4377 29865 4387
rect 29940 4403 29984 4419
rect 29940 4383 29949 4403
rect 29969 4383 29984 4403
rect 29940 4377 29984 4383
rect 30034 4407 30083 4419
rect 30034 4387 30052 4407
rect 30072 4387 30083 4407
rect 30034 4377 30083 4387
rect 26980 4337 26998 4357
rect 27018 4337 27029 4357
rect 26980 4325 27029 4337
rect 869 3876 918 3888
rect 4708 3921 4757 3931
rect 4708 3901 4719 3921
rect 4739 3901 4757 3921
rect 4708 3889 4757 3901
rect 4807 3925 4851 3931
rect 4807 3905 4822 3925
rect 4842 3905 4851 3925
rect 4807 3889 4851 3905
rect 4926 3921 4975 3931
rect 4926 3901 4937 3921
rect 4957 3901 4975 3921
rect 4926 3889 4975 3901
rect 5025 3925 5069 3931
rect 5025 3905 5040 3925
rect 5060 3905 5069 3925
rect 5025 3889 5069 3905
rect 5139 3925 5183 3931
rect 5139 3905 5148 3925
rect 5168 3905 5183 3925
rect 5139 3889 5183 3905
rect 5233 3921 5282 3931
rect 5233 3901 5251 3921
rect 5271 3901 5282 3921
rect 18512 4148 18561 4158
rect 18512 4128 18523 4148
rect 18543 4128 18561 4148
rect 18512 4116 18561 4128
rect 18611 4152 18655 4158
rect 18611 4132 18626 4152
rect 18646 4132 18655 4152
rect 18611 4116 18655 4132
rect 18730 4148 18779 4158
rect 18730 4128 18741 4148
rect 18761 4128 18779 4148
rect 18730 4116 18779 4128
rect 18829 4152 18873 4158
rect 18829 4132 18844 4152
rect 18864 4132 18873 4152
rect 18829 4116 18873 4132
rect 18943 4152 18987 4158
rect 18943 4132 18952 4152
rect 18972 4132 18987 4152
rect 18943 4116 18987 4132
rect 19037 4148 19086 4158
rect 19037 4128 19055 4148
rect 19075 4128 19086 4148
rect 19037 4116 19086 4128
rect 19871 4156 19920 4168
rect 19871 4136 19882 4156
rect 19902 4136 19920 4156
rect 19871 4126 19920 4136
rect 19970 4152 20014 4168
rect 19970 4132 19985 4152
rect 20005 4132 20014 4152
rect 19970 4126 20014 4132
rect 20084 4152 20128 4168
rect 20084 4132 20093 4152
rect 20113 4132 20128 4152
rect 20084 4126 20128 4132
rect 20178 4156 20227 4168
rect 20178 4136 20196 4156
rect 20216 4136 20227 4156
rect 20178 4126 20227 4136
rect 20302 4152 20346 4168
rect 20302 4132 20311 4152
rect 20331 4132 20346 4152
rect 20302 4126 20346 4132
rect 20396 4156 20445 4168
rect 33873 4420 33922 4432
rect 33873 4400 33884 4420
rect 33904 4400 33922 4420
rect 30819 4370 30868 4380
rect 30819 4350 30830 4370
rect 30850 4350 30868 4370
rect 30819 4338 30868 4350
rect 30918 4374 30962 4380
rect 30918 4354 30933 4374
rect 30953 4354 30962 4374
rect 30918 4338 30962 4354
rect 31037 4370 31086 4380
rect 31037 4350 31048 4370
rect 31068 4350 31086 4370
rect 31037 4338 31086 4350
rect 31136 4374 31180 4380
rect 31136 4354 31151 4374
rect 31171 4354 31180 4374
rect 31136 4338 31180 4354
rect 31250 4374 31294 4380
rect 31250 4354 31259 4374
rect 31279 4354 31294 4374
rect 31250 4338 31294 4354
rect 31344 4370 31393 4380
rect 33873 4390 33922 4400
rect 33972 4416 34016 4432
rect 33972 4396 33987 4416
rect 34007 4396 34016 4416
rect 33972 4390 34016 4396
rect 34086 4416 34130 4432
rect 34086 4396 34095 4416
rect 34115 4396 34130 4416
rect 34086 4390 34130 4396
rect 34180 4420 34229 4432
rect 34180 4400 34198 4420
rect 34218 4400 34229 4420
rect 34180 4390 34229 4400
rect 34304 4416 34348 4432
rect 34304 4396 34313 4416
rect 34333 4396 34348 4416
rect 34304 4390 34348 4396
rect 34398 4420 34447 4432
rect 34398 4400 34416 4420
rect 34436 4400 34447 4420
rect 34398 4390 34447 4400
rect 31344 4350 31362 4370
rect 31382 4350 31393 4370
rect 31344 4338 31393 4350
rect 20396 4136 20414 4156
rect 20434 4136 20445 4156
rect 20396 4126 20445 4136
rect 22876 4161 22925 4171
rect 22876 4141 22887 4161
rect 22907 4141 22925 4161
rect 5233 3889 5282 3901
rect 9085 3933 9134 3943
rect 9085 3913 9096 3933
rect 9116 3913 9134 3933
rect 9085 3901 9134 3913
rect 9184 3937 9228 3943
rect 9184 3917 9199 3937
rect 9219 3917 9228 3937
rect 9184 3901 9228 3917
rect 9303 3933 9352 3943
rect 9303 3913 9314 3933
rect 9334 3913 9352 3933
rect 9303 3901 9352 3913
rect 9402 3937 9446 3943
rect 9402 3917 9417 3937
rect 9437 3917 9446 3937
rect 9402 3901 9446 3917
rect 9516 3937 9560 3943
rect 9516 3917 9525 3937
rect 9545 3917 9560 3937
rect 9516 3901 9560 3917
rect 9610 3933 9659 3943
rect 9610 3913 9628 3933
rect 9648 3913 9659 3933
rect 22876 4129 22925 4141
rect 22975 4165 23019 4171
rect 22975 4145 22990 4165
rect 23010 4145 23019 4165
rect 22975 4129 23019 4145
rect 23094 4161 23143 4171
rect 23094 4141 23105 4161
rect 23125 4141 23143 4161
rect 23094 4129 23143 4141
rect 23193 4165 23237 4171
rect 23193 4145 23208 4165
rect 23228 4145 23237 4165
rect 23193 4129 23237 4145
rect 23307 4165 23351 4171
rect 23307 4145 23316 4165
rect 23336 4145 23351 4165
rect 23307 4129 23351 4145
rect 23401 4161 23450 4171
rect 23401 4141 23419 4161
rect 23439 4141 23450 4161
rect 23401 4129 23450 4141
rect 24235 4169 24284 4181
rect 24235 4149 24246 4169
rect 24266 4149 24284 4169
rect 24235 4139 24284 4149
rect 24334 4165 24378 4181
rect 24334 4145 24349 4165
rect 24369 4145 24378 4165
rect 24334 4139 24378 4145
rect 24448 4165 24492 4181
rect 24448 4145 24457 4165
rect 24477 4145 24492 4165
rect 24448 4139 24492 4145
rect 24542 4169 24591 4181
rect 24542 4149 24560 4169
rect 24580 4149 24591 4169
rect 24542 4139 24591 4149
rect 24666 4165 24710 4181
rect 24666 4145 24675 4165
rect 24695 4145 24710 4165
rect 24666 4139 24710 4145
rect 24760 4169 24809 4181
rect 24760 4149 24778 4169
rect 24798 4149 24809 4169
rect 24760 4139 24809 4149
rect 9610 3901 9659 3913
rect 13449 3946 13498 3956
rect 13449 3926 13460 3946
rect 13480 3926 13498 3946
rect 13449 3914 13498 3926
rect 13548 3950 13592 3956
rect 13548 3930 13563 3950
rect 13583 3930 13592 3950
rect 13548 3914 13592 3930
rect 13667 3946 13716 3956
rect 13667 3926 13678 3946
rect 13698 3926 13716 3946
rect 13667 3914 13716 3926
rect 13766 3950 13810 3956
rect 13766 3930 13781 3950
rect 13801 3930 13810 3950
rect 13766 3914 13810 3930
rect 13880 3950 13924 3956
rect 13880 3930 13889 3950
rect 13909 3930 13924 3950
rect 13880 3914 13924 3930
rect 13974 3946 14023 3956
rect 13974 3926 13992 3946
rect 14012 3926 14023 3946
rect 13974 3914 14023 3926
rect 27253 4173 27302 4183
rect 27253 4153 27264 4173
rect 27284 4153 27302 4173
rect 27253 4141 27302 4153
rect 27352 4177 27396 4183
rect 27352 4157 27367 4177
rect 27387 4157 27396 4177
rect 27352 4141 27396 4157
rect 27471 4173 27520 4183
rect 27471 4153 27482 4173
rect 27502 4153 27520 4173
rect 27471 4141 27520 4153
rect 27570 4177 27614 4183
rect 27570 4157 27585 4177
rect 27605 4157 27614 4177
rect 27570 4141 27614 4157
rect 27684 4177 27728 4183
rect 27684 4157 27693 4177
rect 27713 4157 27728 4177
rect 27684 4141 27728 4157
rect 27778 4173 27827 4183
rect 27778 4153 27796 4173
rect 27816 4153 27827 4173
rect 27778 4141 27827 4153
rect 28612 4181 28661 4193
rect 28612 4161 28623 4181
rect 28643 4161 28661 4181
rect 28612 4151 28661 4161
rect 28711 4177 28755 4193
rect 28711 4157 28726 4177
rect 28746 4157 28755 4177
rect 28711 4151 28755 4157
rect 28825 4177 28869 4193
rect 28825 4157 28834 4177
rect 28854 4157 28869 4177
rect 28825 4151 28869 4157
rect 28919 4181 28968 4193
rect 28919 4161 28937 4181
rect 28957 4161 28968 4181
rect 28919 4151 28968 4161
rect 29043 4177 29087 4193
rect 29043 4157 29052 4177
rect 29072 4157 29087 4177
rect 29043 4151 29087 4157
rect 29137 4181 29186 4193
rect 29137 4161 29155 4181
rect 29175 4161 29186 4181
rect 29137 4151 29186 4161
rect 31617 4186 31666 4196
rect 31617 4166 31628 4186
rect 31648 4166 31666 4186
rect 17715 3920 17764 3930
rect 17715 3900 17726 3920
rect 17746 3900 17764 3920
rect 17715 3888 17764 3900
rect 17814 3924 17858 3930
rect 17814 3904 17829 3924
rect 17849 3904 17858 3924
rect 17814 3888 17858 3904
rect 17933 3920 17982 3930
rect 17933 3900 17944 3920
rect 17964 3900 17982 3920
rect 17933 3888 17982 3900
rect 18032 3924 18076 3930
rect 18032 3904 18047 3924
rect 18067 3904 18076 3924
rect 18032 3888 18076 3904
rect 18146 3924 18190 3930
rect 18146 3904 18155 3924
rect 18175 3904 18190 3924
rect 18146 3888 18190 3904
rect 18240 3920 18289 3930
rect 18240 3900 18258 3920
rect 18278 3900 18289 3920
rect 31617 4154 31666 4166
rect 31716 4190 31760 4196
rect 31716 4170 31731 4190
rect 31751 4170 31760 4190
rect 31716 4154 31760 4170
rect 31835 4186 31884 4196
rect 31835 4166 31846 4186
rect 31866 4166 31884 4186
rect 31835 4154 31884 4166
rect 31934 4190 31978 4196
rect 31934 4170 31949 4190
rect 31969 4170 31978 4190
rect 31934 4154 31978 4170
rect 32048 4190 32092 4196
rect 32048 4170 32057 4190
rect 32077 4170 32092 4190
rect 32048 4154 32092 4170
rect 32142 4186 32191 4196
rect 32142 4166 32160 4186
rect 32180 4166 32191 4186
rect 32142 4154 32191 4166
rect 32976 4194 33025 4206
rect 32976 4174 32987 4194
rect 33007 4174 33025 4194
rect 32976 4164 33025 4174
rect 33075 4190 33119 4206
rect 33075 4170 33090 4190
rect 33110 4170 33119 4190
rect 33075 4164 33119 4170
rect 33189 4190 33233 4206
rect 33189 4170 33198 4190
rect 33218 4170 33233 4190
rect 33189 4164 33233 4170
rect 33283 4194 33332 4206
rect 33283 4174 33301 4194
rect 33321 4174 33332 4194
rect 33283 4164 33332 4174
rect 33407 4190 33451 4206
rect 33407 4170 33416 4190
rect 33436 4170 33451 4190
rect 33407 4164 33451 4170
rect 33501 4194 33550 4206
rect 33501 4174 33519 4194
rect 33539 4174 33550 4194
rect 33501 4164 33550 4174
rect 18240 3888 18289 3900
rect 22079 3933 22128 3943
rect 22079 3913 22090 3933
rect 22110 3913 22128 3933
rect 22079 3901 22128 3913
rect 22178 3937 22222 3943
rect 22178 3917 22193 3937
rect 22213 3917 22222 3937
rect 22178 3901 22222 3917
rect 22297 3933 22346 3943
rect 22297 3913 22308 3933
rect 22328 3913 22346 3933
rect 22297 3901 22346 3913
rect 22396 3937 22440 3943
rect 22396 3917 22411 3937
rect 22431 3917 22440 3937
rect 22396 3901 22440 3917
rect 22510 3937 22554 3943
rect 22510 3917 22519 3937
rect 22539 3917 22554 3937
rect 22510 3901 22554 3917
rect 22604 3933 22653 3943
rect 22604 3913 22622 3933
rect 22642 3913 22653 3933
rect 22604 3901 22653 3913
rect 26456 3945 26505 3955
rect 26456 3925 26467 3945
rect 26487 3925 26505 3945
rect 26456 3913 26505 3925
rect 26555 3949 26599 3955
rect 26555 3929 26570 3949
rect 26590 3929 26599 3949
rect 26555 3913 26599 3929
rect 26674 3945 26723 3955
rect 26674 3925 26685 3945
rect 26705 3925 26723 3945
rect 26674 3913 26723 3925
rect 26773 3949 26817 3955
rect 26773 3929 26788 3949
rect 26808 3929 26817 3949
rect 26773 3913 26817 3929
rect 26887 3949 26931 3955
rect 26887 3929 26896 3949
rect 26916 3929 26931 3949
rect 26887 3913 26931 3929
rect 26981 3945 27030 3955
rect 26981 3925 26999 3945
rect 27019 3925 27030 3945
rect 26981 3913 27030 3925
rect 30820 3958 30869 3968
rect 30820 3938 30831 3958
rect 30851 3938 30869 3958
rect 30820 3926 30869 3938
rect 30919 3962 30963 3968
rect 30919 3942 30934 3962
rect 30954 3942 30963 3962
rect 30919 3926 30963 3942
rect 31038 3958 31087 3968
rect 31038 3938 31049 3958
rect 31069 3938 31087 3958
rect 31038 3926 31087 3938
rect 31137 3962 31181 3968
rect 31137 3942 31152 3962
rect 31172 3942 31181 3962
rect 31137 3926 31181 3942
rect 31251 3962 31295 3968
rect 31251 3942 31260 3962
rect 31280 3942 31295 3962
rect 31251 3926 31295 3942
rect 31345 3958 31394 3968
rect 31345 3938 31363 3958
rect 31383 3938 31394 3958
rect 31345 3926 31394 3938
rect 3379 3764 3428 3776
rect 3379 3744 3390 3764
rect 3410 3744 3428 3764
rect 3379 3734 3428 3744
rect 3478 3760 3522 3776
rect 3478 3740 3493 3760
rect 3513 3740 3522 3760
rect 3478 3734 3522 3740
rect 3592 3760 3636 3776
rect 3592 3740 3601 3760
rect 3621 3740 3636 3760
rect 3592 3734 3636 3740
rect 3686 3764 3735 3776
rect 3686 3744 3704 3764
rect 3724 3744 3735 3764
rect 3686 3734 3735 3744
rect 3810 3760 3854 3776
rect 3810 3740 3819 3760
rect 3839 3740 3854 3760
rect 3810 3734 3854 3740
rect 3904 3764 3953 3776
rect 3904 3744 3922 3764
rect 3942 3744 3953 3764
rect 3904 3734 3953 3744
rect 7743 3777 7792 3789
rect 7743 3757 7754 3777
rect 7774 3757 7792 3777
rect 7743 3747 7792 3757
rect 7842 3773 7886 3789
rect 7842 3753 7857 3773
rect 7877 3753 7886 3773
rect 7842 3747 7886 3753
rect 7956 3773 8000 3789
rect 7956 3753 7965 3773
rect 7985 3753 8000 3773
rect 7956 3747 8000 3753
rect 8050 3777 8099 3789
rect 8050 3757 8068 3777
rect 8088 3757 8099 3777
rect 8050 3747 8099 3757
rect 8174 3773 8218 3789
rect 8174 3753 8183 3773
rect 8203 3753 8218 3773
rect 8174 3747 8218 3753
rect 8268 3777 8317 3789
rect 8268 3757 8286 3777
rect 8306 3757 8317 3777
rect 8268 3747 8317 3757
rect 12120 3789 12169 3801
rect 12120 3769 12131 3789
rect 12151 3769 12169 3789
rect 12120 3759 12169 3769
rect 12219 3785 12263 3801
rect 12219 3765 12234 3785
rect 12254 3765 12263 3785
rect 12219 3759 12263 3765
rect 12333 3785 12377 3801
rect 12333 3765 12342 3785
rect 12362 3765 12377 3785
rect 12333 3759 12377 3765
rect 12427 3789 12476 3801
rect 12427 3769 12445 3789
rect 12465 3769 12476 3789
rect 12427 3759 12476 3769
rect 12551 3785 12595 3801
rect 12551 3765 12560 3785
rect 12580 3765 12595 3785
rect 12551 3759 12595 3765
rect 12645 3789 12694 3801
rect 12645 3769 12663 3789
rect 12683 3769 12694 3789
rect 12645 3759 12694 3769
rect 16484 3802 16533 3814
rect 1223 3528 1272 3538
rect 1223 3508 1234 3528
rect 1254 3508 1272 3528
rect 1223 3496 1272 3508
rect 1322 3532 1366 3538
rect 1322 3512 1337 3532
rect 1357 3512 1366 3532
rect 1322 3496 1366 3512
rect 1441 3528 1490 3538
rect 1441 3508 1452 3528
rect 1472 3508 1490 3528
rect 1441 3496 1490 3508
rect 1540 3532 1584 3538
rect 1540 3512 1555 3532
rect 1575 3512 1584 3532
rect 1540 3496 1584 3512
rect 1654 3532 1698 3538
rect 1654 3512 1663 3532
rect 1683 3512 1698 3532
rect 1654 3496 1698 3512
rect 1748 3528 1797 3538
rect 1748 3508 1766 3528
rect 1786 3508 1797 3528
rect 1748 3496 1797 3508
rect 2582 3536 2631 3548
rect 2582 3516 2593 3536
rect 2613 3516 2631 3536
rect 2582 3506 2631 3516
rect 2681 3532 2725 3548
rect 2681 3512 2696 3532
rect 2716 3512 2725 3532
rect 2681 3506 2725 3512
rect 2795 3532 2839 3548
rect 2795 3512 2804 3532
rect 2824 3512 2839 3532
rect 2795 3506 2839 3512
rect 2889 3536 2938 3548
rect 2889 3516 2907 3536
rect 2927 3516 2938 3536
rect 2889 3506 2938 3516
rect 3013 3532 3057 3548
rect 3013 3512 3022 3532
rect 3042 3512 3057 3532
rect 3013 3506 3057 3512
rect 3107 3536 3156 3548
rect 16484 3782 16495 3802
rect 16515 3782 16533 3802
rect 16484 3772 16533 3782
rect 16583 3798 16627 3814
rect 16583 3778 16598 3798
rect 16618 3778 16627 3798
rect 16583 3772 16627 3778
rect 16697 3798 16741 3814
rect 16697 3778 16706 3798
rect 16726 3778 16741 3798
rect 16697 3772 16741 3778
rect 16791 3802 16840 3814
rect 16791 3782 16809 3802
rect 16829 3782 16840 3802
rect 16791 3772 16840 3782
rect 16915 3798 16959 3814
rect 16915 3778 16924 3798
rect 16944 3778 16959 3798
rect 16915 3772 16959 3778
rect 17009 3802 17058 3814
rect 17009 3782 17027 3802
rect 17047 3782 17058 3802
rect 17009 3772 17058 3782
rect 3107 3516 3125 3536
rect 3145 3516 3156 3536
rect 3107 3506 3156 3516
rect 5587 3541 5636 3551
rect 5587 3521 5598 3541
rect 5618 3521 5636 3541
rect 5587 3509 5636 3521
rect 5686 3545 5730 3551
rect 5686 3525 5701 3545
rect 5721 3525 5730 3545
rect 5686 3509 5730 3525
rect 5805 3541 5854 3551
rect 5805 3521 5816 3541
rect 5836 3521 5854 3541
rect 5805 3509 5854 3521
rect 5904 3545 5948 3551
rect 5904 3525 5919 3545
rect 5939 3525 5948 3545
rect 5904 3509 5948 3525
rect 6018 3545 6062 3551
rect 6018 3525 6027 3545
rect 6047 3525 6062 3545
rect 6018 3509 6062 3525
rect 6112 3541 6161 3551
rect 6112 3521 6130 3541
rect 6150 3521 6161 3541
rect 6112 3509 6161 3521
rect 6946 3549 6995 3561
rect 6946 3529 6957 3549
rect 6977 3529 6995 3549
rect 6946 3519 6995 3529
rect 7045 3545 7089 3561
rect 7045 3525 7060 3545
rect 7080 3525 7089 3545
rect 7045 3519 7089 3525
rect 7159 3545 7203 3561
rect 7159 3525 7168 3545
rect 7188 3525 7203 3545
rect 7159 3519 7203 3525
rect 7253 3549 7302 3561
rect 7253 3529 7271 3549
rect 7291 3529 7302 3549
rect 7253 3519 7302 3529
rect 7377 3545 7421 3561
rect 7377 3525 7386 3545
rect 7406 3525 7421 3545
rect 7377 3519 7421 3525
rect 7471 3549 7520 3561
rect 7471 3529 7489 3549
rect 7509 3529 7520 3549
rect 7471 3519 7520 3529
rect 20750 3776 20799 3788
rect 20750 3756 20761 3776
rect 20781 3756 20799 3776
rect 20750 3746 20799 3756
rect 20849 3772 20893 3788
rect 20849 3752 20864 3772
rect 20884 3752 20893 3772
rect 20849 3746 20893 3752
rect 20963 3772 21007 3788
rect 20963 3752 20972 3772
rect 20992 3752 21007 3772
rect 20963 3746 21007 3752
rect 21057 3776 21106 3788
rect 21057 3756 21075 3776
rect 21095 3756 21106 3776
rect 21057 3746 21106 3756
rect 21181 3772 21225 3788
rect 21181 3752 21190 3772
rect 21210 3752 21225 3772
rect 21181 3746 21225 3752
rect 21275 3776 21324 3788
rect 21275 3756 21293 3776
rect 21313 3756 21324 3776
rect 21275 3746 21324 3756
rect 25114 3789 25163 3801
rect 9964 3553 10013 3563
rect 9964 3533 9975 3553
rect 9995 3533 10013 3553
rect 9964 3521 10013 3533
rect 10063 3557 10107 3563
rect 10063 3537 10078 3557
rect 10098 3537 10107 3557
rect 10063 3521 10107 3537
rect 10182 3553 10231 3563
rect 10182 3533 10193 3553
rect 10213 3533 10231 3553
rect 10182 3521 10231 3533
rect 10281 3557 10325 3563
rect 10281 3537 10296 3557
rect 10316 3537 10325 3557
rect 10281 3521 10325 3537
rect 10395 3557 10439 3563
rect 10395 3537 10404 3557
rect 10424 3537 10439 3557
rect 10395 3521 10439 3537
rect 10489 3553 10538 3563
rect 10489 3533 10507 3553
rect 10527 3533 10538 3553
rect 10489 3521 10538 3533
rect 11323 3561 11372 3573
rect 11323 3541 11334 3561
rect 11354 3541 11372 3561
rect 11323 3531 11372 3541
rect 11422 3557 11466 3573
rect 11422 3537 11437 3557
rect 11457 3537 11466 3557
rect 11422 3531 11466 3537
rect 11536 3557 11580 3573
rect 11536 3537 11545 3557
rect 11565 3537 11580 3557
rect 11536 3531 11580 3537
rect 11630 3561 11679 3573
rect 11630 3541 11648 3561
rect 11668 3541 11679 3561
rect 11630 3531 11679 3541
rect 11754 3557 11798 3573
rect 11754 3537 11763 3557
rect 11783 3537 11798 3557
rect 11754 3531 11798 3537
rect 11848 3561 11897 3573
rect 25114 3769 25125 3789
rect 25145 3769 25163 3789
rect 25114 3759 25163 3769
rect 25213 3785 25257 3801
rect 25213 3765 25228 3785
rect 25248 3765 25257 3785
rect 25213 3759 25257 3765
rect 25327 3785 25371 3801
rect 25327 3765 25336 3785
rect 25356 3765 25371 3785
rect 25327 3759 25371 3765
rect 25421 3789 25470 3801
rect 25421 3769 25439 3789
rect 25459 3769 25470 3789
rect 25421 3759 25470 3769
rect 25545 3785 25589 3801
rect 25545 3765 25554 3785
rect 25574 3765 25589 3785
rect 25545 3759 25589 3765
rect 25639 3789 25688 3801
rect 25639 3769 25657 3789
rect 25677 3769 25688 3789
rect 25639 3759 25688 3769
rect 29491 3801 29540 3813
rect 11848 3541 11866 3561
rect 11886 3541 11897 3561
rect 11848 3531 11897 3541
rect 14328 3566 14377 3576
rect 14328 3546 14339 3566
rect 14359 3546 14377 3566
rect 3380 3352 3429 3364
rect 3380 3332 3391 3352
rect 3411 3332 3429 3352
rect 326 3302 375 3312
rect 326 3282 337 3302
rect 357 3282 375 3302
rect 326 3270 375 3282
rect 425 3306 469 3312
rect 425 3286 440 3306
rect 460 3286 469 3306
rect 425 3270 469 3286
rect 544 3302 593 3312
rect 544 3282 555 3302
rect 575 3282 593 3302
rect 544 3270 593 3282
rect 643 3306 687 3312
rect 643 3286 658 3306
rect 678 3286 687 3306
rect 643 3270 687 3286
rect 757 3306 801 3312
rect 757 3286 766 3306
rect 786 3286 801 3306
rect 757 3270 801 3286
rect 851 3302 900 3312
rect 3380 3322 3429 3332
rect 3479 3348 3523 3364
rect 3479 3328 3494 3348
rect 3514 3328 3523 3348
rect 3479 3322 3523 3328
rect 3593 3348 3637 3364
rect 3593 3328 3602 3348
rect 3622 3328 3637 3348
rect 3593 3322 3637 3328
rect 3687 3352 3736 3364
rect 3687 3332 3705 3352
rect 3725 3332 3736 3352
rect 3687 3322 3736 3332
rect 3811 3348 3855 3364
rect 3811 3328 3820 3348
rect 3840 3328 3855 3348
rect 3811 3322 3855 3328
rect 3905 3352 3954 3364
rect 3905 3332 3923 3352
rect 3943 3332 3954 3352
rect 3905 3322 3954 3332
rect 851 3282 869 3302
rect 889 3282 900 3302
rect 851 3270 900 3282
rect 14328 3534 14377 3546
rect 14427 3570 14471 3576
rect 14427 3550 14442 3570
rect 14462 3550 14471 3570
rect 14427 3534 14471 3550
rect 14546 3566 14595 3576
rect 14546 3546 14557 3566
rect 14577 3546 14595 3566
rect 14546 3534 14595 3546
rect 14645 3570 14689 3576
rect 14645 3550 14660 3570
rect 14680 3550 14689 3570
rect 14645 3534 14689 3550
rect 14759 3570 14803 3576
rect 14759 3550 14768 3570
rect 14788 3550 14803 3570
rect 14759 3534 14803 3550
rect 14853 3566 14902 3576
rect 14853 3546 14871 3566
rect 14891 3546 14902 3566
rect 14853 3534 14902 3546
rect 15687 3574 15736 3586
rect 15687 3554 15698 3574
rect 15718 3554 15736 3574
rect 15687 3544 15736 3554
rect 15786 3570 15830 3586
rect 15786 3550 15801 3570
rect 15821 3550 15830 3570
rect 15786 3544 15830 3550
rect 15900 3570 15944 3586
rect 15900 3550 15909 3570
rect 15929 3550 15944 3570
rect 15900 3544 15944 3550
rect 15994 3574 16043 3586
rect 15994 3554 16012 3574
rect 16032 3554 16043 3574
rect 15994 3544 16043 3554
rect 16118 3570 16162 3586
rect 16118 3550 16127 3570
rect 16147 3550 16162 3570
rect 16118 3544 16162 3550
rect 16212 3574 16261 3586
rect 16212 3554 16230 3574
rect 16250 3554 16261 3574
rect 16212 3544 16261 3554
rect 29491 3781 29502 3801
rect 29522 3781 29540 3801
rect 29491 3771 29540 3781
rect 29590 3797 29634 3813
rect 29590 3777 29605 3797
rect 29625 3777 29634 3797
rect 29590 3771 29634 3777
rect 29704 3797 29748 3813
rect 29704 3777 29713 3797
rect 29733 3777 29748 3797
rect 29704 3771 29748 3777
rect 29798 3801 29847 3813
rect 29798 3781 29816 3801
rect 29836 3781 29847 3801
rect 29798 3771 29847 3781
rect 29922 3797 29966 3813
rect 29922 3777 29931 3797
rect 29951 3777 29966 3797
rect 29922 3771 29966 3777
rect 30016 3801 30065 3813
rect 30016 3781 30034 3801
rect 30054 3781 30065 3801
rect 30016 3771 30065 3781
rect 33855 3814 33904 3826
rect 7744 3365 7793 3377
rect 7744 3345 7755 3365
rect 7775 3345 7793 3365
rect 4690 3315 4739 3325
rect 4690 3295 4701 3315
rect 4721 3295 4739 3315
rect 4690 3283 4739 3295
rect 4789 3319 4833 3325
rect 4789 3299 4804 3319
rect 4824 3299 4833 3319
rect 4789 3283 4833 3299
rect 4908 3315 4957 3325
rect 4908 3295 4919 3315
rect 4939 3295 4957 3315
rect 4908 3283 4957 3295
rect 5007 3319 5051 3325
rect 5007 3299 5022 3319
rect 5042 3299 5051 3319
rect 5007 3283 5051 3299
rect 5121 3319 5165 3325
rect 5121 3299 5130 3319
rect 5150 3299 5165 3319
rect 5121 3283 5165 3299
rect 5215 3315 5264 3325
rect 7744 3335 7793 3345
rect 7843 3361 7887 3377
rect 7843 3341 7858 3361
rect 7878 3341 7887 3361
rect 7843 3335 7887 3341
rect 7957 3361 8001 3377
rect 7957 3341 7966 3361
rect 7986 3341 8001 3361
rect 7957 3335 8001 3341
rect 8051 3365 8100 3377
rect 8051 3345 8069 3365
rect 8089 3345 8100 3365
rect 8051 3335 8100 3345
rect 8175 3361 8219 3377
rect 8175 3341 8184 3361
rect 8204 3341 8219 3361
rect 8175 3335 8219 3341
rect 8269 3365 8318 3377
rect 8269 3345 8287 3365
rect 8307 3345 8318 3365
rect 8269 3335 8318 3345
rect 5215 3295 5233 3315
rect 5253 3295 5264 3315
rect 5215 3283 5264 3295
rect 18594 3540 18643 3550
rect 18594 3520 18605 3540
rect 18625 3520 18643 3540
rect 18594 3508 18643 3520
rect 18693 3544 18737 3550
rect 18693 3524 18708 3544
rect 18728 3524 18737 3544
rect 18693 3508 18737 3524
rect 18812 3540 18861 3550
rect 18812 3520 18823 3540
rect 18843 3520 18861 3540
rect 18812 3508 18861 3520
rect 18911 3544 18955 3550
rect 18911 3524 18926 3544
rect 18946 3524 18955 3544
rect 18911 3508 18955 3524
rect 19025 3544 19069 3550
rect 19025 3524 19034 3544
rect 19054 3524 19069 3544
rect 19025 3508 19069 3524
rect 19119 3540 19168 3550
rect 19119 3520 19137 3540
rect 19157 3520 19168 3540
rect 19119 3508 19168 3520
rect 19953 3548 20002 3560
rect 19953 3528 19964 3548
rect 19984 3528 20002 3548
rect 19953 3518 20002 3528
rect 20052 3544 20096 3560
rect 20052 3524 20067 3544
rect 20087 3524 20096 3544
rect 20052 3518 20096 3524
rect 20166 3544 20210 3560
rect 20166 3524 20175 3544
rect 20195 3524 20210 3544
rect 20166 3518 20210 3524
rect 20260 3548 20309 3560
rect 20260 3528 20278 3548
rect 20298 3528 20309 3548
rect 20260 3518 20309 3528
rect 20384 3544 20428 3560
rect 20384 3524 20393 3544
rect 20413 3524 20428 3544
rect 20384 3518 20428 3524
rect 20478 3548 20527 3560
rect 33855 3794 33866 3814
rect 33886 3794 33904 3814
rect 33855 3784 33904 3794
rect 33954 3810 33998 3826
rect 33954 3790 33969 3810
rect 33989 3790 33998 3810
rect 33954 3784 33998 3790
rect 34068 3810 34112 3826
rect 34068 3790 34077 3810
rect 34097 3790 34112 3810
rect 34068 3784 34112 3790
rect 34162 3814 34211 3826
rect 34162 3794 34180 3814
rect 34200 3794 34211 3814
rect 34162 3784 34211 3794
rect 34286 3810 34330 3826
rect 34286 3790 34295 3810
rect 34315 3790 34330 3810
rect 34286 3784 34330 3790
rect 34380 3814 34429 3826
rect 34380 3794 34398 3814
rect 34418 3794 34429 3814
rect 34380 3784 34429 3794
rect 20478 3528 20496 3548
rect 20516 3528 20527 3548
rect 20478 3518 20527 3528
rect 22958 3553 23007 3563
rect 22958 3533 22969 3553
rect 22989 3533 23007 3553
rect 12121 3377 12170 3389
rect 12121 3357 12132 3377
rect 12152 3357 12170 3377
rect 9067 3327 9116 3337
rect 9067 3307 9078 3327
rect 9098 3307 9116 3327
rect 9067 3295 9116 3307
rect 9166 3331 9210 3337
rect 9166 3311 9181 3331
rect 9201 3311 9210 3331
rect 9166 3295 9210 3311
rect 9285 3327 9334 3337
rect 9285 3307 9296 3327
rect 9316 3307 9334 3327
rect 9285 3295 9334 3307
rect 9384 3331 9428 3337
rect 9384 3311 9399 3331
rect 9419 3311 9428 3331
rect 9384 3295 9428 3311
rect 9498 3331 9542 3337
rect 9498 3311 9507 3331
rect 9527 3311 9542 3331
rect 9498 3295 9542 3311
rect 9592 3327 9641 3337
rect 12121 3347 12170 3357
rect 12220 3373 12264 3389
rect 12220 3353 12235 3373
rect 12255 3353 12264 3373
rect 12220 3347 12264 3353
rect 12334 3373 12378 3389
rect 12334 3353 12343 3373
rect 12363 3353 12378 3373
rect 12334 3347 12378 3353
rect 12428 3377 12477 3389
rect 12428 3357 12446 3377
rect 12466 3357 12477 3377
rect 12428 3347 12477 3357
rect 12552 3373 12596 3389
rect 12552 3353 12561 3373
rect 12581 3353 12596 3373
rect 12552 3347 12596 3353
rect 12646 3377 12695 3389
rect 12646 3357 12664 3377
rect 12684 3357 12695 3377
rect 12646 3347 12695 3357
rect 9592 3307 9610 3327
rect 9630 3307 9641 3327
rect 9592 3295 9641 3307
rect 2417 3128 2466 3140
rect 1124 3118 1173 3128
rect 1124 3098 1135 3118
rect 1155 3098 1173 3118
rect 1124 3086 1173 3098
rect 1223 3122 1267 3128
rect 1223 3102 1238 3122
rect 1258 3102 1267 3122
rect 1223 3086 1267 3102
rect 1342 3118 1391 3128
rect 1342 3098 1353 3118
rect 1373 3098 1391 3118
rect 1342 3086 1391 3098
rect 1441 3122 1485 3128
rect 1441 3102 1456 3122
rect 1476 3102 1485 3122
rect 1441 3086 1485 3102
rect 1555 3122 1599 3128
rect 1555 3102 1564 3122
rect 1584 3102 1599 3122
rect 1555 3086 1599 3102
rect 1649 3118 1698 3128
rect 1649 3098 1667 3118
rect 1687 3098 1698 3118
rect 2417 3108 2428 3128
rect 2448 3108 2466 3128
rect 2417 3098 2466 3108
rect 2516 3124 2560 3140
rect 2516 3104 2531 3124
rect 2551 3104 2560 3124
rect 2516 3098 2560 3104
rect 2630 3124 2674 3140
rect 2630 3104 2639 3124
rect 2659 3104 2674 3124
rect 2630 3098 2674 3104
rect 2724 3128 2773 3140
rect 2724 3108 2742 3128
rect 2762 3108 2773 3128
rect 2724 3098 2773 3108
rect 2848 3124 2892 3140
rect 2848 3104 2857 3124
rect 2877 3104 2892 3124
rect 2848 3098 2892 3104
rect 2942 3128 2991 3140
rect 16485 3390 16534 3402
rect 16485 3370 16496 3390
rect 16516 3370 16534 3390
rect 13431 3340 13480 3350
rect 13431 3320 13442 3340
rect 13462 3320 13480 3340
rect 13431 3308 13480 3320
rect 13530 3344 13574 3350
rect 13530 3324 13545 3344
rect 13565 3324 13574 3344
rect 13530 3308 13574 3324
rect 13649 3340 13698 3350
rect 13649 3320 13660 3340
rect 13680 3320 13698 3340
rect 13649 3308 13698 3320
rect 13748 3344 13792 3350
rect 13748 3324 13763 3344
rect 13783 3324 13792 3344
rect 13748 3308 13792 3324
rect 13862 3344 13906 3350
rect 13862 3324 13871 3344
rect 13891 3324 13906 3344
rect 13862 3308 13906 3324
rect 13956 3340 14005 3350
rect 16485 3360 16534 3370
rect 16584 3386 16628 3402
rect 16584 3366 16599 3386
rect 16619 3366 16628 3386
rect 16584 3360 16628 3366
rect 16698 3386 16742 3402
rect 16698 3366 16707 3386
rect 16727 3366 16742 3386
rect 16698 3360 16742 3366
rect 16792 3390 16841 3402
rect 16792 3370 16810 3390
rect 16830 3370 16841 3390
rect 16792 3360 16841 3370
rect 16916 3386 16960 3402
rect 16916 3366 16925 3386
rect 16945 3366 16960 3386
rect 16916 3360 16960 3366
rect 17010 3390 17059 3402
rect 17010 3370 17028 3390
rect 17048 3370 17059 3390
rect 17010 3360 17059 3370
rect 22958 3521 23007 3533
rect 23057 3557 23101 3563
rect 23057 3537 23072 3557
rect 23092 3537 23101 3557
rect 23057 3521 23101 3537
rect 23176 3553 23225 3563
rect 23176 3533 23187 3553
rect 23207 3533 23225 3553
rect 23176 3521 23225 3533
rect 23275 3557 23319 3563
rect 23275 3537 23290 3557
rect 23310 3537 23319 3557
rect 23275 3521 23319 3537
rect 23389 3557 23433 3563
rect 23389 3537 23398 3557
rect 23418 3537 23433 3557
rect 23389 3521 23433 3537
rect 23483 3553 23532 3563
rect 23483 3533 23501 3553
rect 23521 3533 23532 3553
rect 23483 3521 23532 3533
rect 24317 3561 24366 3573
rect 24317 3541 24328 3561
rect 24348 3541 24366 3561
rect 24317 3531 24366 3541
rect 24416 3557 24460 3573
rect 24416 3537 24431 3557
rect 24451 3537 24460 3557
rect 24416 3531 24460 3537
rect 24530 3557 24574 3573
rect 24530 3537 24539 3557
rect 24559 3537 24574 3557
rect 24530 3531 24574 3537
rect 24624 3561 24673 3573
rect 24624 3541 24642 3561
rect 24662 3541 24673 3561
rect 24624 3531 24673 3541
rect 24748 3557 24792 3573
rect 24748 3537 24757 3557
rect 24777 3537 24792 3557
rect 24748 3531 24792 3537
rect 24842 3561 24891 3573
rect 24842 3541 24860 3561
rect 24880 3541 24891 3561
rect 24842 3531 24891 3541
rect 27335 3565 27384 3575
rect 27335 3545 27346 3565
rect 27366 3545 27384 3565
rect 13956 3320 13974 3340
rect 13994 3320 14005 3340
rect 13956 3308 14005 3320
rect 6781 3141 6830 3153
rect 2942 3108 2960 3128
rect 2980 3108 2991 3128
rect 2942 3098 2991 3108
rect 1649 3086 1698 3098
rect 5488 3131 5537 3141
rect 5488 3111 5499 3131
rect 5519 3111 5537 3131
rect 5488 3099 5537 3111
rect 5587 3135 5631 3141
rect 5587 3115 5602 3135
rect 5622 3115 5631 3135
rect 5587 3099 5631 3115
rect 5706 3131 5755 3141
rect 5706 3111 5717 3131
rect 5737 3111 5755 3131
rect 5706 3099 5755 3111
rect 5805 3135 5849 3141
rect 5805 3115 5820 3135
rect 5840 3115 5849 3135
rect 5805 3099 5849 3115
rect 5919 3135 5963 3141
rect 5919 3115 5928 3135
rect 5948 3115 5963 3135
rect 5919 3099 5963 3115
rect 6013 3131 6062 3141
rect 6013 3111 6031 3131
rect 6051 3111 6062 3131
rect 6781 3121 6792 3141
rect 6812 3121 6830 3141
rect 6781 3111 6830 3121
rect 6880 3137 6924 3153
rect 6880 3117 6895 3137
rect 6915 3117 6924 3137
rect 6880 3111 6924 3117
rect 6994 3137 7038 3153
rect 6994 3117 7003 3137
rect 7023 3117 7038 3137
rect 6994 3111 7038 3117
rect 7088 3141 7137 3153
rect 7088 3121 7106 3141
rect 7126 3121 7137 3141
rect 7088 3111 7137 3121
rect 7212 3137 7256 3153
rect 7212 3117 7221 3137
rect 7241 3117 7256 3137
rect 7212 3111 7256 3117
rect 7306 3141 7355 3153
rect 27335 3533 27384 3545
rect 27434 3569 27478 3575
rect 27434 3549 27449 3569
rect 27469 3549 27478 3569
rect 27434 3533 27478 3549
rect 27553 3565 27602 3575
rect 27553 3545 27564 3565
rect 27584 3545 27602 3565
rect 27553 3533 27602 3545
rect 27652 3569 27696 3575
rect 27652 3549 27667 3569
rect 27687 3549 27696 3569
rect 27652 3533 27696 3549
rect 27766 3569 27810 3575
rect 27766 3549 27775 3569
rect 27795 3549 27810 3569
rect 27766 3533 27810 3549
rect 27860 3565 27909 3575
rect 27860 3545 27878 3565
rect 27898 3545 27909 3565
rect 27860 3533 27909 3545
rect 28694 3573 28743 3585
rect 28694 3553 28705 3573
rect 28725 3553 28743 3573
rect 28694 3543 28743 3553
rect 28793 3569 28837 3585
rect 28793 3549 28808 3569
rect 28828 3549 28837 3569
rect 28793 3543 28837 3549
rect 28907 3569 28951 3585
rect 28907 3549 28916 3569
rect 28936 3549 28951 3569
rect 28907 3543 28951 3549
rect 29001 3573 29050 3585
rect 29001 3553 29019 3573
rect 29039 3553 29050 3573
rect 29001 3543 29050 3553
rect 29125 3569 29169 3585
rect 29125 3549 29134 3569
rect 29154 3549 29169 3569
rect 29125 3543 29169 3549
rect 29219 3573 29268 3585
rect 29219 3553 29237 3573
rect 29257 3553 29268 3573
rect 29219 3543 29268 3553
rect 31699 3578 31748 3588
rect 31699 3558 31710 3578
rect 31730 3558 31748 3578
rect 20751 3364 20800 3376
rect 20751 3344 20762 3364
rect 20782 3344 20800 3364
rect 11158 3153 11207 3165
rect 7306 3121 7324 3141
rect 7344 3121 7355 3141
rect 7306 3111 7355 3121
rect 6013 3099 6062 3111
rect 9865 3143 9914 3153
rect 9865 3123 9876 3143
rect 9896 3123 9914 3143
rect 9865 3111 9914 3123
rect 9964 3147 10008 3153
rect 9964 3127 9979 3147
rect 9999 3127 10008 3147
rect 9964 3111 10008 3127
rect 10083 3143 10132 3153
rect 10083 3123 10094 3143
rect 10114 3123 10132 3143
rect 10083 3111 10132 3123
rect 10182 3147 10226 3153
rect 10182 3127 10197 3147
rect 10217 3127 10226 3147
rect 10182 3111 10226 3127
rect 10296 3147 10340 3153
rect 10296 3127 10305 3147
rect 10325 3127 10340 3147
rect 10296 3111 10340 3127
rect 10390 3143 10439 3153
rect 10390 3123 10408 3143
rect 10428 3123 10439 3143
rect 11158 3133 11169 3153
rect 11189 3133 11207 3153
rect 11158 3123 11207 3133
rect 11257 3149 11301 3165
rect 11257 3129 11272 3149
rect 11292 3129 11301 3149
rect 11257 3123 11301 3129
rect 11371 3149 11415 3165
rect 11371 3129 11380 3149
rect 11400 3129 11415 3149
rect 11371 3123 11415 3129
rect 11465 3153 11514 3165
rect 11465 3133 11483 3153
rect 11503 3133 11514 3153
rect 11465 3123 11514 3133
rect 11589 3149 11633 3165
rect 11589 3129 11598 3149
rect 11618 3129 11633 3149
rect 11589 3123 11633 3129
rect 11683 3153 11732 3165
rect 17697 3314 17746 3324
rect 17697 3294 17708 3314
rect 17728 3294 17746 3314
rect 17697 3282 17746 3294
rect 17796 3318 17840 3324
rect 17796 3298 17811 3318
rect 17831 3298 17840 3318
rect 17796 3282 17840 3298
rect 17915 3314 17964 3324
rect 17915 3294 17926 3314
rect 17946 3294 17964 3314
rect 17915 3282 17964 3294
rect 18014 3318 18058 3324
rect 18014 3298 18029 3318
rect 18049 3298 18058 3318
rect 18014 3282 18058 3298
rect 18128 3318 18172 3324
rect 18128 3298 18137 3318
rect 18157 3298 18172 3318
rect 18128 3282 18172 3298
rect 18222 3314 18271 3324
rect 20751 3334 20800 3344
rect 20850 3360 20894 3376
rect 20850 3340 20865 3360
rect 20885 3340 20894 3360
rect 20850 3334 20894 3340
rect 20964 3360 21008 3376
rect 20964 3340 20973 3360
rect 20993 3340 21008 3360
rect 20964 3334 21008 3340
rect 21058 3364 21107 3376
rect 21058 3344 21076 3364
rect 21096 3344 21107 3364
rect 21058 3334 21107 3344
rect 21182 3360 21226 3376
rect 21182 3340 21191 3360
rect 21211 3340 21226 3360
rect 21182 3334 21226 3340
rect 21276 3364 21325 3376
rect 21276 3344 21294 3364
rect 21314 3344 21325 3364
rect 21276 3334 21325 3344
rect 18222 3294 18240 3314
rect 18260 3294 18271 3314
rect 18222 3282 18271 3294
rect 31699 3546 31748 3558
rect 31798 3582 31842 3588
rect 31798 3562 31813 3582
rect 31833 3562 31842 3582
rect 31798 3546 31842 3562
rect 31917 3578 31966 3588
rect 31917 3558 31928 3578
rect 31948 3558 31966 3578
rect 31917 3546 31966 3558
rect 32016 3582 32060 3588
rect 32016 3562 32031 3582
rect 32051 3562 32060 3582
rect 32016 3546 32060 3562
rect 32130 3582 32174 3588
rect 32130 3562 32139 3582
rect 32159 3562 32174 3582
rect 32130 3546 32174 3562
rect 32224 3578 32273 3588
rect 32224 3558 32242 3578
rect 32262 3558 32273 3578
rect 32224 3546 32273 3558
rect 33058 3586 33107 3598
rect 33058 3566 33069 3586
rect 33089 3566 33107 3586
rect 33058 3556 33107 3566
rect 33157 3582 33201 3598
rect 33157 3562 33172 3582
rect 33192 3562 33201 3582
rect 33157 3556 33201 3562
rect 33271 3582 33315 3598
rect 33271 3562 33280 3582
rect 33300 3562 33315 3582
rect 33271 3556 33315 3562
rect 33365 3586 33414 3598
rect 33365 3566 33383 3586
rect 33403 3566 33414 3586
rect 33365 3556 33414 3566
rect 33489 3582 33533 3598
rect 33489 3562 33498 3582
rect 33518 3562 33533 3582
rect 33489 3556 33533 3562
rect 33583 3586 33632 3598
rect 33583 3566 33601 3586
rect 33621 3566 33632 3586
rect 33583 3556 33632 3566
rect 25115 3377 25164 3389
rect 25115 3357 25126 3377
rect 25146 3357 25164 3377
rect 22061 3327 22110 3337
rect 22061 3307 22072 3327
rect 22092 3307 22110 3327
rect 22061 3295 22110 3307
rect 22160 3331 22204 3337
rect 22160 3311 22175 3331
rect 22195 3311 22204 3331
rect 22160 3295 22204 3311
rect 22279 3327 22328 3337
rect 22279 3307 22290 3327
rect 22310 3307 22328 3327
rect 22279 3295 22328 3307
rect 22378 3331 22422 3337
rect 22378 3311 22393 3331
rect 22413 3311 22422 3331
rect 22378 3295 22422 3311
rect 22492 3331 22536 3337
rect 22492 3311 22501 3331
rect 22521 3311 22536 3331
rect 22492 3295 22536 3311
rect 22586 3327 22635 3337
rect 25115 3347 25164 3357
rect 25214 3373 25258 3389
rect 25214 3353 25229 3373
rect 25249 3353 25258 3373
rect 25214 3347 25258 3353
rect 25328 3373 25372 3389
rect 25328 3353 25337 3373
rect 25357 3353 25372 3373
rect 25328 3347 25372 3353
rect 25422 3377 25471 3389
rect 25422 3357 25440 3377
rect 25460 3357 25471 3377
rect 25422 3347 25471 3357
rect 25546 3373 25590 3389
rect 25546 3353 25555 3373
rect 25575 3353 25590 3373
rect 25546 3347 25590 3353
rect 25640 3377 25689 3389
rect 25640 3357 25658 3377
rect 25678 3357 25689 3377
rect 25640 3347 25689 3357
rect 22586 3307 22604 3327
rect 22624 3307 22635 3327
rect 22586 3295 22635 3307
rect 15522 3166 15571 3178
rect 11683 3133 11701 3153
rect 11721 3133 11732 3153
rect 11683 3123 11732 3133
rect 10390 3111 10439 3123
rect 327 2890 376 2900
rect 327 2870 338 2890
rect 358 2870 376 2890
rect 327 2858 376 2870
rect 426 2894 470 2900
rect 426 2874 441 2894
rect 461 2874 470 2894
rect 426 2858 470 2874
rect 545 2890 594 2900
rect 545 2870 556 2890
rect 576 2870 594 2890
rect 545 2858 594 2870
rect 644 2894 688 2900
rect 644 2874 659 2894
rect 679 2874 688 2894
rect 644 2858 688 2874
rect 758 2894 802 2900
rect 758 2874 767 2894
rect 787 2874 802 2894
rect 758 2858 802 2874
rect 852 2890 901 2900
rect 852 2870 870 2890
rect 890 2870 901 2890
rect 14229 3156 14278 3166
rect 14229 3136 14240 3156
rect 14260 3136 14278 3156
rect 14229 3124 14278 3136
rect 14328 3160 14372 3166
rect 14328 3140 14343 3160
rect 14363 3140 14372 3160
rect 14328 3124 14372 3140
rect 14447 3156 14496 3166
rect 14447 3136 14458 3156
rect 14478 3136 14496 3156
rect 14447 3124 14496 3136
rect 14546 3160 14590 3166
rect 14546 3140 14561 3160
rect 14581 3140 14590 3160
rect 14546 3124 14590 3140
rect 14660 3160 14704 3166
rect 14660 3140 14669 3160
rect 14689 3140 14704 3160
rect 14660 3124 14704 3140
rect 14754 3156 14803 3166
rect 14754 3136 14772 3156
rect 14792 3136 14803 3156
rect 15522 3146 15533 3166
rect 15553 3146 15571 3166
rect 15522 3136 15571 3146
rect 15621 3162 15665 3178
rect 15621 3142 15636 3162
rect 15656 3142 15665 3162
rect 15621 3136 15665 3142
rect 15735 3162 15779 3178
rect 15735 3142 15744 3162
rect 15764 3142 15779 3162
rect 15735 3136 15779 3142
rect 15829 3166 15878 3178
rect 15829 3146 15847 3166
rect 15867 3146 15878 3166
rect 15829 3136 15878 3146
rect 15953 3162 15997 3178
rect 15953 3142 15962 3162
rect 15982 3142 15997 3162
rect 15953 3136 15997 3142
rect 16047 3166 16096 3178
rect 16047 3146 16065 3166
rect 16085 3146 16096 3166
rect 16047 3136 16096 3146
rect 29492 3389 29541 3401
rect 29492 3369 29503 3389
rect 29523 3369 29541 3389
rect 26438 3339 26487 3349
rect 26438 3319 26449 3339
rect 26469 3319 26487 3339
rect 26438 3307 26487 3319
rect 26537 3343 26581 3349
rect 26537 3323 26552 3343
rect 26572 3323 26581 3343
rect 26537 3307 26581 3323
rect 26656 3339 26705 3349
rect 26656 3319 26667 3339
rect 26687 3319 26705 3339
rect 26656 3307 26705 3319
rect 26755 3343 26799 3349
rect 26755 3323 26770 3343
rect 26790 3323 26799 3343
rect 26755 3307 26799 3323
rect 26869 3343 26913 3349
rect 26869 3323 26878 3343
rect 26898 3323 26913 3343
rect 26869 3307 26913 3323
rect 26963 3339 27012 3349
rect 29492 3359 29541 3369
rect 29591 3385 29635 3401
rect 29591 3365 29606 3385
rect 29626 3365 29635 3385
rect 29591 3359 29635 3365
rect 29705 3385 29749 3401
rect 29705 3365 29714 3385
rect 29734 3365 29749 3385
rect 29705 3359 29749 3365
rect 29799 3389 29848 3401
rect 29799 3369 29817 3389
rect 29837 3369 29848 3389
rect 29799 3359 29848 3369
rect 29923 3385 29967 3401
rect 29923 3365 29932 3385
rect 29952 3365 29967 3385
rect 29923 3359 29967 3365
rect 30017 3389 30066 3401
rect 30017 3369 30035 3389
rect 30055 3369 30066 3389
rect 30017 3359 30066 3369
rect 26963 3319 26981 3339
rect 27001 3319 27012 3339
rect 26963 3307 27012 3319
rect 19788 3140 19837 3152
rect 14754 3124 14803 3136
rect 852 2858 901 2870
rect 4691 2903 4740 2913
rect 4691 2883 4702 2903
rect 4722 2883 4740 2903
rect 4691 2871 4740 2883
rect 4790 2907 4834 2913
rect 4790 2887 4805 2907
rect 4825 2887 4834 2907
rect 4790 2871 4834 2887
rect 4909 2903 4958 2913
rect 4909 2883 4920 2903
rect 4940 2883 4958 2903
rect 4909 2871 4958 2883
rect 5008 2907 5052 2913
rect 5008 2887 5023 2907
rect 5043 2887 5052 2907
rect 5008 2871 5052 2887
rect 5122 2907 5166 2913
rect 5122 2887 5131 2907
rect 5151 2887 5166 2907
rect 5122 2871 5166 2887
rect 5216 2903 5265 2913
rect 5216 2883 5234 2903
rect 5254 2883 5265 2903
rect 18495 3130 18544 3140
rect 18495 3110 18506 3130
rect 18526 3110 18544 3130
rect 18495 3098 18544 3110
rect 18594 3134 18638 3140
rect 18594 3114 18609 3134
rect 18629 3114 18638 3134
rect 18594 3098 18638 3114
rect 18713 3130 18762 3140
rect 18713 3110 18724 3130
rect 18744 3110 18762 3130
rect 18713 3098 18762 3110
rect 18812 3134 18856 3140
rect 18812 3114 18827 3134
rect 18847 3114 18856 3134
rect 18812 3098 18856 3114
rect 18926 3134 18970 3140
rect 18926 3114 18935 3134
rect 18955 3114 18970 3134
rect 18926 3098 18970 3114
rect 19020 3130 19069 3140
rect 19020 3110 19038 3130
rect 19058 3110 19069 3130
rect 19788 3120 19799 3140
rect 19819 3120 19837 3140
rect 19788 3110 19837 3120
rect 19887 3136 19931 3152
rect 19887 3116 19902 3136
rect 19922 3116 19931 3136
rect 19887 3110 19931 3116
rect 20001 3136 20045 3152
rect 20001 3116 20010 3136
rect 20030 3116 20045 3136
rect 20001 3110 20045 3116
rect 20095 3140 20144 3152
rect 20095 3120 20113 3140
rect 20133 3120 20144 3140
rect 20095 3110 20144 3120
rect 20219 3136 20263 3152
rect 20219 3116 20228 3136
rect 20248 3116 20263 3136
rect 20219 3110 20263 3116
rect 20313 3140 20362 3152
rect 33856 3402 33905 3414
rect 33856 3382 33867 3402
rect 33887 3382 33905 3402
rect 30802 3352 30851 3362
rect 30802 3332 30813 3352
rect 30833 3332 30851 3352
rect 30802 3320 30851 3332
rect 30901 3356 30945 3362
rect 30901 3336 30916 3356
rect 30936 3336 30945 3356
rect 30901 3320 30945 3336
rect 31020 3352 31069 3362
rect 31020 3332 31031 3352
rect 31051 3332 31069 3352
rect 31020 3320 31069 3332
rect 31119 3356 31163 3362
rect 31119 3336 31134 3356
rect 31154 3336 31163 3356
rect 31119 3320 31163 3336
rect 31233 3356 31277 3362
rect 31233 3336 31242 3356
rect 31262 3336 31277 3356
rect 31233 3320 31277 3336
rect 31327 3352 31376 3362
rect 33856 3372 33905 3382
rect 33955 3398 33999 3414
rect 33955 3378 33970 3398
rect 33990 3378 33999 3398
rect 33955 3372 33999 3378
rect 34069 3398 34113 3414
rect 34069 3378 34078 3398
rect 34098 3378 34113 3398
rect 34069 3372 34113 3378
rect 34163 3402 34212 3414
rect 34163 3382 34181 3402
rect 34201 3382 34212 3402
rect 34163 3372 34212 3382
rect 34287 3398 34331 3414
rect 34287 3378 34296 3398
rect 34316 3378 34331 3398
rect 34287 3372 34331 3378
rect 34381 3402 34430 3414
rect 34381 3382 34399 3402
rect 34419 3382 34430 3402
rect 34381 3372 34430 3382
rect 31327 3332 31345 3352
rect 31365 3332 31376 3352
rect 31327 3320 31376 3332
rect 24152 3153 24201 3165
rect 20313 3120 20331 3140
rect 20351 3120 20362 3140
rect 20313 3110 20362 3120
rect 19020 3098 19069 3110
rect 5216 2871 5265 2883
rect 9068 2915 9117 2925
rect 9068 2895 9079 2915
rect 9099 2895 9117 2915
rect 9068 2883 9117 2895
rect 9167 2919 9211 2925
rect 9167 2899 9182 2919
rect 9202 2899 9211 2919
rect 9167 2883 9211 2899
rect 9286 2915 9335 2925
rect 9286 2895 9297 2915
rect 9317 2895 9335 2915
rect 9286 2883 9335 2895
rect 9385 2919 9429 2925
rect 9385 2899 9400 2919
rect 9420 2899 9429 2919
rect 9385 2883 9429 2899
rect 9499 2919 9543 2925
rect 9499 2899 9508 2919
rect 9528 2899 9543 2919
rect 9499 2883 9543 2899
rect 9593 2915 9642 2925
rect 9593 2895 9611 2915
rect 9631 2895 9642 2915
rect 22859 3143 22908 3153
rect 22859 3123 22870 3143
rect 22890 3123 22908 3143
rect 22859 3111 22908 3123
rect 22958 3147 23002 3153
rect 22958 3127 22973 3147
rect 22993 3127 23002 3147
rect 22958 3111 23002 3127
rect 23077 3143 23126 3153
rect 23077 3123 23088 3143
rect 23108 3123 23126 3143
rect 23077 3111 23126 3123
rect 23176 3147 23220 3153
rect 23176 3127 23191 3147
rect 23211 3127 23220 3147
rect 23176 3111 23220 3127
rect 23290 3147 23334 3153
rect 23290 3127 23299 3147
rect 23319 3127 23334 3147
rect 23290 3111 23334 3127
rect 23384 3143 23433 3153
rect 23384 3123 23402 3143
rect 23422 3123 23433 3143
rect 24152 3133 24163 3153
rect 24183 3133 24201 3153
rect 24152 3123 24201 3133
rect 24251 3149 24295 3165
rect 24251 3129 24266 3149
rect 24286 3129 24295 3149
rect 24251 3123 24295 3129
rect 24365 3149 24409 3165
rect 24365 3129 24374 3149
rect 24394 3129 24409 3149
rect 24365 3123 24409 3129
rect 24459 3153 24508 3165
rect 24459 3133 24477 3153
rect 24497 3133 24508 3153
rect 24459 3123 24508 3133
rect 24583 3149 24627 3165
rect 24583 3129 24592 3149
rect 24612 3129 24627 3149
rect 24583 3123 24627 3129
rect 24677 3153 24726 3165
rect 28529 3165 28578 3177
rect 24677 3133 24695 3153
rect 24715 3133 24726 3153
rect 24677 3123 24726 3133
rect 23384 3111 23433 3123
rect 9593 2883 9642 2895
rect 13432 2928 13481 2938
rect 13432 2908 13443 2928
rect 13463 2908 13481 2928
rect 13432 2896 13481 2908
rect 13531 2932 13575 2938
rect 13531 2912 13546 2932
rect 13566 2912 13575 2932
rect 13531 2896 13575 2912
rect 13650 2928 13699 2938
rect 13650 2908 13661 2928
rect 13681 2908 13699 2928
rect 13650 2896 13699 2908
rect 13749 2932 13793 2938
rect 13749 2912 13764 2932
rect 13784 2912 13793 2932
rect 13749 2896 13793 2912
rect 13863 2932 13907 2938
rect 13863 2912 13872 2932
rect 13892 2912 13907 2932
rect 13863 2896 13907 2912
rect 13957 2928 14006 2938
rect 13957 2908 13975 2928
rect 13995 2908 14006 2928
rect 13957 2896 14006 2908
rect 27236 3155 27285 3165
rect 27236 3135 27247 3155
rect 27267 3135 27285 3155
rect 27236 3123 27285 3135
rect 27335 3159 27379 3165
rect 27335 3139 27350 3159
rect 27370 3139 27379 3159
rect 27335 3123 27379 3139
rect 27454 3155 27503 3165
rect 27454 3135 27465 3155
rect 27485 3135 27503 3155
rect 27454 3123 27503 3135
rect 27553 3159 27597 3165
rect 27553 3139 27568 3159
rect 27588 3139 27597 3159
rect 27553 3123 27597 3139
rect 27667 3159 27711 3165
rect 27667 3139 27676 3159
rect 27696 3139 27711 3159
rect 27667 3123 27711 3139
rect 27761 3155 27810 3165
rect 27761 3135 27779 3155
rect 27799 3135 27810 3155
rect 28529 3145 28540 3165
rect 28560 3145 28578 3165
rect 28529 3135 28578 3145
rect 28628 3161 28672 3177
rect 28628 3141 28643 3161
rect 28663 3141 28672 3161
rect 28628 3135 28672 3141
rect 28742 3161 28786 3177
rect 28742 3141 28751 3161
rect 28771 3141 28786 3161
rect 28742 3135 28786 3141
rect 28836 3165 28885 3177
rect 28836 3145 28854 3165
rect 28874 3145 28885 3165
rect 28836 3135 28885 3145
rect 28960 3161 29004 3177
rect 28960 3141 28969 3161
rect 28989 3141 29004 3161
rect 28960 3135 29004 3141
rect 29054 3165 29103 3177
rect 32893 3178 32942 3190
rect 29054 3145 29072 3165
rect 29092 3145 29103 3165
rect 29054 3135 29103 3145
rect 27761 3123 27810 3135
rect 17698 2902 17747 2912
rect 17698 2882 17709 2902
rect 17729 2882 17747 2902
rect 17698 2870 17747 2882
rect 17797 2906 17841 2912
rect 17797 2886 17812 2906
rect 17832 2886 17841 2906
rect 17797 2870 17841 2886
rect 17916 2902 17965 2912
rect 17916 2882 17927 2902
rect 17947 2882 17965 2902
rect 17916 2870 17965 2882
rect 18015 2906 18059 2912
rect 18015 2886 18030 2906
rect 18050 2886 18059 2906
rect 18015 2870 18059 2886
rect 18129 2906 18173 2912
rect 18129 2886 18138 2906
rect 18158 2886 18173 2906
rect 18129 2870 18173 2886
rect 18223 2902 18272 2912
rect 18223 2882 18241 2902
rect 18261 2882 18272 2902
rect 31600 3168 31649 3178
rect 31600 3148 31611 3168
rect 31631 3148 31649 3168
rect 31600 3136 31649 3148
rect 31699 3172 31743 3178
rect 31699 3152 31714 3172
rect 31734 3152 31743 3172
rect 31699 3136 31743 3152
rect 31818 3168 31867 3178
rect 31818 3148 31829 3168
rect 31849 3148 31867 3168
rect 31818 3136 31867 3148
rect 31917 3172 31961 3178
rect 31917 3152 31932 3172
rect 31952 3152 31961 3172
rect 31917 3136 31961 3152
rect 32031 3172 32075 3178
rect 32031 3152 32040 3172
rect 32060 3152 32075 3172
rect 32031 3136 32075 3152
rect 32125 3168 32174 3178
rect 32125 3148 32143 3168
rect 32163 3148 32174 3168
rect 32893 3158 32904 3178
rect 32924 3158 32942 3178
rect 32893 3148 32942 3158
rect 32992 3174 33036 3190
rect 32992 3154 33007 3174
rect 33027 3154 33036 3174
rect 32992 3148 33036 3154
rect 33106 3174 33150 3190
rect 33106 3154 33115 3174
rect 33135 3154 33150 3174
rect 33106 3148 33150 3154
rect 33200 3178 33249 3190
rect 33200 3158 33218 3178
rect 33238 3158 33249 3178
rect 33200 3148 33249 3158
rect 33324 3174 33368 3190
rect 33324 3154 33333 3174
rect 33353 3154 33368 3174
rect 33324 3148 33368 3154
rect 33418 3178 33467 3190
rect 33418 3158 33436 3178
rect 33456 3158 33467 3178
rect 33418 3148 33467 3158
rect 32125 3136 32174 3148
rect 18223 2870 18272 2882
rect 22062 2915 22111 2925
rect 22062 2895 22073 2915
rect 22093 2895 22111 2915
rect 22062 2883 22111 2895
rect 22161 2919 22205 2925
rect 22161 2899 22176 2919
rect 22196 2899 22205 2919
rect 22161 2883 22205 2899
rect 22280 2915 22329 2925
rect 22280 2895 22291 2915
rect 22311 2895 22329 2915
rect 22280 2883 22329 2895
rect 22379 2919 22423 2925
rect 22379 2899 22394 2919
rect 22414 2899 22423 2919
rect 22379 2883 22423 2899
rect 22493 2919 22537 2925
rect 22493 2899 22502 2919
rect 22522 2899 22537 2919
rect 22493 2883 22537 2899
rect 22587 2915 22636 2925
rect 22587 2895 22605 2915
rect 22625 2895 22636 2915
rect 22587 2883 22636 2895
rect 26439 2927 26488 2937
rect 26439 2907 26450 2927
rect 26470 2907 26488 2927
rect 26439 2895 26488 2907
rect 26538 2931 26582 2937
rect 26538 2911 26553 2931
rect 26573 2911 26582 2931
rect 26538 2895 26582 2911
rect 26657 2927 26706 2937
rect 26657 2907 26668 2927
rect 26688 2907 26706 2927
rect 26657 2895 26706 2907
rect 26756 2931 26800 2937
rect 26756 2911 26771 2931
rect 26791 2911 26800 2931
rect 26756 2895 26800 2911
rect 26870 2931 26914 2937
rect 26870 2911 26879 2931
rect 26899 2911 26914 2931
rect 26870 2895 26914 2911
rect 26964 2927 27013 2937
rect 26964 2907 26982 2927
rect 27002 2907 27013 2927
rect 26964 2895 27013 2907
rect 30803 2940 30852 2950
rect 30803 2920 30814 2940
rect 30834 2920 30852 2940
rect 30803 2908 30852 2920
rect 30902 2944 30946 2950
rect 30902 2924 30917 2944
rect 30937 2924 30946 2944
rect 30902 2908 30946 2924
rect 31021 2940 31070 2950
rect 31021 2920 31032 2940
rect 31052 2920 31070 2940
rect 31021 2908 31070 2920
rect 31120 2944 31164 2950
rect 31120 2924 31135 2944
rect 31155 2924 31164 2944
rect 31120 2908 31164 2924
rect 31234 2944 31278 2950
rect 31234 2924 31243 2944
rect 31263 2924 31278 2944
rect 31234 2908 31278 2924
rect 31328 2940 31377 2950
rect 31328 2920 31346 2940
rect 31366 2920 31377 2940
rect 31328 2908 31377 2920
rect 3359 2746 3408 2758
rect 3359 2726 3370 2746
rect 3390 2726 3408 2746
rect 3359 2716 3408 2726
rect 3458 2742 3502 2758
rect 3458 2722 3473 2742
rect 3493 2722 3502 2742
rect 3458 2716 3502 2722
rect 3572 2742 3616 2758
rect 3572 2722 3581 2742
rect 3601 2722 3616 2742
rect 3572 2716 3616 2722
rect 3666 2746 3715 2758
rect 3666 2726 3684 2746
rect 3704 2726 3715 2746
rect 3666 2716 3715 2726
rect 3790 2742 3834 2758
rect 3790 2722 3799 2742
rect 3819 2722 3834 2742
rect 3790 2716 3834 2722
rect 3884 2746 3933 2758
rect 3884 2726 3902 2746
rect 3922 2726 3933 2746
rect 3884 2716 3933 2726
rect 7723 2759 7772 2771
rect 7723 2739 7734 2759
rect 7754 2739 7772 2759
rect 7723 2729 7772 2739
rect 7822 2755 7866 2771
rect 7822 2735 7837 2755
rect 7857 2735 7866 2755
rect 7822 2729 7866 2735
rect 7936 2755 7980 2771
rect 7936 2735 7945 2755
rect 7965 2735 7980 2755
rect 7936 2729 7980 2735
rect 8030 2759 8079 2771
rect 8030 2739 8048 2759
rect 8068 2739 8079 2759
rect 8030 2729 8079 2739
rect 8154 2755 8198 2771
rect 8154 2735 8163 2755
rect 8183 2735 8198 2755
rect 8154 2729 8198 2735
rect 8248 2759 8297 2771
rect 8248 2739 8266 2759
rect 8286 2739 8297 2759
rect 8248 2729 8297 2739
rect 12100 2771 12149 2783
rect 12100 2751 12111 2771
rect 12131 2751 12149 2771
rect 12100 2741 12149 2751
rect 12199 2767 12243 2783
rect 12199 2747 12214 2767
rect 12234 2747 12243 2767
rect 12199 2741 12243 2747
rect 12313 2767 12357 2783
rect 12313 2747 12322 2767
rect 12342 2747 12357 2767
rect 12313 2741 12357 2747
rect 12407 2771 12456 2783
rect 12407 2751 12425 2771
rect 12445 2751 12456 2771
rect 12407 2741 12456 2751
rect 12531 2767 12575 2783
rect 12531 2747 12540 2767
rect 12560 2747 12575 2767
rect 12531 2741 12575 2747
rect 12625 2771 12674 2783
rect 12625 2751 12643 2771
rect 12663 2751 12674 2771
rect 12625 2741 12674 2751
rect 16464 2784 16513 2796
rect 2562 2518 2611 2530
rect 1269 2508 1318 2518
rect 1269 2488 1280 2508
rect 1300 2488 1318 2508
rect 1269 2476 1318 2488
rect 1368 2512 1412 2518
rect 1368 2492 1383 2512
rect 1403 2492 1412 2512
rect 1368 2476 1412 2492
rect 1487 2508 1536 2518
rect 1487 2488 1498 2508
rect 1518 2488 1536 2508
rect 1487 2476 1536 2488
rect 1586 2512 1630 2518
rect 1586 2492 1601 2512
rect 1621 2492 1630 2512
rect 1586 2476 1630 2492
rect 1700 2512 1744 2518
rect 1700 2492 1709 2512
rect 1729 2492 1744 2512
rect 1700 2476 1744 2492
rect 1794 2508 1843 2518
rect 1794 2488 1812 2508
rect 1832 2488 1843 2508
rect 2562 2498 2573 2518
rect 2593 2498 2611 2518
rect 2562 2488 2611 2498
rect 2661 2514 2705 2530
rect 2661 2494 2676 2514
rect 2696 2494 2705 2514
rect 2661 2488 2705 2494
rect 2775 2514 2819 2530
rect 2775 2494 2784 2514
rect 2804 2494 2819 2514
rect 2775 2488 2819 2494
rect 2869 2518 2918 2530
rect 2869 2498 2887 2518
rect 2907 2498 2918 2518
rect 2869 2488 2918 2498
rect 2993 2514 3037 2530
rect 2993 2494 3002 2514
rect 3022 2494 3037 2514
rect 2993 2488 3037 2494
rect 3087 2518 3136 2530
rect 3087 2498 3105 2518
rect 3125 2498 3136 2518
rect 3087 2488 3136 2498
rect 16464 2764 16475 2784
rect 16495 2764 16513 2784
rect 16464 2754 16513 2764
rect 16563 2780 16607 2796
rect 16563 2760 16578 2780
rect 16598 2760 16607 2780
rect 16563 2754 16607 2760
rect 16677 2780 16721 2796
rect 16677 2760 16686 2780
rect 16706 2760 16721 2780
rect 16677 2754 16721 2760
rect 16771 2784 16820 2796
rect 16771 2764 16789 2784
rect 16809 2764 16820 2784
rect 16771 2754 16820 2764
rect 16895 2780 16939 2796
rect 16895 2760 16904 2780
rect 16924 2760 16939 2780
rect 16895 2754 16939 2760
rect 16989 2784 17038 2796
rect 16989 2764 17007 2784
rect 17027 2764 17038 2784
rect 16989 2754 17038 2764
rect 6926 2531 6975 2543
rect 5633 2521 5682 2531
rect 5633 2501 5644 2521
rect 5664 2501 5682 2521
rect 1794 2476 1843 2488
rect 5633 2489 5682 2501
rect 5732 2525 5776 2531
rect 5732 2505 5747 2525
rect 5767 2505 5776 2525
rect 5732 2489 5776 2505
rect 5851 2521 5900 2531
rect 5851 2501 5862 2521
rect 5882 2501 5900 2521
rect 5851 2489 5900 2501
rect 5950 2525 5994 2531
rect 5950 2505 5965 2525
rect 5985 2505 5994 2525
rect 5950 2489 5994 2505
rect 6064 2525 6108 2531
rect 6064 2505 6073 2525
rect 6093 2505 6108 2525
rect 6064 2489 6108 2505
rect 6158 2521 6207 2531
rect 6158 2501 6176 2521
rect 6196 2501 6207 2521
rect 6926 2511 6937 2531
rect 6957 2511 6975 2531
rect 6926 2501 6975 2511
rect 7025 2527 7069 2543
rect 7025 2507 7040 2527
rect 7060 2507 7069 2527
rect 7025 2501 7069 2507
rect 7139 2527 7183 2543
rect 7139 2507 7148 2527
rect 7168 2507 7183 2527
rect 7139 2501 7183 2507
rect 7233 2531 7282 2543
rect 7233 2511 7251 2531
rect 7271 2511 7282 2531
rect 7233 2501 7282 2511
rect 7357 2527 7401 2543
rect 7357 2507 7366 2527
rect 7386 2507 7401 2527
rect 7357 2501 7401 2507
rect 7451 2531 7500 2543
rect 7451 2511 7469 2531
rect 7489 2511 7500 2531
rect 7451 2501 7500 2511
rect 20730 2758 20779 2770
rect 20730 2738 20741 2758
rect 20761 2738 20779 2758
rect 20730 2728 20779 2738
rect 20829 2754 20873 2770
rect 20829 2734 20844 2754
rect 20864 2734 20873 2754
rect 20829 2728 20873 2734
rect 20943 2754 20987 2770
rect 20943 2734 20952 2754
rect 20972 2734 20987 2754
rect 20943 2728 20987 2734
rect 21037 2758 21086 2770
rect 21037 2738 21055 2758
rect 21075 2738 21086 2758
rect 21037 2728 21086 2738
rect 21161 2754 21205 2770
rect 21161 2734 21170 2754
rect 21190 2734 21205 2754
rect 21161 2728 21205 2734
rect 21255 2758 21304 2770
rect 21255 2738 21273 2758
rect 21293 2738 21304 2758
rect 21255 2728 21304 2738
rect 25094 2771 25143 2783
rect 11303 2543 11352 2555
rect 10010 2533 10059 2543
rect 10010 2513 10021 2533
rect 10041 2513 10059 2533
rect 6158 2489 6207 2501
rect 10010 2501 10059 2513
rect 10109 2537 10153 2543
rect 10109 2517 10124 2537
rect 10144 2517 10153 2537
rect 10109 2501 10153 2517
rect 10228 2533 10277 2543
rect 10228 2513 10239 2533
rect 10259 2513 10277 2533
rect 10228 2501 10277 2513
rect 10327 2537 10371 2543
rect 10327 2517 10342 2537
rect 10362 2517 10371 2537
rect 10327 2501 10371 2517
rect 10441 2537 10485 2543
rect 10441 2517 10450 2537
rect 10470 2517 10485 2537
rect 10441 2501 10485 2517
rect 10535 2533 10584 2543
rect 10535 2513 10553 2533
rect 10573 2513 10584 2533
rect 11303 2523 11314 2543
rect 11334 2523 11352 2543
rect 11303 2513 11352 2523
rect 11402 2539 11446 2555
rect 11402 2519 11417 2539
rect 11437 2519 11446 2539
rect 11402 2513 11446 2519
rect 11516 2539 11560 2555
rect 11516 2519 11525 2539
rect 11545 2519 11560 2539
rect 11516 2513 11560 2519
rect 11610 2543 11659 2555
rect 11610 2523 11628 2543
rect 11648 2523 11659 2543
rect 11610 2513 11659 2523
rect 11734 2539 11778 2555
rect 11734 2519 11743 2539
rect 11763 2519 11778 2539
rect 11734 2513 11778 2519
rect 11828 2543 11877 2555
rect 11828 2523 11846 2543
rect 11866 2523 11877 2543
rect 11828 2513 11877 2523
rect 25094 2751 25105 2771
rect 25125 2751 25143 2771
rect 25094 2741 25143 2751
rect 25193 2767 25237 2783
rect 25193 2747 25208 2767
rect 25228 2747 25237 2767
rect 25193 2741 25237 2747
rect 25307 2767 25351 2783
rect 25307 2747 25316 2767
rect 25336 2747 25351 2767
rect 25307 2741 25351 2747
rect 25401 2771 25450 2783
rect 25401 2751 25419 2771
rect 25439 2751 25450 2771
rect 25401 2741 25450 2751
rect 25525 2767 25569 2783
rect 25525 2747 25534 2767
rect 25554 2747 25569 2767
rect 25525 2741 25569 2747
rect 25619 2771 25668 2783
rect 25619 2751 25637 2771
rect 25657 2751 25668 2771
rect 25619 2741 25668 2751
rect 29471 2783 29520 2795
rect 15667 2556 15716 2568
rect 14374 2546 14423 2556
rect 14374 2526 14385 2546
rect 14405 2526 14423 2546
rect 10535 2501 10584 2513
rect 3360 2334 3409 2346
rect 3360 2314 3371 2334
rect 3391 2314 3409 2334
rect 306 2284 355 2294
rect 306 2264 317 2284
rect 337 2264 355 2284
rect 306 2252 355 2264
rect 405 2288 449 2294
rect 405 2268 420 2288
rect 440 2268 449 2288
rect 405 2252 449 2268
rect 524 2284 573 2294
rect 524 2264 535 2284
rect 555 2264 573 2284
rect 524 2252 573 2264
rect 623 2288 667 2294
rect 623 2268 638 2288
rect 658 2268 667 2288
rect 623 2252 667 2268
rect 737 2288 781 2294
rect 737 2268 746 2288
rect 766 2268 781 2288
rect 737 2252 781 2268
rect 831 2284 880 2294
rect 3360 2304 3409 2314
rect 3459 2330 3503 2346
rect 3459 2310 3474 2330
rect 3494 2310 3503 2330
rect 3459 2304 3503 2310
rect 3573 2330 3617 2346
rect 3573 2310 3582 2330
rect 3602 2310 3617 2330
rect 3573 2304 3617 2310
rect 3667 2334 3716 2346
rect 3667 2314 3685 2334
rect 3705 2314 3716 2334
rect 3667 2304 3716 2314
rect 3791 2330 3835 2346
rect 3791 2310 3800 2330
rect 3820 2310 3835 2330
rect 3791 2304 3835 2310
rect 3885 2334 3934 2346
rect 3885 2314 3903 2334
rect 3923 2314 3934 2334
rect 3885 2304 3934 2314
rect 831 2264 849 2284
rect 869 2264 880 2284
rect 831 2252 880 2264
rect 14374 2514 14423 2526
rect 14473 2550 14517 2556
rect 14473 2530 14488 2550
rect 14508 2530 14517 2550
rect 14473 2514 14517 2530
rect 14592 2546 14641 2556
rect 14592 2526 14603 2546
rect 14623 2526 14641 2546
rect 14592 2514 14641 2526
rect 14691 2550 14735 2556
rect 14691 2530 14706 2550
rect 14726 2530 14735 2550
rect 14691 2514 14735 2530
rect 14805 2550 14849 2556
rect 14805 2530 14814 2550
rect 14834 2530 14849 2550
rect 14805 2514 14849 2530
rect 14899 2546 14948 2556
rect 14899 2526 14917 2546
rect 14937 2526 14948 2546
rect 15667 2536 15678 2556
rect 15698 2536 15716 2556
rect 15667 2526 15716 2536
rect 15766 2552 15810 2568
rect 15766 2532 15781 2552
rect 15801 2532 15810 2552
rect 15766 2526 15810 2532
rect 15880 2552 15924 2568
rect 15880 2532 15889 2552
rect 15909 2532 15924 2552
rect 15880 2526 15924 2532
rect 15974 2556 16023 2568
rect 15974 2536 15992 2556
rect 16012 2536 16023 2556
rect 15974 2526 16023 2536
rect 16098 2552 16142 2568
rect 16098 2532 16107 2552
rect 16127 2532 16142 2552
rect 16098 2526 16142 2532
rect 16192 2556 16241 2568
rect 16192 2536 16210 2556
rect 16230 2536 16241 2556
rect 16192 2526 16241 2536
rect 29471 2763 29482 2783
rect 29502 2763 29520 2783
rect 29471 2753 29520 2763
rect 29570 2779 29614 2795
rect 29570 2759 29585 2779
rect 29605 2759 29614 2779
rect 29570 2753 29614 2759
rect 29684 2779 29728 2795
rect 29684 2759 29693 2779
rect 29713 2759 29728 2779
rect 29684 2753 29728 2759
rect 29778 2783 29827 2795
rect 29778 2763 29796 2783
rect 29816 2763 29827 2783
rect 29778 2753 29827 2763
rect 29902 2779 29946 2795
rect 29902 2759 29911 2779
rect 29931 2759 29946 2779
rect 29902 2753 29946 2759
rect 29996 2783 30045 2795
rect 29996 2763 30014 2783
rect 30034 2763 30045 2783
rect 29996 2753 30045 2763
rect 33835 2796 33884 2808
rect 19933 2530 19982 2542
rect 14899 2514 14948 2526
rect 7724 2347 7773 2359
rect 7724 2327 7735 2347
rect 7755 2327 7773 2347
rect 4670 2297 4719 2307
rect 4670 2277 4681 2297
rect 4701 2277 4719 2297
rect 4670 2265 4719 2277
rect 4769 2301 4813 2307
rect 4769 2281 4784 2301
rect 4804 2281 4813 2301
rect 4769 2265 4813 2281
rect 4888 2297 4937 2307
rect 4888 2277 4899 2297
rect 4919 2277 4937 2297
rect 4888 2265 4937 2277
rect 4987 2301 5031 2307
rect 4987 2281 5002 2301
rect 5022 2281 5031 2301
rect 4987 2265 5031 2281
rect 5101 2301 5145 2307
rect 5101 2281 5110 2301
rect 5130 2281 5145 2301
rect 5101 2265 5145 2281
rect 5195 2297 5244 2307
rect 7724 2317 7773 2327
rect 7823 2343 7867 2359
rect 7823 2323 7838 2343
rect 7858 2323 7867 2343
rect 7823 2317 7867 2323
rect 7937 2343 7981 2359
rect 7937 2323 7946 2343
rect 7966 2323 7981 2343
rect 7937 2317 7981 2323
rect 8031 2347 8080 2359
rect 8031 2327 8049 2347
rect 8069 2327 8080 2347
rect 8031 2317 8080 2327
rect 8155 2343 8199 2359
rect 8155 2323 8164 2343
rect 8184 2323 8199 2343
rect 8155 2317 8199 2323
rect 8249 2347 8298 2359
rect 8249 2327 8267 2347
rect 8287 2327 8298 2347
rect 8249 2317 8298 2327
rect 5195 2277 5213 2297
rect 5233 2277 5244 2297
rect 5195 2265 5244 2277
rect 18640 2520 18689 2530
rect 18640 2500 18651 2520
rect 18671 2500 18689 2520
rect 18640 2488 18689 2500
rect 18739 2524 18783 2530
rect 18739 2504 18754 2524
rect 18774 2504 18783 2524
rect 18739 2488 18783 2504
rect 18858 2520 18907 2530
rect 18858 2500 18869 2520
rect 18889 2500 18907 2520
rect 18858 2488 18907 2500
rect 18957 2524 19001 2530
rect 18957 2504 18972 2524
rect 18992 2504 19001 2524
rect 18957 2488 19001 2504
rect 19071 2524 19115 2530
rect 19071 2504 19080 2524
rect 19100 2504 19115 2524
rect 19071 2488 19115 2504
rect 19165 2520 19214 2530
rect 19165 2500 19183 2520
rect 19203 2500 19214 2520
rect 19933 2510 19944 2530
rect 19964 2510 19982 2530
rect 19933 2500 19982 2510
rect 20032 2526 20076 2542
rect 20032 2506 20047 2526
rect 20067 2506 20076 2526
rect 20032 2500 20076 2506
rect 20146 2526 20190 2542
rect 20146 2506 20155 2526
rect 20175 2506 20190 2526
rect 20146 2500 20190 2506
rect 20240 2530 20289 2542
rect 20240 2510 20258 2530
rect 20278 2510 20289 2530
rect 20240 2500 20289 2510
rect 20364 2526 20408 2542
rect 20364 2506 20373 2526
rect 20393 2506 20408 2526
rect 20364 2500 20408 2506
rect 20458 2530 20507 2542
rect 20458 2510 20476 2530
rect 20496 2510 20507 2530
rect 20458 2500 20507 2510
rect 33835 2776 33846 2796
rect 33866 2776 33884 2796
rect 33835 2766 33884 2776
rect 33934 2792 33978 2808
rect 33934 2772 33949 2792
rect 33969 2772 33978 2792
rect 33934 2766 33978 2772
rect 34048 2792 34092 2808
rect 34048 2772 34057 2792
rect 34077 2772 34092 2792
rect 34048 2766 34092 2772
rect 34142 2796 34191 2808
rect 34142 2776 34160 2796
rect 34180 2776 34191 2796
rect 34142 2766 34191 2776
rect 34266 2792 34310 2808
rect 34266 2772 34275 2792
rect 34295 2772 34310 2792
rect 34266 2766 34310 2772
rect 34360 2796 34409 2808
rect 34360 2776 34378 2796
rect 34398 2776 34409 2796
rect 34360 2766 34409 2776
rect 24297 2543 24346 2555
rect 23004 2533 23053 2543
rect 23004 2513 23015 2533
rect 23035 2513 23053 2533
rect 19165 2488 19214 2500
rect 12101 2359 12150 2371
rect 12101 2339 12112 2359
rect 12132 2339 12150 2359
rect 9047 2309 9096 2319
rect 9047 2289 9058 2309
rect 9078 2289 9096 2309
rect 9047 2277 9096 2289
rect 9146 2313 9190 2319
rect 9146 2293 9161 2313
rect 9181 2293 9190 2313
rect 9146 2277 9190 2293
rect 9265 2309 9314 2319
rect 9265 2289 9276 2309
rect 9296 2289 9314 2309
rect 9265 2277 9314 2289
rect 9364 2313 9408 2319
rect 9364 2293 9379 2313
rect 9399 2293 9408 2313
rect 9364 2277 9408 2293
rect 9478 2313 9522 2319
rect 9478 2293 9487 2313
rect 9507 2293 9522 2313
rect 9478 2277 9522 2293
rect 9572 2309 9621 2319
rect 12101 2329 12150 2339
rect 12200 2355 12244 2371
rect 12200 2335 12215 2355
rect 12235 2335 12244 2355
rect 12200 2329 12244 2335
rect 12314 2355 12358 2371
rect 12314 2335 12323 2355
rect 12343 2335 12358 2355
rect 12314 2329 12358 2335
rect 12408 2359 12457 2371
rect 12408 2339 12426 2359
rect 12446 2339 12457 2359
rect 12408 2329 12457 2339
rect 12532 2355 12576 2371
rect 12532 2335 12541 2355
rect 12561 2335 12576 2355
rect 12532 2329 12576 2335
rect 12626 2359 12675 2371
rect 12626 2339 12644 2359
rect 12664 2339 12675 2359
rect 12626 2329 12675 2339
rect 9572 2289 9590 2309
rect 9610 2289 9621 2309
rect 9572 2277 9621 2289
rect 1104 2100 1153 2110
rect 1104 2080 1115 2100
rect 1135 2080 1153 2100
rect 1104 2068 1153 2080
rect 1203 2104 1247 2110
rect 1203 2084 1218 2104
rect 1238 2084 1247 2104
rect 1203 2068 1247 2084
rect 1322 2100 1371 2110
rect 1322 2080 1333 2100
rect 1353 2080 1371 2100
rect 1322 2068 1371 2080
rect 1421 2104 1465 2110
rect 1421 2084 1436 2104
rect 1456 2084 1465 2104
rect 1421 2068 1465 2084
rect 1535 2104 1579 2110
rect 1535 2084 1544 2104
rect 1564 2084 1579 2104
rect 1535 2068 1579 2084
rect 1629 2100 1678 2110
rect 1629 2080 1647 2100
rect 1667 2080 1678 2100
rect 1629 2068 1678 2080
rect 2463 2108 2512 2120
rect 2463 2088 2474 2108
rect 2494 2088 2512 2108
rect 2463 2078 2512 2088
rect 2562 2104 2606 2120
rect 2562 2084 2577 2104
rect 2597 2084 2606 2104
rect 2562 2078 2606 2084
rect 2676 2104 2720 2120
rect 2676 2084 2685 2104
rect 2705 2084 2720 2104
rect 2676 2078 2720 2084
rect 2770 2108 2819 2120
rect 2770 2088 2788 2108
rect 2808 2088 2819 2108
rect 2770 2078 2819 2088
rect 2894 2104 2938 2120
rect 2894 2084 2903 2104
rect 2923 2084 2938 2104
rect 2894 2078 2938 2084
rect 2988 2108 3037 2120
rect 16465 2372 16514 2384
rect 16465 2352 16476 2372
rect 16496 2352 16514 2372
rect 13411 2322 13460 2332
rect 13411 2302 13422 2322
rect 13442 2302 13460 2322
rect 13411 2290 13460 2302
rect 13510 2326 13554 2332
rect 13510 2306 13525 2326
rect 13545 2306 13554 2326
rect 13510 2290 13554 2306
rect 13629 2322 13678 2332
rect 13629 2302 13640 2322
rect 13660 2302 13678 2322
rect 13629 2290 13678 2302
rect 13728 2326 13772 2332
rect 13728 2306 13743 2326
rect 13763 2306 13772 2326
rect 13728 2290 13772 2306
rect 13842 2326 13886 2332
rect 13842 2306 13851 2326
rect 13871 2306 13886 2326
rect 13842 2290 13886 2306
rect 13936 2322 13985 2332
rect 16465 2342 16514 2352
rect 16564 2368 16608 2384
rect 16564 2348 16579 2368
rect 16599 2348 16608 2368
rect 16564 2342 16608 2348
rect 16678 2368 16722 2384
rect 16678 2348 16687 2368
rect 16707 2348 16722 2368
rect 16678 2342 16722 2348
rect 16772 2372 16821 2384
rect 16772 2352 16790 2372
rect 16810 2352 16821 2372
rect 16772 2342 16821 2352
rect 16896 2368 16940 2384
rect 16896 2348 16905 2368
rect 16925 2348 16940 2368
rect 16896 2342 16940 2348
rect 16990 2372 17039 2384
rect 16990 2352 17008 2372
rect 17028 2352 17039 2372
rect 16990 2342 17039 2352
rect 23004 2501 23053 2513
rect 23103 2537 23147 2543
rect 23103 2517 23118 2537
rect 23138 2517 23147 2537
rect 23103 2501 23147 2517
rect 23222 2533 23271 2543
rect 23222 2513 23233 2533
rect 23253 2513 23271 2533
rect 23222 2501 23271 2513
rect 23321 2537 23365 2543
rect 23321 2517 23336 2537
rect 23356 2517 23365 2537
rect 23321 2501 23365 2517
rect 23435 2537 23479 2543
rect 23435 2517 23444 2537
rect 23464 2517 23479 2537
rect 23435 2501 23479 2517
rect 23529 2533 23578 2543
rect 23529 2513 23547 2533
rect 23567 2513 23578 2533
rect 24297 2523 24308 2543
rect 24328 2523 24346 2543
rect 24297 2513 24346 2523
rect 24396 2539 24440 2555
rect 24396 2519 24411 2539
rect 24431 2519 24440 2539
rect 24396 2513 24440 2519
rect 24510 2539 24554 2555
rect 24510 2519 24519 2539
rect 24539 2519 24554 2539
rect 24510 2513 24554 2519
rect 24604 2543 24653 2555
rect 24604 2523 24622 2543
rect 24642 2523 24653 2543
rect 24604 2513 24653 2523
rect 24728 2539 24772 2555
rect 24728 2519 24737 2539
rect 24757 2519 24772 2539
rect 24728 2513 24772 2519
rect 24822 2543 24871 2555
rect 24822 2523 24840 2543
rect 24860 2523 24871 2543
rect 24822 2513 24871 2523
rect 28674 2555 28723 2567
rect 27381 2545 27430 2555
rect 27381 2525 27392 2545
rect 27412 2525 27430 2545
rect 23529 2501 23578 2513
rect 13936 2302 13954 2322
rect 13974 2302 13985 2322
rect 13936 2290 13985 2302
rect 2988 2088 3006 2108
rect 3026 2088 3037 2108
rect 2988 2078 3037 2088
rect 5468 2113 5517 2123
rect 5468 2093 5479 2113
rect 5499 2093 5517 2113
rect 5468 2081 5517 2093
rect 5567 2117 5611 2123
rect 5567 2097 5582 2117
rect 5602 2097 5611 2117
rect 5567 2081 5611 2097
rect 5686 2113 5735 2123
rect 5686 2093 5697 2113
rect 5717 2093 5735 2113
rect 5686 2081 5735 2093
rect 5785 2117 5829 2123
rect 5785 2097 5800 2117
rect 5820 2097 5829 2117
rect 5785 2081 5829 2097
rect 5899 2117 5943 2123
rect 5899 2097 5908 2117
rect 5928 2097 5943 2117
rect 5899 2081 5943 2097
rect 5993 2113 6042 2123
rect 5993 2093 6011 2113
rect 6031 2093 6042 2113
rect 5993 2081 6042 2093
rect 6827 2121 6876 2133
rect 6827 2101 6838 2121
rect 6858 2101 6876 2121
rect 6827 2091 6876 2101
rect 6926 2117 6970 2133
rect 6926 2097 6941 2117
rect 6961 2097 6970 2117
rect 6926 2091 6970 2097
rect 7040 2117 7084 2133
rect 7040 2097 7049 2117
rect 7069 2097 7084 2117
rect 7040 2091 7084 2097
rect 7134 2121 7183 2133
rect 7134 2101 7152 2121
rect 7172 2101 7183 2121
rect 7134 2091 7183 2101
rect 7258 2117 7302 2133
rect 7258 2097 7267 2117
rect 7287 2097 7302 2117
rect 7258 2091 7302 2097
rect 7352 2121 7401 2133
rect 27381 2513 27430 2525
rect 27480 2549 27524 2555
rect 27480 2529 27495 2549
rect 27515 2529 27524 2549
rect 27480 2513 27524 2529
rect 27599 2545 27648 2555
rect 27599 2525 27610 2545
rect 27630 2525 27648 2545
rect 27599 2513 27648 2525
rect 27698 2549 27742 2555
rect 27698 2529 27713 2549
rect 27733 2529 27742 2549
rect 27698 2513 27742 2529
rect 27812 2549 27856 2555
rect 27812 2529 27821 2549
rect 27841 2529 27856 2549
rect 27812 2513 27856 2529
rect 27906 2545 27955 2555
rect 27906 2525 27924 2545
rect 27944 2525 27955 2545
rect 28674 2535 28685 2555
rect 28705 2535 28723 2555
rect 28674 2525 28723 2535
rect 28773 2551 28817 2567
rect 28773 2531 28788 2551
rect 28808 2531 28817 2551
rect 28773 2525 28817 2531
rect 28887 2551 28931 2567
rect 28887 2531 28896 2551
rect 28916 2531 28931 2551
rect 28887 2525 28931 2531
rect 28981 2555 29030 2567
rect 28981 2535 28999 2555
rect 29019 2535 29030 2555
rect 28981 2525 29030 2535
rect 29105 2551 29149 2567
rect 29105 2531 29114 2551
rect 29134 2531 29149 2551
rect 29105 2525 29149 2531
rect 29199 2555 29248 2567
rect 29199 2535 29217 2555
rect 29237 2535 29248 2555
rect 29199 2525 29248 2535
rect 33038 2568 33087 2580
rect 31745 2558 31794 2568
rect 31745 2538 31756 2558
rect 31776 2538 31794 2558
rect 27906 2513 27955 2525
rect 20731 2346 20780 2358
rect 20731 2326 20742 2346
rect 20762 2326 20780 2346
rect 7352 2101 7370 2121
rect 7390 2101 7401 2121
rect 7352 2091 7401 2101
rect 9845 2125 9894 2135
rect 9845 2105 9856 2125
rect 9876 2105 9894 2125
rect 9845 2093 9894 2105
rect 9944 2129 9988 2135
rect 9944 2109 9959 2129
rect 9979 2109 9988 2129
rect 9944 2093 9988 2109
rect 10063 2125 10112 2135
rect 10063 2105 10074 2125
rect 10094 2105 10112 2125
rect 10063 2093 10112 2105
rect 10162 2129 10206 2135
rect 10162 2109 10177 2129
rect 10197 2109 10206 2129
rect 10162 2093 10206 2109
rect 10276 2129 10320 2135
rect 10276 2109 10285 2129
rect 10305 2109 10320 2129
rect 10276 2093 10320 2109
rect 10370 2125 10419 2135
rect 10370 2105 10388 2125
rect 10408 2105 10419 2125
rect 10370 2093 10419 2105
rect 11204 2133 11253 2145
rect 11204 2113 11215 2133
rect 11235 2113 11253 2133
rect 11204 2103 11253 2113
rect 11303 2129 11347 2145
rect 11303 2109 11318 2129
rect 11338 2109 11347 2129
rect 11303 2103 11347 2109
rect 11417 2129 11461 2145
rect 11417 2109 11426 2129
rect 11446 2109 11461 2129
rect 11417 2103 11461 2109
rect 11511 2133 11560 2145
rect 11511 2113 11529 2133
rect 11549 2113 11560 2133
rect 11511 2103 11560 2113
rect 11635 2129 11679 2145
rect 11635 2109 11644 2129
rect 11664 2109 11679 2129
rect 11635 2103 11679 2109
rect 11729 2133 11778 2145
rect 17677 2296 17726 2306
rect 17677 2276 17688 2296
rect 17708 2276 17726 2296
rect 17677 2264 17726 2276
rect 17776 2300 17820 2306
rect 17776 2280 17791 2300
rect 17811 2280 17820 2300
rect 17776 2264 17820 2280
rect 17895 2296 17944 2306
rect 17895 2276 17906 2296
rect 17926 2276 17944 2296
rect 17895 2264 17944 2276
rect 17994 2300 18038 2306
rect 17994 2280 18009 2300
rect 18029 2280 18038 2300
rect 17994 2264 18038 2280
rect 18108 2300 18152 2306
rect 18108 2280 18117 2300
rect 18137 2280 18152 2300
rect 18108 2264 18152 2280
rect 18202 2296 18251 2306
rect 20731 2316 20780 2326
rect 20830 2342 20874 2358
rect 20830 2322 20845 2342
rect 20865 2322 20874 2342
rect 20830 2316 20874 2322
rect 20944 2342 20988 2358
rect 20944 2322 20953 2342
rect 20973 2322 20988 2342
rect 20944 2316 20988 2322
rect 21038 2346 21087 2358
rect 21038 2326 21056 2346
rect 21076 2326 21087 2346
rect 21038 2316 21087 2326
rect 21162 2342 21206 2358
rect 21162 2322 21171 2342
rect 21191 2322 21206 2342
rect 21162 2316 21206 2322
rect 21256 2346 21305 2358
rect 21256 2326 21274 2346
rect 21294 2326 21305 2346
rect 21256 2316 21305 2326
rect 18202 2276 18220 2296
rect 18240 2276 18251 2296
rect 18202 2264 18251 2276
rect 31745 2526 31794 2538
rect 31844 2562 31888 2568
rect 31844 2542 31859 2562
rect 31879 2542 31888 2562
rect 31844 2526 31888 2542
rect 31963 2558 32012 2568
rect 31963 2538 31974 2558
rect 31994 2538 32012 2558
rect 31963 2526 32012 2538
rect 32062 2562 32106 2568
rect 32062 2542 32077 2562
rect 32097 2542 32106 2562
rect 32062 2526 32106 2542
rect 32176 2562 32220 2568
rect 32176 2542 32185 2562
rect 32205 2542 32220 2562
rect 32176 2526 32220 2542
rect 32270 2558 32319 2568
rect 32270 2538 32288 2558
rect 32308 2538 32319 2558
rect 33038 2548 33049 2568
rect 33069 2548 33087 2568
rect 33038 2538 33087 2548
rect 33137 2564 33181 2580
rect 33137 2544 33152 2564
rect 33172 2544 33181 2564
rect 33137 2538 33181 2544
rect 33251 2564 33295 2580
rect 33251 2544 33260 2564
rect 33280 2544 33295 2564
rect 33251 2538 33295 2544
rect 33345 2568 33394 2580
rect 33345 2548 33363 2568
rect 33383 2548 33394 2568
rect 33345 2538 33394 2548
rect 33469 2564 33513 2580
rect 33469 2544 33478 2564
rect 33498 2544 33513 2564
rect 33469 2538 33513 2544
rect 33563 2568 33612 2580
rect 33563 2548 33581 2568
rect 33601 2548 33612 2568
rect 33563 2538 33612 2548
rect 32270 2526 32319 2538
rect 25095 2359 25144 2371
rect 25095 2339 25106 2359
rect 25126 2339 25144 2359
rect 22041 2309 22090 2319
rect 22041 2289 22052 2309
rect 22072 2289 22090 2309
rect 22041 2277 22090 2289
rect 22140 2313 22184 2319
rect 22140 2293 22155 2313
rect 22175 2293 22184 2313
rect 22140 2277 22184 2293
rect 22259 2309 22308 2319
rect 22259 2289 22270 2309
rect 22290 2289 22308 2309
rect 22259 2277 22308 2289
rect 22358 2313 22402 2319
rect 22358 2293 22373 2313
rect 22393 2293 22402 2313
rect 22358 2277 22402 2293
rect 22472 2313 22516 2319
rect 22472 2293 22481 2313
rect 22501 2293 22516 2313
rect 22472 2277 22516 2293
rect 22566 2309 22615 2319
rect 25095 2329 25144 2339
rect 25194 2355 25238 2371
rect 25194 2335 25209 2355
rect 25229 2335 25238 2355
rect 25194 2329 25238 2335
rect 25308 2355 25352 2371
rect 25308 2335 25317 2355
rect 25337 2335 25352 2355
rect 25308 2329 25352 2335
rect 25402 2359 25451 2371
rect 25402 2339 25420 2359
rect 25440 2339 25451 2359
rect 25402 2329 25451 2339
rect 25526 2355 25570 2371
rect 25526 2335 25535 2355
rect 25555 2335 25570 2355
rect 25526 2329 25570 2335
rect 25620 2359 25669 2371
rect 25620 2339 25638 2359
rect 25658 2339 25669 2359
rect 25620 2329 25669 2339
rect 22566 2289 22584 2309
rect 22604 2289 22615 2309
rect 22566 2277 22615 2289
rect 11729 2113 11747 2133
rect 11767 2113 11778 2133
rect 11729 2103 11778 2113
rect 14209 2138 14258 2148
rect 14209 2118 14220 2138
rect 14240 2118 14258 2138
rect 307 1872 356 1882
rect 307 1852 318 1872
rect 338 1852 356 1872
rect 307 1840 356 1852
rect 406 1876 450 1882
rect 406 1856 421 1876
rect 441 1856 450 1876
rect 406 1840 450 1856
rect 525 1872 574 1882
rect 525 1852 536 1872
rect 556 1852 574 1872
rect 525 1840 574 1852
rect 624 1876 668 1882
rect 624 1856 639 1876
rect 659 1856 668 1876
rect 624 1840 668 1856
rect 738 1876 782 1882
rect 738 1856 747 1876
rect 767 1856 782 1876
rect 738 1840 782 1856
rect 832 1872 881 1882
rect 832 1852 850 1872
rect 870 1852 881 1872
rect 14209 2106 14258 2118
rect 14308 2142 14352 2148
rect 14308 2122 14323 2142
rect 14343 2122 14352 2142
rect 14308 2106 14352 2122
rect 14427 2138 14476 2148
rect 14427 2118 14438 2138
rect 14458 2118 14476 2138
rect 14427 2106 14476 2118
rect 14526 2142 14570 2148
rect 14526 2122 14541 2142
rect 14561 2122 14570 2142
rect 14526 2106 14570 2122
rect 14640 2142 14684 2148
rect 14640 2122 14649 2142
rect 14669 2122 14684 2142
rect 14640 2106 14684 2122
rect 14734 2138 14783 2148
rect 14734 2118 14752 2138
rect 14772 2118 14783 2138
rect 14734 2106 14783 2118
rect 15568 2146 15617 2158
rect 15568 2126 15579 2146
rect 15599 2126 15617 2146
rect 15568 2116 15617 2126
rect 15667 2142 15711 2158
rect 15667 2122 15682 2142
rect 15702 2122 15711 2142
rect 15667 2116 15711 2122
rect 15781 2142 15825 2158
rect 15781 2122 15790 2142
rect 15810 2122 15825 2142
rect 15781 2116 15825 2122
rect 15875 2146 15924 2158
rect 15875 2126 15893 2146
rect 15913 2126 15924 2146
rect 15875 2116 15924 2126
rect 15999 2142 16043 2158
rect 15999 2122 16008 2142
rect 16028 2122 16043 2142
rect 15999 2116 16043 2122
rect 16093 2146 16142 2158
rect 16093 2126 16111 2146
rect 16131 2126 16142 2146
rect 16093 2116 16142 2126
rect 29472 2371 29521 2383
rect 29472 2351 29483 2371
rect 29503 2351 29521 2371
rect 26418 2321 26467 2331
rect 26418 2301 26429 2321
rect 26449 2301 26467 2321
rect 26418 2289 26467 2301
rect 26517 2325 26561 2331
rect 26517 2305 26532 2325
rect 26552 2305 26561 2325
rect 26517 2289 26561 2305
rect 26636 2321 26685 2331
rect 26636 2301 26647 2321
rect 26667 2301 26685 2321
rect 26636 2289 26685 2301
rect 26735 2325 26779 2331
rect 26735 2305 26750 2325
rect 26770 2305 26779 2325
rect 26735 2289 26779 2305
rect 26849 2325 26893 2331
rect 26849 2305 26858 2325
rect 26878 2305 26893 2325
rect 26849 2289 26893 2305
rect 26943 2321 26992 2331
rect 29472 2341 29521 2351
rect 29571 2367 29615 2383
rect 29571 2347 29586 2367
rect 29606 2347 29615 2367
rect 29571 2341 29615 2347
rect 29685 2367 29729 2383
rect 29685 2347 29694 2367
rect 29714 2347 29729 2367
rect 29685 2341 29729 2347
rect 29779 2371 29828 2383
rect 29779 2351 29797 2371
rect 29817 2351 29828 2371
rect 29779 2341 29828 2351
rect 29903 2367 29947 2383
rect 29903 2347 29912 2367
rect 29932 2347 29947 2367
rect 29903 2341 29947 2347
rect 29997 2371 30046 2383
rect 29997 2351 30015 2371
rect 30035 2351 30046 2371
rect 29997 2341 30046 2351
rect 26943 2301 26961 2321
rect 26981 2301 26992 2321
rect 26943 2289 26992 2301
rect 832 1840 881 1852
rect 4671 1885 4720 1895
rect 4671 1865 4682 1885
rect 4702 1865 4720 1885
rect 4671 1853 4720 1865
rect 4770 1889 4814 1895
rect 4770 1869 4785 1889
rect 4805 1869 4814 1889
rect 4770 1853 4814 1869
rect 4889 1885 4938 1895
rect 4889 1865 4900 1885
rect 4920 1865 4938 1885
rect 4889 1853 4938 1865
rect 4988 1889 5032 1895
rect 4988 1869 5003 1889
rect 5023 1869 5032 1889
rect 4988 1853 5032 1869
rect 5102 1889 5146 1895
rect 5102 1869 5111 1889
rect 5131 1869 5146 1889
rect 5102 1853 5146 1869
rect 5196 1885 5245 1895
rect 5196 1865 5214 1885
rect 5234 1865 5245 1885
rect 18475 2112 18524 2122
rect 18475 2092 18486 2112
rect 18506 2092 18524 2112
rect 18475 2080 18524 2092
rect 18574 2116 18618 2122
rect 18574 2096 18589 2116
rect 18609 2096 18618 2116
rect 18574 2080 18618 2096
rect 18693 2112 18742 2122
rect 18693 2092 18704 2112
rect 18724 2092 18742 2112
rect 18693 2080 18742 2092
rect 18792 2116 18836 2122
rect 18792 2096 18807 2116
rect 18827 2096 18836 2116
rect 18792 2080 18836 2096
rect 18906 2116 18950 2122
rect 18906 2096 18915 2116
rect 18935 2096 18950 2116
rect 18906 2080 18950 2096
rect 19000 2112 19049 2122
rect 19000 2092 19018 2112
rect 19038 2092 19049 2112
rect 19000 2080 19049 2092
rect 19834 2120 19883 2132
rect 19834 2100 19845 2120
rect 19865 2100 19883 2120
rect 19834 2090 19883 2100
rect 19933 2116 19977 2132
rect 19933 2096 19948 2116
rect 19968 2096 19977 2116
rect 19933 2090 19977 2096
rect 20047 2116 20091 2132
rect 20047 2096 20056 2116
rect 20076 2096 20091 2116
rect 20047 2090 20091 2096
rect 20141 2120 20190 2132
rect 20141 2100 20159 2120
rect 20179 2100 20190 2120
rect 20141 2090 20190 2100
rect 20265 2116 20309 2132
rect 20265 2096 20274 2116
rect 20294 2096 20309 2116
rect 20265 2090 20309 2096
rect 20359 2120 20408 2132
rect 33836 2384 33885 2396
rect 33836 2364 33847 2384
rect 33867 2364 33885 2384
rect 30782 2334 30831 2344
rect 30782 2314 30793 2334
rect 30813 2314 30831 2334
rect 30782 2302 30831 2314
rect 30881 2338 30925 2344
rect 30881 2318 30896 2338
rect 30916 2318 30925 2338
rect 30881 2302 30925 2318
rect 31000 2334 31049 2344
rect 31000 2314 31011 2334
rect 31031 2314 31049 2334
rect 31000 2302 31049 2314
rect 31099 2338 31143 2344
rect 31099 2318 31114 2338
rect 31134 2318 31143 2338
rect 31099 2302 31143 2318
rect 31213 2338 31257 2344
rect 31213 2318 31222 2338
rect 31242 2318 31257 2338
rect 31213 2302 31257 2318
rect 31307 2334 31356 2344
rect 33836 2354 33885 2364
rect 33935 2380 33979 2396
rect 33935 2360 33950 2380
rect 33970 2360 33979 2380
rect 33935 2354 33979 2360
rect 34049 2380 34093 2396
rect 34049 2360 34058 2380
rect 34078 2360 34093 2380
rect 34049 2354 34093 2360
rect 34143 2384 34192 2396
rect 34143 2364 34161 2384
rect 34181 2364 34192 2384
rect 34143 2354 34192 2364
rect 34267 2380 34311 2396
rect 34267 2360 34276 2380
rect 34296 2360 34311 2380
rect 34267 2354 34311 2360
rect 34361 2384 34410 2396
rect 34361 2364 34379 2384
rect 34399 2364 34410 2384
rect 34361 2354 34410 2364
rect 31307 2314 31325 2334
rect 31345 2314 31356 2334
rect 31307 2302 31356 2314
rect 20359 2100 20377 2120
rect 20397 2100 20408 2120
rect 20359 2090 20408 2100
rect 22839 2125 22888 2135
rect 22839 2105 22850 2125
rect 22870 2105 22888 2125
rect 5196 1853 5245 1865
rect 9048 1897 9097 1907
rect 9048 1877 9059 1897
rect 9079 1877 9097 1897
rect 9048 1865 9097 1877
rect 9147 1901 9191 1907
rect 9147 1881 9162 1901
rect 9182 1881 9191 1901
rect 9147 1865 9191 1881
rect 9266 1897 9315 1907
rect 9266 1877 9277 1897
rect 9297 1877 9315 1897
rect 9266 1865 9315 1877
rect 9365 1901 9409 1907
rect 9365 1881 9380 1901
rect 9400 1881 9409 1901
rect 9365 1865 9409 1881
rect 9479 1901 9523 1907
rect 9479 1881 9488 1901
rect 9508 1881 9523 1901
rect 9479 1865 9523 1881
rect 9573 1897 9622 1907
rect 9573 1877 9591 1897
rect 9611 1877 9622 1897
rect 22839 2093 22888 2105
rect 22938 2129 22982 2135
rect 22938 2109 22953 2129
rect 22973 2109 22982 2129
rect 22938 2093 22982 2109
rect 23057 2125 23106 2135
rect 23057 2105 23068 2125
rect 23088 2105 23106 2125
rect 23057 2093 23106 2105
rect 23156 2129 23200 2135
rect 23156 2109 23171 2129
rect 23191 2109 23200 2129
rect 23156 2093 23200 2109
rect 23270 2129 23314 2135
rect 23270 2109 23279 2129
rect 23299 2109 23314 2129
rect 23270 2093 23314 2109
rect 23364 2125 23413 2135
rect 23364 2105 23382 2125
rect 23402 2105 23413 2125
rect 23364 2093 23413 2105
rect 24198 2133 24247 2145
rect 24198 2113 24209 2133
rect 24229 2113 24247 2133
rect 24198 2103 24247 2113
rect 24297 2129 24341 2145
rect 24297 2109 24312 2129
rect 24332 2109 24341 2129
rect 24297 2103 24341 2109
rect 24411 2129 24455 2145
rect 24411 2109 24420 2129
rect 24440 2109 24455 2129
rect 24411 2103 24455 2109
rect 24505 2133 24554 2145
rect 24505 2113 24523 2133
rect 24543 2113 24554 2133
rect 24505 2103 24554 2113
rect 24629 2129 24673 2145
rect 24629 2109 24638 2129
rect 24658 2109 24673 2129
rect 24629 2103 24673 2109
rect 24723 2133 24772 2145
rect 24723 2113 24741 2133
rect 24761 2113 24772 2133
rect 24723 2103 24772 2113
rect 9573 1865 9622 1877
rect 13412 1910 13461 1920
rect 13412 1890 13423 1910
rect 13443 1890 13461 1910
rect 13412 1878 13461 1890
rect 13511 1914 13555 1920
rect 13511 1894 13526 1914
rect 13546 1894 13555 1914
rect 13511 1878 13555 1894
rect 13630 1910 13679 1920
rect 13630 1890 13641 1910
rect 13661 1890 13679 1910
rect 13630 1878 13679 1890
rect 13729 1914 13773 1920
rect 13729 1894 13744 1914
rect 13764 1894 13773 1914
rect 13729 1878 13773 1894
rect 13843 1914 13887 1920
rect 13843 1894 13852 1914
rect 13872 1894 13887 1914
rect 13843 1878 13887 1894
rect 13937 1910 13986 1920
rect 13937 1890 13955 1910
rect 13975 1890 13986 1910
rect 13937 1878 13986 1890
rect 27216 2137 27265 2147
rect 27216 2117 27227 2137
rect 27247 2117 27265 2137
rect 27216 2105 27265 2117
rect 27315 2141 27359 2147
rect 27315 2121 27330 2141
rect 27350 2121 27359 2141
rect 27315 2105 27359 2121
rect 27434 2137 27483 2147
rect 27434 2117 27445 2137
rect 27465 2117 27483 2137
rect 27434 2105 27483 2117
rect 27533 2141 27577 2147
rect 27533 2121 27548 2141
rect 27568 2121 27577 2141
rect 27533 2105 27577 2121
rect 27647 2141 27691 2147
rect 27647 2121 27656 2141
rect 27676 2121 27691 2141
rect 27647 2105 27691 2121
rect 27741 2137 27790 2147
rect 27741 2117 27759 2137
rect 27779 2117 27790 2137
rect 27741 2105 27790 2117
rect 28575 2145 28624 2157
rect 28575 2125 28586 2145
rect 28606 2125 28624 2145
rect 28575 2115 28624 2125
rect 28674 2141 28718 2157
rect 28674 2121 28689 2141
rect 28709 2121 28718 2141
rect 28674 2115 28718 2121
rect 28788 2141 28832 2157
rect 28788 2121 28797 2141
rect 28817 2121 28832 2141
rect 28788 2115 28832 2121
rect 28882 2145 28931 2157
rect 28882 2125 28900 2145
rect 28920 2125 28931 2145
rect 28882 2115 28931 2125
rect 29006 2141 29050 2157
rect 29006 2121 29015 2141
rect 29035 2121 29050 2141
rect 29006 2115 29050 2121
rect 29100 2145 29149 2157
rect 29100 2125 29118 2145
rect 29138 2125 29149 2145
rect 29100 2115 29149 2125
rect 31580 2150 31629 2160
rect 31580 2130 31591 2150
rect 31611 2130 31629 2150
rect 17678 1884 17727 1894
rect 17678 1864 17689 1884
rect 17709 1864 17727 1884
rect 17678 1852 17727 1864
rect 17777 1888 17821 1894
rect 17777 1868 17792 1888
rect 17812 1868 17821 1888
rect 17777 1852 17821 1868
rect 17896 1884 17945 1894
rect 17896 1864 17907 1884
rect 17927 1864 17945 1884
rect 17896 1852 17945 1864
rect 17995 1888 18039 1894
rect 17995 1868 18010 1888
rect 18030 1868 18039 1888
rect 17995 1852 18039 1868
rect 18109 1888 18153 1894
rect 18109 1868 18118 1888
rect 18138 1868 18153 1888
rect 18109 1852 18153 1868
rect 18203 1884 18252 1894
rect 18203 1864 18221 1884
rect 18241 1864 18252 1884
rect 31580 2118 31629 2130
rect 31679 2154 31723 2160
rect 31679 2134 31694 2154
rect 31714 2134 31723 2154
rect 31679 2118 31723 2134
rect 31798 2150 31847 2160
rect 31798 2130 31809 2150
rect 31829 2130 31847 2150
rect 31798 2118 31847 2130
rect 31897 2154 31941 2160
rect 31897 2134 31912 2154
rect 31932 2134 31941 2154
rect 31897 2118 31941 2134
rect 32011 2154 32055 2160
rect 32011 2134 32020 2154
rect 32040 2134 32055 2154
rect 32011 2118 32055 2134
rect 32105 2150 32154 2160
rect 32105 2130 32123 2150
rect 32143 2130 32154 2150
rect 32105 2118 32154 2130
rect 32939 2158 32988 2170
rect 32939 2138 32950 2158
rect 32970 2138 32988 2158
rect 32939 2128 32988 2138
rect 33038 2154 33082 2170
rect 33038 2134 33053 2154
rect 33073 2134 33082 2154
rect 33038 2128 33082 2134
rect 33152 2154 33196 2170
rect 33152 2134 33161 2154
rect 33181 2134 33196 2154
rect 33152 2128 33196 2134
rect 33246 2158 33295 2170
rect 33246 2138 33264 2158
rect 33284 2138 33295 2158
rect 33246 2128 33295 2138
rect 33370 2154 33414 2170
rect 33370 2134 33379 2154
rect 33399 2134 33414 2154
rect 33370 2128 33414 2134
rect 33464 2158 33513 2170
rect 33464 2138 33482 2158
rect 33502 2138 33513 2158
rect 33464 2128 33513 2138
rect 18203 1852 18252 1864
rect 22042 1897 22091 1907
rect 22042 1877 22053 1897
rect 22073 1877 22091 1897
rect 22042 1865 22091 1877
rect 22141 1901 22185 1907
rect 22141 1881 22156 1901
rect 22176 1881 22185 1901
rect 22141 1865 22185 1881
rect 22260 1897 22309 1907
rect 22260 1877 22271 1897
rect 22291 1877 22309 1897
rect 22260 1865 22309 1877
rect 22359 1901 22403 1907
rect 22359 1881 22374 1901
rect 22394 1881 22403 1901
rect 22359 1865 22403 1881
rect 22473 1901 22517 1907
rect 22473 1881 22482 1901
rect 22502 1881 22517 1901
rect 22473 1865 22517 1881
rect 22567 1897 22616 1907
rect 22567 1877 22585 1897
rect 22605 1877 22616 1897
rect 22567 1865 22616 1877
rect 26419 1909 26468 1919
rect 26419 1889 26430 1909
rect 26450 1889 26468 1909
rect 26419 1877 26468 1889
rect 26518 1913 26562 1919
rect 26518 1893 26533 1913
rect 26553 1893 26562 1913
rect 26518 1877 26562 1893
rect 26637 1909 26686 1919
rect 26637 1889 26648 1909
rect 26668 1889 26686 1909
rect 26637 1877 26686 1889
rect 26736 1913 26780 1919
rect 26736 1893 26751 1913
rect 26771 1893 26780 1913
rect 26736 1877 26780 1893
rect 26850 1913 26894 1919
rect 26850 1893 26859 1913
rect 26879 1893 26894 1913
rect 26850 1877 26894 1893
rect 26944 1909 26993 1919
rect 26944 1889 26962 1909
rect 26982 1889 26993 1909
rect 26944 1877 26993 1889
rect 30783 1922 30832 1932
rect 30783 1902 30794 1922
rect 30814 1902 30832 1922
rect 30783 1890 30832 1902
rect 30882 1926 30926 1932
rect 30882 1906 30897 1926
rect 30917 1906 30926 1926
rect 30882 1890 30926 1906
rect 31001 1922 31050 1932
rect 31001 1902 31012 1922
rect 31032 1902 31050 1922
rect 31001 1890 31050 1902
rect 31100 1926 31144 1932
rect 31100 1906 31115 1926
rect 31135 1906 31144 1926
rect 31100 1890 31144 1906
rect 31214 1926 31258 1932
rect 31214 1906 31223 1926
rect 31243 1906 31258 1926
rect 31214 1890 31258 1906
rect 31308 1922 31357 1932
rect 31308 1902 31326 1922
rect 31346 1902 31357 1922
rect 31308 1890 31357 1902
rect 3342 1728 3391 1740
rect 3342 1708 3353 1728
rect 3373 1708 3391 1728
rect 3342 1698 3391 1708
rect 3441 1724 3485 1740
rect 3441 1704 3456 1724
rect 3476 1704 3485 1724
rect 3441 1698 3485 1704
rect 3555 1724 3599 1740
rect 3555 1704 3564 1724
rect 3584 1704 3599 1724
rect 3555 1698 3599 1704
rect 3649 1728 3698 1740
rect 3649 1708 3667 1728
rect 3687 1708 3698 1728
rect 3649 1698 3698 1708
rect 3773 1724 3817 1740
rect 3773 1704 3782 1724
rect 3802 1704 3817 1724
rect 3773 1698 3817 1704
rect 3867 1728 3916 1740
rect 3867 1708 3885 1728
rect 3905 1708 3916 1728
rect 3867 1698 3916 1708
rect 7706 1741 7755 1753
rect 7706 1721 7717 1741
rect 7737 1721 7755 1741
rect 7706 1711 7755 1721
rect 7805 1737 7849 1753
rect 7805 1717 7820 1737
rect 7840 1717 7849 1737
rect 7805 1711 7849 1717
rect 7919 1737 7963 1753
rect 7919 1717 7928 1737
rect 7948 1717 7963 1737
rect 7919 1711 7963 1717
rect 8013 1741 8062 1753
rect 8013 1721 8031 1741
rect 8051 1721 8062 1741
rect 8013 1711 8062 1721
rect 8137 1737 8181 1753
rect 8137 1717 8146 1737
rect 8166 1717 8181 1737
rect 8137 1711 8181 1717
rect 8231 1741 8280 1753
rect 8231 1721 8249 1741
rect 8269 1721 8280 1741
rect 8231 1711 8280 1721
rect 12083 1753 12132 1765
rect 12083 1733 12094 1753
rect 12114 1733 12132 1753
rect 12083 1723 12132 1733
rect 12182 1749 12226 1765
rect 12182 1729 12197 1749
rect 12217 1729 12226 1749
rect 12182 1723 12226 1729
rect 12296 1749 12340 1765
rect 12296 1729 12305 1749
rect 12325 1729 12340 1749
rect 12296 1723 12340 1729
rect 12390 1753 12439 1765
rect 12390 1733 12408 1753
rect 12428 1733 12439 1753
rect 12390 1723 12439 1733
rect 12514 1749 12558 1765
rect 12514 1729 12523 1749
rect 12543 1729 12558 1749
rect 12514 1723 12558 1729
rect 12608 1753 12657 1765
rect 12608 1733 12626 1753
rect 12646 1733 12657 1753
rect 12608 1723 12657 1733
rect 16447 1766 16496 1778
rect 1186 1492 1235 1502
rect 1186 1472 1197 1492
rect 1217 1472 1235 1492
rect 1186 1460 1235 1472
rect 1285 1496 1329 1502
rect 1285 1476 1300 1496
rect 1320 1476 1329 1496
rect 1285 1460 1329 1476
rect 1404 1492 1453 1502
rect 1404 1472 1415 1492
rect 1435 1472 1453 1492
rect 1404 1460 1453 1472
rect 1503 1496 1547 1502
rect 1503 1476 1518 1496
rect 1538 1476 1547 1496
rect 1503 1460 1547 1476
rect 1617 1496 1661 1502
rect 1617 1476 1626 1496
rect 1646 1476 1661 1496
rect 1617 1460 1661 1476
rect 1711 1492 1760 1502
rect 1711 1472 1729 1492
rect 1749 1472 1760 1492
rect 1711 1460 1760 1472
rect 2545 1500 2594 1512
rect 2545 1480 2556 1500
rect 2576 1480 2594 1500
rect 2545 1470 2594 1480
rect 2644 1496 2688 1512
rect 2644 1476 2659 1496
rect 2679 1476 2688 1496
rect 2644 1470 2688 1476
rect 2758 1496 2802 1512
rect 2758 1476 2767 1496
rect 2787 1476 2802 1496
rect 2758 1470 2802 1476
rect 2852 1500 2901 1512
rect 2852 1480 2870 1500
rect 2890 1480 2901 1500
rect 2852 1470 2901 1480
rect 2976 1496 3020 1512
rect 2976 1476 2985 1496
rect 3005 1476 3020 1496
rect 2976 1470 3020 1476
rect 3070 1500 3119 1512
rect 16447 1746 16458 1766
rect 16478 1746 16496 1766
rect 16447 1736 16496 1746
rect 16546 1762 16590 1778
rect 16546 1742 16561 1762
rect 16581 1742 16590 1762
rect 16546 1736 16590 1742
rect 16660 1762 16704 1778
rect 16660 1742 16669 1762
rect 16689 1742 16704 1762
rect 16660 1736 16704 1742
rect 16754 1766 16803 1778
rect 16754 1746 16772 1766
rect 16792 1746 16803 1766
rect 16754 1736 16803 1746
rect 16878 1762 16922 1778
rect 16878 1742 16887 1762
rect 16907 1742 16922 1762
rect 16878 1736 16922 1742
rect 16972 1766 17021 1778
rect 16972 1746 16990 1766
rect 17010 1746 17021 1766
rect 16972 1736 17021 1746
rect 3070 1480 3088 1500
rect 3108 1480 3119 1500
rect 3070 1470 3119 1480
rect 5550 1505 5599 1515
rect 5550 1485 5561 1505
rect 5581 1485 5599 1505
rect 5550 1473 5599 1485
rect 5649 1509 5693 1515
rect 5649 1489 5664 1509
rect 5684 1489 5693 1509
rect 5649 1473 5693 1489
rect 5768 1505 5817 1515
rect 5768 1485 5779 1505
rect 5799 1485 5817 1505
rect 5768 1473 5817 1485
rect 5867 1509 5911 1515
rect 5867 1489 5882 1509
rect 5902 1489 5911 1509
rect 5867 1473 5911 1489
rect 5981 1509 6025 1515
rect 5981 1489 5990 1509
rect 6010 1489 6025 1509
rect 5981 1473 6025 1489
rect 6075 1505 6124 1515
rect 6075 1485 6093 1505
rect 6113 1485 6124 1505
rect 6075 1473 6124 1485
rect 6909 1513 6958 1525
rect 6909 1493 6920 1513
rect 6940 1493 6958 1513
rect 6909 1483 6958 1493
rect 7008 1509 7052 1525
rect 7008 1489 7023 1509
rect 7043 1489 7052 1509
rect 7008 1483 7052 1489
rect 7122 1509 7166 1525
rect 7122 1489 7131 1509
rect 7151 1489 7166 1509
rect 7122 1483 7166 1489
rect 7216 1513 7265 1525
rect 7216 1493 7234 1513
rect 7254 1493 7265 1513
rect 7216 1483 7265 1493
rect 7340 1509 7384 1525
rect 7340 1489 7349 1509
rect 7369 1489 7384 1509
rect 7340 1483 7384 1489
rect 7434 1513 7483 1525
rect 7434 1493 7452 1513
rect 7472 1493 7483 1513
rect 7434 1483 7483 1493
rect 20713 1740 20762 1752
rect 20713 1720 20724 1740
rect 20744 1720 20762 1740
rect 20713 1710 20762 1720
rect 20812 1736 20856 1752
rect 20812 1716 20827 1736
rect 20847 1716 20856 1736
rect 20812 1710 20856 1716
rect 20926 1736 20970 1752
rect 20926 1716 20935 1736
rect 20955 1716 20970 1736
rect 20926 1710 20970 1716
rect 21020 1740 21069 1752
rect 21020 1720 21038 1740
rect 21058 1720 21069 1740
rect 21020 1710 21069 1720
rect 21144 1736 21188 1752
rect 21144 1716 21153 1736
rect 21173 1716 21188 1736
rect 21144 1710 21188 1716
rect 21238 1740 21287 1752
rect 21238 1720 21256 1740
rect 21276 1720 21287 1740
rect 21238 1710 21287 1720
rect 25077 1753 25126 1765
rect 9927 1517 9976 1527
rect 9927 1497 9938 1517
rect 9958 1497 9976 1517
rect 9927 1485 9976 1497
rect 10026 1521 10070 1527
rect 10026 1501 10041 1521
rect 10061 1501 10070 1521
rect 10026 1485 10070 1501
rect 10145 1517 10194 1527
rect 10145 1497 10156 1517
rect 10176 1497 10194 1517
rect 10145 1485 10194 1497
rect 10244 1521 10288 1527
rect 10244 1501 10259 1521
rect 10279 1501 10288 1521
rect 10244 1485 10288 1501
rect 10358 1521 10402 1527
rect 10358 1501 10367 1521
rect 10387 1501 10402 1521
rect 10358 1485 10402 1501
rect 10452 1517 10501 1527
rect 10452 1497 10470 1517
rect 10490 1497 10501 1517
rect 10452 1485 10501 1497
rect 11286 1525 11335 1537
rect 11286 1505 11297 1525
rect 11317 1505 11335 1525
rect 11286 1495 11335 1505
rect 11385 1521 11429 1537
rect 11385 1501 11400 1521
rect 11420 1501 11429 1521
rect 11385 1495 11429 1501
rect 11499 1521 11543 1537
rect 11499 1501 11508 1521
rect 11528 1501 11543 1521
rect 11499 1495 11543 1501
rect 11593 1525 11642 1537
rect 11593 1505 11611 1525
rect 11631 1505 11642 1525
rect 11593 1495 11642 1505
rect 11717 1521 11761 1537
rect 11717 1501 11726 1521
rect 11746 1501 11761 1521
rect 11717 1495 11761 1501
rect 11811 1525 11860 1537
rect 25077 1733 25088 1753
rect 25108 1733 25126 1753
rect 25077 1723 25126 1733
rect 25176 1749 25220 1765
rect 25176 1729 25191 1749
rect 25211 1729 25220 1749
rect 25176 1723 25220 1729
rect 25290 1749 25334 1765
rect 25290 1729 25299 1749
rect 25319 1729 25334 1749
rect 25290 1723 25334 1729
rect 25384 1753 25433 1765
rect 25384 1733 25402 1753
rect 25422 1733 25433 1753
rect 25384 1723 25433 1733
rect 25508 1749 25552 1765
rect 25508 1729 25517 1749
rect 25537 1729 25552 1749
rect 25508 1723 25552 1729
rect 25602 1753 25651 1765
rect 25602 1733 25620 1753
rect 25640 1733 25651 1753
rect 25602 1723 25651 1733
rect 29454 1765 29503 1777
rect 11811 1505 11829 1525
rect 11849 1505 11860 1525
rect 11811 1495 11860 1505
rect 14291 1530 14340 1540
rect 14291 1510 14302 1530
rect 14322 1510 14340 1530
rect 3343 1316 3392 1328
rect 3343 1296 3354 1316
rect 3374 1296 3392 1316
rect 289 1266 338 1276
rect 289 1246 300 1266
rect 320 1246 338 1266
rect 289 1234 338 1246
rect 388 1270 432 1276
rect 388 1250 403 1270
rect 423 1250 432 1270
rect 388 1234 432 1250
rect 507 1266 556 1276
rect 507 1246 518 1266
rect 538 1246 556 1266
rect 507 1234 556 1246
rect 606 1270 650 1276
rect 606 1250 621 1270
rect 641 1250 650 1270
rect 606 1234 650 1250
rect 720 1270 764 1276
rect 720 1250 729 1270
rect 749 1250 764 1270
rect 720 1234 764 1250
rect 814 1266 863 1276
rect 3343 1286 3392 1296
rect 3442 1312 3486 1328
rect 3442 1292 3457 1312
rect 3477 1292 3486 1312
rect 3442 1286 3486 1292
rect 3556 1312 3600 1328
rect 3556 1292 3565 1312
rect 3585 1292 3600 1312
rect 3556 1286 3600 1292
rect 3650 1316 3699 1328
rect 3650 1296 3668 1316
rect 3688 1296 3699 1316
rect 3650 1286 3699 1296
rect 3774 1312 3818 1328
rect 3774 1292 3783 1312
rect 3803 1292 3818 1312
rect 3774 1286 3818 1292
rect 3868 1316 3917 1328
rect 3868 1296 3886 1316
rect 3906 1296 3917 1316
rect 3868 1286 3917 1296
rect 814 1246 832 1266
rect 852 1246 863 1266
rect 814 1234 863 1246
rect 14291 1498 14340 1510
rect 14390 1534 14434 1540
rect 14390 1514 14405 1534
rect 14425 1514 14434 1534
rect 14390 1498 14434 1514
rect 14509 1530 14558 1540
rect 14509 1510 14520 1530
rect 14540 1510 14558 1530
rect 14509 1498 14558 1510
rect 14608 1534 14652 1540
rect 14608 1514 14623 1534
rect 14643 1514 14652 1534
rect 14608 1498 14652 1514
rect 14722 1534 14766 1540
rect 14722 1514 14731 1534
rect 14751 1514 14766 1534
rect 14722 1498 14766 1514
rect 14816 1530 14865 1540
rect 14816 1510 14834 1530
rect 14854 1510 14865 1530
rect 14816 1498 14865 1510
rect 15650 1538 15699 1550
rect 15650 1518 15661 1538
rect 15681 1518 15699 1538
rect 15650 1508 15699 1518
rect 15749 1534 15793 1550
rect 15749 1514 15764 1534
rect 15784 1514 15793 1534
rect 15749 1508 15793 1514
rect 15863 1534 15907 1550
rect 15863 1514 15872 1534
rect 15892 1514 15907 1534
rect 15863 1508 15907 1514
rect 15957 1538 16006 1550
rect 15957 1518 15975 1538
rect 15995 1518 16006 1538
rect 15957 1508 16006 1518
rect 16081 1534 16125 1550
rect 16081 1514 16090 1534
rect 16110 1514 16125 1534
rect 16081 1508 16125 1514
rect 16175 1538 16224 1550
rect 16175 1518 16193 1538
rect 16213 1518 16224 1538
rect 16175 1508 16224 1518
rect 29454 1745 29465 1765
rect 29485 1745 29503 1765
rect 29454 1735 29503 1745
rect 29553 1761 29597 1777
rect 29553 1741 29568 1761
rect 29588 1741 29597 1761
rect 29553 1735 29597 1741
rect 29667 1761 29711 1777
rect 29667 1741 29676 1761
rect 29696 1741 29711 1761
rect 29667 1735 29711 1741
rect 29761 1765 29810 1777
rect 29761 1745 29779 1765
rect 29799 1745 29810 1765
rect 29761 1735 29810 1745
rect 29885 1761 29929 1777
rect 29885 1741 29894 1761
rect 29914 1741 29929 1761
rect 29885 1735 29929 1741
rect 29979 1765 30028 1777
rect 29979 1745 29997 1765
rect 30017 1745 30028 1765
rect 29979 1735 30028 1745
rect 33818 1778 33867 1790
rect 7707 1329 7756 1341
rect 7707 1309 7718 1329
rect 7738 1309 7756 1329
rect 4653 1279 4702 1289
rect 4653 1259 4664 1279
rect 4684 1259 4702 1279
rect 4653 1247 4702 1259
rect 4752 1283 4796 1289
rect 4752 1263 4767 1283
rect 4787 1263 4796 1283
rect 4752 1247 4796 1263
rect 4871 1279 4920 1289
rect 4871 1259 4882 1279
rect 4902 1259 4920 1279
rect 4871 1247 4920 1259
rect 4970 1283 5014 1289
rect 4970 1263 4985 1283
rect 5005 1263 5014 1283
rect 4970 1247 5014 1263
rect 5084 1283 5128 1289
rect 5084 1263 5093 1283
rect 5113 1263 5128 1283
rect 5084 1247 5128 1263
rect 5178 1279 5227 1289
rect 7707 1299 7756 1309
rect 7806 1325 7850 1341
rect 7806 1305 7821 1325
rect 7841 1305 7850 1325
rect 7806 1299 7850 1305
rect 7920 1325 7964 1341
rect 7920 1305 7929 1325
rect 7949 1305 7964 1325
rect 7920 1299 7964 1305
rect 8014 1329 8063 1341
rect 8014 1309 8032 1329
rect 8052 1309 8063 1329
rect 8014 1299 8063 1309
rect 8138 1325 8182 1341
rect 8138 1305 8147 1325
rect 8167 1305 8182 1325
rect 8138 1299 8182 1305
rect 8232 1329 8281 1341
rect 8232 1309 8250 1329
rect 8270 1309 8281 1329
rect 8232 1299 8281 1309
rect 5178 1259 5196 1279
rect 5216 1259 5227 1279
rect 5178 1247 5227 1259
rect 18557 1504 18606 1514
rect 18557 1484 18568 1504
rect 18588 1484 18606 1504
rect 18557 1472 18606 1484
rect 18656 1508 18700 1514
rect 18656 1488 18671 1508
rect 18691 1488 18700 1508
rect 18656 1472 18700 1488
rect 18775 1504 18824 1514
rect 18775 1484 18786 1504
rect 18806 1484 18824 1504
rect 18775 1472 18824 1484
rect 18874 1508 18918 1514
rect 18874 1488 18889 1508
rect 18909 1488 18918 1508
rect 18874 1472 18918 1488
rect 18988 1508 19032 1514
rect 18988 1488 18997 1508
rect 19017 1488 19032 1508
rect 18988 1472 19032 1488
rect 19082 1504 19131 1514
rect 19082 1484 19100 1504
rect 19120 1484 19131 1504
rect 19082 1472 19131 1484
rect 19916 1512 19965 1524
rect 19916 1492 19927 1512
rect 19947 1492 19965 1512
rect 19916 1482 19965 1492
rect 20015 1508 20059 1524
rect 20015 1488 20030 1508
rect 20050 1488 20059 1508
rect 20015 1482 20059 1488
rect 20129 1508 20173 1524
rect 20129 1488 20138 1508
rect 20158 1488 20173 1508
rect 20129 1482 20173 1488
rect 20223 1512 20272 1524
rect 20223 1492 20241 1512
rect 20261 1492 20272 1512
rect 20223 1482 20272 1492
rect 20347 1508 20391 1524
rect 20347 1488 20356 1508
rect 20376 1488 20391 1508
rect 20347 1482 20391 1488
rect 20441 1512 20490 1524
rect 33818 1758 33829 1778
rect 33849 1758 33867 1778
rect 33818 1748 33867 1758
rect 33917 1774 33961 1790
rect 33917 1754 33932 1774
rect 33952 1754 33961 1774
rect 33917 1748 33961 1754
rect 34031 1774 34075 1790
rect 34031 1754 34040 1774
rect 34060 1754 34075 1774
rect 34031 1748 34075 1754
rect 34125 1778 34174 1790
rect 34125 1758 34143 1778
rect 34163 1758 34174 1778
rect 34125 1748 34174 1758
rect 34249 1774 34293 1790
rect 34249 1754 34258 1774
rect 34278 1754 34293 1774
rect 34249 1748 34293 1754
rect 34343 1778 34392 1790
rect 34343 1758 34361 1778
rect 34381 1758 34392 1778
rect 34343 1748 34392 1758
rect 20441 1492 20459 1512
rect 20479 1492 20490 1512
rect 20441 1482 20490 1492
rect 22921 1517 22970 1527
rect 22921 1497 22932 1517
rect 22952 1497 22970 1517
rect 12084 1341 12133 1353
rect 12084 1321 12095 1341
rect 12115 1321 12133 1341
rect 9030 1291 9079 1301
rect 9030 1271 9041 1291
rect 9061 1271 9079 1291
rect 9030 1259 9079 1271
rect 9129 1295 9173 1301
rect 9129 1275 9144 1295
rect 9164 1275 9173 1295
rect 9129 1259 9173 1275
rect 9248 1291 9297 1301
rect 9248 1271 9259 1291
rect 9279 1271 9297 1291
rect 9248 1259 9297 1271
rect 9347 1295 9391 1301
rect 9347 1275 9362 1295
rect 9382 1275 9391 1295
rect 9347 1259 9391 1275
rect 9461 1295 9505 1301
rect 9461 1275 9470 1295
rect 9490 1275 9505 1295
rect 9461 1259 9505 1275
rect 9555 1291 9604 1301
rect 12084 1311 12133 1321
rect 12183 1337 12227 1353
rect 12183 1317 12198 1337
rect 12218 1317 12227 1337
rect 12183 1311 12227 1317
rect 12297 1337 12341 1353
rect 12297 1317 12306 1337
rect 12326 1317 12341 1337
rect 12297 1311 12341 1317
rect 12391 1341 12440 1353
rect 12391 1321 12409 1341
rect 12429 1321 12440 1341
rect 12391 1311 12440 1321
rect 12515 1337 12559 1353
rect 12515 1317 12524 1337
rect 12544 1317 12559 1337
rect 12515 1311 12559 1317
rect 12609 1341 12658 1353
rect 12609 1321 12627 1341
rect 12647 1321 12658 1341
rect 12609 1311 12658 1321
rect 9555 1271 9573 1291
rect 9593 1271 9604 1291
rect 9555 1259 9604 1271
rect 16448 1354 16497 1366
rect 16448 1334 16459 1354
rect 16479 1334 16497 1354
rect 13394 1304 13443 1314
rect 13394 1284 13405 1304
rect 13425 1284 13443 1304
rect 13394 1272 13443 1284
rect 13493 1308 13537 1314
rect 13493 1288 13508 1308
rect 13528 1288 13537 1308
rect 13493 1272 13537 1288
rect 13612 1304 13661 1314
rect 13612 1284 13623 1304
rect 13643 1284 13661 1304
rect 13612 1272 13661 1284
rect 13711 1308 13755 1314
rect 13711 1288 13726 1308
rect 13746 1288 13755 1308
rect 13711 1272 13755 1288
rect 13825 1308 13869 1314
rect 13825 1288 13834 1308
rect 13854 1288 13869 1308
rect 13825 1272 13869 1288
rect 13919 1304 13968 1314
rect 16448 1324 16497 1334
rect 16547 1350 16591 1366
rect 16547 1330 16562 1350
rect 16582 1330 16591 1350
rect 16547 1324 16591 1330
rect 16661 1350 16705 1366
rect 16661 1330 16670 1350
rect 16690 1330 16705 1350
rect 16661 1324 16705 1330
rect 16755 1354 16804 1366
rect 16755 1334 16773 1354
rect 16793 1334 16804 1354
rect 16755 1324 16804 1334
rect 16879 1350 16923 1366
rect 16879 1330 16888 1350
rect 16908 1330 16923 1350
rect 16879 1324 16923 1330
rect 16973 1354 17022 1366
rect 16973 1334 16991 1354
rect 17011 1334 17022 1354
rect 16973 1324 17022 1334
rect 22921 1485 22970 1497
rect 23020 1521 23064 1527
rect 23020 1501 23035 1521
rect 23055 1501 23064 1521
rect 23020 1485 23064 1501
rect 23139 1517 23188 1527
rect 23139 1497 23150 1517
rect 23170 1497 23188 1517
rect 23139 1485 23188 1497
rect 23238 1521 23282 1527
rect 23238 1501 23253 1521
rect 23273 1501 23282 1521
rect 23238 1485 23282 1501
rect 23352 1521 23396 1527
rect 23352 1501 23361 1521
rect 23381 1501 23396 1521
rect 23352 1485 23396 1501
rect 23446 1517 23495 1527
rect 23446 1497 23464 1517
rect 23484 1497 23495 1517
rect 23446 1485 23495 1497
rect 24280 1525 24329 1537
rect 24280 1505 24291 1525
rect 24311 1505 24329 1525
rect 24280 1495 24329 1505
rect 24379 1521 24423 1537
rect 24379 1501 24394 1521
rect 24414 1501 24423 1521
rect 24379 1495 24423 1501
rect 24493 1521 24537 1537
rect 24493 1501 24502 1521
rect 24522 1501 24537 1521
rect 24493 1495 24537 1501
rect 24587 1525 24636 1537
rect 24587 1505 24605 1525
rect 24625 1505 24636 1525
rect 24587 1495 24636 1505
rect 24711 1521 24755 1537
rect 24711 1501 24720 1521
rect 24740 1501 24755 1521
rect 24711 1495 24755 1501
rect 24805 1525 24854 1537
rect 24805 1505 24823 1525
rect 24843 1505 24854 1525
rect 24805 1495 24854 1505
rect 27298 1529 27347 1539
rect 27298 1509 27309 1529
rect 27329 1509 27347 1529
rect 13919 1284 13937 1304
rect 13957 1284 13968 1304
rect 13919 1272 13968 1284
rect 27298 1497 27347 1509
rect 27397 1533 27441 1539
rect 27397 1513 27412 1533
rect 27432 1513 27441 1533
rect 27397 1497 27441 1513
rect 27516 1529 27565 1539
rect 27516 1509 27527 1529
rect 27547 1509 27565 1529
rect 27516 1497 27565 1509
rect 27615 1533 27659 1539
rect 27615 1513 27630 1533
rect 27650 1513 27659 1533
rect 27615 1497 27659 1513
rect 27729 1533 27773 1539
rect 27729 1513 27738 1533
rect 27758 1513 27773 1533
rect 27729 1497 27773 1513
rect 27823 1529 27872 1539
rect 27823 1509 27841 1529
rect 27861 1509 27872 1529
rect 27823 1497 27872 1509
rect 28657 1537 28706 1549
rect 28657 1517 28668 1537
rect 28688 1517 28706 1537
rect 28657 1507 28706 1517
rect 28756 1533 28800 1549
rect 28756 1513 28771 1533
rect 28791 1513 28800 1533
rect 28756 1507 28800 1513
rect 28870 1533 28914 1549
rect 28870 1513 28879 1533
rect 28899 1513 28914 1533
rect 28870 1507 28914 1513
rect 28964 1537 29013 1549
rect 28964 1517 28982 1537
rect 29002 1517 29013 1537
rect 28964 1507 29013 1517
rect 29088 1533 29132 1549
rect 29088 1513 29097 1533
rect 29117 1513 29132 1533
rect 29088 1507 29132 1513
rect 29182 1537 29231 1549
rect 29182 1517 29200 1537
rect 29220 1517 29231 1537
rect 29182 1507 29231 1517
rect 31662 1542 31711 1552
rect 31662 1522 31673 1542
rect 31693 1522 31711 1542
rect 20714 1328 20763 1340
rect 20714 1308 20725 1328
rect 20745 1308 20763 1328
rect 17660 1278 17709 1288
rect 17660 1258 17671 1278
rect 17691 1258 17709 1278
rect 17660 1246 17709 1258
rect 17759 1282 17803 1288
rect 17759 1262 17774 1282
rect 17794 1262 17803 1282
rect 17759 1246 17803 1262
rect 17878 1278 17927 1288
rect 17878 1258 17889 1278
rect 17909 1258 17927 1278
rect 17878 1246 17927 1258
rect 17977 1282 18021 1288
rect 17977 1262 17992 1282
rect 18012 1262 18021 1282
rect 17977 1246 18021 1262
rect 18091 1282 18135 1288
rect 18091 1262 18100 1282
rect 18120 1262 18135 1282
rect 18091 1246 18135 1262
rect 18185 1278 18234 1288
rect 20714 1298 20763 1308
rect 20813 1324 20857 1340
rect 20813 1304 20828 1324
rect 20848 1304 20857 1324
rect 20813 1298 20857 1304
rect 20927 1324 20971 1340
rect 20927 1304 20936 1324
rect 20956 1304 20971 1324
rect 20927 1298 20971 1304
rect 21021 1328 21070 1340
rect 21021 1308 21039 1328
rect 21059 1308 21070 1328
rect 21021 1298 21070 1308
rect 21145 1324 21189 1340
rect 21145 1304 21154 1324
rect 21174 1304 21189 1324
rect 21145 1298 21189 1304
rect 21239 1328 21288 1340
rect 21239 1308 21257 1328
rect 21277 1308 21288 1328
rect 21239 1298 21288 1308
rect 18185 1258 18203 1278
rect 18223 1258 18234 1278
rect 18185 1246 18234 1258
rect 31662 1510 31711 1522
rect 31761 1546 31805 1552
rect 31761 1526 31776 1546
rect 31796 1526 31805 1546
rect 31761 1510 31805 1526
rect 31880 1542 31929 1552
rect 31880 1522 31891 1542
rect 31911 1522 31929 1542
rect 31880 1510 31929 1522
rect 31979 1546 32023 1552
rect 31979 1526 31994 1546
rect 32014 1526 32023 1546
rect 31979 1510 32023 1526
rect 32093 1546 32137 1552
rect 32093 1526 32102 1546
rect 32122 1526 32137 1546
rect 32093 1510 32137 1526
rect 32187 1542 32236 1552
rect 32187 1522 32205 1542
rect 32225 1522 32236 1542
rect 32187 1510 32236 1522
rect 33021 1550 33070 1562
rect 33021 1530 33032 1550
rect 33052 1530 33070 1550
rect 33021 1520 33070 1530
rect 33120 1546 33164 1562
rect 33120 1526 33135 1546
rect 33155 1526 33164 1546
rect 33120 1520 33164 1526
rect 33234 1546 33278 1562
rect 33234 1526 33243 1546
rect 33263 1526 33278 1546
rect 33234 1520 33278 1526
rect 33328 1550 33377 1562
rect 33328 1530 33346 1550
rect 33366 1530 33377 1550
rect 33328 1520 33377 1530
rect 33452 1546 33496 1562
rect 33452 1526 33461 1546
rect 33481 1526 33496 1546
rect 33452 1520 33496 1526
rect 33546 1550 33595 1562
rect 33546 1530 33564 1550
rect 33584 1530 33595 1550
rect 33546 1520 33595 1530
rect 25078 1341 25127 1353
rect 25078 1321 25089 1341
rect 25109 1321 25127 1341
rect 22024 1291 22073 1301
rect 22024 1271 22035 1291
rect 22055 1271 22073 1291
rect 22024 1259 22073 1271
rect 22123 1295 22167 1301
rect 22123 1275 22138 1295
rect 22158 1275 22167 1295
rect 22123 1259 22167 1275
rect 22242 1291 22291 1301
rect 22242 1271 22253 1291
rect 22273 1271 22291 1291
rect 22242 1259 22291 1271
rect 22341 1295 22385 1301
rect 22341 1275 22356 1295
rect 22376 1275 22385 1295
rect 22341 1259 22385 1275
rect 22455 1295 22499 1301
rect 22455 1275 22464 1295
rect 22484 1275 22499 1295
rect 22455 1259 22499 1275
rect 22549 1291 22598 1301
rect 25078 1311 25127 1321
rect 25177 1337 25221 1353
rect 25177 1317 25192 1337
rect 25212 1317 25221 1337
rect 25177 1311 25221 1317
rect 25291 1337 25335 1353
rect 25291 1317 25300 1337
rect 25320 1317 25335 1337
rect 25291 1311 25335 1317
rect 25385 1341 25434 1353
rect 25385 1321 25403 1341
rect 25423 1321 25434 1341
rect 25385 1311 25434 1321
rect 25509 1337 25553 1353
rect 25509 1317 25518 1337
rect 25538 1317 25553 1337
rect 25509 1311 25553 1317
rect 25603 1341 25652 1353
rect 25603 1321 25621 1341
rect 25641 1321 25652 1341
rect 25603 1311 25652 1321
rect 22549 1271 22567 1291
rect 22587 1271 22598 1291
rect 22549 1259 22598 1271
rect 1087 1082 1136 1092
rect 1087 1062 1098 1082
rect 1118 1062 1136 1082
rect 1087 1050 1136 1062
rect 1186 1086 1230 1092
rect 1186 1066 1201 1086
rect 1221 1066 1230 1086
rect 1186 1050 1230 1066
rect 1305 1082 1354 1092
rect 1305 1062 1316 1082
rect 1336 1062 1354 1082
rect 1305 1050 1354 1062
rect 1404 1086 1448 1092
rect 1404 1066 1419 1086
rect 1439 1066 1448 1086
rect 1404 1050 1448 1066
rect 1518 1086 1562 1092
rect 1518 1066 1527 1086
rect 1547 1066 1562 1086
rect 1518 1050 1562 1066
rect 1612 1082 1661 1092
rect 1612 1062 1630 1082
rect 1650 1062 1661 1082
rect 1612 1050 1661 1062
rect 5451 1095 5500 1105
rect 5451 1075 5462 1095
rect 5482 1075 5500 1095
rect 5451 1063 5500 1075
rect 5550 1099 5594 1105
rect 5550 1079 5565 1099
rect 5585 1079 5594 1099
rect 5550 1063 5594 1079
rect 5669 1095 5718 1105
rect 5669 1075 5680 1095
rect 5700 1075 5718 1095
rect 5669 1063 5718 1075
rect 5768 1099 5812 1105
rect 5768 1079 5783 1099
rect 5803 1079 5812 1099
rect 5768 1063 5812 1079
rect 5882 1099 5926 1105
rect 5882 1079 5891 1099
rect 5911 1079 5926 1099
rect 5882 1063 5926 1079
rect 5976 1095 6025 1105
rect 5976 1075 5994 1095
rect 6014 1075 6025 1095
rect 5976 1063 6025 1075
rect 9828 1107 9877 1117
rect 9828 1087 9839 1107
rect 9859 1087 9877 1107
rect 9828 1075 9877 1087
rect 9927 1111 9971 1117
rect 9927 1091 9942 1111
rect 9962 1091 9971 1111
rect 9927 1075 9971 1091
rect 10046 1107 10095 1117
rect 10046 1087 10057 1107
rect 10077 1087 10095 1107
rect 10046 1075 10095 1087
rect 10145 1111 10189 1117
rect 10145 1091 10160 1111
rect 10180 1091 10189 1111
rect 10145 1075 10189 1091
rect 10259 1111 10303 1117
rect 10259 1091 10268 1111
rect 10288 1091 10303 1111
rect 10259 1075 10303 1091
rect 10353 1107 10402 1117
rect 10353 1087 10371 1107
rect 10391 1087 10402 1107
rect 10353 1075 10402 1087
rect 14192 1120 14241 1130
rect 14192 1100 14203 1120
rect 14223 1100 14241 1120
rect 290 854 339 864
rect 290 834 301 854
rect 321 834 339 854
rect 290 822 339 834
rect 389 858 433 864
rect 389 838 404 858
rect 424 838 433 858
rect 389 822 433 838
rect 508 854 557 864
rect 508 834 519 854
rect 539 834 557 854
rect 508 822 557 834
rect 607 858 651 864
rect 607 838 622 858
rect 642 838 651 858
rect 607 822 651 838
rect 721 858 765 864
rect 721 838 730 858
rect 750 838 765 858
rect 721 822 765 838
rect 815 854 864 864
rect 815 834 833 854
rect 853 834 864 854
rect 14192 1088 14241 1100
rect 14291 1124 14335 1130
rect 14291 1104 14306 1124
rect 14326 1104 14335 1124
rect 14291 1088 14335 1104
rect 14410 1120 14459 1130
rect 14410 1100 14421 1120
rect 14441 1100 14459 1120
rect 14410 1088 14459 1100
rect 14509 1124 14553 1130
rect 14509 1104 14524 1124
rect 14544 1104 14553 1124
rect 14509 1088 14553 1104
rect 14623 1124 14667 1130
rect 14623 1104 14632 1124
rect 14652 1104 14667 1124
rect 14623 1088 14667 1104
rect 14717 1120 14766 1130
rect 14717 1100 14735 1120
rect 14755 1100 14766 1120
rect 14717 1088 14766 1100
rect 29455 1353 29504 1365
rect 29455 1333 29466 1353
rect 29486 1333 29504 1353
rect 26401 1303 26450 1313
rect 26401 1283 26412 1303
rect 26432 1283 26450 1303
rect 26401 1271 26450 1283
rect 26500 1307 26544 1313
rect 26500 1287 26515 1307
rect 26535 1287 26544 1307
rect 26500 1271 26544 1287
rect 26619 1303 26668 1313
rect 26619 1283 26630 1303
rect 26650 1283 26668 1303
rect 26619 1271 26668 1283
rect 26718 1307 26762 1313
rect 26718 1287 26733 1307
rect 26753 1287 26762 1307
rect 26718 1271 26762 1287
rect 26832 1307 26876 1313
rect 26832 1287 26841 1307
rect 26861 1287 26876 1307
rect 26832 1271 26876 1287
rect 26926 1303 26975 1313
rect 29455 1323 29504 1333
rect 29554 1349 29598 1365
rect 29554 1329 29569 1349
rect 29589 1329 29598 1349
rect 29554 1323 29598 1329
rect 29668 1349 29712 1365
rect 29668 1329 29677 1349
rect 29697 1329 29712 1349
rect 29668 1323 29712 1329
rect 29762 1353 29811 1365
rect 29762 1333 29780 1353
rect 29800 1333 29811 1353
rect 29762 1323 29811 1333
rect 29886 1349 29930 1365
rect 29886 1329 29895 1349
rect 29915 1329 29930 1349
rect 29886 1323 29930 1329
rect 29980 1353 30029 1365
rect 29980 1333 29998 1353
rect 30018 1333 30029 1353
rect 29980 1323 30029 1333
rect 26926 1283 26944 1303
rect 26964 1283 26975 1303
rect 26926 1271 26975 1283
rect 33819 1366 33868 1378
rect 33819 1346 33830 1366
rect 33850 1346 33868 1366
rect 30765 1316 30814 1326
rect 30765 1296 30776 1316
rect 30796 1296 30814 1316
rect 30765 1284 30814 1296
rect 30864 1320 30908 1326
rect 30864 1300 30879 1320
rect 30899 1300 30908 1320
rect 30864 1284 30908 1300
rect 30983 1316 31032 1326
rect 30983 1296 30994 1316
rect 31014 1296 31032 1316
rect 30983 1284 31032 1296
rect 31082 1320 31126 1326
rect 31082 1300 31097 1320
rect 31117 1300 31126 1320
rect 31082 1284 31126 1300
rect 31196 1320 31240 1326
rect 31196 1300 31205 1320
rect 31225 1300 31240 1320
rect 31196 1284 31240 1300
rect 31290 1316 31339 1326
rect 33819 1336 33868 1346
rect 33918 1362 33962 1378
rect 33918 1342 33933 1362
rect 33953 1342 33962 1362
rect 33918 1336 33962 1342
rect 34032 1362 34076 1378
rect 34032 1342 34041 1362
rect 34061 1342 34076 1362
rect 34032 1336 34076 1342
rect 34126 1366 34175 1378
rect 34126 1346 34144 1366
rect 34164 1346 34175 1366
rect 34126 1336 34175 1346
rect 34250 1362 34294 1378
rect 34250 1342 34259 1362
rect 34279 1342 34294 1362
rect 34250 1336 34294 1342
rect 34344 1366 34393 1378
rect 34344 1346 34362 1366
rect 34382 1346 34393 1366
rect 34344 1336 34393 1346
rect 31290 1296 31308 1316
rect 31328 1296 31339 1316
rect 31290 1284 31339 1296
rect 815 822 864 834
rect 4654 867 4703 877
rect 4654 847 4665 867
rect 4685 847 4703 867
rect 4654 835 4703 847
rect 4753 871 4797 877
rect 4753 851 4768 871
rect 4788 851 4797 871
rect 4753 835 4797 851
rect 4872 867 4921 877
rect 4872 847 4883 867
rect 4903 847 4921 867
rect 4872 835 4921 847
rect 4971 871 5015 877
rect 4971 851 4986 871
rect 5006 851 5015 871
rect 4971 835 5015 851
rect 5085 871 5129 877
rect 5085 851 5094 871
rect 5114 851 5129 871
rect 5085 835 5129 851
rect 5179 867 5228 877
rect 5179 847 5197 867
rect 5217 847 5228 867
rect 18458 1094 18507 1104
rect 18458 1074 18469 1094
rect 18489 1074 18507 1094
rect 18458 1062 18507 1074
rect 18557 1098 18601 1104
rect 18557 1078 18572 1098
rect 18592 1078 18601 1098
rect 18557 1062 18601 1078
rect 18676 1094 18725 1104
rect 18676 1074 18687 1094
rect 18707 1074 18725 1094
rect 18676 1062 18725 1074
rect 18775 1098 18819 1104
rect 18775 1078 18790 1098
rect 18810 1078 18819 1098
rect 18775 1062 18819 1078
rect 18889 1098 18933 1104
rect 18889 1078 18898 1098
rect 18918 1078 18933 1098
rect 18889 1062 18933 1078
rect 18983 1094 19032 1104
rect 18983 1074 19001 1094
rect 19021 1074 19032 1094
rect 18983 1062 19032 1074
rect 22822 1107 22871 1117
rect 22822 1087 22833 1107
rect 22853 1087 22871 1107
rect 5179 835 5228 847
rect 9031 879 9080 889
rect 9031 859 9042 879
rect 9062 859 9080 879
rect 9031 847 9080 859
rect 9130 883 9174 889
rect 9130 863 9145 883
rect 9165 863 9174 883
rect 9130 847 9174 863
rect 9249 879 9298 889
rect 9249 859 9260 879
rect 9280 859 9298 879
rect 9249 847 9298 859
rect 9348 883 9392 889
rect 9348 863 9363 883
rect 9383 863 9392 883
rect 9348 847 9392 863
rect 9462 883 9506 889
rect 9462 863 9471 883
rect 9491 863 9506 883
rect 9462 847 9506 863
rect 9556 879 9605 889
rect 9556 859 9574 879
rect 9594 859 9605 879
rect 22822 1075 22871 1087
rect 22921 1111 22965 1117
rect 22921 1091 22936 1111
rect 22956 1091 22965 1111
rect 22921 1075 22965 1091
rect 23040 1107 23089 1117
rect 23040 1087 23051 1107
rect 23071 1087 23089 1107
rect 23040 1075 23089 1087
rect 23139 1111 23183 1117
rect 23139 1091 23154 1111
rect 23174 1091 23183 1111
rect 23139 1075 23183 1091
rect 23253 1111 23297 1117
rect 23253 1091 23262 1111
rect 23282 1091 23297 1111
rect 23253 1075 23297 1091
rect 23347 1107 23396 1117
rect 23347 1087 23365 1107
rect 23385 1087 23396 1107
rect 23347 1075 23396 1087
rect 27199 1119 27248 1129
rect 27199 1099 27210 1119
rect 27230 1099 27248 1119
rect 9556 847 9605 859
rect 13395 892 13444 902
rect 13395 872 13406 892
rect 13426 872 13444 892
rect 13395 860 13444 872
rect 13494 896 13538 902
rect 13494 876 13509 896
rect 13529 876 13538 896
rect 13494 860 13538 876
rect 13613 892 13662 902
rect 13613 872 13624 892
rect 13644 872 13662 892
rect 13613 860 13662 872
rect 13712 896 13756 902
rect 13712 876 13727 896
rect 13747 876 13756 896
rect 13712 860 13756 876
rect 13826 896 13870 902
rect 13826 876 13835 896
rect 13855 876 13870 896
rect 13826 860 13870 876
rect 13920 892 13969 902
rect 13920 872 13938 892
rect 13958 872 13969 892
rect 13920 860 13969 872
rect 27199 1087 27248 1099
rect 27298 1123 27342 1129
rect 27298 1103 27313 1123
rect 27333 1103 27342 1123
rect 27298 1087 27342 1103
rect 27417 1119 27466 1129
rect 27417 1099 27428 1119
rect 27448 1099 27466 1119
rect 27417 1087 27466 1099
rect 27516 1123 27560 1129
rect 27516 1103 27531 1123
rect 27551 1103 27560 1123
rect 27516 1087 27560 1103
rect 27630 1123 27674 1129
rect 27630 1103 27639 1123
rect 27659 1103 27674 1123
rect 27630 1087 27674 1103
rect 27724 1119 27773 1129
rect 27724 1099 27742 1119
rect 27762 1099 27773 1119
rect 27724 1087 27773 1099
rect 31563 1132 31612 1142
rect 31563 1112 31574 1132
rect 31594 1112 31612 1132
rect 17661 866 17710 876
rect 17661 846 17672 866
rect 17692 846 17710 866
rect 17661 834 17710 846
rect 17760 870 17804 876
rect 17760 850 17775 870
rect 17795 850 17804 870
rect 17760 834 17804 850
rect 17879 866 17928 876
rect 17879 846 17890 866
rect 17910 846 17928 866
rect 17879 834 17928 846
rect 17978 870 18022 876
rect 17978 850 17993 870
rect 18013 850 18022 870
rect 17978 834 18022 850
rect 18092 870 18136 876
rect 18092 850 18101 870
rect 18121 850 18136 870
rect 18092 834 18136 850
rect 18186 866 18235 876
rect 18186 846 18204 866
rect 18224 846 18235 866
rect 31563 1100 31612 1112
rect 31662 1136 31706 1142
rect 31662 1116 31677 1136
rect 31697 1116 31706 1136
rect 31662 1100 31706 1116
rect 31781 1132 31830 1142
rect 31781 1112 31792 1132
rect 31812 1112 31830 1132
rect 31781 1100 31830 1112
rect 31880 1136 31924 1142
rect 31880 1116 31895 1136
rect 31915 1116 31924 1136
rect 31880 1100 31924 1116
rect 31994 1136 32038 1142
rect 31994 1116 32003 1136
rect 32023 1116 32038 1136
rect 31994 1100 32038 1116
rect 32088 1132 32137 1142
rect 32088 1112 32106 1132
rect 32126 1112 32137 1132
rect 32088 1100 32137 1112
rect 18186 834 18235 846
rect 22025 879 22074 889
rect 22025 859 22036 879
rect 22056 859 22074 879
rect 22025 847 22074 859
rect 22124 883 22168 889
rect 22124 863 22139 883
rect 22159 863 22168 883
rect 22124 847 22168 863
rect 22243 879 22292 889
rect 22243 859 22254 879
rect 22274 859 22292 879
rect 22243 847 22292 859
rect 22342 883 22386 889
rect 22342 863 22357 883
rect 22377 863 22386 883
rect 22342 847 22386 863
rect 22456 883 22500 889
rect 22456 863 22465 883
rect 22485 863 22500 883
rect 22456 847 22500 863
rect 22550 879 22599 889
rect 22550 859 22568 879
rect 22588 859 22599 879
rect 22550 847 22599 859
rect 26402 891 26451 901
rect 26402 871 26413 891
rect 26433 871 26451 891
rect 26402 859 26451 871
rect 26501 895 26545 901
rect 26501 875 26516 895
rect 26536 875 26545 895
rect 26501 859 26545 875
rect 26620 891 26669 901
rect 26620 871 26631 891
rect 26651 871 26669 891
rect 26620 859 26669 871
rect 26719 895 26763 901
rect 26719 875 26734 895
rect 26754 875 26763 895
rect 26719 859 26763 875
rect 26833 895 26877 901
rect 26833 875 26842 895
rect 26862 875 26877 895
rect 26833 859 26877 875
rect 26927 891 26976 901
rect 26927 871 26945 891
rect 26965 871 26976 891
rect 26927 859 26976 871
rect 30766 904 30815 914
rect 30766 884 30777 904
rect 30797 884 30815 904
rect 30766 872 30815 884
rect 30865 908 30909 914
rect 30865 888 30880 908
rect 30900 888 30909 908
rect 30865 872 30909 888
rect 30984 904 31033 914
rect 30984 884 30995 904
rect 31015 884 31033 904
rect 30984 872 31033 884
rect 31083 908 31127 914
rect 31083 888 31098 908
rect 31118 888 31127 908
rect 31083 872 31127 888
rect 31197 908 31241 914
rect 31197 888 31206 908
rect 31226 888 31241 908
rect 31197 872 31241 888
rect 31291 904 31340 914
rect 31291 884 31309 904
rect 31329 884 31340 904
rect 31291 872 31340 884
rect 5867 291 5916 301
rect 1503 278 1552 288
rect 1503 258 1514 278
rect 1534 258 1552 278
rect 1503 246 1552 258
rect 1602 282 1646 288
rect 1602 262 1617 282
rect 1637 262 1646 282
rect 1602 246 1646 262
rect 1721 278 1770 288
rect 1721 258 1732 278
rect 1752 258 1770 278
rect 1721 246 1770 258
rect 1820 282 1864 288
rect 1820 262 1835 282
rect 1855 262 1864 282
rect 1820 246 1864 262
rect 1934 282 1978 288
rect 1934 262 1943 282
rect 1963 262 1978 282
rect 1934 246 1978 262
rect 2028 278 2077 288
rect 2028 258 2046 278
rect 2066 258 2077 278
rect 2028 246 2077 258
rect 5867 271 5878 291
rect 5898 271 5916 291
rect 5867 259 5916 271
rect 5966 295 6010 301
rect 5966 275 5981 295
rect 6001 275 6010 295
rect 5966 259 6010 275
rect 6085 291 6134 301
rect 6085 271 6096 291
rect 6116 271 6134 291
rect 6085 259 6134 271
rect 6184 295 6228 301
rect 6184 275 6199 295
rect 6219 275 6228 295
rect 6184 259 6228 275
rect 6298 295 6342 301
rect 6298 275 6307 295
rect 6327 275 6342 295
rect 6298 259 6342 275
rect 6392 291 6441 301
rect 6392 271 6410 291
rect 6430 271 6441 291
rect 6392 259 6441 271
rect 14608 316 14657 326
rect 10244 303 10293 313
rect 10244 283 10255 303
rect 10275 283 10293 303
rect 10244 271 10293 283
rect 10343 307 10387 313
rect 10343 287 10358 307
rect 10378 287 10387 307
rect 10343 271 10387 287
rect 10462 303 10511 313
rect 10462 283 10473 303
rect 10493 283 10511 303
rect 10462 271 10511 283
rect 10561 307 10605 313
rect 10561 287 10576 307
rect 10596 287 10605 307
rect 10561 271 10605 287
rect 10675 307 10719 313
rect 10675 287 10684 307
rect 10704 287 10719 307
rect 10675 271 10719 287
rect 10769 303 10818 313
rect 10769 283 10787 303
rect 10807 283 10818 303
rect 10769 271 10818 283
rect 14608 296 14619 316
rect 14639 296 14657 316
rect 14608 284 14657 296
rect 14707 320 14751 326
rect 14707 300 14722 320
rect 14742 300 14751 320
rect 14707 284 14751 300
rect 14826 316 14875 326
rect 14826 296 14837 316
rect 14857 296 14875 316
rect 14826 284 14875 296
rect 14925 320 14969 326
rect 14925 300 14940 320
rect 14960 300 14969 320
rect 14925 284 14969 300
rect 15039 320 15083 326
rect 15039 300 15048 320
rect 15068 300 15083 320
rect 15039 284 15083 300
rect 15133 316 15182 326
rect 15133 296 15151 316
rect 15171 296 15182 316
rect 15133 284 15182 296
rect 23238 303 23287 313
rect 18874 290 18923 300
rect 18874 270 18885 290
rect 18905 270 18923 290
rect 18874 258 18923 270
rect 18973 294 19017 300
rect 18973 274 18988 294
rect 19008 274 19017 294
rect 18973 258 19017 274
rect 19092 290 19141 300
rect 19092 270 19103 290
rect 19123 270 19141 290
rect 19092 258 19141 270
rect 19191 294 19235 300
rect 19191 274 19206 294
rect 19226 274 19235 294
rect 19191 258 19235 274
rect 19305 294 19349 300
rect 19305 274 19314 294
rect 19334 274 19349 294
rect 19305 258 19349 274
rect 19399 290 19448 300
rect 19399 270 19417 290
rect 19437 270 19448 290
rect 19399 258 19448 270
rect 8440 228 8489 238
rect 3992 204 4041 214
rect 3992 184 4003 204
rect 4023 184 4041 204
rect 3992 172 4041 184
rect 4091 208 4135 214
rect 4091 188 4106 208
rect 4126 188 4135 208
rect 4091 172 4135 188
rect 4210 204 4259 214
rect 4210 184 4221 204
rect 4241 184 4259 204
rect 4210 172 4259 184
rect 4309 208 4353 214
rect 4309 188 4324 208
rect 4344 188 4353 208
rect 4309 172 4353 188
rect 4423 208 4467 214
rect 4423 188 4432 208
rect 4452 188 4467 208
rect 4423 172 4467 188
rect 4517 204 4566 214
rect 4517 184 4535 204
rect 4555 184 4566 204
rect 8440 208 8451 228
rect 8471 208 8489 228
rect 8440 196 8489 208
rect 8539 232 8583 238
rect 8539 212 8554 232
rect 8574 212 8583 232
rect 8539 196 8583 212
rect 8658 228 8707 238
rect 8658 208 8669 228
rect 8689 208 8707 228
rect 8658 196 8707 208
rect 8757 232 8801 238
rect 8757 212 8772 232
rect 8792 212 8801 232
rect 8757 196 8801 212
rect 8871 232 8915 238
rect 8871 212 8880 232
rect 8900 212 8915 232
rect 8871 196 8915 212
rect 8965 228 9014 238
rect 8965 208 8983 228
rect 9003 208 9014 228
rect 8965 196 9014 208
rect 12733 229 12782 239
rect 12733 209 12744 229
rect 12764 209 12782 229
rect 12733 197 12782 209
rect 12832 233 12876 239
rect 12832 213 12847 233
rect 12867 213 12876 233
rect 12832 197 12876 213
rect 12951 229 13000 239
rect 12951 209 12962 229
rect 12982 209 13000 229
rect 12951 197 13000 209
rect 13050 233 13094 239
rect 13050 213 13065 233
rect 13085 213 13094 233
rect 13050 197 13094 213
rect 13164 233 13208 239
rect 13164 213 13173 233
rect 13193 213 13208 233
rect 13164 197 13208 213
rect 13258 229 13307 239
rect 13258 209 13276 229
rect 13296 209 13307 229
rect 13258 197 13307 209
rect 4517 172 4566 184
rect 23238 283 23249 303
rect 23269 283 23287 303
rect 23238 271 23287 283
rect 23337 307 23381 313
rect 23337 287 23352 307
rect 23372 287 23381 307
rect 23337 271 23381 287
rect 23456 303 23505 313
rect 23456 283 23467 303
rect 23487 283 23505 303
rect 23456 271 23505 283
rect 23555 307 23599 313
rect 23555 287 23570 307
rect 23590 287 23599 307
rect 23555 271 23599 287
rect 23669 307 23713 313
rect 23669 287 23678 307
rect 23698 287 23713 307
rect 23669 271 23713 287
rect 23763 303 23812 313
rect 23763 283 23781 303
rect 23801 283 23812 303
rect 23763 271 23812 283
rect 31979 328 32028 338
rect 27615 315 27664 325
rect 27615 295 27626 315
rect 27646 295 27664 315
rect 27615 283 27664 295
rect 27714 319 27758 325
rect 27714 299 27729 319
rect 27749 299 27758 319
rect 27714 283 27758 299
rect 27833 315 27882 325
rect 27833 295 27844 315
rect 27864 295 27882 315
rect 27833 283 27882 295
rect 27932 319 27976 325
rect 27932 299 27947 319
rect 27967 299 27976 319
rect 27932 283 27976 299
rect 28046 319 28090 325
rect 28046 299 28055 319
rect 28075 299 28090 319
rect 28046 283 28090 299
rect 28140 315 28189 325
rect 28140 295 28158 315
rect 28178 295 28189 315
rect 28140 283 28189 295
rect 31979 308 31990 328
rect 32010 308 32028 328
rect 31979 296 32028 308
rect 32078 332 32122 338
rect 32078 312 32093 332
rect 32113 312 32122 332
rect 32078 296 32122 312
rect 32197 328 32246 338
rect 32197 308 32208 328
rect 32228 308 32246 328
rect 32197 296 32246 308
rect 32296 332 32340 338
rect 32296 312 32311 332
rect 32331 312 32340 332
rect 32296 296 32340 312
rect 32410 332 32454 338
rect 32410 312 32419 332
rect 32439 312 32454 332
rect 32410 296 32454 312
rect 32504 328 32553 338
rect 32504 308 32522 328
rect 32542 308 32553 328
rect 32504 296 32553 308
rect 25811 240 25860 250
rect 21363 216 21412 226
rect 21363 196 21374 216
rect 21394 196 21412 216
rect 21363 184 21412 196
rect 21462 220 21506 226
rect 21462 200 21477 220
rect 21497 200 21506 220
rect 21462 184 21506 200
rect 21581 216 21630 226
rect 21581 196 21592 216
rect 21612 196 21630 216
rect 21581 184 21630 196
rect 21680 220 21724 226
rect 21680 200 21695 220
rect 21715 200 21724 220
rect 21680 184 21724 200
rect 21794 220 21838 226
rect 21794 200 21803 220
rect 21823 200 21838 220
rect 21794 184 21838 200
rect 21888 216 21937 226
rect 21888 196 21906 216
rect 21926 196 21937 216
rect 25811 220 25822 240
rect 25842 220 25860 240
rect 25811 208 25860 220
rect 25910 244 25954 250
rect 25910 224 25925 244
rect 25945 224 25954 244
rect 25910 208 25954 224
rect 26029 240 26078 250
rect 26029 220 26040 240
rect 26060 220 26078 240
rect 26029 208 26078 220
rect 26128 244 26172 250
rect 26128 224 26143 244
rect 26163 224 26172 244
rect 26128 208 26172 224
rect 26242 244 26286 250
rect 26242 224 26251 244
rect 26271 224 26286 244
rect 26242 208 26286 224
rect 26336 240 26385 250
rect 26336 220 26354 240
rect 26374 220 26385 240
rect 26336 208 26385 220
rect 30104 241 30153 251
rect 30104 221 30115 241
rect 30135 221 30153 241
rect 30104 209 30153 221
rect 30203 245 30247 251
rect 30203 225 30218 245
rect 30238 225 30247 245
rect 30203 209 30247 225
rect 30322 241 30371 251
rect 30322 221 30333 241
rect 30353 221 30371 241
rect 30322 209 30371 221
rect 30421 245 30465 251
rect 30421 225 30436 245
rect 30456 225 30465 245
rect 30421 209 30465 225
rect 30535 245 30579 251
rect 30535 225 30544 245
rect 30564 225 30579 245
rect 30535 209 30579 225
rect 30629 241 30678 251
rect 30629 221 30647 241
rect 30667 221 30678 241
rect 30629 209 30678 221
rect 21888 184 21937 196
rect 16930 165 16979 175
rect 16930 145 16941 165
rect 16961 145 16979 165
rect 16930 133 16979 145
rect 17029 169 17073 175
rect 17029 149 17044 169
rect 17064 149 17073 169
rect 17029 133 17073 149
rect 17148 165 17197 175
rect 17148 145 17159 165
rect 17179 145 17197 165
rect 17148 133 17197 145
rect 17247 169 17291 175
rect 17247 149 17262 169
rect 17282 149 17291 169
rect 17247 133 17291 149
rect 17361 169 17405 175
rect 17361 149 17370 169
rect 17390 149 17405 169
rect 17361 133 17405 149
rect 17455 165 17504 175
rect 17455 145 17473 165
rect 17493 145 17504 165
rect 17455 133 17504 145
<< pdiff >>
rect 3474 8705 3518 8747
rect 3474 8685 3486 8705
rect 3506 8685 3518 8705
rect 3474 8678 3518 8685
rect 3473 8647 3518 8678
rect 3568 8705 3610 8747
rect 3568 8685 3582 8705
rect 3602 8685 3610 8705
rect 3568 8647 3610 8685
rect 3684 8705 3726 8747
rect 3684 8685 3692 8705
rect 3712 8685 3726 8705
rect 3684 8647 3726 8685
rect 3776 8705 3820 8747
rect 3776 8685 3788 8705
rect 3808 8685 3820 8705
rect 3776 8647 3820 8685
rect 3902 8705 3944 8747
rect 3902 8685 3910 8705
rect 3930 8685 3944 8705
rect 3902 8647 3944 8685
rect 3994 8705 4038 8747
rect 3994 8685 4006 8705
rect 4026 8685 4038 8705
rect 3994 8647 4038 8685
rect 7838 8718 7882 8760
rect 7838 8698 7850 8718
rect 7870 8698 7882 8718
rect 7838 8691 7882 8698
rect 7837 8660 7882 8691
rect 7932 8718 7974 8760
rect 7932 8698 7946 8718
rect 7966 8698 7974 8718
rect 7932 8660 7974 8698
rect 8048 8718 8090 8760
rect 8048 8698 8056 8718
rect 8076 8698 8090 8718
rect 8048 8660 8090 8698
rect 8140 8718 8184 8760
rect 8140 8698 8152 8718
rect 8172 8698 8184 8718
rect 8140 8660 8184 8698
rect 8266 8718 8308 8760
rect 8266 8698 8274 8718
rect 8294 8698 8308 8718
rect 8266 8660 8308 8698
rect 8358 8718 8402 8760
rect 8358 8698 8370 8718
rect 8390 8698 8402 8718
rect 8358 8660 8402 8698
rect 12215 8730 12259 8772
rect 12215 8710 12227 8730
rect 12247 8710 12259 8730
rect 12215 8703 12259 8710
rect 12214 8672 12259 8703
rect 12309 8730 12351 8772
rect 12309 8710 12323 8730
rect 12343 8710 12351 8730
rect 12309 8672 12351 8710
rect 12425 8730 12467 8772
rect 12425 8710 12433 8730
rect 12453 8710 12467 8730
rect 12425 8672 12467 8710
rect 12517 8730 12561 8772
rect 12517 8710 12529 8730
rect 12549 8710 12561 8730
rect 12517 8672 12561 8710
rect 12643 8730 12685 8772
rect 12643 8710 12651 8730
rect 12671 8710 12685 8730
rect 12643 8672 12685 8710
rect 12735 8730 12779 8772
rect 12735 8710 12747 8730
rect 12767 8710 12779 8730
rect 12735 8672 12779 8710
rect 16579 8743 16623 8785
rect 16579 8723 16591 8743
rect 16611 8723 16623 8743
rect 16579 8716 16623 8723
rect 16578 8685 16623 8716
rect 16673 8743 16715 8785
rect 16673 8723 16687 8743
rect 16707 8723 16715 8743
rect 16673 8685 16715 8723
rect 16789 8743 16831 8785
rect 16789 8723 16797 8743
rect 16817 8723 16831 8743
rect 16789 8685 16831 8723
rect 16881 8743 16925 8785
rect 16881 8723 16893 8743
rect 16913 8723 16925 8743
rect 16881 8685 16925 8723
rect 17007 8743 17049 8785
rect 17007 8723 17015 8743
rect 17035 8723 17049 8743
rect 17007 8685 17049 8723
rect 17099 8743 17143 8785
rect 17099 8723 17111 8743
rect 17131 8723 17143 8743
rect 17099 8685 17143 8723
rect 20845 8717 20889 8759
rect 20845 8697 20857 8717
rect 20877 8697 20889 8717
rect 20845 8690 20889 8697
rect 20844 8659 20889 8690
rect 20939 8717 20981 8759
rect 20939 8697 20953 8717
rect 20973 8697 20981 8717
rect 20939 8659 20981 8697
rect 21055 8717 21097 8759
rect 21055 8697 21063 8717
rect 21083 8697 21097 8717
rect 21055 8659 21097 8697
rect 21147 8717 21191 8759
rect 21147 8697 21159 8717
rect 21179 8697 21191 8717
rect 21147 8659 21191 8697
rect 21273 8717 21315 8759
rect 21273 8697 21281 8717
rect 21301 8697 21315 8717
rect 21273 8659 21315 8697
rect 21365 8717 21409 8759
rect 21365 8697 21377 8717
rect 21397 8697 21409 8717
rect 21365 8659 21409 8697
rect 25209 8730 25253 8772
rect 25209 8710 25221 8730
rect 25241 8710 25253 8730
rect 25209 8703 25253 8710
rect 421 8541 465 8579
rect 421 8521 433 8541
rect 453 8521 465 8541
rect 421 8479 465 8521
rect 515 8541 557 8579
rect 515 8521 529 8541
rect 549 8521 557 8541
rect 515 8479 557 8521
rect 639 8541 683 8579
rect 639 8521 651 8541
rect 671 8521 683 8541
rect 639 8479 683 8521
rect 733 8541 775 8579
rect 733 8521 747 8541
rect 767 8521 775 8541
rect 733 8479 775 8521
rect 849 8541 891 8579
rect 849 8521 857 8541
rect 877 8521 891 8541
rect 849 8479 891 8521
rect 941 8548 986 8579
rect 941 8541 985 8548
rect 941 8521 953 8541
rect 973 8521 985 8541
rect 941 8479 985 8521
rect 4785 8554 4829 8592
rect 4785 8534 4797 8554
rect 4817 8534 4829 8554
rect 2677 8477 2721 8519
rect 2677 8457 2689 8477
rect 2709 8457 2721 8477
rect 2677 8450 2721 8457
rect 2676 8419 2721 8450
rect 2771 8477 2813 8519
rect 2771 8457 2785 8477
rect 2805 8457 2813 8477
rect 2771 8419 2813 8457
rect 2887 8477 2929 8519
rect 2887 8457 2895 8477
rect 2915 8457 2929 8477
rect 2887 8419 2929 8457
rect 2979 8477 3023 8519
rect 2979 8457 2991 8477
rect 3011 8457 3023 8477
rect 2979 8419 3023 8457
rect 3105 8477 3147 8519
rect 3105 8457 3113 8477
rect 3133 8457 3147 8477
rect 3105 8419 3147 8457
rect 3197 8477 3241 8519
rect 4785 8492 4829 8534
rect 4879 8554 4921 8592
rect 4879 8534 4893 8554
rect 4913 8534 4921 8554
rect 4879 8492 4921 8534
rect 5003 8554 5047 8592
rect 5003 8534 5015 8554
rect 5035 8534 5047 8554
rect 5003 8492 5047 8534
rect 5097 8554 5139 8592
rect 5097 8534 5111 8554
rect 5131 8534 5139 8554
rect 5097 8492 5139 8534
rect 5213 8554 5255 8592
rect 5213 8534 5221 8554
rect 5241 8534 5255 8554
rect 5213 8492 5255 8534
rect 5305 8561 5350 8592
rect 5305 8554 5349 8561
rect 5305 8534 5317 8554
rect 5337 8534 5349 8554
rect 5305 8492 5349 8534
rect 9162 8566 9206 8604
rect 9162 8546 9174 8566
rect 9194 8546 9206 8566
rect 3197 8457 3209 8477
rect 3229 8457 3241 8477
rect 3197 8419 3241 8457
rect 1219 8357 1263 8395
rect 1219 8337 1231 8357
rect 1251 8337 1263 8357
rect 1219 8295 1263 8337
rect 1313 8357 1355 8395
rect 1313 8337 1327 8357
rect 1347 8337 1355 8357
rect 1313 8295 1355 8337
rect 1437 8357 1481 8395
rect 1437 8337 1449 8357
rect 1469 8337 1481 8357
rect 1437 8295 1481 8337
rect 1531 8357 1573 8395
rect 1531 8337 1545 8357
rect 1565 8337 1573 8357
rect 1531 8295 1573 8337
rect 1647 8357 1689 8395
rect 1647 8337 1655 8357
rect 1675 8337 1689 8357
rect 1647 8295 1689 8337
rect 1739 8364 1784 8395
rect 1739 8357 1783 8364
rect 1739 8337 1751 8357
rect 1771 8337 1783 8357
rect 1739 8295 1783 8337
rect 7041 8490 7085 8532
rect 7041 8470 7053 8490
rect 7073 8470 7085 8490
rect 7041 8463 7085 8470
rect 7040 8432 7085 8463
rect 7135 8490 7177 8532
rect 7135 8470 7149 8490
rect 7169 8470 7177 8490
rect 7135 8432 7177 8470
rect 7251 8490 7293 8532
rect 7251 8470 7259 8490
rect 7279 8470 7293 8490
rect 7251 8432 7293 8470
rect 7343 8490 7387 8532
rect 7343 8470 7355 8490
rect 7375 8470 7387 8490
rect 7343 8432 7387 8470
rect 7469 8490 7511 8532
rect 7469 8470 7477 8490
rect 7497 8470 7511 8490
rect 7469 8432 7511 8470
rect 7561 8490 7605 8532
rect 9162 8504 9206 8546
rect 9256 8566 9298 8604
rect 9256 8546 9270 8566
rect 9290 8546 9298 8566
rect 9256 8504 9298 8546
rect 9380 8566 9424 8604
rect 9380 8546 9392 8566
rect 9412 8546 9424 8566
rect 9380 8504 9424 8546
rect 9474 8566 9516 8604
rect 9474 8546 9488 8566
rect 9508 8546 9516 8566
rect 9474 8504 9516 8546
rect 9590 8566 9632 8604
rect 9590 8546 9598 8566
rect 9618 8546 9632 8566
rect 9590 8504 9632 8546
rect 9682 8573 9727 8604
rect 9682 8566 9726 8573
rect 9682 8546 9694 8566
rect 9714 8546 9726 8566
rect 9682 8504 9726 8546
rect 13526 8579 13570 8617
rect 13526 8559 13538 8579
rect 13558 8559 13570 8579
rect 7561 8470 7573 8490
rect 7593 8470 7605 8490
rect 7561 8432 7605 8470
rect 5583 8370 5627 8408
rect 5583 8350 5595 8370
rect 5615 8350 5627 8370
rect 3475 8293 3519 8335
rect 3475 8273 3487 8293
rect 3507 8273 3519 8293
rect 3475 8266 3519 8273
rect 3474 8235 3519 8266
rect 3569 8293 3611 8335
rect 3569 8273 3583 8293
rect 3603 8273 3611 8293
rect 3569 8235 3611 8273
rect 3685 8293 3727 8335
rect 3685 8273 3693 8293
rect 3713 8273 3727 8293
rect 3685 8235 3727 8273
rect 3777 8293 3821 8335
rect 3777 8273 3789 8293
rect 3809 8273 3821 8293
rect 3777 8235 3821 8273
rect 3903 8293 3945 8335
rect 3903 8273 3911 8293
rect 3931 8273 3945 8293
rect 3903 8235 3945 8273
rect 3995 8293 4039 8335
rect 5583 8308 5627 8350
rect 5677 8370 5719 8408
rect 5677 8350 5691 8370
rect 5711 8350 5719 8370
rect 5677 8308 5719 8350
rect 5801 8370 5845 8408
rect 5801 8350 5813 8370
rect 5833 8350 5845 8370
rect 5801 8308 5845 8350
rect 5895 8370 5937 8408
rect 5895 8350 5909 8370
rect 5929 8350 5937 8370
rect 5895 8308 5937 8350
rect 6011 8370 6053 8408
rect 6011 8350 6019 8370
rect 6039 8350 6053 8370
rect 6011 8308 6053 8350
rect 6103 8377 6148 8408
rect 6103 8370 6147 8377
rect 6103 8350 6115 8370
rect 6135 8350 6147 8370
rect 6103 8308 6147 8350
rect 11418 8502 11462 8544
rect 11418 8482 11430 8502
rect 11450 8482 11462 8502
rect 11418 8475 11462 8482
rect 11417 8444 11462 8475
rect 11512 8502 11554 8544
rect 11512 8482 11526 8502
rect 11546 8482 11554 8502
rect 11512 8444 11554 8482
rect 11628 8502 11670 8544
rect 11628 8482 11636 8502
rect 11656 8482 11670 8502
rect 11628 8444 11670 8482
rect 11720 8502 11764 8544
rect 11720 8482 11732 8502
rect 11752 8482 11764 8502
rect 11720 8444 11764 8482
rect 11846 8502 11888 8544
rect 11846 8482 11854 8502
rect 11874 8482 11888 8502
rect 11846 8444 11888 8482
rect 11938 8502 11982 8544
rect 13526 8517 13570 8559
rect 13620 8579 13662 8617
rect 13620 8559 13634 8579
rect 13654 8559 13662 8579
rect 13620 8517 13662 8559
rect 13744 8579 13788 8617
rect 13744 8559 13756 8579
rect 13776 8559 13788 8579
rect 13744 8517 13788 8559
rect 13838 8579 13880 8617
rect 13838 8559 13852 8579
rect 13872 8559 13880 8579
rect 13838 8517 13880 8559
rect 13954 8579 13996 8617
rect 13954 8559 13962 8579
rect 13982 8559 13996 8579
rect 13954 8517 13996 8559
rect 14046 8586 14091 8617
rect 14046 8579 14090 8586
rect 14046 8559 14058 8579
rect 14078 8559 14090 8579
rect 14046 8517 14090 8559
rect 25208 8672 25253 8703
rect 25303 8730 25345 8772
rect 25303 8710 25317 8730
rect 25337 8710 25345 8730
rect 25303 8672 25345 8710
rect 25419 8730 25461 8772
rect 25419 8710 25427 8730
rect 25447 8710 25461 8730
rect 25419 8672 25461 8710
rect 25511 8730 25555 8772
rect 25511 8710 25523 8730
rect 25543 8710 25555 8730
rect 25511 8672 25555 8710
rect 25637 8730 25679 8772
rect 25637 8710 25645 8730
rect 25665 8710 25679 8730
rect 25637 8672 25679 8710
rect 25729 8730 25773 8772
rect 25729 8710 25741 8730
rect 25761 8710 25773 8730
rect 25729 8672 25773 8710
rect 29586 8742 29630 8784
rect 29586 8722 29598 8742
rect 29618 8722 29630 8742
rect 29586 8715 29630 8722
rect 29585 8684 29630 8715
rect 29680 8742 29722 8784
rect 29680 8722 29694 8742
rect 29714 8722 29722 8742
rect 29680 8684 29722 8722
rect 29796 8742 29838 8784
rect 29796 8722 29804 8742
rect 29824 8722 29838 8742
rect 29796 8684 29838 8722
rect 29888 8742 29932 8784
rect 29888 8722 29900 8742
rect 29920 8722 29932 8742
rect 29888 8684 29932 8722
rect 30014 8742 30056 8784
rect 30014 8722 30022 8742
rect 30042 8722 30056 8742
rect 30014 8684 30056 8722
rect 30106 8742 30150 8784
rect 30106 8722 30118 8742
rect 30138 8722 30150 8742
rect 30106 8684 30150 8722
rect 33950 8755 33994 8797
rect 33950 8735 33962 8755
rect 33982 8735 33994 8755
rect 33950 8728 33994 8735
rect 33949 8697 33994 8728
rect 34044 8755 34086 8797
rect 34044 8735 34058 8755
rect 34078 8735 34086 8755
rect 34044 8697 34086 8735
rect 34160 8755 34202 8797
rect 34160 8735 34168 8755
rect 34188 8735 34202 8755
rect 34160 8697 34202 8735
rect 34252 8755 34296 8797
rect 34252 8735 34264 8755
rect 34284 8735 34296 8755
rect 34252 8697 34296 8735
rect 34378 8755 34420 8797
rect 34378 8735 34386 8755
rect 34406 8735 34420 8755
rect 34378 8697 34420 8735
rect 34470 8755 34514 8797
rect 34470 8735 34482 8755
rect 34502 8735 34514 8755
rect 34470 8697 34514 8735
rect 11938 8482 11950 8502
rect 11970 8482 11982 8502
rect 11938 8444 11982 8482
rect 9960 8382 10004 8420
rect 9960 8362 9972 8382
rect 9992 8362 10004 8382
rect 3995 8273 4007 8293
rect 4027 8273 4039 8293
rect 3995 8235 4039 8273
rect 7839 8306 7883 8348
rect 7839 8286 7851 8306
rect 7871 8286 7883 8306
rect 7839 8279 7883 8286
rect 7838 8248 7883 8279
rect 7933 8306 7975 8348
rect 7933 8286 7947 8306
rect 7967 8286 7975 8306
rect 7933 8248 7975 8286
rect 8049 8306 8091 8348
rect 8049 8286 8057 8306
rect 8077 8286 8091 8306
rect 8049 8248 8091 8286
rect 8141 8306 8185 8348
rect 8141 8286 8153 8306
rect 8173 8286 8185 8306
rect 8141 8248 8185 8286
rect 8267 8306 8309 8348
rect 8267 8286 8275 8306
rect 8295 8286 8309 8306
rect 8267 8248 8309 8286
rect 8359 8306 8403 8348
rect 9960 8320 10004 8362
rect 10054 8382 10096 8420
rect 10054 8362 10068 8382
rect 10088 8362 10096 8382
rect 10054 8320 10096 8362
rect 10178 8382 10222 8420
rect 10178 8362 10190 8382
rect 10210 8362 10222 8382
rect 10178 8320 10222 8362
rect 10272 8382 10314 8420
rect 10272 8362 10286 8382
rect 10306 8362 10314 8382
rect 10272 8320 10314 8362
rect 10388 8382 10430 8420
rect 10388 8362 10396 8382
rect 10416 8362 10430 8382
rect 10388 8320 10430 8362
rect 10480 8389 10525 8420
rect 10480 8382 10524 8389
rect 10480 8362 10492 8382
rect 10512 8362 10524 8382
rect 10480 8320 10524 8362
rect 15782 8515 15826 8557
rect 15782 8495 15794 8515
rect 15814 8495 15826 8515
rect 15782 8488 15826 8495
rect 15781 8457 15826 8488
rect 15876 8515 15918 8557
rect 15876 8495 15890 8515
rect 15910 8495 15918 8515
rect 15876 8457 15918 8495
rect 15992 8515 16034 8557
rect 15992 8495 16000 8515
rect 16020 8495 16034 8515
rect 15992 8457 16034 8495
rect 16084 8515 16128 8557
rect 16084 8495 16096 8515
rect 16116 8495 16128 8515
rect 16084 8457 16128 8495
rect 16210 8515 16252 8557
rect 16210 8495 16218 8515
rect 16238 8495 16252 8515
rect 16210 8457 16252 8495
rect 16302 8515 16346 8557
rect 17792 8553 17836 8591
rect 17792 8533 17804 8553
rect 17824 8533 17836 8553
rect 16302 8495 16314 8515
rect 16334 8495 16346 8515
rect 16302 8457 16346 8495
rect 17792 8491 17836 8533
rect 17886 8553 17928 8591
rect 17886 8533 17900 8553
rect 17920 8533 17928 8553
rect 17886 8491 17928 8533
rect 18010 8553 18054 8591
rect 18010 8533 18022 8553
rect 18042 8533 18054 8553
rect 18010 8491 18054 8533
rect 18104 8553 18146 8591
rect 18104 8533 18118 8553
rect 18138 8533 18146 8553
rect 18104 8491 18146 8533
rect 18220 8553 18262 8591
rect 18220 8533 18228 8553
rect 18248 8533 18262 8553
rect 18220 8491 18262 8533
rect 18312 8560 18357 8591
rect 18312 8553 18356 8560
rect 18312 8533 18324 8553
rect 18344 8533 18356 8553
rect 18312 8491 18356 8533
rect 22156 8566 22200 8604
rect 22156 8546 22168 8566
rect 22188 8546 22200 8566
rect 14324 8395 14368 8433
rect 14324 8375 14336 8395
rect 14356 8375 14368 8395
rect 8359 8286 8371 8306
rect 8391 8286 8403 8306
rect 8359 8248 8403 8286
rect 422 8129 466 8167
rect 422 8109 434 8129
rect 454 8109 466 8129
rect 422 8067 466 8109
rect 516 8129 558 8167
rect 516 8109 530 8129
rect 550 8109 558 8129
rect 516 8067 558 8109
rect 640 8129 684 8167
rect 640 8109 652 8129
rect 672 8109 684 8129
rect 640 8067 684 8109
rect 734 8129 776 8167
rect 734 8109 748 8129
rect 768 8109 776 8129
rect 734 8067 776 8109
rect 850 8129 892 8167
rect 850 8109 858 8129
rect 878 8109 892 8129
rect 850 8067 892 8109
rect 942 8136 987 8167
rect 942 8129 986 8136
rect 942 8109 954 8129
rect 974 8109 986 8129
rect 12216 8318 12260 8360
rect 12216 8298 12228 8318
rect 12248 8298 12260 8318
rect 12216 8291 12260 8298
rect 12215 8260 12260 8291
rect 12310 8318 12352 8360
rect 12310 8298 12324 8318
rect 12344 8298 12352 8318
rect 12310 8260 12352 8298
rect 12426 8318 12468 8360
rect 12426 8298 12434 8318
rect 12454 8298 12468 8318
rect 12426 8260 12468 8298
rect 12518 8318 12562 8360
rect 12518 8298 12530 8318
rect 12550 8298 12562 8318
rect 12518 8260 12562 8298
rect 12644 8318 12686 8360
rect 12644 8298 12652 8318
rect 12672 8298 12686 8318
rect 12644 8260 12686 8298
rect 12736 8318 12780 8360
rect 14324 8333 14368 8375
rect 14418 8395 14460 8433
rect 14418 8375 14432 8395
rect 14452 8375 14460 8395
rect 14418 8333 14460 8375
rect 14542 8395 14586 8433
rect 14542 8375 14554 8395
rect 14574 8375 14586 8395
rect 14542 8333 14586 8375
rect 14636 8395 14678 8433
rect 14636 8375 14650 8395
rect 14670 8375 14678 8395
rect 14636 8333 14678 8375
rect 14752 8395 14794 8433
rect 14752 8375 14760 8395
rect 14780 8375 14794 8395
rect 14752 8333 14794 8375
rect 14844 8402 14889 8433
rect 14844 8395 14888 8402
rect 14844 8375 14856 8395
rect 14876 8375 14888 8395
rect 14844 8333 14888 8375
rect 20048 8489 20092 8531
rect 20048 8469 20060 8489
rect 20080 8469 20092 8489
rect 20048 8462 20092 8469
rect 20047 8431 20092 8462
rect 20142 8489 20184 8531
rect 20142 8469 20156 8489
rect 20176 8469 20184 8489
rect 20142 8431 20184 8469
rect 20258 8489 20300 8531
rect 20258 8469 20266 8489
rect 20286 8469 20300 8489
rect 20258 8431 20300 8469
rect 20350 8489 20394 8531
rect 20350 8469 20362 8489
rect 20382 8469 20394 8489
rect 20350 8431 20394 8469
rect 20476 8489 20518 8531
rect 20476 8469 20484 8489
rect 20504 8469 20518 8489
rect 20476 8431 20518 8469
rect 20568 8489 20612 8531
rect 22156 8504 22200 8546
rect 22250 8566 22292 8604
rect 22250 8546 22264 8566
rect 22284 8546 22292 8566
rect 22250 8504 22292 8546
rect 22374 8566 22418 8604
rect 22374 8546 22386 8566
rect 22406 8546 22418 8566
rect 22374 8504 22418 8546
rect 22468 8566 22510 8604
rect 22468 8546 22482 8566
rect 22502 8546 22510 8566
rect 22468 8504 22510 8546
rect 22584 8566 22626 8604
rect 22584 8546 22592 8566
rect 22612 8546 22626 8566
rect 22584 8504 22626 8546
rect 22676 8573 22721 8604
rect 22676 8566 22720 8573
rect 22676 8546 22688 8566
rect 22708 8546 22720 8566
rect 22676 8504 22720 8546
rect 26533 8578 26577 8616
rect 26533 8558 26545 8578
rect 26565 8558 26577 8578
rect 20568 8469 20580 8489
rect 20600 8469 20612 8489
rect 20568 8431 20612 8469
rect 12736 8298 12748 8318
rect 12768 8298 12780 8318
rect 12736 8260 12780 8298
rect 4786 8142 4830 8180
rect 942 8067 986 8109
rect 2578 8067 2622 8109
rect 2578 8047 2590 8067
rect 2610 8047 2622 8067
rect 2578 8040 2622 8047
rect 2577 8009 2622 8040
rect 2672 8067 2714 8109
rect 2672 8047 2686 8067
rect 2706 8047 2714 8067
rect 2672 8009 2714 8047
rect 2788 8067 2830 8109
rect 2788 8047 2796 8067
rect 2816 8047 2830 8067
rect 2788 8009 2830 8047
rect 2880 8067 2924 8109
rect 2880 8047 2892 8067
rect 2912 8047 2924 8067
rect 2880 8009 2924 8047
rect 3006 8067 3048 8109
rect 3006 8047 3014 8067
rect 3034 8047 3048 8067
rect 3006 8009 3048 8047
rect 3098 8067 3142 8109
rect 4786 8122 4798 8142
rect 4818 8122 4830 8142
rect 3098 8047 3110 8067
rect 3130 8047 3142 8067
rect 4786 8080 4830 8122
rect 4880 8142 4922 8180
rect 4880 8122 4894 8142
rect 4914 8122 4922 8142
rect 4880 8080 4922 8122
rect 5004 8142 5048 8180
rect 5004 8122 5016 8142
rect 5036 8122 5048 8142
rect 5004 8080 5048 8122
rect 5098 8142 5140 8180
rect 5098 8122 5112 8142
rect 5132 8122 5140 8142
rect 5098 8080 5140 8122
rect 5214 8142 5256 8180
rect 5214 8122 5222 8142
rect 5242 8122 5256 8142
rect 5214 8080 5256 8122
rect 5306 8149 5351 8180
rect 5306 8142 5350 8149
rect 5306 8122 5318 8142
rect 5338 8122 5350 8142
rect 16580 8331 16624 8373
rect 16580 8311 16592 8331
rect 16612 8311 16624 8331
rect 16580 8304 16624 8311
rect 16579 8273 16624 8304
rect 16674 8331 16716 8373
rect 16674 8311 16688 8331
rect 16708 8311 16716 8331
rect 16674 8273 16716 8311
rect 16790 8331 16832 8373
rect 16790 8311 16798 8331
rect 16818 8311 16832 8331
rect 16790 8273 16832 8311
rect 16882 8331 16926 8373
rect 16882 8311 16894 8331
rect 16914 8311 16926 8331
rect 16882 8273 16926 8311
rect 17008 8331 17050 8373
rect 17008 8311 17016 8331
rect 17036 8311 17050 8331
rect 17008 8273 17050 8311
rect 17100 8331 17144 8373
rect 18590 8369 18634 8407
rect 18590 8349 18602 8369
rect 18622 8349 18634 8369
rect 17100 8311 17112 8331
rect 17132 8311 17144 8331
rect 17100 8273 17144 8311
rect 18590 8307 18634 8349
rect 18684 8369 18726 8407
rect 18684 8349 18698 8369
rect 18718 8349 18726 8369
rect 18684 8307 18726 8349
rect 18808 8369 18852 8407
rect 18808 8349 18820 8369
rect 18840 8349 18852 8369
rect 18808 8307 18852 8349
rect 18902 8369 18944 8407
rect 18902 8349 18916 8369
rect 18936 8349 18944 8369
rect 18902 8307 18944 8349
rect 19018 8369 19060 8407
rect 19018 8349 19026 8369
rect 19046 8349 19060 8369
rect 19018 8307 19060 8349
rect 19110 8376 19155 8407
rect 19110 8369 19154 8376
rect 19110 8349 19122 8369
rect 19142 8349 19154 8369
rect 19110 8307 19154 8349
rect 24412 8502 24456 8544
rect 24412 8482 24424 8502
rect 24444 8482 24456 8502
rect 24412 8475 24456 8482
rect 24411 8444 24456 8475
rect 24506 8502 24548 8544
rect 24506 8482 24520 8502
rect 24540 8482 24548 8502
rect 24506 8444 24548 8482
rect 24622 8502 24664 8544
rect 24622 8482 24630 8502
rect 24650 8482 24664 8502
rect 24622 8444 24664 8482
rect 24714 8502 24758 8544
rect 24714 8482 24726 8502
rect 24746 8482 24758 8502
rect 24714 8444 24758 8482
rect 24840 8502 24882 8544
rect 24840 8482 24848 8502
rect 24868 8482 24882 8502
rect 24840 8444 24882 8482
rect 24932 8502 24976 8544
rect 26533 8516 26577 8558
rect 26627 8578 26669 8616
rect 26627 8558 26641 8578
rect 26661 8558 26669 8578
rect 26627 8516 26669 8558
rect 26751 8578 26795 8616
rect 26751 8558 26763 8578
rect 26783 8558 26795 8578
rect 26751 8516 26795 8558
rect 26845 8578 26887 8616
rect 26845 8558 26859 8578
rect 26879 8558 26887 8578
rect 26845 8516 26887 8558
rect 26961 8578 27003 8616
rect 26961 8558 26969 8578
rect 26989 8558 27003 8578
rect 26961 8516 27003 8558
rect 27053 8585 27098 8616
rect 27053 8578 27097 8585
rect 27053 8558 27065 8578
rect 27085 8558 27097 8578
rect 27053 8516 27097 8558
rect 30897 8591 30941 8629
rect 30897 8571 30909 8591
rect 30929 8571 30941 8591
rect 24932 8482 24944 8502
rect 24964 8482 24976 8502
rect 24932 8444 24976 8482
rect 22954 8382 22998 8420
rect 22954 8362 22966 8382
rect 22986 8362 22998 8382
rect 9163 8154 9207 8192
rect 5306 8080 5350 8122
rect 6942 8080 6986 8122
rect 3098 8009 3142 8047
rect 6942 8060 6954 8080
rect 6974 8060 6986 8080
rect 6942 8053 6986 8060
rect 6941 8022 6986 8053
rect 7036 8080 7078 8122
rect 7036 8060 7050 8080
rect 7070 8060 7078 8080
rect 7036 8022 7078 8060
rect 7152 8080 7194 8122
rect 7152 8060 7160 8080
rect 7180 8060 7194 8080
rect 7152 8022 7194 8060
rect 7244 8080 7288 8122
rect 7244 8060 7256 8080
rect 7276 8060 7288 8080
rect 7244 8022 7288 8060
rect 7370 8080 7412 8122
rect 7370 8060 7378 8080
rect 7398 8060 7412 8080
rect 7370 8022 7412 8060
rect 7462 8080 7506 8122
rect 9163 8134 9175 8154
rect 9195 8134 9207 8154
rect 7462 8060 7474 8080
rect 7494 8060 7506 8080
rect 9163 8092 9207 8134
rect 9257 8154 9299 8192
rect 9257 8134 9271 8154
rect 9291 8134 9299 8154
rect 9257 8092 9299 8134
rect 9381 8154 9425 8192
rect 9381 8134 9393 8154
rect 9413 8134 9425 8154
rect 9381 8092 9425 8134
rect 9475 8154 9517 8192
rect 9475 8134 9489 8154
rect 9509 8134 9517 8154
rect 9475 8092 9517 8134
rect 9591 8154 9633 8192
rect 9591 8134 9599 8154
rect 9619 8134 9633 8154
rect 9591 8092 9633 8134
rect 9683 8161 9728 8192
rect 9683 8154 9727 8161
rect 9683 8134 9695 8154
rect 9715 8134 9727 8154
rect 20846 8305 20890 8347
rect 20846 8285 20858 8305
rect 20878 8285 20890 8305
rect 20846 8278 20890 8285
rect 20845 8247 20890 8278
rect 20940 8305 20982 8347
rect 20940 8285 20954 8305
rect 20974 8285 20982 8305
rect 20940 8247 20982 8285
rect 21056 8305 21098 8347
rect 21056 8285 21064 8305
rect 21084 8285 21098 8305
rect 21056 8247 21098 8285
rect 21148 8305 21192 8347
rect 21148 8285 21160 8305
rect 21180 8285 21192 8305
rect 21148 8247 21192 8285
rect 21274 8305 21316 8347
rect 21274 8285 21282 8305
rect 21302 8285 21316 8305
rect 21274 8247 21316 8285
rect 21366 8305 21410 8347
rect 22954 8320 22998 8362
rect 23048 8382 23090 8420
rect 23048 8362 23062 8382
rect 23082 8362 23090 8382
rect 23048 8320 23090 8362
rect 23172 8382 23216 8420
rect 23172 8362 23184 8382
rect 23204 8362 23216 8382
rect 23172 8320 23216 8362
rect 23266 8382 23308 8420
rect 23266 8362 23280 8382
rect 23300 8362 23308 8382
rect 23266 8320 23308 8362
rect 23382 8382 23424 8420
rect 23382 8362 23390 8382
rect 23410 8362 23424 8382
rect 23382 8320 23424 8362
rect 23474 8389 23519 8420
rect 23474 8382 23518 8389
rect 23474 8362 23486 8382
rect 23506 8362 23518 8382
rect 23474 8320 23518 8362
rect 28789 8514 28833 8556
rect 28789 8494 28801 8514
rect 28821 8494 28833 8514
rect 28789 8487 28833 8494
rect 28788 8456 28833 8487
rect 28883 8514 28925 8556
rect 28883 8494 28897 8514
rect 28917 8494 28925 8514
rect 28883 8456 28925 8494
rect 28999 8514 29041 8556
rect 28999 8494 29007 8514
rect 29027 8494 29041 8514
rect 28999 8456 29041 8494
rect 29091 8514 29135 8556
rect 29091 8494 29103 8514
rect 29123 8494 29135 8514
rect 29091 8456 29135 8494
rect 29217 8514 29259 8556
rect 29217 8494 29225 8514
rect 29245 8494 29259 8514
rect 29217 8456 29259 8494
rect 29309 8514 29353 8556
rect 30897 8529 30941 8571
rect 30991 8591 31033 8629
rect 30991 8571 31005 8591
rect 31025 8571 31033 8591
rect 30991 8529 31033 8571
rect 31115 8591 31159 8629
rect 31115 8571 31127 8591
rect 31147 8571 31159 8591
rect 31115 8529 31159 8571
rect 31209 8591 31251 8629
rect 31209 8571 31223 8591
rect 31243 8571 31251 8591
rect 31209 8529 31251 8571
rect 31325 8591 31367 8629
rect 31325 8571 31333 8591
rect 31353 8571 31367 8591
rect 31325 8529 31367 8571
rect 31417 8598 31462 8629
rect 31417 8591 31461 8598
rect 31417 8571 31429 8591
rect 31449 8571 31461 8591
rect 31417 8529 31461 8571
rect 29309 8494 29321 8514
rect 29341 8494 29353 8514
rect 29309 8456 29353 8494
rect 27331 8394 27375 8432
rect 27331 8374 27343 8394
rect 27363 8374 27375 8394
rect 21366 8285 21378 8305
rect 21398 8285 21410 8305
rect 21366 8247 21410 8285
rect 13527 8167 13571 8205
rect 9683 8092 9727 8134
rect 11319 8092 11363 8134
rect 7462 8022 7506 8060
rect 11319 8072 11331 8092
rect 11351 8072 11363 8092
rect 11319 8065 11363 8072
rect 11318 8034 11363 8065
rect 11413 8092 11455 8134
rect 11413 8072 11427 8092
rect 11447 8072 11455 8092
rect 11413 8034 11455 8072
rect 11529 8092 11571 8134
rect 11529 8072 11537 8092
rect 11557 8072 11571 8092
rect 11529 8034 11571 8072
rect 11621 8092 11665 8134
rect 11621 8072 11633 8092
rect 11653 8072 11665 8092
rect 11621 8034 11665 8072
rect 11747 8092 11789 8134
rect 11747 8072 11755 8092
rect 11775 8072 11789 8092
rect 11747 8034 11789 8072
rect 11839 8092 11883 8134
rect 13527 8147 13539 8167
rect 13559 8147 13571 8167
rect 11839 8072 11851 8092
rect 11871 8072 11883 8092
rect 13527 8105 13571 8147
rect 13621 8167 13663 8205
rect 13621 8147 13635 8167
rect 13655 8147 13663 8167
rect 13621 8105 13663 8147
rect 13745 8167 13789 8205
rect 13745 8147 13757 8167
rect 13777 8147 13789 8167
rect 13745 8105 13789 8147
rect 13839 8167 13881 8205
rect 13839 8147 13853 8167
rect 13873 8147 13881 8167
rect 13839 8105 13881 8147
rect 13955 8167 13997 8205
rect 13955 8147 13963 8167
rect 13983 8147 13997 8167
rect 13955 8105 13997 8147
rect 14047 8174 14092 8205
rect 14047 8167 14091 8174
rect 14047 8147 14059 8167
rect 14079 8147 14091 8167
rect 25210 8318 25254 8360
rect 25210 8298 25222 8318
rect 25242 8298 25254 8318
rect 25210 8291 25254 8298
rect 25209 8260 25254 8291
rect 25304 8318 25346 8360
rect 25304 8298 25318 8318
rect 25338 8298 25346 8318
rect 25304 8260 25346 8298
rect 25420 8318 25462 8360
rect 25420 8298 25428 8318
rect 25448 8298 25462 8318
rect 25420 8260 25462 8298
rect 25512 8318 25556 8360
rect 25512 8298 25524 8318
rect 25544 8298 25556 8318
rect 25512 8260 25556 8298
rect 25638 8318 25680 8360
rect 25638 8298 25646 8318
rect 25666 8298 25680 8318
rect 25638 8260 25680 8298
rect 25730 8318 25774 8360
rect 27331 8332 27375 8374
rect 27425 8394 27467 8432
rect 27425 8374 27439 8394
rect 27459 8374 27467 8394
rect 27425 8332 27467 8374
rect 27549 8394 27593 8432
rect 27549 8374 27561 8394
rect 27581 8374 27593 8394
rect 27549 8332 27593 8374
rect 27643 8394 27685 8432
rect 27643 8374 27657 8394
rect 27677 8374 27685 8394
rect 27643 8332 27685 8374
rect 27759 8394 27801 8432
rect 27759 8374 27767 8394
rect 27787 8374 27801 8394
rect 27759 8332 27801 8374
rect 27851 8401 27896 8432
rect 27851 8394 27895 8401
rect 27851 8374 27863 8394
rect 27883 8374 27895 8394
rect 27851 8332 27895 8374
rect 33153 8527 33197 8569
rect 33153 8507 33165 8527
rect 33185 8507 33197 8527
rect 33153 8500 33197 8507
rect 33152 8469 33197 8500
rect 33247 8527 33289 8569
rect 33247 8507 33261 8527
rect 33281 8507 33289 8527
rect 33247 8469 33289 8507
rect 33363 8527 33405 8569
rect 33363 8507 33371 8527
rect 33391 8507 33405 8527
rect 33363 8469 33405 8507
rect 33455 8527 33499 8569
rect 33455 8507 33467 8527
rect 33487 8507 33499 8527
rect 33455 8469 33499 8507
rect 33581 8527 33623 8569
rect 33581 8507 33589 8527
rect 33609 8507 33623 8527
rect 33581 8469 33623 8507
rect 33673 8527 33717 8569
rect 33673 8507 33685 8527
rect 33705 8507 33717 8527
rect 33673 8469 33717 8507
rect 31695 8407 31739 8445
rect 31695 8387 31707 8407
rect 31727 8387 31739 8407
rect 25730 8298 25742 8318
rect 25762 8298 25774 8318
rect 25730 8260 25774 8298
rect 14047 8105 14091 8147
rect 15683 8105 15727 8147
rect 11839 8034 11883 8072
rect 15683 8085 15695 8105
rect 15715 8085 15727 8105
rect 15683 8078 15727 8085
rect 15682 8047 15727 8078
rect 15777 8105 15819 8147
rect 15777 8085 15791 8105
rect 15811 8085 15819 8105
rect 15777 8047 15819 8085
rect 15893 8105 15935 8147
rect 15893 8085 15901 8105
rect 15921 8085 15935 8105
rect 15893 8047 15935 8085
rect 15985 8105 16029 8147
rect 15985 8085 15997 8105
rect 16017 8085 16029 8105
rect 15985 8047 16029 8085
rect 16111 8105 16153 8147
rect 16111 8085 16119 8105
rect 16139 8085 16153 8105
rect 16111 8047 16153 8085
rect 16203 8105 16247 8147
rect 16203 8085 16215 8105
rect 16235 8085 16247 8105
rect 17793 8141 17837 8179
rect 17793 8121 17805 8141
rect 17825 8121 17837 8141
rect 16203 8047 16247 8085
rect 17793 8079 17837 8121
rect 17887 8141 17929 8179
rect 17887 8121 17901 8141
rect 17921 8121 17929 8141
rect 17887 8079 17929 8121
rect 18011 8141 18055 8179
rect 18011 8121 18023 8141
rect 18043 8121 18055 8141
rect 18011 8079 18055 8121
rect 18105 8141 18147 8179
rect 18105 8121 18119 8141
rect 18139 8121 18147 8141
rect 18105 8079 18147 8121
rect 18221 8141 18263 8179
rect 18221 8121 18229 8141
rect 18249 8121 18263 8141
rect 18221 8079 18263 8121
rect 18313 8148 18358 8179
rect 18313 8141 18357 8148
rect 18313 8121 18325 8141
rect 18345 8121 18357 8141
rect 29587 8330 29631 8372
rect 29587 8310 29599 8330
rect 29619 8310 29631 8330
rect 29587 8303 29631 8310
rect 29586 8272 29631 8303
rect 29681 8330 29723 8372
rect 29681 8310 29695 8330
rect 29715 8310 29723 8330
rect 29681 8272 29723 8310
rect 29797 8330 29839 8372
rect 29797 8310 29805 8330
rect 29825 8310 29839 8330
rect 29797 8272 29839 8310
rect 29889 8330 29933 8372
rect 29889 8310 29901 8330
rect 29921 8310 29933 8330
rect 29889 8272 29933 8310
rect 30015 8330 30057 8372
rect 30015 8310 30023 8330
rect 30043 8310 30057 8330
rect 30015 8272 30057 8310
rect 30107 8330 30151 8372
rect 31695 8345 31739 8387
rect 31789 8407 31831 8445
rect 31789 8387 31803 8407
rect 31823 8387 31831 8407
rect 31789 8345 31831 8387
rect 31913 8407 31957 8445
rect 31913 8387 31925 8407
rect 31945 8387 31957 8407
rect 31913 8345 31957 8387
rect 32007 8407 32049 8445
rect 32007 8387 32021 8407
rect 32041 8387 32049 8407
rect 32007 8345 32049 8387
rect 32123 8407 32165 8445
rect 32123 8387 32131 8407
rect 32151 8387 32165 8407
rect 32123 8345 32165 8387
rect 32215 8414 32260 8445
rect 32215 8407 32259 8414
rect 32215 8387 32227 8407
rect 32247 8387 32259 8407
rect 32215 8345 32259 8387
rect 30107 8310 30119 8330
rect 30139 8310 30151 8330
rect 30107 8272 30151 8310
rect 22157 8154 22201 8192
rect 18313 8079 18357 8121
rect 19949 8079 19993 8121
rect 19949 8059 19961 8079
rect 19981 8059 19993 8079
rect 19949 8052 19993 8059
rect 19948 8021 19993 8052
rect 20043 8079 20085 8121
rect 20043 8059 20057 8079
rect 20077 8059 20085 8079
rect 20043 8021 20085 8059
rect 20159 8079 20201 8121
rect 20159 8059 20167 8079
rect 20187 8059 20201 8079
rect 20159 8021 20201 8059
rect 20251 8079 20295 8121
rect 20251 8059 20263 8079
rect 20283 8059 20295 8079
rect 20251 8021 20295 8059
rect 20377 8079 20419 8121
rect 20377 8059 20385 8079
rect 20405 8059 20419 8079
rect 20377 8021 20419 8059
rect 20469 8079 20513 8121
rect 22157 8134 22169 8154
rect 22189 8134 22201 8154
rect 20469 8059 20481 8079
rect 20501 8059 20513 8079
rect 22157 8092 22201 8134
rect 22251 8154 22293 8192
rect 22251 8134 22265 8154
rect 22285 8134 22293 8154
rect 22251 8092 22293 8134
rect 22375 8154 22419 8192
rect 22375 8134 22387 8154
rect 22407 8134 22419 8154
rect 22375 8092 22419 8134
rect 22469 8154 22511 8192
rect 22469 8134 22483 8154
rect 22503 8134 22511 8154
rect 22469 8092 22511 8134
rect 22585 8154 22627 8192
rect 22585 8134 22593 8154
rect 22613 8134 22627 8154
rect 22585 8092 22627 8134
rect 22677 8161 22722 8192
rect 22677 8154 22721 8161
rect 22677 8134 22689 8154
rect 22709 8134 22721 8154
rect 33951 8343 33995 8385
rect 33951 8323 33963 8343
rect 33983 8323 33995 8343
rect 33951 8316 33995 8323
rect 33950 8285 33995 8316
rect 34045 8343 34087 8385
rect 34045 8323 34059 8343
rect 34079 8323 34087 8343
rect 34045 8285 34087 8323
rect 34161 8343 34203 8385
rect 34161 8323 34169 8343
rect 34189 8323 34203 8343
rect 34161 8285 34203 8323
rect 34253 8343 34297 8385
rect 34253 8323 34265 8343
rect 34285 8323 34297 8343
rect 34253 8285 34297 8323
rect 34379 8343 34421 8385
rect 34379 8323 34387 8343
rect 34407 8323 34421 8343
rect 34379 8285 34421 8323
rect 34471 8343 34515 8385
rect 34471 8323 34483 8343
rect 34503 8323 34515 8343
rect 34471 8285 34515 8323
rect 26534 8166 26578 8204
rect 22677 8092 22721 8134
rect 24313 8092 24357 8134
rect 20469 8021 20513 8059
rect 24313 8072 24325 8092
rect 24345 8072 24357 8092
rect 24313 8065 24357 8072
rect 24312 8034 24357 8065
rect 24407 8092 24449 8134
rect 24407 8072 24421 8092
rect 24441 8072 24449 8092
rect 24407 8034 24449 8072
rect 24523 8092 24565 8134
rect 24523 8072 24531 8092
rect 24551 8072 24565 8092
rect 24523 8034 24565 8072
rect 24615 8092 24659 8134
rect 24615 8072 24627 8092
rect 24647 8072 24659 8092
rect 24615 8034 24659 8072
rect 24741 8092 24783 8134
rect 24741 8072 24749 8092
rect 24769 8072 24783 8092
rect 24741 8034 24783 8072
rect 24833 8092 24877 8134
rect 26534 8146 26546 8166
rect 26566 8146 26578 8166
rect 24833 8072 24845 8092
rect 24865 8072 24877 8092
rect 26534 8104 26578 8146
rect 26628 8166 26670 8204
rect 26628 8146 26642 8166
rect 26662 8146 26670 8166
rect 26628 8104 26670 8146
rect 26752 8166 26796 8204
rect 26752 8146 26764 8166
rect 26784 8146 26796 8166
rect 26752 8104 26796 8146
rect 26846 8166 26888 8204
rect 26846 8146 26860 8166
rect 26880 8146 26888 8166
rect 26846 8104 26888 8146
rect 26962 8166 27004 8204
rect 26962 8146 26970 8166
rect 26990 8146 27004 8166
rect 26962 8104 27004 8146
rect 27054 8173 27099 8204
rect 27054 8166 27098 8173
rect 27054 8146 27066 8166
rect 27086 8146 27098 8166
rect 30898 8179 30942 8217
rect 27054 8104 27098 8146
rect 28690 8104 28734 8146
rect 24833 8034 24877 8072
rect 28690 8084 28702 8104
rect 28722 8084 28734 8104
rect 28690 8077 28734 8084
rect 28689 8046 28734 8077
rect 28784 8104 28826 8146
rect 28784 8084 28798 8104
rect 28818 8084 28826 8104
rect 28784 8046 28826 8084
rect 28900 8104 28942 8146
rect 28900 8084 28908 8104
rect 28928 8084 28942 8104
rect 28900 8046 28942 8084
rect 28992 8104 29036 8146
rect 28992 8084 29004 8104
rect 29024 8084 29036 8104
rect 28992 8046 29036 8084
rect 29118 8104 29160 8146
rect 29118 8084 29126 8104
rect 29146 8084 29160 8104
rect 29118 8046 29160 8084
rect 29210 8104 29254 8146
rect 30898 8159 30910 8179
rect 30930 8159 30942 8179
rect 29210 8084 29222 8104
rect 29242 8084 29254 8104
rect 30898 8117 30942 8159
rect 30992 8179 31034 8217
rect 30992 8159 31006 8179
rect 31026 8159 31034 8179
rect 30992 8117 31034 8159
rect 31116 8179 31160 8217
rect 31116 8159 31128 8179
rect 31148 8159 31160 8179
rect 31116 8117 31160 8159
rect 31210 8179 31252 8217
rect 31210 8159 31224 8179
rect 31244 8159 31252 8179
rect 31210 8117 31252 8159
rect 31326 8179 31368 8217
rect 31326 8159 31334 8179
rect 31354 8159 31368 8179
rect 31326 8117 31368 8159
rect 31418 8186 31463 8217
rect 31418 8179 31462 8186
rect 31418 8159 31430 8179
rect 31450 8159 31462 8179
rect 31418 8117 31462 8159
rect 33054 8117 33098 8159
rect 29210 8046 29254 8084
rect 33054 8097 33066 8117
rect 33086 8097 33098 8117
rect 33054 8090 33098 8097
rect 33053 8059 33098 8090
rect 33148 8117 33190 8159
rect 33148 8097 33162 8117
rect 33182 8097 33190 8117
rect 33148 8059 33190 8097
rect 33264 8117 33306 8159
rect 33264 8097 33272 8117
rect 33292 8097 33306 8117
rect 33264 8059 33306 8097
rect 33356 8117 33400 8159
rect 33356 8097 33368 8117
rect 33388 8097 33400 8117
rect 33356 8059 33400 8097
rect 33482 8117 33524 8159
rect 33482 8097 33490 8117
rect 33510 8097 33524 8117
rect 33482 8059 33524 8097
rect 33574 8117 33618 8159
rect 33574 8097 33586 8117
rect 33606 8097 33618 8117
rect 33574 8059 33618 8097
rect 1301 7749 1345 7787
rect 1301 7729 1313 7749
rect 1333 7729 1345 7749
rect 1301 7687 1345 7729
rect 1395 7749 1437 7787
rect 1395 7729 1409 7749
rect 1429 7729 1437 7749
rect 1395 7687 1437 7729
rect 1519 7749 1563 7787
rect 1519 7729 1531 7749
rect 1551 7729 1563 7749
rect 1519 7687 1563 7729
rect 1613 7749 1655 7787
rect 1613 7729 1627 7749
rect 1647 7729 1655 7749
rect 1613 7687 1655 7729
rect 1729 7749 1771 7787
rect 1729 7729 1737 7749
rect 1757 7729 1771 7749
rect 1729 7687 1771 7729
rect 1821 7756 1866 7787
rect 1821 7749 1865 7756
rect 1821 7729 1833 7749
rect 1853 7729 1865 7749
rect 5665 7762 5709 7800
rect 1821 7687 1865 7729
rect 3457 7687 3501 7729
rect 3457 7667 3469 7687
rect 3489 7667 3501 7687
rect 3457 7660 3501 7667
rect 3456 7629 3501 7660
rect 3551 7687 3593 7729
rect 3551 7667 3565 7687
rect 3585 7667 3593 7687
rect 3551 7629 3593 7667
rect 3667 7687 3709 7729
rect 3667 7667 3675 7687
rect 3695 7667 3709 7687
rect 3667 7629 3709 7667
rect 3759 7687 3803 7729
rect 3759 7667 3771 7687
rect 3791 7667 3803 7687
rect 3759 7629 3803 7667
rect 3885 7687 3927 7729
rect 3885 7667 3893 7687
rect 3913 7667 3927 7687
rect 3885 7629 3927 7667
rect 3977 7687 4021 7729
rect 5665 7742 5677 7762
rect 5697 7742 5709 7762
rect 3977 7667 3989 7687
rect 4009 7667 4021 7687
rect 5665 7700 5709 7742
rect 5759 7762 5801 7800
rect 5759 7742 5773 7762
rect 5793 7742 5801 7762
rect 5759 7700 5801 7742
rect 5883 7762 5927 7800
rect 5883 7742 5895 7762
rect 5915 7742 5927 7762
rect 5883 7700 5927 7742
rect 5977 7762 6019 7800
rect 5977 7742 5991 7762
rect 6011 7742 6019 7762
rect 5977 7700 6019 7742
rect 6093 7762 6135 7800
rect 6093 7742 6101 7762
rect 6121 7742 6135 7762
rect 6093 7700 6135 7742
rect 6185 7769 6230 7800
rect 6185 7762 6229 7769
rect 6185 7742 6197 7762
rect 6217 7742 6229 7762
rect 10042 7774 10086 7812
rect 6185 7700 6229 7742
rect 7821 7700 7865 7742
rect 3977 7629 4021 7667
rect 7821 7680 7833 7700
rect 7853 7680 7865 7700
rect 7821 7673 7865 7680
rect 7820 7642 7865 7673
rect 7915 7700 7957 7742
rect 7915 7680 7929 7700
rect 7949 7680 7957 7700
rect 7915 7642 7957 7680
rect 8031 7700 8073 7742
rect 8031 7680 8039 7700
rect 8059 7680 8073 7700
rect 8031 7642 8073 7680
rect 8123 7700 8167 7742
rect 8123 7680 8135 7700
rect 8155 7680 8167 7700
rect 8123 7642 8167 7680
rect 8249 7700 8291 7742
rect 8249 7680 8257 7700
rect 8277 7680 8291 7700
rect 8249 7642 8291 7680
rect 8341 7700 8385 7742
rect 10042 7754 10054 7774
rect 10074 7754 10086 7774
rect 8341 7680 8353 7700
rect 8373 7680 8385 7700
rect 10042 7712 10086 7754
rect 10136 7774 10178 7812
rect 10136 7754 10150 7774
rect 10170 7754 10178 7774
rect 10136 7712 10178 7754
rect 10260 7774 10304 7812
rect 10260 7754 10272 7774
rect 10292 7754 10304 7774
rect 10260 7712 10304 7754
rect 10354 7774 10396 7812
rect 10354 7754 10368 7774
rect 10388 7754 10396 7774
rect 10354 7712 10396 7754
rect 10470 7774 10512 7812
rect 10470 7754 10478 7774
rect 10498 7754 10512 7774
rect 10470 7712 10512 7754
rect 10562 7781 10607 7812
rect 10562 7774 10606 7781
rect 10562 7754 10574 7774
rect 10594 7754 10606 7774
rect 14406 7787 14450 7825
rect 10562 7712 10606 7754
rect 12198 7712 12242 7754
rect 8341 7642 8385 7680
rect 404 7523 448 7561
rect 404 7503 416 7523
rect 436 7503 448 7523
rect 404 7461 448 7503
rect 498 7523 540 7561
rect 498 7503 512 7523
rect 532 7503 540 7523
rect 498 7461 540 7503
rect 622 7523 666 7561
rect 622 7503 634 7523
rect 654 7503 666 7523
rect 622 7461 666 7503
rect 716 7523 758 7561
rect 716 7503 730 7523
rect 750 7503 758 7523
rect 716 7461 758 7503
rect 832 7523 874 7561
rect 832 7503 840 7523
rect 860 7503 874 7523
rect 832 7461 874 7503
rect 924 7530 969 7561
rect 924 7523 968 7530
rect 924 7503 936 7523
rect 956 7503 968 7523
rect 924 7461 968 7503
rect 12198 7692 12210 7712
rect 12230 7692 12242 7712
rect 12198 7685 12242 7692
rect 12197 7654 12242 7685
rect 12292 7712 12334 7754
rect 12292 7692 12306 7712
rect 12326 7692 12334 7712
rect 12292 7654 12334 7692
rect 12408 7712 12450 7754
rect 12408 7692 12416 7712
rect 12436 7692 12450 7712
rect 12408 7654 12450 7692
rect 12500 7712 12544 7754
rect 12500 7692 12512 7712
rect 12532 7692 12544 7712
rect 12500 7654 12544 7692
rect 12626 7712 12668 7754
rect 12626 7692 12634 7712
rect 12654 7692 12668 7712
rect 12626 7654 12668 7692
rect 12718 7712 12762 7754
rect 14406 7767 14418 7787
rect 14438 7767 14450 7787
rect 12718 7692 12730 7712
rect 12750 7692 12762 7712
rect 14406 7725 14450 7767
rect 14500 7787 14542 7825
rect 14500 7767 14514 7787
rect 14534 7767 14542 7787
rect 14500 7725 14542 7767
rect 14624 7787 14668 7825
rect 14624 7767 14636 7787
rect 14656 7767 14668 7787
rect 14624 7725 14668 7767
rect 14718 7787 14760 7825
rect 14718 7767 14732 7787
rect 14752 7767 14760 7787
rect 14718 7725 14760 7767
rect 14834 7787 14876 7825
rect 14834 7767 14842 7787
rect 14862 7767 14876 7787
rect 14834 7725 14876 7767
rect 14926 7794 14971 7825
rect 14926 7787 14970 7794
rect 14926 7767 14938 7787
rect 14958 7767 14970 7787
rect 14926 7725 14970 7767
rect 16562 7725 16606 7767
rect 12718 7654 12762 7692
rect 4768 7536 4812 7574
rect 4768 7516 4780 7536
rect 4800 7516 4812 7536
rect 2660 7459 2704 7501
rect 2660 7439 2672 7459
rect 2692 7439 2704 7459
rect 2660 7432 2704 7439
rect 2659 7401 2704 7432
rect 2754 7459 2796 7501
rect 2754 7439 2768 7459
rect 2788 7439 2796 7459
rect 2754 7401 2796 7439
rect 2870 7459 2912 7501
rect 2870 7439 2878 7459
rect 2898 7439 2912 7459
rect 2870 7401 2912 7439
rect 2962 7459 3006 7501
rect 2962 7439 2974 7459
rect 2994 7439 3006 7459
rect 2962 7401 3006 7439
rect 3088 7459 3130 7501
rect 3088 7439 3096 7459
rect 3116 7439 3130 7459
rect 3088 7401 3130 7439
rect 3180 7459 3224 7501
rect 4768 7474 4812 7516
rect 4862 7536 4904 7574
rect 4862 7516 4876 7536
rect 4896 7516 4904 7536
rect 4862 7474 4904 7516
rect 4986 7536 5030 7574
rect 4986 7516 4998 7536
rect 5018 7516 5030 7536
rect 4986 7474 5030 7516
rect 5080 7536 5122 7574
rect 5080 7516 5094 7536
rect 5114 7516 5122 7536
rect 5080 7474 5122 7516
rect 5196 7536 5238 7574
rect 5196 7516 5204 7536
rect 5224 7516 5238 7536
rect 5196 7474 5238 7516
rect 5288 7543 5333 7574
rect 5288 7536 5332 7543
rect 5288 7516 5300 7536
rect 5320 7516 5332 7536
rect 5288 7474 5332 7516
rect 16562 7705 16574 7725
rect 16594 7705 16606 7725
rect 16562 7698 16606 7705
rect 16561 7667 16606 7698
rect 16656 7725 16698 7767
rect 16656 7705 16670 7725
rect 16690 7705 16698 7725
rect 16656 7667 16698 7705
rect 16772 7725 16814 7767
rect 16772 7705 16780 7725
rect 16800 7705 16814 7725
rect 16772 7667 16814 7705
rect 16864 7725 16908 7767
rect 16864 7705 16876 7725
rect 16896 7705 16908 7725
rect 16864 7667 16908 7705
rect 16990 7725 17032 7767
rect 16990 7705 16998 7725
rect 17018 7705 17032 7725
rect 16990 7667 17032 7705
rect 17082 7725 17126 7767
rect 18672 7761 18716 7799
rect 17082 7705 17094 7725
rect 17114 7705 17126 7725
rect 17082 7667 17126 7705
rect 18672 7741 18684 7761
rect 18704 7741 18716 7761
rect 18672 7699 18716 7741
rect 18766 7761 18808 7799
rect 18766 7741 18780 7761
rect 18800 7741 18808 7761
rect 18766 7699 18808 7741
rect 18890 7761 18934 7799
rect 18890 7741 18902 7761
rect 18922 7741 18934 7761
rect 18890 7699 18934 7741
rect 18984 7761 19026 7799
rect 18984 7741 18998 7761
rect 19018 7741 19026 7761
rect 18984 7699 19026 7741
rect 19100 7761 19142 7799
rect 19100 7741 19108 7761
rect 19128 7741 19142 7761
rect 19100 7699 19142 7741
rect 19192 7768 19237 7799
rect 19192 7761 19236 7768
rect 19192 7741 19204 7761
rect 19224 7741 19236 7761
rect 23036 7774 23080 7812
rect 19192 7699 19236 7741
rect 20828 7699 20872 7741
rect 9145 7548 9189 7586
rect 9145 7528 9157 7548
rect 9177 7528 9189 7548
rect 3180 7439 3192 7459
rect 3212 7439 3224 7459
rect 3180 7401 3224 7439
rect 1202 7339 1246 7377
rect 1202 7319 1214 7339
rect 1234 7319 1246 7339
rect 1202 7277 1246 7319
rect 1296 7339 1338 7377
rect 1296 7319 1310 7339
rect 1330 7319 1338 7339
rect 1296 7277 1338 7319
rect 1420 7339 1464 7377
rect 1420 7319 1432 7339
rect 1452 7319 1464 7339
rect 1420 7277 1464 7319
rect 1514 7339 1556 7377
rect 1514 7319 1528 7339
rect 1548 7319 1556 7339
rect 1514 7277 1556 7319
rect 1630 7339 1672 7377
rect 1630 7319 1638 7339
rect 1658 7319 1672 7339
rect 1630 7277 1672 7319
rect 1722 7346 1767 7377
rect 1722 7339 1766 7346
rect 1722 7319 1734 7339
rect 1754 7319 1766 7339
rect 1722 7277 1766 7319
rect 7024 7472 7068 7514
rect 7024 7452 7036 7472
rect 7056 7452 7068 7472
rect 7024 7445 7068 7452
rect 7023 7414 7068 7445
rect 7118 7472 7160 7514
rect 7118 7452 7132 7472
rect 7152 7452 7160 7472
rect 7118 7414 7160 7452
rect 7234 7472 7276 7514
rect 7234 7452 7242 7472
rect 7262 7452 7276 7472
rect 7234 7414 7276 7452
rect 7326 7472 7370 7514
rect 7326 7452 7338 7472
rect 7358 7452 7370 7472
rect 7326 7414 7370 7452
rect 7452 7472 7494 7514
rect 7452 7452 7460 7472
rect 7480 7452 7494 7472
rect 7452 7414 7494 7452
rect 7544 7472 7588 7514
rect 9145 7486 9189 7528
rect 9239 7548 9281 7586
rect 9239 7528 9253 7548
rect 9273 7528 9281 7548
rect 9239 7486 9281 7528
rect 9363 7548 9407 7586
rect 9363 7528 9375 7548
rect 9395 7528 9407 7548
rect 9363 7486 9407 7528
rect 9457 7548 9499 7586
rect 9457 7528 9471 7548
rect 9491 7528 9499 7548
rect 9457 7486 9499 7528
rect 9573 7548 9615 7586
rect 9573 7528 9581 7548
rect 9601 7528 9615 7548
rect 9573 7486 9615 7528
rect 9665 7555 9710 7586
rect 9665 7548 9709 7555
rect 9665 7528 9677 7548
rect 9697 7528 9709 7548
rect 9665 7486 9709 7528
rect 20828 7679 20840 7699
rect 20860 7679 20872 7699
rect 20828 7672 20872 7679
rect 20827 7641 20872 7672
rect 20922 7699 20964 7741
rect 20922 7679 20936 7699
rect 20956 7679 20964 7699
rect 20922 7641 20964 7679
rect 21038 7699 21080 7741
rect 21038 7679 21046 7699
rect 21066 7679 21080 7699
rect 21038 7641 21080 7679
rect 21130 7699 21174 7741
rect 21130 7679 21142 7699
rect 21162 7679 21174 7699
rect 21130 7641 21174 7679
rect 21256 7699 21298 7741
rect 21256 7679 21264 7699
rect 21284 7679 21298 7699
rect 21256 7641 21298 7679
rect 21348 7699 21392 7741
rect 23036 7754 23048 7774
rect 23068 7754 23080 7774
rect 21348 7679 21360 7699
rect 21380 7679 21392 7699
rect 23036 7712 23080 7754
rect 23130 7774 23172 7812
rect 23130 7754 23144 7774
rect 23164 7754 23172 7774
rect 23130 7712 23172 7754
rect 23254 7774 23298 7812
rect 23254 7754 23266 7774
rect 23286 7754 23298 7774
rect 23254 7712 23298 7754
rect 23348 7774 23390 7812
rect 23348 7754 23362 7774
rect 23382 7754 23390 7774
rect 23348 7712 23390 7754
rect 23464 7774 23506 7812
rect 23464 7754 23472 7774
rect 23492 7754 23506 7774
rect 23464 7712 23506 7754
rect 23556 7781 23601 7812
rect 23556 7774 23600 7781
rect 23556 7754 23568 7774
rect 23588 7754 23600 7774
rect 27413 7786 27457 7824
rect 23556 7712 23600 7754
rect 25192 7712 25236 7754
rect 21348 7641 21392 7679
rect 13509 7561 13553 7599
rect 13509 7541 13521 7561
rect 13541 7541 13553 7561
rect 7544 7452 7556 7472
rect 7576 7452 7588 7472
rect 7544 7414 7588 7452
rect 5566 7352 5610 7390
rect 5566 7332 5578 7352
rect 5598 7332 5610 7352
rect 3458 7275 3502 7317
rect 3458 7255 3470 7275
rect 3490 7255 3502 7275
rect 3458 7248 3502 7255
rect 3457 7217 3502 7248
rect 3552 7275 3594 7317
rect 3552 7255 3566 7275
rect 3586 7255 3594 7275
rect 3552 7217 3594 7255
rect 3668 7275 3710 7317
rect 3668 7255 3676 7275
rect 3696 7255 3710 7275
rect 3668 7217 3710 7255
rect 3760 7275 3804 7317
rect 3760 7255 3772 7275
rect 3792 7255 3804 7275
rect 3760 7217 3804 7255
rect 3886 7275 3928 7317
rect 3886 7255 3894 7275
rect 3914 7255 3928 7275
rect 3886 7217 3928 7255
rect 3978 7275 4022 7317
rect 5566 7290 5610 7332
rect 5660 7352 5702 7390
rect 5660 7332 5674 7352
rect 5694 7332 5702 7352
rect 5660 7290 5702 7332
rect 5784 7352 5828 7390
rect 5784 7332 5796 7352
rect 5816 7332 5828 7352
rect 5784 7290 5828 7332
rect 5878 7352 5920 7390
rect 5878 7332 5892 7352
rect 5912 7332 5920 7352
rect 5878 7290 5920 7332
rect 5994 7352 6036 7390
rect 5994 7332 6002 7352
rect 6022 7332 6036 7352
rect 5994 7290 6036 7332
rect 6086 7359 6131 7390
rect 6086 7352 6130 7359
rect 6086 7332 6098 7352
rect 6118 7332 6130 7352
rect 6086 7290 6130 7332
rect 11401 7484 11445 7526
rect 11401 7464 11413 7484
rect 11433 7464 11445 7484
rect 11401 7457 11445 7464
rect 11400 7426 11445 7457
rect 11495 7484 11537 7526
rect 11495 7464 11509 7484
rect 11529 7464 11537 7484
rect 11495 7426 11537 7464
rect 11611 7484 11653 7526
rect 11611 7464 11619 7484
rect 11639 7464 11653 7484
rect 11611 7426 11653 7464
rect 11703 7484 11747 7526
rect 11703 7464 11715 7484
rect 11735 7464 11747 7484
rect 11703 7426 11747 7464
rect 11829 7484 11871 7526
rect 11829 7464 11837 7484
rect 11857 7464 11871 7484
rect 11829 7426 11871 7464
rect 11921 7484 11965 7526
rect 13509 7499 13553 7541
rect 13603 7561 13645 7599
rect 13603 7541 13617 7561
rect 13637 7541 13645 7561
rect 13603 7499 13645 7541
rect 13727 7561 13771 7599
rect 13727 7541 13739 7561
rect 13759 7541 13771 7561
rect 13727 7499 13771 7541
rect 13821 7561 13863 7599
rect 13821 7541 13835 7561
rect 13855 7541 13863 7561
rect 13821 7499 13863 7541
rect 13937 7561 13979 7599
rect 13937 7541 13945 7561
rect 13965 7541 13979 7561
rect 13937 7499 13979 7541
rect 14029 7568 14074 7599
rect 14029 7561 14073 7568
rect 14029 7541 14041 7561
rect 14061 7541 14073 7561
rect 14029 7499 14073 7541
rect 25192 7692 25204 7712
rect 25224 7692 25236 7712
rect 25192 7685 25236 7692
rect 25191 7654 25236 7685
rect 25286 7712 25328 7754
rect 25286 7692 25300 7712
rect 25320 7692 25328 7712
rect 25286 7654 25328 7692
rect 25402 7712 25444 7754
rect 25402 7692 25410 7712
rect 25430 7692 25444 7712
rect 25402 7654 25444 7692
rect 25494 7712 25538 7754
rect 25494 7692 25506 7712
rect 25526 7692 25538 7712
rect 25494 7654 25538 7692
rect 25620 7712 25662 7754
rect 25620 7692 25628 7712
rect 25648 7692 25662 7712
rect 25620 7654 25662 7692
rect 25712 7712 25756 7754
rect 27413 7766 27425 7786
rect 27445 7766 27457 7786
rect 25712 7692 25724 7712
rect 25744 7692 25756 7712
rect 27413 7724 27457 7766
rect 27507 7786 27549 7824
rect 27507 7766 27521 7786
rect 27541 7766 27549 7786
rect 27507 7724 27549 7766
rect 27631 7786 27675 7824
rect 27631 7766 27643 7786
rect 27663 7766 27675 7786
rect 27631 7724 27675 7766
rect 27725 7786 27767 7824
rect 27725 7766 27739 7786
rect 27759 7766 27767 7786
rect 27725 7724 27767 7766
rect 27841 7786 27883 7824
rect 27841 7766 27849 7786
rect 27869 7766 27883 7786
rect 27841 7724 27883 7766
rect 27933 7793 27978 7824
rect 27933 7786 27977 7793
rect 27933 7766 27945 7786
rect 27965 7766 27977 7786
rect 31777 7799 31821 7837
rect 27933 7724 27977 7766
rect 29569 7724 29613 7766
rect 25712 7654 25756 7692
rect 11921 7464 11933 7484
rect 11953 7464 11965 7484
rect 11921 7426 11965 7464
rect 9943 7364 9987 7402
rect 9943 7344 9955 7364
rect 9975 7344 9987 7364
rect 3978 7255 3990 7275
rect 4010 7255 4022 7275
rect 3978 7217 4022 7255
rect 7822 7288 7866 7330
rect 7822 7268 7834 7288
rect 7854 7268 7866 7288
rect 7822 7261 7866 7268
rect 7821 7230 7866 7261
rect 7916 7288 7958 7330
rect 7916 7268 7930 7288
rect 7950 7268 7958 7288
rect 7916 7230 7958 7268
rect 8032 7288 8074 7330
rect 8032 7268 8040 7288
rect 8060 7268 8074 7288
rect 8032 7230 8074 7268
rect 8124 7288 8168 7330
rect 8124 7268 8136 7288
rect 8156 7268 8168 7288
rect 8124 7230 8168 7268
rect 8250 7288 8292 7330
rect 8250 7268 8258 7288
rect 8278 7268 8292 7288
rect 8250 7230 8292 7268
rect 8342 7288 8386 7330
rect 9943 7302 9987 7344
rect 10037 7364 10079 7402
rect 10037 7344 10051 7364
rect 10071 7344 10079 7364
rect 10037 7302 10079 7344
rect 10161 7364 10205 7402
rect 10161 7344 10173 7364
rect 10193 7344 10205 7364
rect 10161 7302 10205 7344
rect 10255 7364 10297 7402
rect 10255 7344 10269 7364
rect 10289 7344 10297 7364
rect 10255 7302 10297 7344
rect 10371 7364 10413 7402
rect 10371 7344 10379 7364
rect 10399 7344 10413 7364
rect 10371 7302 10413 7344
rect 10463 7371 10508 7402
rect 10463 7364 10507 7371
rect 10463 7344 10475 7364
rect 10495 7344 10507 7364
rect 10463 7302 10507 7344
rect 15765 7497 15809 7539
rect 15765 7477 15777 7497
rect 15797 7477 15809 7497
rect 15765 7470 15809 7477
rect 15764 7439 15809 7470
rect 15859 7497 15901 7539
rect 15859 7477 15873 7497
rect 15893 7477 15901 7497
rect 15859 7439 15901 7477
rect 15975 7497 16017 7539
rect 15975 7477 15983 7497
rect 16003 7477 16017 7497
rect 15975 7439 16017 7477
rect 16067 7497 16111 7539
rect 16067 7477 16079 7497
rect 16099 7477 16111 7497
rect 16067 7439 16111 7477
rect 16193 7497 16235 7539
rect 16193 7477 16201 7497
rect 16221 7477 16235 7497
rect 16193 7439 16235 7477
rect 16285 7497 16329 7539
rect 17775 7535 17819 7573
rect 17775 7515 17787 7535
rect 17807 7515 17819 7535
rect 16285 7477 16297 7497
rect 16317 7477 16329 7497
rect 16285 7439 16329 7477
rect 17775 7473 17819 7515
rect 17869 7535 17911 7573
rect 17869 7515 17883 7535
rect 17903 7515 17911 7535
rect 17869 7473 17911 7515
rect 17993 7535 18037 7573
rect 17993 7515 18005 7535
rect 18025 7515 18037 7535
rect 17993 7473 18037 7515
rect 18087 7535 18129 7573
rect 18087 7515 18101 7535
rect 18121 7515 18129 7535
rect 18087 7473 18129 7515
rect 18203 7535 18245 7573
rect 18203 7515 18211 7535
rect 18231 7515 18245 7535
rect 18203 7473 18245 7515
rect 18295 7542 18340 7573
rect 18295 7535 18339 7542
rect 18295 7515 18307 7535
rect 18327 7515 18339 7535
rect 18295 7473 18339 7515
rect 29569 7704 29581 7724
rect 29601 7704 29613 7724
rect 29569 7697 29613 7704
rect 29568 7666 29613 7697
rect 29663 7724 29705 7766
rect 29663 7704 29677 7724
rect 29697 7704 29705 7724
rect 29663 7666 29705 7704
rect 29779 7724 29821 7766
rect 29779 7704 29787 7724
rect 29807 7704 29821 7724
rect 29779 7666 29821 7704
rect 29871 7724 29915 7766
rect 29871 7704 29883 7724
rect 29903 7704 29915 7724
rect 29871 7666 29915 7704
rect 29997 7724 30039 7766
rect 29997 7704 30005 7724
rect 30025 7704 30039 7724
rect 29997 7666 30039 7704
rect 30089 7724 30133 7766
rect 31777 7779 31789 7799
rect 31809 7779 31821 7799
rect 30089 7704 30101 7724
rect 30121 7704 30133 7724
rect 31777 7737 31821 7779
rect 31871 7799 31913 7837
rect 31871 7779 31885 7799
rect 31905 7779 31913 7799
rect 31871 7737 31913 7779
rect 31995 7799 32039 7837
rect 31995 7779 32007 7799
rect 32027 7779 32039 7799
rect 31995 7737 32039 7779
rect 32089 7799 32131 7837
rect 32089 7779 32103 7799
rect 32123 7779 32131 7799
rect 32089 7737 32131 7779
rect 32205 7799 32247 7837
rect 32205 7779 32213 7799
rect 32233 7779 32247 7799
rect 32205 7737 32247 7779
rect 32297 7806 32342 7837
rect 32297 7799 32341 7806
rect 32297 7779 32309 7799
rect 32329 7779 32341 7799
rect 32297 7737 32341 7779
rect 33933 7737 33977 7779
rect 30089 7666 30133 7704
rect 22139 7548 22183 7586
rect 22139 7528 22151 7548
rect 22171 7528 22183 7548
rect 14307 7377 14351 7415
rect 14307 7357 14319 7377
rect 14339 7357 14351 7377
rect 8342 7268 8354 7288
rect 8374 7268 8386 7288
rect 8342 7230 8386 7268
rect 405 7111 449 7149
rect 405 7091 417 7111
rect 437 7091 449 7111
rect 405 7049 449 7091
rect 499 7111 541 7149
rect 499 7091 513 7111
rect 533 7091 541 7111
rect 499 7049 541 7091
rect 623 7111 667 7149
rect 623 7091 635 7111
rect 655 7091 667 7111
rect 623 7049 667 7091
rect 717 7111 759 7149
rect 717 7091 731 7111
rect 751 7091 759 7111
rect 717 7049 759 7091
rect 833 7111 875 7149
rect 833 7091 841 7111
rect 861 7091 875 7111
rect 833 7049 875 7091
rect 925 7118 970 7149
rect 925 7111 969 7118
rect 925 7091 937 7111
rect 957 7091 969 7111
rect 12199 7300 12243 7342
rect 12199 7280 12211 7300
rect 12231 7280 12243 7300
rect 12199 7273 12243 7280
rect 12198 7242 12243 7273
rect 12293 7300 12335 7342
rect 12293 7280 12307 7300
rect 12327 7280 12335 7300
rect 12293 7242 12335 7280
rect 12409 7300 12451 7342
rect 12409 7280 12417 7300
rect 12437 7280 12451 7300
rect 12409 7242 12451 7280
rect 12501 7300 12545 7342
rect 12501 7280 12513 7300
rect 12533 7280 12545 7300
rect 12501 7242 12545 7280
rect 12627 7300 12669 7342
rect 12627 7280 12635 7300
rect 12655 7280 12669 7300
rect 12627 7242 12669 7280
rect 12719 7300 12763 7342
rect 14307 7315 14351 7357
rect 14401 7377 14443 7415
rect 14401 7357 14415 7377
rect 14435 7357 14443 7377
rect 14401 7315 14443 7357
rect 14525 7377 14569 7415
rect 14525 7357 14537 7377
rect 14557 7357 14569 7377
rect 14525 7315 14569 7357
rect 14619 7377 14661 7415
rect 14619 7357 14633 7377
rect 14653 7357 14661 7377
rect 14619 7315 14661 7357
rect 14735 7377 14777 7415
rect 14735 7357 14743 7377
rect 14763 7357 14777 7377
rect 14735 7315 14777 7357
rect 14827 7384 14872 7415
rect 14827 7377 14871 7384
rect 14827 7357 14839 7377
rect 14859 7357 14871 7377
rect 14827 7315 14871 7357
rect 20031 7471 20075 7513
rect 20031 7451 20043 7471
rect 20063 7451 20075 7471
rect 20031 7444 20075 7451
rect 20030 7413 20075 7444
rect 20125 7471 20167 7513
rect 20125 7451 20139 7471
rect 20159 7451 20167 7471
rect 20125 7413 20167 7451
rect 20241 7471 20283 7513
rect 20241 7451 20249 7471
rect 20269 7451 20283 7471
rect 20241 7413 20283 7451
rect 20333 7471 20377 7513
rect 20333 7451 20345 7471
rect 20365 7451 20377 7471
rect 20333 7413 20377 7451
rect 20459 7471 20501 7513
rect 20459 7451 20467 7471
rect 20487 7451 20501 7471
rect 20459 7413 20501 7451
rect 20551 7471 20595 7513
rect 22139 7486 22183 7528
rect 22233 7548 22275 7586
rect 22233 7528 22247 7548
rect 22267 7528 22275 7548
rect 22233 7486 22275 7528
rect 22357 7548 22401 7586
rect 22357 7528 22369 7548
rect 22389 7528 22401 7548
rect 22357 7486 22401 7528
rect 22451 7548 22493 7586
rect 22451 7528 22465 7548
rect 22485 7528 22493 7548
rect 22451 7486 22493 7528
rect 22567 7548 22609 7586
rect 22567 7528 22575 7548
rect 22595 7528 22609 7548
rect 22567 7486 22609 7528
rect 22659 7555 22704 7586
rect 22659 7548 22703 7555
rect 22659 7528 22671 7548
rect 22691 7528 22703 7548
rect 22659 7486 22703 7528
rect 33933 7717 33945 7737
rect 33965 7717 33977 7737
rect 33933 7710 33977 7717
rect 33932 7679 33977 7710
rect 34027 7737 34069 7779
rect 34027 7717 34041 7737
rect 34061 7717 34069 7737
rect 34027 7679 34069 7717
rect 34143 7737 34185 7779
rect 34143 7717 34151 7737
rect 34171 7717 34185 7737
rect 34143 7679 34185 7717
rect 34235 7737 34279 7779
rect 34235 7717 34247 7737
rect 34267 7717 34279 7737
rect 34235 7679 34279 7717
rect 34361 7737 34403 7779
rect 34361 7717 34369 7737
rect 34389 7717 34403 7737
rect 34361 7679 34403 7717
rect 34453 7737 34497 7779
rect 34453 7717 34465 7737
rect 34485 7717 34497 7737
rect 34453 7679 34497 7717
rect 26516 7560 26560 7598
rect 26516 7540 26528 7560
rect 26548 7540 26560 7560
rect 20551 7451 20563 7471
rect 20583 7451 20595 7471
rect 20551 7413 20595 7451
rect 12719 7280 12731 7300
rect 12751 7280 12763 7300
rect 12719 7242 12763 7280
rect 4769 7124 4813 7162
rect 925 7049 969 7091
rect 2495 7051 2539 7093
rect 2495 7031 2507 7051
rect 2527 7031 2539 7051
rect 2495 7024 2539 7031
rect 2494 6993 2539 7024
rect 2589 7051 2631 7093
rect 2589 7031 2603 7051
rect 2623 7031 2631 7051
rect 2589 6993 2631 7031
rect 2705 7051 2747 7093
rect 2705 7031 2713 7051
rect 2733 7031 2747 7051
rect 2705 6993 2747 7031
rect 2797 7051 2841 7093
rect 2797 7031 2809 7051
rect 2829 7031 2841 7051
rect 2797 6993 2841 7031
rect 2923 7051 2965 7093
rect 2923 7031 2931 7051
rect 2951 7031 2965 7051
rect 2923 6993 2965 7031
rect 3015 7051 3059 7093
rect 4769 7104 4781 7124
rect 4801 7104 4813 7124
rect 3015 7031 3027 7051
rect 3047 7031 3059 7051
rect 4769 7062 4813 7104
rect 4863 7124 4905 7162
rect 4863 7104 4877 7124
rect 4897 7104 4905 7124
rect 4863 7062 4905 7104
rect 4987 7124 5031 7162
rect 4987 7104 4999 7124
rect 5019 7104 5031 7124
rect 4987 7062 5031 7104
rect 5081 7124 5123 7162
rect 5081 7104 5095 7124
rect 5115 7104 5123 7124
rect 5081 7062 5123 7104
rect 5197 7124 5239 7162
rect 5197 7104 5205 7124
rect 5225 7104 5239 7124
rect 5197 7062 5239 7104
rect 5289 7131 5334 7162
rect 5289 7124 5333 7131
rect 5289 7104 5301 7124
rect 5321 7104 5333 7124
rect 16563 7313 16607 7355
rect 16563 7293 16575 7313
rect 16595 7293 16607 7313
rect 16563 7286 16607 7293
rect 16562 7255 16607 7286
rect 16657 7313 16699 7355
rect 16657 7293 16671 7313
rect 16691 7293 16699 7313
rect 16657 7255 16699 7293
rect 16773 7313 16815 7355
rect 16773 7293 16781 7313
rect 16801 7293 16815 7313
rect 16773 7255 16815 7293
rect 16865 7313 16909 7355
rect 16865 7293 16877 7313
rect 16897 7293 16909 7313
rect 16865 7255 16909 7293
rect 16991 7313 17033 7355
rect 16991 7293 16999 7313
rect 17019 7293 17033 7313
rect 16991 7255 17033 7293
rect 17083 7313 17127 7355
rect 18573 7351 18617 7389
rect 18573 7331 18585 7351
rect 18605 7331 18617 7351
rect 17083 7293 17095 7313
rect 17115 7293 17127 7313
rect 17083 7255 17127 7293
rect 18573 7289 18617 7331
rect 18667 7351 18709 7389
rect 18667 7331 18681 7351
rect 18701 7331 18709 7351
rect 18667 7289 18709 7331
rect 18791 7351 18835 7389
rect 18791 7331 18803 7351
rect 18823 7331 18835 7351
rect 18791 7289 18835 7331
rect 18885 7351 18927 7389
rect 18885 7331 18899 7351
rect 18919 7331 18927 7351
rect 18885 7289 18927 7331
rect 19001 7351 19043 7389
rect 19001 7331 19009 7351
rect 19029 7331 19043 7351
rect 19001 7289 19043 7331
rect 19093 7358 19138 7389
rect 19093 7351 19137 7358
rect 19093 7331 19105 7351
rect 19125 7331 19137 7351
rect 19093 7289 19137 7331
rect 24395 7484 24439 7526
rect 24395 7464 24407 7484
rect 24427 7464 24439 7484
rect 24395 7457 24439 7464
rect 24394 7426 24439 7457
rect 24489 7484 24531 7526
rect 24489 7464 24503 7484
rect 24523 7464 24531 7484
rect 24489 7426 24531 7464
rect 24605 7484 24647 7526
rect 24605 7464 24613 7484
rect 24633 7464 24647 7484
rect 24605 7426 24647 7464
rect 24697 7484 24741 7526
rect 24697 7464 24709 7484
rect 24729 7464 24741 7484
rect 24697 7426 24741 7464
rect 24823 7484 24865 7526
rect 24823 7464 24831 7484
rect 24851 7464 24865 7484
rect 24823 7426 24865 7464
rect 24915 7484 24959 7526
rect 26516 7498 26560 7540
rect 26610 7560 26652 7598
rect 26610 7540 26624 7560
rect 26644 7540 26652 7560
rect 26610 7498 26652 7540
rect 26734 7560 26778 7598
rect 26734 7540 26746 7560
rect 26766 7540 26778 7560
rect 26734 7498 26778 7540
rect 26828 7560 26870 7598
rect 26828 7540 26842 7560
rect 26862 7540 26870 7560
rect 26828 7498 26870 7540
rect 26944 7560 26986 7598
rect 26944 7540 26952 7560
rect 26972 7540 26986 7560
rect 26944 7498 26986 7540
rect 27036 7567 27081 7598
rect 27036 7560 27080 7567
rect 27036 7540 27048 7560
rect 27068 7540 27080 7560
rect 27036 7498 27080 7540
rect 30880 7573 30924 7611
rect 30880 7553 30892 7573
rect 30912 7553 30924 7573
rect 24915 7464 24927 7484
rect 24947 7464 24959 7484
rect 24915 7426 24959 7464
rect 22937 7364 22981 7402
rect 22937 7344 22949 7364
rect 22969 7344 22981 7364
rect 9146 7136 9190 7174
rect 5289 7062 5333 7104
rect 6859 7064 6903 7106
rect 3015 6993 3059 7031
rect 6859 7044 6871 7064
rect 6891 7044 6903 7064
rect 6859 7037 6903 7044
rect 6858 7006 6903 7037
rect 6953 7064 6995 7106
rect 6953 7044 6967 7064
rect 6987 7044 6995 7064
rect 6953 7006 6995 7044
rect 7069 7064 7111 7106
rect 7069 7044 7077 7064
rect 7097 7044 7111 7064
rect 7069 7006 7111 7044
rect 7161 7064 7205 7106
rect 7161 7044 7173 7064
rect 7193 7044 7205 7064
rect 7161 7006 7205 7044
rect 7287 7064 7329 7106
rect 7287 7044 7295 7064
rect 7315 7044 7329 7064
rect 7287 7006 7329 7044
rect 7379 7064 7423 7106
rect 9146 7116 9158 7136
rect 9178 7116 9190 7136
rect 7379 7044 7391 7064
rect 7411 7044 7423 7064
rect 9146 7074 9190 7116
rect 9240 7136 9282 7174
rect 9240 7116 9254 7136
rect 9274 7116 9282 7136
rect 9240 7074 9282 7116
rect 9364 7136 9408 7174
rect 9364 7116 9376 7136
rect 9396 7116 9408 7136
rect 9364 7074 9408 7116
rect 9458 7136 9500 7174
rect 9458 7116 9472 7136
rect 9492 7116 9500 7136
rect 9458 7074 9500 7116
rect 9574 7136 9616 7174
rect 9574 7116 9582 7136
rect 9602 7116 9616 7136
rect 9574 7074 9616 7116
rect 9666 7143 9711 7174
rect 9666 7136 9710 7143
rect 9666 7116 9678 7136
rect 9698 7116 9710 7136
rect 20829 7287 20873 7329
rect 20829 7267 20841 7287
rect 20861 7267 20873 7287
rect 20829 7260 20873 7267
rect 20828 7229 20873 7260
rect 20923 7287 20965 7329
rect 20923 7267 20937 7287
rect 20957 7267 20965 7287
rect 20923 7229 20965 7267
rect 21039 7287 21081 7329
rect 21039 7267 21047 7287
rect 21067 7267 21081 7287
rect 21039 7229 21081 7267
rect 21131 7287 21175 7329
rect 21131 7267 21143 7287
rect 21163 7267 21175 7287
rect 21131 7229 21175 7267
rect 21257 7287 21299 7329
rect 21257 7267 21265 7287
rect 21285 7267 21299 7287
rect 21257 7229 21299 7267
rect 21349 7287 21393 7329
rect 22937 7302 22981 7344
rect 23031 7364 23073 7402
rect 23031 7344 23045 7364
rect 23065 7344 23073 7364
rect 23031 7302 23073 7344
rect 23155 7364 23199 7402
rect 23155 7344 23167 7364
rect 23187 7344 23199 7364
rect 23155 7302 23199 7344
rect 23249 7364 23291 7402
rect 23249 7344 23263 7364
rect 23283 7344 23291 7364
rect 23249 7302 23291 7344
rect 23365 7364 23407 7402
rect 23365 7344 23373 7364
rect 23393 7344 23407 7364
rect 23365 7302 23407 7344
rect 23457 7371 23502 7402
rect 23457 7364 23501 7371
rect 23457 7344 23469 7364
rect 23489 7344 23501 7364
rect 23457 7302 23501 7344
rect 28772 7496 28816 7538
rect 28772 7476 28784 7496
rect 28804 7476 28816 7496
rect 28772 7469 28816 7476
rect 28771 7438 28816 7469
rect 28866 7496 28908 7538
rect 28866 7476 28880 7496
rect 28900 7476 28908 7496
rect 28866 7438 28908 7476
rect 28982 7496 29024 7538
rect 28982 7476 28990 7496
rect 29010 7476 29024 7496
rect 28982 7438 29024 7476
rect 29074 7496 29118 7538
rect 29074 7476 29086 7496
rect 29106 7476 29118 7496
rect 29074 7438 29118 7476
rect 29200 7496 29242 7538
rect 29200 7476 29208 7496
rect 29228 7476 29242 7496
rect 29200 7438 29242 7476
rect 29292 7496 29336 7538
rect 30880 7511 30924 7553
rect 30974 7573 31016 7611
rect 30974 7553 30988 7573
rect 31008 7553 31016 7573
rect 30974 7511 31016 7553
rect 31098 7573 31142 7611
rect 31098 7553 31110 7573
rect 31130 7553 31142 7573
rect 31098 7511 31142 7553
rect 31192 7573 31234 7611
rect 31192 7553 31206 7573
rect 31226 7553 31234 7573
rect 31192 7511 31234 7553
rect 31308 7573 31350 7611
rect 31308 7553 31316 7573
rect 31336 7553 31350 7573
rect 31308 7511 31350 7553
rect 31400 7580 31445 7611
rect 31400 7573 31444 7580
rect 31400 7553 31412 7573
rect 31432 7553 31444 7573
rect 31400 7511 31444 7553
rect 29292 7476 29304 7496
rect 29324 7476 29336 7496
rect 29292 7438 29336 7476
rect 27314 7376 27358 7414
rect 27314 7356 27326 7376
rect 27346 7356 27358 7376
rect 21349 7267 21361 7287
rect 21381 7267 21393 7287
rect 21349 7229 21393 7267
rect 13510 7149 13554 7187
rect 9666 7074 9710 7116
rect 11236 7076 11280 7118
rect 7379 7006 7423 7044
rect 11236 7056 11248 7076
rect 11268 7056 11280 7076
rect 11236 7049 11280 7056
rect 11235 7018 11280 7049
rect 11330 7076 11372 7118
rect 11330 7056 11344 7076
rect 11364 7056 11372 7076
rect 11330 7018 11372 7056
rect 11446 7076 11488 7118
rect 11446 7056 11454 7076
rect 11474 7056 11488 7076
rect 11446 7018 11488 7056
rect 11538 7076 11582 7118
rect 11538 7056 11550 7076
rect 11570 7056 11582 7076
rect 11538 7018 11582 7056
rect 11664 7076 11706 7118
rect 11664 7056 11672 7076
rect 11692 7056 11706 7076
rect 11664 7018 11706 7056
rect 11756 7076 11800 7118
rect 13510 7129 13522 7149
rect 13542 7129 13554 7149
rect 11756 7056 11768 7076
rect 11788 7056 11800 7076
rect 13510 7087 13554 7129
rect 13604 7149 13646 7187
rect 13604 7129 13618 7149
rect 13638 7129 13646 7149
rect 13604 7087 13646 7129
rect 13728 7149 13772 7187
rect 13728 7129 13740 7149
rect 13760 7129 13772 7149
rect 13728 7087 13772 7129
rect 13822 7149 13864 7187
rect 13822 7129 13836 7149
rect 13856 7129 13864 7149
rect 13822 7087 13864 7129
rect 13938 7149 13980 7187
rect 13938 7129 13946 7149
rect 13966 7129 13980 7149
rect 13938 7087 13980 7129
rect 14030 7156 14075 7187
rect 14030 7149 14074 7156
rect 14030 7129 14042 7149
rect 14062 7129 14074 7149
rect 25193 7300 25237 7342
rect 25193 7280 25205 7300
rect 25225 7280 25237 7300
rect 25193 7273 25237 7280
rect 25192 7242 25237 7273
rect 25287 7300 25329 7342
rect 25287 7280 25301 7300
rect 25321 7280 25329 7300
rect 25287 7242 25329 7280
rect 25403 7300 25445 7342
rect 25403 7280 25411 7300
rect 25431 7280 25445 7300
rect 25403 7242 25445 7280
rect 25495 7300 25539 7342
rect 25495 7280 25507 7300
rect 25527 7280 25539 7300
rect 25495 7242 25539 7280
rect 25621 7300 25663 7342
rect 25621 7280 25629 7300
rect 25649 7280 25663 7300
rect 25621 7242 25663 7280
rect 25713 7300 25757 7342
rect 27314 7314 27358 7356
rect 27408 7376 27450 7414
rect 27408 7356 27422 7376
rect 27442 7356 27450 7376
rect 27408 7314 27450 7356
rect 27532 7376 27576 7414
rect 27532 7356 27544 7376
rect 27564 7356 27576 7376
rect 27532 7314 27576 7356
rect 27626 7376 27668 7414
rect 27626 7356 27640 7376
rect 27660 7356 27668 7376
rect 27626 7314 27668 7356
rect 27742 7376 27784 7414
rect 27742 7356 27750 7376
rect 27770 7356 27784 7376
rect 27742 7314 27784 7356
rect 27834 7383 27879 7414
rect 27834 7376 27878 7383
rect 27834 7356 27846 7376
rect 27866 7356 27878 7376
rect 27834 7314 27878 7356
rect 33136 7509 33180 7551
rect 33136 7489 33148 7509
rect 33168 7489 33180 7509
rect 33136 7482 33180 7489
rect 33135 7451 33180 7482
rect 33230 7509 33272 7551
rect 33230 7489 33244 7509
rect 33264 7489 33272 7509
rect 33230 7451 33272 7489
rect 33346 7509 33388 7551
rect 33346 7489 33354 7509
rect 33374 7489 33388 7509
rect 33346 7451 33388 7489
rect 33438 7509 33482 7551
rect 33438 7489 33450 7509
rect 33470 7489 33482 7509
rect 33438 7451 33482 7489
rect 33564 7509 33606 7551
rect 33564 7489 33572 7509
rect 33592 7489 33606 7509
rect 33564 7451 33606 7489
rect 33656 7509 33700 7551
rect 33656 7489 33668 7509
rect 33688 7489 33700 7509
rect 33656 7451 33700 7489
rect 31678 7389 31722 7427
rect 31678 7369 31690 7389
rect 31710 7369 31722 7389
rect 25713 7280 25725 7300
rect 25745 7280 25757 7300
rect 25713 7242 25757 7280
rect 14030 7087 14074 7129
rect 15600 7089 15644 7131
rect 11756 7018 11800 7056
rect 15600 7069 15612 7089
rect 15632 7069 15644 7089
rect 15600 7062 15644 7069
rect 15599 7031 15644 7062
rect 15694 7089 15736 7131
rect 15694 7069 15708 7089
rect 15728 7069 15736 7089
rect 15694 7031 15736 7069
rect 15810 7089 15852 7131
rect 15810 7069 15818 7089
rect 15838 7069 15852 7089
rect 15810 7031 15852 7069
rect 15902 7089 15946 7131
rect 15902 7069 15914 7089
rect 15934 7069 15946 7089
rect 15902 7031 15946 7069
rect 16028 7089 16070 7131
rect 16028 7069 16036 7089
rect 16056 7069 16070 7089
rect 16028 7031 16070 7069
rect 16120 7089 16164 7131
rect 16120 7069 16132 7089
rect 16152 7069 16164 7089
rect 17776 7123 17820 7161
rect 17776 7103 17788 7123
rect 17808 7103 17820 7123
rect 16120 7031 16164 7069
rect 17776 7061 17820 7103
rect 17870 7123 17912 7161
rect 17870 7103 17884 7123
rect 17904 7103 17912 7123
rect 17870 7061 17912 7103
rect 17994 7123 18038 7161
rect 17994 7103 18006 7123
rect 18026 7103 18038 7123
rect 17994 7061 18038 7103
rect 18088 7123 18130 7161
rect 18088 7103 18102 7123
rect 18122 7103 18130 7123
rect 18088 7061 18130 7103
rect 18204 7123 18246 7161
rect 18204 7103 18212 7123
rect 18232 7103 18246 7123
rect 18204 7061 18246 7103
rect 18296 7130 18341 7161
rect 18296 7123 18340 7130
rect 18296 7103 18308 7123
rect 18328 7103 18340 7123
rect 29570 7312 29614 7354
rect 29570 7292 29582 7312
rect 29602 7292 29614 7312
rect 29570 7285 29614 7292
rect 29569 7254 29614 7285
rect 29664 7312 29706 7354
rect 29664 7292 29678 7312
rect 29698 7292 29706 7312
rect 29664 7254 29706 7292
rect 29780 7312 29822 7354
rect 29780 7292 29788 7312
rect 29808 7292 29822 7312
rect 29780 7254 29822 7292
rect 29872 7312 29916 7354
rect 29872 7292 29884 7312
rect 29904 7292 29916 7312
rect 29872 7254 29916 7292
rect 29998 7312 30040 7354
rect 29998 7292 30006 7312
rect 30026 7292 30040 7312
rect 29998 7254 30040 7292
rect 30090 7312 30134 7354
rect 31678 7327 31722 7369
rect 31772 7389 31814 7427
rect 31772 7369 31786 7389
rect 31806 7369 31814 7389
rect 31772 7327 31814 7369
rect 31896 7389 31940 7427
rect 31896 7369 31908 7389
rect 31928 7369 31940 7389
rect 31896 7327 31940 7369
rect 31990 7389 32032 7427
rect 31990 7369 32004 7389
rect 32024 7369 32032 7389
rect 31990 7327 32032 7369
rect 32106 7389 32148 7427
rect 32106 7369 32114 7389
rect 32134 7369 32148 7389
rect 32106 7327 32148 7369
rect 32198 7396 32243 7427
rect 32198 7389 32242 7396
rect 32198 7369 32210 7389
rect 32230 7369 32242 7389
rect 32198 7327 32242 7369
rect 30090 7292 30102 7312
rect 30122 7292 30134 7312
rect 30090 7254 30134 7292
rect 22140 7136 22184 7174
rect 18296 7061 18340 7103
rect 19866 7063 19910 7105
rect 19866 7043 19878 7063
rect 19898 7043 19910 7063
rect 19866 7036 19910 7043
rect 19865 7005 19910 7036
rect 19960 7063 20002 7105
rect 19960 7043 19974 7063
rect 19994 7043 20002 7063
rect 19960 7005 20002 7043
rect 20076 7063 20118 7105
rect 20076 7043 20084 7063
rect 20104 7043 20118 7063
rect 20076 7005 20118 7043
rect 20168 7063 20212 7105
rect 20168 7043 20180 7063
rect 20200 7043 20212 7063
rect 20168 7005 20212 7043
rect 20294 7063 20336 7105
rect 20294 7043 20302 7063
rect 20322 7043 20336 7063
rect 20294 7005 20336 7043
rect 20386 7063 20430 7105
rect 22140 7116 22152 7136
rect 22172 7116 22184 7136
rect 20386 7043 20398 7063
rect 20418 7043 20430 7063
rect 22140 7074 22184 7116
rect 22234 7136 22276 7174
rect 22234 7116 22248 7136
rect 22268 7116 22276 7136
rect 22234 7074 22276 7116
rect 22358 7136 22402 7174
rect 22358 7116 22370 7136
rect 22390 7116 22402 7136
rect 22358 7074 22402 7116
rect 22452 7136 22494 7174
rect 22452 7116 22466 7136
rect 22486 7116 22494 7136
rect 22452 7074 22494 7116
rect 22568 7136 22610 7174
rect 22568 7116 22576 7136
rect 22596 7116 22610 7136
rect 22568 7074 22610 7116
rect 22660 7143 22705 7174
rect 22660 7136 22704 7143
rect 22660 7116 22672 7136
rect 22692 7116 22704 7136
rect 33934 7325 33978 7367
rect 33934 7305 33946 7325
rect 33966 7305 33978 7325
rect 33934 7298 33978 7305
rect 33933 7267 33978 7298
rect 34028 7325 34070 7367
rect 34028 7305 34042 7325
rect 34062 7305 34070 7325
rect 34028 7267 34070 7305
rect 34144 7325 34186 7367
rect 34144 7305 34152 7325
rect 34172 7305 34186 7325
rect 34144 7267 34186 7305
rect 34236 7325 34280 7367
rect 34236 7305 34248 7325
rect 34268 7305 34280 7325
rect 34236 7267 34280 7305
rect 34362 7325 34404 7367
rect 34362 7305 34370 7325
rect 34390 7305 34404 7325
rect 34362 7267 34404 7305
rect 34454 7325 34498 7367
rect 34454 7305 34466 7325
rect 34486 7305 34498 7325
rect 34454 7267 34498 7305
rect 26517 7148 26561 7186
rect 22660 7074 22704 7116
rect 24230 7076 24274 7118
rect 20386 7005 20430 7043
rect 24230 7056 24242 7076
rect 24262 7056 24274 7076
rect 24230 7049 24274 7056
rect 24229 7018 24274 7049
rect 24324 7076 24366 7118
rect 24324 7056 24338 7076
rect 24358 7056 24366 7076
rect 24324 7018 24366 7056
rect 24440 7076 24482 7118
rect 24440 7056 24448 7076
rect 24468 7056 24482 7076
rect 24440 7018 24482 7056
rect 24532 7076 24576 7118
rect 24532 7056 24544 7076
rect 24564 7056 24576 7076
rect 24532 7018 24576 7056
rect 24658 7076 24700 7118
rect 24658 7056 24666 7076
rect 24686 7056 24700 7076
rect 24658 7018 24700 7056
rect 24750 7076 24794 7118
rect 26517 7128 26529 7148
rect 26549 7128 26561 7148
rect 24750 7056 24762 7076
rect 24782 7056 24794 7076
rect 26517 7086 26561 7128
rect 26611 7148 26653 7186
rect 26611 7128 26625 7148
rect 26645 7128 26653 7148
rect 26611 7086 26653 7128
rect 26735 7148 26779 7186
rect 26735 7128 26747 7148
rect 26767 7128 26779 7148
rect 26735 7086 26779 7128
rect 26829 7148 26871 7186
rect 26829 7128 26843 7148
rect 26863 7128 26871 7148
rect 26829 7086 26871 7128
rect 26945 7148 26987 7186
rect 26945 7128 26953 7148
rect 26973 7128 26987 7148
rect 26945 7086 26987 7128
rect 27037 7155 27082 7186
rect 27037 7148 27081 7155
rect 27037 7128 27049 7148
rect 27069 7128 27081 7148
rect 30881 7161 30925 7199
rect 27037 7086 27081 7128
rect 28607 7088 28651 7130
rect 24750 7018 24794 7056
rect 28607 7068 28619 7088
rect 28639 7068 28651 7088
rect 28607 7061 28651 7068
rect 28606 7030 28651 7061
rect 28701 7088 28743 7130
rect 28701 7068 28715 7088
rect 28735 7068 28743 7088
rect 28701 7030 28743 7068
rect 28817 7088 28859 7130
rect 28817 7068 28825 7088
rect 28845 7068 28859 7088
rect 28817 7030 28859 7068
rect 28909 7088 28953 7130
rect 28909 7068 28921 7088
rect 28941 7068 28953 7088
rect 28909 7030 28953 7068
rect 29035 7088 29077 7130
rect 29035 7068 29043 7088
rect 29063 7068 29077 7088
rect 29035 7030 29077 7068
rect 29127 7088 29171 7130
rect 30881 7141 30893 7161
rect 30913 7141 30925 7161
rect 29127 7068 29139 7088
rect 29159 7068 29171 7088
rect 30881 7099 30925 7141
rect 30975 7161 31017 7199
rect 30975 7141 30989 7161
rect 31009 7141 31017 7161
rect 30975 7099 31017 7141
rect 31099 7161 31143 7199
rect 31099 7141 31111 7161
rect 31131 7141 31143 7161
rect 31099 7099 31143 7141
rect 31193 7161 31235 7199
rect 31193 7141 31207 7161
rect 31227 7141 31235 7161
rect 31193 7099 31235 7141
rect 31309 7161 31351 7199
rect 31309 7141 31317 7161
rect 31337 7141 31351 7161
rect 31309 7099 31351 7141
rect 31401 7168 31446 7199
rect 31401 7161 31445 7168
rect 31401 7141 31413 7161
rect 31433 7141 31445 7161
rect 31401 7099 31445 7141
rect 32971 7101 33015 7143
rect 29127 7030 29171 7068
rect 32971 7081 32983 7101
rect 33003 7081 33015 7101
rect 32971 7074 33015 7081
rect 32970 7043 33015 7074
rect 33065 7101 33107 7143
rect 33065 7081 33079 7101
rect 33099 7081 33107 7101
rect 33065 7043 33107 7081
rect 33181 7101 33223 7143
rect 33181 7081 33189 7101
rect 33209 7081 33223 7101
rect 33181 7043 33223 7081
rect 33273 7101 33317 7143
rect 33273 7081 33285 7101
rect 33305 7081 33317 7101
rect 33273 7043 33317 7081
rect 33399 7101 33441 7143
rect 33399 7081 33407 7101
rect 33427 7081 33441 7101
rect 33399 7043 33441 7081
rect 33491 7101 33535 7143
rect 33491 7081 33503 7101
rect 33523 7081 33535 7101
rect 33491 7043 33535 7081
rect 1347 6729 1391 6767
rect 1347 6709 1359 6729
rect 1379 6709 1391 6729
rect 1347 6667 1391 6709
rect 1441 6729 1483 6767
rect 1441 6709 1455 6729
rect 1475 6709 1483 6729
rect 1441 6667 1483 6709
rect 1565 6729 1609 6767
rect 1565 6709 1577 6729
rect 1597 6709 1609 6729
rect 1565 6667 1609 6709
rect 1659 6729 1701 6767
rect 1659 6709 1673 6729
rect 1693 6709 1701 6729
rect 1659 6667 1701 6709
rect 1775 6729 1817 6767
rect 1775 6709 1783 6729
rect 1803 6709 1817 6729
rect 1775 6667 1817 6709
rect 1867 6736 1912 6767
rect 1867 6729 1911 6736
rect 1867 6709 1879 6729
rect 1899 6709 1911 6729
rect 5711 6742 5755 6780
rect 1867 6667 1911 6709
rect 3437 6669 3481 6711
rect 3437 6649 3449 6669
rect 3469 6649 3481 6669
rect 3437 6642 3481 6649
rect 3436 6611 3481 6642
rect 3531 6669 3573 6711
rect 3531 6649 3545 6669
rect 3565 6649 3573 6669
rect 3531 6611 3573 6649
rect 3647 6669 3689 6711
rect 3647 6649 3655 6669
rect 3675 6649 3689 6669
rect 3647 6611 3689 6649
rect 3739 6669 3783 6711
rect 3739 6649 3751 6669
rect 3771 6649 3783 6669
rect 3739 6611 3783 6649
rect 3865 6669 3907 6711
rect 3865 6649 3873 6669
rect 3893 6649 3907 6669
rect 3865 6611 3907 6649
rect 3957 6669 4001 6711
rect 5711 6722 5723 6742
rect 5743 6722 5755 6742
rect 3957 6649 3969 6669
rect 3989 6649 4001 6669
rect 5711 6680 5755 6722
rect 5805 6742 5847 6780
rect 5805 6722 5819 6742
rect 5839 6722 5847 6742
rect 5805 6680 5847 6722
rect 5929 6742 5973 6780
rect 5929 6722 5941 6742
rect 5961 6722 5973 6742
rect 5929 6680 5973 6722
rect 6023 6742 6065 6780
rect 6023 6722 6037 6742
rect 6057 6722 6065 6742
rect 6023 6680 6065 6722
rect 6139 6742 6181 6780
rect 6139 6722 6147 6742
rect 6167 6722 6181 6742
rect 6139 6680 6181 6722
rect 6231 6749 6276 6780
rect 6231 6742 6275 6749
rect 6231 6722 6243 6742
rect 6263 6722 6275 6742
rect 10088 6754 10132 6792
rect 6231 6680 6275 6722
rect 7801 6682 7845 6724
rect 3957 6611 4001 6649
rect 7801 6662 7813 6682
rect 7833 6662 7845 6682
rect 7801 6655 7845 6662
rect 7800 6624 7845 6655
rect 7895 6682 7937 6724
rect 7895 6662 7909 6682
rect 7929 6662 7937 6682
rect 7895 6624 7937 6662
rect 8011 6682 8053 6724
rect 8011 6662 8019 6682
rect 8039 6662 8053 6682
rect 8011 6624 8053 6662
rect 8103 6682 8147 6724
rect 8103 6662 8115 6682
rect 8135 6662 8147 6682
rect 8103 6624 8147 6662
rect 8229 6682 8271 6724
rect 8229 6662 8237 6682
rect 8257 6662 8271 6682
rect 8229 6624 8271 6662
rect 8321 6682 8365 6724
rect 10088 6734 10100 6754
rect 10120 6734 10132 6754
rect 8321 6662 8333 6682
rect 8353 6662 8365 6682
rect 10088 6692 10132 6734
rect 10182 6754 10224 6792
rect 10182 6734 10196 6754
rect 10216 6734 10224 6754
rect 10182 6692 10224 6734
rect 10306 6754 10350 6792
rect 10306 6734 10318 6754
rect 10338 6734 10350 6754
rect 10306 6692 10350 6734
rect 10400 6754 10442 6792
rect 10400 6734 10414 6754
rect 10434 6734 10442 6754
rect 10400 6692 10442 6734
rect 10516 6754 10558 6792
rect 10516 6734 10524 6754
rect 10544 6734 10558 6754
rect 10516 6692 10558 6734
rect 10608 6761 10653 6792
rect 10608 6754 10652 6761
rect 10608 6734 10620 6754
rect 10640 6734 10652 6754
rect 14452 6767 14496 6805
rect 10608 6692 10652 6734
rect 12178 6694 12222 6736
rect 8321 6624 8365 6662
rect 384 6505 428 6543
rect 384 6485 396 6505
rect 416 6485 428 6505
rect 384 6443 428 6485
rect 478 6505 520 6543
rect 478 6485 492 6505
rect 512 6485 520 6505
rect 478 6443 520 6485
rect 602 6505 646 6543
rect 602 6485 614 6505
rect 634 6485 646 6505
rect 602 6443 646 6485
rect 696 6505 738 6543
rect 696 6485 710 6505
rect 730 6485 738 6505
rect 696 6443 738 6485
rect 812 6505 854 6543
rect 812 6485 820 6505
rect 840 6485 854 6505
rect 812 6443 854 6485
rect 904 6512 949 6543
rect 904 6505 948 6512
rect 904 6485 916 6505
rect 936 6485 948 6505
rect 904 6443 948 6485
rect 12178 6674 12190 6694
rect 12210 6674 12222 6694
rect 12178 6667 12222 6674
rect 12177 6636 12222 6667
rect 12272 6694 12314 6736
rect 12272 6674 12286 6694
rect 12306 6674 12314 6694
rect 12272 6636 12314 6674
rect 12388 6694 12430 6736
rect 12388 6674 12396 6694
rect 12416 6674 12430 6694
rect 12388 6636 12430 6674
rect 12480 6694 12524 6736
rect 12480 6674 12492 6694
rect 12512 6674 12524 6694
rect 12480 6636 12524 6674
rect 12606 6694 12648 6736
rect 12606 6674 12614 6694
rect 12634 6674 12648 6694
rect 12606 6636 12648 6674
rect 12698 6694 12742 6736
rect 14452 6747 14464 6767
rect 14484 6747 14496 6767
rect 12698 6674 12710 6694
rect 12730 6674 12742 6694
rect 14452 6705 14496 6747
rect 14546 6767 14588 6805
rect 14546 6747 14560 6767
rect 14580 6747 14588 6767
rect 14546 6705 14588 6747
rect 14670 6767 14714 6805
rect 14670 6747 14682 6767
rect 14702 6747 14714 6767
rect 14670 6705 14714 6747
rect 14764 6767 14806 6805
rect 14764 6747 14778 6767
rect 14798 6747 14806 6767
rect 14764 6705 14806 6747
rect 14880 6767 14922 6805
rect 14880 6747 14888 6767
rect 14908 6747 14922 6767
rect 14880 6705 14922 6747
rect 14972 6774 15017 6805
rect 14972 6767 15016 6774
rect 14972 6747 14984 6767
rect 15004 6747 15016 6767
rect 14972 6705 15016 6747
rect 16542 6707 16586 6749
rect 12698 6636 12742 6674
rect 4748 6518 4792 6556
rect 4748 6498 4760 6518
rect 4780 6498 4792 6518
rect 2640 6441 2684 6483
rect 2640 6421 2652 6441
rect 2672 6421 2684 6441
rect 2640 6414 2684 6421
rect 2639 6383 2684 6414
rect 2734 6441 2776 6483
rect 2734 6421 2748 6441
rect 2768 6421 2776 6441
rect 2734 6383 2776 6421
rect 2850 6441 2892 6483
rect 2850 6421 2858 6441
rect 2878 6421 2892 6441
rect 2850 6383 2892 6421
rect 2942 6441 2986 6483
rect 2942 6421 2954 6441
rect 2974 6421 2986 6441
rect 2942 6383 2986 6421
rect 3068 6441 3110 6483
rect 3068 6421 3076 6441
rect 3096 6421 3110 6441
rect 3068 6383 3110 6421
rect 3160 6441 3204 6483
rect 4748 6456 4792 6498
rect 4842 6518 4884 6556
rect 4842 6498 4856 6518
rect 4876 6498 4884 6518
rect 4842 6456 4884 6498
rect 4966 6518 5010 6556
rect 4966 6498 4978 6518
rect 4998 6498 5010 6518
rect 4966 6456 5010 6498
rect 5060 6518 5102 6556
rect 5060 6498 5074 6518
rect 5094 6498 5102 6518
rect 5060 6456 5102 6498
rect 5176 6518 5218 6556
rect 5176 6498 5184 6518
rect 5204 6498 5218 6518
rect 5176 6456 5218 6498
rect 5268 6525 5313 6556
rect 5268 6518 5312 6525
rect 5268 6498 5280 6518
rect 5300 6498 5312 6518
rect 5268 6456 5312 6498
rect 16542 6687 16554 6707
rect 16574 6687 16586 6707
rect 16542 6680 16586 6687
rect 16541 6649 16586 6680
rect 16636 6707 16678 6749
rect 16636 6687 16650 6707
rect 16670 6687 16678 6707
rect 16636 6649 16678 6687
rect 16752 6707 16794 6749
rect 16752 6687 16760 6707
rect 16780 6687 16794 6707
rect 16752 6649 16794 6687
rect 16844 6707 16888 6749
rect 16844 6687 16856 6707
rect 16876 6687 16888 6707
rect 16844 6649 16888 6687
rect 16970 6707 17012 6749
rect 16970 6687 16978 6707
rect 16998 6687 17012 6707
rect 16970 6649 17012 6687
rect 17062 6707 17106 6749
rect 18718 6741 18762 6779
rect 17062 6687 17074 6707
rect 17094 6687 17106 6707
rect 17062 6649 17106 6687
rect 18718 6721 18730 6741
rect 18750 6721 18762 6741
rect 18718 6679 18762 6721
rect 18812 6741 18854 6779
rect 18812 6721 18826 6741
rect 18846 6721 18854 6741
rect 18812 6679 18854 6721
rect 18936 6741 18980 6779
rect 18936 6721 18948 6741
rect 18968 6721 18980 6741
rect 18936 6679 18980 6721
rect 19030 6741 19072 6779
rect 19030 6721 19044 6741
rect 19064 6721 19072 6741
rect 19030 6679 19072 6721
rect 19146 6741 19188 6779
rect 19146 6721 19154 6741
rect 19174 6721 19188 6741
rect 19146 6679 19188 6721
rect 19238 6748 19283 6779
rect 19238 6741 19282 6748
rect 19238 6721 19250 6741
rect 19270 6721 19282 6741
rect 23082 6754 23126 6792
rect 19238 6679 19282 6721
rect 20808 6681 20852 6723
rect 9125 6530 9169 6568
rect 9125 6510 9137 6530
rect 9157 6510 9169 6530
rect 3160 6421 3172 6441
rect 3192 6421 3204 6441
rect 3160 6383 3204 6421
rect 1182 6321 1226 6359
rect 1182 6301 1194 6321
rect 1214 6301 1226 6321
rect 1182 6259 1226 6301
rect 1276 6321 1318 6359
rect 1276 6301 1290 6321
rect 1310 6301 1318 6321
rect 1276 6259 1318 6301
rect 1400 6321 1444 6359
rect 1400 6301 1412 6321
rect 1432 6301 1444 6321
rect 1400 6259 1444 6301
rect 1494 6321 1536 6359
rect 1494 6301 1508 6321
rect 1528 6301 1536 6321
rect 1494 6259 1536 6301
rect 1610 6321 1652 6359
rect 1610 6301 1618 6321
rect 1638 6301 1652 6321
rect 1610 6259 1652 6301
rect 1702 6328 1747 6359
rect 1702 6321 1746 6328
rect 1702 6301 1714 6321
rect 1734 6301 1746 6321
rect 1702 6259 1746 6301
rect 7004 6454 7048 6496
rect 7004 6434 7016 6454
rect 7036 6434 7048 6454
rect 7004 6427 7048 6434
rect 7003 6396 7048 6427
rect 7098 6454 7140 6496
rect 7098 6434 7112 6454
rect 7132 6434 7140 6454
rect 7098 6396 7140 6434
rect 7214 6454 7256 6496
rect 7214 6434 7222 6454
rect 7242 6434 7256 6454
rect 7214 6396 7256 6434
rect 7306 6454 7350 6496
rect 7306 6434 7318 6454
rect 7338 6434 7350 6454
rect 7306 6396 7350 6434
rect 7432 6454 7474 6496
rect 7432 6434 7440 6454
rect 7460 6434 7474 6454
rect 7432 6396 7474 6434
rect 7524 6454 7568 6496
rect 9125 6468 9169 6510
rect 9219 6530 9261 6568
rect 9219 6510 9233 6530
rect 9253 6510 9261 6530
rect 9219 6468 9261 6510
rect 9343 6530 9387 6568
rect 9343 6510 9355 6530
rect 9375 6510 9387 6530
rect 9343 6468 9387 6510
rect 9437 6530 9479 6568
rect 9437 6510 9451 6530
rect 9471 6510 9479 6530
rect 9437 6468 9479 6510
rect 9553 6530 9595 6568
rect 9553 6510 9561 6530
rect 9581 6510 9595 6530
rect 9553 6468 9595 6510
rect 9645 6537 9690 6568
rect 9645 6530 9689 6537
rect 9645 6510 9657 6530
rect 9677 6510 9689 6530
rect 9645 6468 9689 6510
rect 20808 6661 20820 6681
rect 20840 6661 20852 6681
rect 20808 6654 20852 6661
rect 20807 6623 20852 6654
rect 20902 6681 20944 6723
rect 20902 6661 20916 6681
rect 20936 6661 20944 6681
rect 20902 6623 20944 6661
rect 21018 6681 21060 6723
rect 21018 6661 21026 6681
rect 21046 6661 21060 6681
rect 21018 6623 21060 6661
rect 21110 6681 21154 6723
rect 21110 6661 21122 6681
rect 21142 6661 21154 6681
rect 21110 6623 21154 6661
rect 21236 6681 21278 6723
rect 21236 6661 21244 6681
rect 21264 6661 21278 6681
rect 21236 6623 21278 6661
rect 21328 6681 21372 6723
rect 23082 6734 23094 6754
rect 23114 6734 23126 6754
rect 21328 6661 21340 6681
rect 21360 6661 21372 6681
rect 23082 6692 23126 6734
rect 23176 6754 23218 6792
rect 23176 6734 23190 6754
rect 23210 6734 23218 6754
rect 23176 6692 23218 6734
rect 23300 6754 23344 6792
rect 23300 6734 23312 6754
rect 23332 6734 23344 6754
rect 23300 6692 23344 6734
rect 23394 6754 23436 6792
rect 23394 6734 23408 6754
rect 23428 6734 23436 6754
rect 23394 6692 23436 6734
rect 23510 6754 23552 6792
rect 23510 6734 23518 6754
rect 23538 6734 23552 6754
rect 23510 6692 23552 6734
rect 23602 6761 23647 6792
rect 23602 6754 23646 6761
rect 23602 6734 23614 6754
rect 23634 6734 23646 6754
rect 27459 6766 27503 6804
rect 23602 6692 23646 6734
rect 25172 6694 25216 6736
rect 21328 6623 21372 6661
rect 13489 6543 13533 6581
rect 13489 6523 13501 6543
rect 13521 6523 13533 6543
rect 7524 6434 7536 6454
rect 7556 6434 7568 6454
rect 7524 6396 7568 6434
rect 5546 6334 5590 6372
rect 5546 6314 5558 6334
rect 5578 6314 5590 6334
rect 3438 6257 3482 6299
rect 3438 6237 3450 6257
rect 3470 6237 3482 6257
rect 3438 6230 3482 6237
rect 3437 6199 3482 6230
rect 3532 6257 3574 6299
rect 3532 6237 3546 6257
rect 3566 6237 3574 6257
rect 3532 6199 3574 6237
rect 3648 6257 3690 6299
rect 3648 6237 3656 6257
rect 3676 6237 3690 6257
rect 3648 6199 3690 6237
rect 3740 6257 3784 6299
rect 3740 6237 3752 6257
rect 3772 6237 3784 6257
rect 3740 6199 3784 6237
rect 3866 6257 3908 6299
rect 3866 6237 3874 6257
rect 3894 6237 3908 6257
rect 3866 6199 3908 6237
rect 3958 6257 4002 6299
rect 5546 6272 5590 6314
rect 5640 6334 5682 6372
rect 5640 6314 5654 6334
rect 5674 6314 5682 6334
rect 5640 6272 5682 6314
rect 5764 6334 5808 6372
rect 5764 6314 5776 6334
rect 5796 6314 5808 6334
rect 5764 6272 5808 6314
rect 5858 6334 5900 6372
rect 5858 6314 5872 6334
rect 5892 6314 5900 6334
rect 5858 6272 5900 6314
rect 5974 6334 6016 6372
rect 5974 6314 5982 6334
rect 6002 6314 6016 6334
rect 5974 6272 6016 6314
rect 6066 6341 6111 6372
rect 6066 6334 6110 6341
rect 6066 6314 6078 6334
rect 6098 6314 6110 6334
rect 6066 6272 6110 6314
rect 11381 6466 11425 6508
rect 11381 6446 11393 6466
rect 11413 6446 11425 6466
rect 11381 6439 11425 6446
rect 11380 6408 11425 6439
rect 11475 6466 11517 6508
rect 11475 6446 11489 6466
rect 11509 6446 11517 6466
rect 11475 6408 11517 6446
rect 11591 6466 11633 6508
rect 11591 6446 11599 6466
rect 11619 6446 11633 6466
rect 11591 6408 11633 6446
rect 11683 6466 11727 6508
rect 11683 6446 11695 6466
rect 11715 6446 11727 6466
rect 11683 6408 11727 6446
rect 11809 6466 11851 6508
rect 11809 6446 11817 6466
rect 11837 6446 11851 6466
rect 11809 6408 11851 6446
rect 11901 6466 11945 6508
rect 13489 6481 13533 6523
rect 13583 6543 13625 6581
rect 13583 6523 13597 6543
rect 13617 6523 13625 6543
rect 13583 6481 13625 6523
rect 13707 6543 13751 6581
rect 13707 6523 13719 6543
rect 13739 6523 13751 6543
rect 13707 6481 13751 6523
rect 13801 6543 13843 6581
rect 13801 6523 13815 6543
rect 13835 6523 13843 6543
rect 13801 6481 13843 6523
rect 13917 6543 13959 6581
rect 13917 6523 13925 6543
rect 13945 6523 13959 6543
rect 13917 6481 13959 6523
rect 14009 6550 14054 6581
rect 14009 6543 14053 6550
rect 14009 6523 14021 6543
rect 14041 6523 14053 6543
rect 14009 6481 14053 6523
rect 25172 6674 25184 6694
rect 25204 6674 25216 6694
rect 25172 6667 25216 6674
rect 25171 6636 25216 6667
rect 25266 6694 25308 6736
rect 25266 6674 25280 6694
rect 25300 6674 25308 6694
rect 25266 6636 25308 6674
rect 25382 6694 25424 6736
rect 25382 6674 25390 6694
rect 25410 6674 25424 6694
rect 25382 6636 25424 6674
rect 25474 6694 25518 6736
rect 25474 6674 25486 6694
rect 25506 6674 25518 6694
rect 25474 6636 25518 6674
rect 25600 6694 25642 6736
rect 25600 6674 25608 6694
rect 25628 6674 25642 6694
rect 25600 6636 25642 6674
rect 25692 6694 25736 6736
rect 27459 6746 27471 6766
rect 27491 6746 27503 6766
rect 25692 6674 25704 6694
rect 25724 6674 25736 6694
rect 27459 6704 27503 6746
rect 27553 6766 27595 6804
rect 27553 6746 27567 6766
rect 27587 6746 27595 6766
rect 27553 6704 27595 6746
rect 27677 6766 27721 6804
rect 27677 6746 27689 6766
rect 27709 6746 27721 6766
rect 27677 6704 27721 6746
rect 27771 6766 27813 6804
rect 27771 6746 27785 6766
rect 27805 6746 27813 6766
rect 27771 6704 27813 6746
rect 27887 6766 27929 6804
rect 27887 6746 27895 6766
rect 27915 6746 27929 6766
rect 27887 6704 27929 6746
rect 27979 6773 28024 6804
rect 27979 6766 28023 6773
rect 27979 6746 27991 6766
rect 28011 6746 28023 6766
rect 31823 6779 31867 6817
rect 27979 6704 28023 6746
rect 29549 6706 29593 6748
rect 25692 6636 25736 6674
rect 11901 6446 11913 6466
rect 11933 6446 11945 6466
rect 11901 6408 11945 6446
rect 9923 6346 9967 6384
rect 9923 6326 9935 6346
rect 9955 6326 9967 6346
rect 3958 6237 3970 6257
rect 3990 6237 4002 6257
rect 3958 6199 4002 6237
rect 7802 6270 7846 6312
rect 7802 6250 7814 6270
rect 7834 6250 7846 6270
rect 7802 6243 7846 6250
rect 7801 6212 7846 6243
rect 7896 6270 7938 6312
rect 7896 6250 7910 6270
rect 7930 6250 7938 6270
rect 7896 6212 7938 6250
rect 8012 6270 8054 6312
rect 8012 6250 8020 6270
rect 8040 6250 8054 6270
rect 8012 6212 8054 6250
rect 8104 6270 8148 6312
rect 8104 6250 8116 6270
rect 8136 6250 8148 6270
rect 8104 6212 8148 6250
rect 8230 6270 8272 6312
rect 8230 6250 8238 6270
rect 8258 6250 8272 6270
rect 8230 6212 8272 6250
rect 8322 6270 8366 6312
rect 9923 6284 9967 6326
rect 10017 6346 10059 6384
rect 10017 6326 10031 6346
rect 10051 6326 10059 6346
rect 10017 6284 10059 6326
rect 10141 6346 10185 6384
rect 10141 6326 10153 6346
rect 10173 6326 10185 6346
rect 10141 6284 10185 6326
rect 10235 6346 10277 6384
rect 10235 6326 10249 6346
rect 10269 6326 10277 6346
rect 10235 6284 10277 6326
rect 10351 6346 10393 6384
rect 10351 6326 10359 6346
rect 10379 6326 10393 6346
rect 10351 6284 10393 6326
rect 10443 6353 10488 6384
rect 10443 6346 10487 6353
rect 10443 6326 10455 6346
rect 10475 6326 10487 6346
rect 10443 6284 10487 6326
rect 15745 6479 15789 6521
rect 15745 6459 15757 6479
rect 15777 6459 15789 6479
rect 15745 6452 15789 6459
rect 15744 6421 15789 6452
rect 15839 6479 15881 6521
rect 15839 6459 15853 6479
rect 15873 6459 15881 6479
rect 15839 6421 15881 6459
rect 15955 6479 15997 6521
rect 15955 6459 15963 6479
rect 15983 6459 15997 6479
rect 15955 6421 15997 6459
rect 16047 6479 16091 6521
rect 16047 6459 16059 6479
rect 16079 6459 16091 6479
rect 16047 6421 16091 6459
rect 16173 6479 16215 6521
rect 16173 6459 16181 6479
rect 16201 6459 16215 6479
rect 16173 6421 16215 6459
rect 16265 6479 16309 6521
rect 17755 6517 17799 6555
rect 17755 6497 17767 6517
rect 17787 6497 17799 6517
rect 16265 6459 16277 6479
rect 16297 6459 16309 6479
rect 16265 6421 16309 6459
rect 17755 6455 17799 6497
rect 17849 6517 17891 6555
rect 17849 6497 17863 6517
rect 17883 6497 17891 6517
rect 17849 6455 17891 6497
rect 17973 6517 18017 6555
rect 17973 6497 17985 6517
rect 18005 6497 18017 6517
rect 17973 6455 18017 6497
rect 18067 6517 18109 6555
rect 18067 6497 18081 6517
rect 18101 6497 18109 6517
rect 18067 6455 18109 6497
rect 18183 6517 18225 6555
rect 18183 6497 18191 6517
rect 18211 6497 18225 6517
rect 18183 6455 18225 6497
rect 18275 6524 18320 6555
rect 18275 6517 18319 6524
rect 18275 6497 18287 6517
rect 18307 6497 18319 6517
rect 18275 6455 18319 6497
rect 29549 6686 29561 6706
rect 29581 6686 29593 6706
rect 29549 6679 29593 6686
rect 29548 6648 29593 6679
rect 29643 6706 29685 6748
rect 29643 6686 29657 6706
rect 29677 6686 29685 6706
rect 29643 6648 29685 6686
rect 29759 6706 29801 6748
rect 29759 6686 29767 6706
rect 29787 6686 29801 6706
rect 29759 6648 29801 6686
rect 29851 6706 29895 6748
rect 29851 6686 29863 6706
rect 29883 6686 29895 6706
rect 29851 6648 29895 6686
rect 29977 6706 30019 6748
rect 29977 6686 29985 6706
rect 30005 6686 30019 6706
rect 29977 6648 30019 6686
rect 30069 6706 30113 6748
rect 31823 6759 31835 6779
rect 31855 6759 31867 6779
rect 30069 6686 30081 6706
rect 30101 6686 30113 6706
rect 31823 6717 31867 6759
rect 31917 6779 31959 6817
rect 31917 6759 31931 6779
rect 31951 6759 31959 6779
rect 31917 6717 31959 6759
rect 32041 6779 32085 6817
rect 32041 6759 32053 6779
rect 32073 6759 32085 6779
rect 32041 6717 32085 6759
rect 32135 6779 32177 6817
rect 32135 6759 32149 6779
rect 32169 6759 32177 6779
rect 32135 6717 32177 6759
rect 32251 6779 32293 6817
rect 32251 6759 32259 6779
rect 32279 6759 32293 6779
rect 32251 6717 32293 6759
rect 32343 6786 32388 6817
rect 32343 6779 32387 6786
rect 32343 6759 32355 6779
rect 32375 6759 32387 6779
rect 32343 6717 32387 6759
rect 33913 6719 33957 6761
rect 30069 6648 30113 6686
rect 22119 6530 22163 6568
rect 22119 6510 22131 6530
rect 22151 6510 22163 6530
rect 14287 6359 14331 6397
rect 14287 6339 14299 6359
rect 14319 6339 14331 6359
rect 8322 6250 8334 6270
rect 8354 6250 8366 6270
rect 8322 6212 8366 6250
rect 385 6093 429 6131
rect 385 6073 397 6093
rect 417 6073 429 6093
rect 385 6031 429 6073
rect 479 6093 521 6131
rect 479 6073 493 6093
rect 513 6073 521 6093
rect 479 6031 521 6073
rect 603 6093 647 6131
rect 603 6073 615 6093
rect 635 6073 647 6093
rect 603 6031 647 6073
rect 697 6093 739 6131
rect 697 6073 711 6093
rect 731 6073 739 6093
rect 697 6031 739 6073
rect 813 6093 855 6131
rect 813 6073 821 6093
rect 841 6073 855 6093
rect 813 6031 855 6073
rect 905 6100 950 6131
rect 905 6093 949 6100
rect 905 6073 917 6093
rect 937 6073 949 6093
rect 12179 6282 12223 6324
rect 12179 6262 12191 6282
rect 12211 6262 12223 6282
rect 12179 6255 12223 6262
rect 12178 6224 12223 6255
rect 12273 6282 12315 6324
rect 12273 6262 12287 6282
rect 12307 6262 12315 6282
rect 12273 6224 12315 6262
rect 12389 6282 12431 6324
rect 12389 6262 12397 6282
rect 12417 6262 12431 6282
rect 12389 6224 12431 6262
rect 12481 6282 12525 6324
rect 12481 6262 12493 6282
rect 12513 6262 12525 6282
rect 12481 6224 12525 6262
rect 12607 6282 12649 6324
rect 12607 6262 12615 6282
rect 12635 6262 12649 6282
rect 12607 6224 12649 6262
rect 12699 6282 12743 6324
rect 14287 6297 14331 6339
rect 14381 6359 14423 6397
rect 14381 6339 14395 6359
rect 14415 6339 14423 6359
rect 14381 6297 14423 6339
rect 14505 6359 14549 6397
rect 14505 6339 14517 6359
rect 14537 6339 14549 6359
rect 14505 6297 14549 6339
rect 14599 6359 14641 6397
rect 14599 6339 14613 6359
rect 14633 6339 14641 6359
rect 14599 6297 14641 6339
rect 14715 6359 14757 6397
rect 14715 6339 14723 6359
rect 14743 6339 14757 6359
rect 14715 6297 14757 6339
rect 14807 6366 14852 6397
rect 14807 6359 14851 6366
rect 14807 6339 14819 6359
rect 14839 6339 14851 6359
rect 14807 6297 14851 6339
rect 20011 6453 20055 6495
rect 20011 6433 20023 6453
rect 20043 6433 20055 6453
rect 20011 6426 20055 6433
rect 20010 6395 20055 6426
rect 20105 6453 20147 6495
rect 20105 6433 20119 6453
rect 20139 6433 20147 6453
rect 20105 6395 20147 6433
rect 20221 6453 20263 6495
rect 20221 6433 20229 6453
rect 20249 6433 20263 6453
rect 20221 6395 20263 6433
rect 20313 6453 20357 6495
rect 20313 6433 20325 6453
rect 20345 6433 20357 6453
rect 20313 6395 20357 6433
rect 20439 6453 20481 6495
rect 20439 6433 20447 6453
rect 20467 6433 20481 6453
rect 20439 6395 20481 6433
rect 20531 6453 20575 6495
rect 22119 6468 22163 6510
rect 22213 6530 22255 6568
rect 22213 6510 22227 6530
rect 22247 6510 22255 6530
rect 22213 6468 22255 6510
rect 22337 6530 22381 6568
rect 22337 6510 22349 6530
rect 22369 6510 22381 6530
rect 22337 6468 22381 6510
rect 22431 6530 22473 6568
rect 22431 6510 22445 6530
rect 22465 6510 22473 6530
rect 22431 6468 22473 6510
rect 22547 6530 22589 6568
rect 22547 6510 22555 6530
rect 22575 6510 22589 6530
rect 22547 6468 22589 6510
rect 22639 6537 22684 6568
rect 22639 6530 22683 6537
rect 22639 6510 22651 6530
rect 22671 6510 22683 6530
rect 22639 6468 22683 6510
rect 33913 6699 33925 6719
rect 33945 6699 33957 6719
rect 33913 6692 33957 6699
rect 33912 6661 33957 6692
rect 34007 6719 34049 6761
rect 34007 6699 34021 6719
rect 34041 6699 34049 6719
rect 34007 6661 34049 6699
rect 34123 6719 34165 6761
rect 34123 6699 34131 6719
rect 34151 6699 34165 6719
rect 34123 6661 34165 6699
rect 34215 6719 34259 6761
rect 34215 6699 34227 6719
rect 34247 6699 34259 6719
rect 34215 6661 34259 6699
rect 34341 6719 34383 6761
rect 34341 6699 34349 6719
rect 34369 6699 34383 6719
rect 34341 6661 34383 6699
rect 34433 6719 34477 6761
rect 34433 6699 34445 6719
rect 34465 6699 34477 6719
rect 34433 6661 34477 6699
rect 26496 6542 26540 6580
rect 26496 6522 26508 6542
rect 26528 6522 26540 6542
rect 20531 6433 20543 6453
rect 20563 6433 20575 6453
rect 20531 6395 20575 6433
rect 12699 6262 12711 6282
rect 12731 6262 12743 6282
rect 12699 6224 12743 6262
rect 4749 6106 4793 6144
rect 905 6031 949 6073
rect 2541 6031 2585 6073
rect 2541 6011 2553 6031
rect 2573 6011 2585 6031
rect 2541 6004 2585 6011
rect 2540 5973 2585 6004
rect 2635 6031 2677 6073
rect 2635 6011 2649 6031
rect 2669 6011 2677 6031
rect 2635 5973 2677 6011
rect 2751 6031 2793 6073
rect 2751 6011 2759 6031
rect 2779 6011 2793 6031
rect 2751 5973 2793 6011
rect 2843 6031 2887 6073
rect 2843 6011 2855 6031
rect 2875 6011 2887 6031
rect 2843 5973 2887 6011
rect 2969 6031 3011 6073
rect 2969 6011 2977 6031
rect 2997 6011 3011 6031
rect 2969 5973 3011 6011
rect 3061 6031 3105 6073
rect 4749 6086 4761 6106
rect 4781 6086 4793 6106
rect 3061 6011 3073 6031
rect 3093 6011 3105 6031
rect 4749 6044 4793 6086
rect 4843 6106 4885 6144
rect 4843 6086 4857 6106
rect 4877 6086 4885 6106
rect 4843 6044 4885 6086
rect 4967 6106 5011 6144
rect 4967 6086 4979 6106
rect 4999 6086 5011 6106
rect 4967 6044 5011 6086
rect 5061 6106 5103 6144
rect 5061 6086 5075 6106
rect 5095 6086 5103 6106
rect 5061 6044 5103 6086
rect 5177 6106 5219 6144
rect 5177 6086 5185 6106
rect 5205 6086 5219 6106
rect 5177 6044 5219 6086
rect 5269 6113 5314 6144
rect 5269 6106 5313 6113
rect 5269 6086 5281 6106
rect 5301 6086 5313 6106
rect 16543 6295 16587 6337
rect 16543 6275 16555 6295
rect 16575 6275 16587 6295
rect 16543 6268 16587 6275
rect 16542 6237 16587 6268
rect 16637 6295 16679 6337
rect 16637 6275 16651 6295
rect 16671 6275 16679 6295
rect 16637 6237 16679 6275
rect 16753 6295 16795 6337
rect 16753 6275 16761 6295
rect 16781 6275 16795 6295
rect 16753 6237 16795 6275
rect 16845 6295 16889 6337
rect 16845 6275 16857 6295
rect 16877 6275 16889 6295
rect 16845 6237 16889 6275
rect 16971 6295 17013 6337
rect 16971 6275 16979 6295
rect 16999 6275 17013 6295
rect 16971 6237 17013 6275
rect 17063 6295 17107 6337
rect 18553 6333 18597 6371
rect 18553 6313 18565 6333
rect 18585 6313 18597 6333
rect 17063 6275 17075 6295
rect 17095 6275 17107 6295
rect 17063 6237 17107 6275
rect 18553 6271 18597 6313
rect 18647 6333 18689 6371
rect 18647 6313 18661 6333
rect 18681 6313 18689 6333
rect 18647 6271 18689 6313
rect 18771 6333 18815 6371
rect 18771 6313 18783 6333
rect 18803 6313 18815 6333
rect 18771 6271 18815 6313
rect 18865 6333 18907 6371
rect 18865 6313 18879 6333
rect 18899 6313 18907 6333
rect 18865 6271 18907 6313
rect 18981 6333 19023 6371
rect 18981 6313 18989 6333
rect 19009 6313 19023 6333
rect 18981 6271 19023 6313
rect 19073 6340 19118 6371
rect 19073 6333 19117 6340
rect 19073 6313 19085 6333
rect 19105 6313 19117 6333
rect 19073 6271 19117 6313
rect 24375 6466 24419 6508
rect 24375 6446 24387 6466
rect 24407 6446 24419 6466
rect 24375 6439 24419 6446
rect 24374 6408 24419 6439
rect 24469 6466 24511 6508
rect 24469 6446 24483 6466
rect 24503 6446 24511 6466
rect 24469 6408 24511 6446
rect 24585 6466 24627 6508
rect 24585 6446 24593 6466
rect 24613 6446 24627 6466
rect 24585 6408 24627 6446
rect 24677 6466 24721 6508
rect 24677 6446 24689 6466
rect 24709 6446 24721 6466
rect 24677 6408 24721 6446
rect 24803 6466 24845 6508
rect 24803 6446 24811 6466
rect 24831 6446 24845 6466
rect 24803 6408 24845 6446
rect 24895 6466 24939 6508
rect 26496 6480 26540 6522
rect 26590 6542 26632 6580
rect 26590 6522 26604 6542
rect 26624 6522 26632 6542
rect 26590 6480 26632 6522
rect 26714 6542 26758 6580
rect 26714 6522 26726 6542
rect 26746 6522 26758 6542
rect 26714 6480 26758 6522
rect 26808 6542 26850 6580
rect 26808 6522 26822 6542
rect 26842 6522 26850 6542
rect 26808 6480 26850 6522
rect 26924 6542 26966 6580
rect 26924 6522 26932 6542
rect 26952 6522 26966 6542
rect 26924 6480 26966 6522
rect 27016 6549 27061 6580
rect 27016 6542 27060 6549
rect 27016 6522 27028 6542
rect 27048 6522 27060 6542
rect 27016 6480 27060 6522
rect 30860 6555 30904 6593
rect 30860 6535 30872 6555
rect 30892 6535 30904 6555
rect 24895 6446 24907 6466
rect 24927 6446 24939 6466
rect 24895 6408 24939 6446
rect 22917 6346 22961 6384
rect 22917 6326 22929 6346
rect 22949 6326 22961 6346
rect 9126 6118 9170 6156
rect 5269 6044 5313 6086
rect 6905 6044 6949 6086
rect 3061 5973 3105 6011
rect 6905 6024 6917 6044
rect 6937 6024 6949 6044
rect 6905 6017 6949 6024
rect 6904 5986 6949 6017
rect 6999 6044 7041 6086
rect 6999 6024 7013 6044
rect 7033 6024 7041 6044
rect 6999 5986 7041 6024
rect 7115 6044 7157 6086
rect 7115 6024 7123 6044
rect 7143 6024 7157 6044
rect 7115 5986 7157 6024
rect 7207 6044 7251 6086
rect 7207 6024 7219 6044
rect 7239 6024 7251 6044
rect 7207 5986 7251 6024
rect 7333 6044 7375 6086
rect 7333 6024 7341 6044
rect 7361 6024 7375 6044
rect 7333 5986 7375 6024
rect 7425 6044 7469 6086
rect 9126 6098 9138 6118
rect 9158 6098 9170 6118
rect 7425 6024 7437 6044
rect 7457 6024 7469 6044
rect 9126 6056 9170 6098
rect 9220 6118 9262 6156
rect 9220 6098 9234 6118
rect 9254 6098 9262 6118
rect 9220 6056 9262 6098
rect 9344 6118 9388 6156
rect 9344 6098 9356 6118
rect 9376 6098 9388 6118
rect 9344 6056 9388 6098
rect 9438 6118 9480 6156
rect 9438 6098 9452 6118
rect 9472 6098 9480 6118
rect 9438 6056 9480 6098
rect 9554 6118 9596 6156
rect 9554 6098 9562 6118
rect 9582 6098 9596 6118
rect 9554 6056 9596 6098
rect 9646 6125 9691 6156
rect 9646 6118 9690 6125
rect 9646 6098 9658 6118
rect 9678 6098 9690 6118
rect 20809 6269 20853 6311
rect 20809 6249 20821 6269
rect 20841 6249 20853 6269
rect 20809 6242 20853 6249
rect 20808 6211 20853 6242
rect 20903 6269 20945 6311
rect 20903 6249 20917 6269
rect 20937 6249 20945 6269
rect 20903 6211 20945 6249
rect 21019 6269 21061 6311
rect 21019 6249 21027 6269
rect 21047 6249 21061 6269
rect 21019 6211 21061 6249
rect 21111 6269 21155 6311
rect 21111 6249 21123 6269
rect 21143 6249 21155 6269
rect 21111 6211 21155 6249
rect 21237 6269 21279 6311
rect 21237 6249 21245 6269
rect 21265 6249 21279 6269
rect 21237 6211 21279 6249
rect 21329 6269 21373 6311
rect 22917 6284 22961 6326
rect 23011 6346 23053 6384
rect 23011 6326 23025 6346
rect 23045 6326 23053 6346
rect 23011 6284 23053 6326
rect 23135 6346 23179 6384
rect 23135 6326 23147 6346
rect 23167 6326 23179 6346
rect 23135 6284 23179 6326
rect 23229 6346 23271 6384
rect 23229 6326 23243 6346
rect 23263 6326 23271 6346
rect 23229 6284 23271 6326
rect 23345 6346 23387 6384
rect 23345 6326 23353 6346
rect 23373 6326 23387 6346
rect 23345 6284 23387 6326
rect 23437 6353 23482 6384
rect 23437 6346 23481 6353
rect 23437 6326 23449 6346
rect 23469 6326 23481 6346
rect 23437 6284 23481 6326
rect 28752 6478 28796 6520
rect 28752 6458 28764 6478
rect 28784 6458 28796 6478
rect 28752 6451 28796 6458
rect 28751 6420 28796 6451
rect 28846 6478 28888 6520
rect 28846 6458 28860 6478
rect 28880 6458 28888 6478
rect 28846 6420 28888 6458
rect 28962 6478 29004 6520
rect 28962 6458 28970 6478
rect 28990 6458 29004 6478
rect 28962 6420 29004 6458
rect 29054 6478 29098 6520
rect 29054 6458 29066 6478
rect 29086 6458 29098 6478
rect 29054 6420 29098 6458
rect 29180 6478 29222 6520
rect 29180 6458 29188 6478
rect 29208 6458 29222 6478
rect 29180 6420 29222 6458
rect 29272 6478 29316 6520
rect 30860 6493 30904 6535
rect 30954 6555 30996 6593
rect 30954 6535 30968 6555
rect 30988 6535 30996 6555
rect 30954 6493 30996 6535
rect 31078 6555 31122 6593
rect 31078 6535 31090 6555
rect 31110 6535 31122 6555
rect 31078 6493 31122 6535
rect 31172 6555 31214 6593
rect 31172 6535 31186 6555
rect 31206 6535 31214 6555
rect 31172 6493 31214 6535
rect 31288 6555 31330 6593
rect 31288 6535 31296 6555
rect 31316 6535 31330 6555
rect 31288 6493 31330 6535
rect 31380 6562 31425 6593
rect 31380 6555 31424 6562
rect 31380 6535 31392 6555
rect 31412 6535 31424 6555
rect 31380 6493 31424 6535
rect 29272 6458 29284 6478
rect 29304 6458 29316 6478
rect 29272 6420 29316 6458
rect 27294 6358 27338 6396
rect 27294 6338 27306 6358
rect 27326 6338 27338 6358
rect 21329 6249 21341 6269
rect 21361 6249 21373 6269
rect 21329 6211 21373 6249
rect 13490 6131 13534 6169
rect 9646 6056 9690 6098
rect 11282 6056 11326 6098
rect 7425 5986 7469 6024
rect 11282 6036 11294 6056
rect 11314 6036 11326 6056
rect 11282 6029 11326 6036
rect 11281 5998 11326 6029
rect 11376 6056 11418 6098
rect 11376 6036 11390 6056
rect 11410 6036 11418 6056
rect 11376 5998 11418 6036
rect 11492 6056 11534 6098
rect 11492 6036 11500 6056
rect 11520 6036 11534 6056
rect 11492 5998 11534 6036
rect 11584 6056 11628 6098
rect 11584 6036 11596 6056
rect 11616 6036 11628 6056
rect 11584 5998 11628 6036
rect 11710 6056 11752 6098
rect 11710 6036 11718 6056
rect 11738 6036 11752 6056
rect 11710 5998 11752 6036
rect 11802 6056 11846 6098
rect 13490 6111 13502 6131
rect 13522 6111 13534 6131
rect 11802 6036 11814 6056
rect 11834 6036 11846 6056
rect 13490 6069 13534 6111
rect 13584 6131 13626 6169
rect 13584 6111 13598 6131
rect 13618 6111 13626 6131
rect 13584 6069 13626 6111
rect 13708 6131 13752 6169
rect 13708 6111 13720 6131
rect 13740 6111 13752 6131
rect 13708 6069 13752 6111
rect 13802 6131 13844 6169
rect 13802 6111 13816 6131
rect 13836 6111 13844 6131
rect 13802 6069 13844 6111
rect 13918 6131 13960 6169
rect 13918 6111 13926 6131
rect 13946 6111 13960 6131
rect 13918 6069 13960 6111
rect 14010 6138 14055 6169
rect 14010 6131 14054 6138
rect 14010 6111 14022 6131
rect 14042 6111 14054 6131
rect 25173 6282 25217 6324
rect 25173 6262 25185 6282
rect 25205 6262 25217 6282
rect 25173 6255 25217 6262
rect 25172 6224 25217 6255
rect 25267 6282 25309 6324
rect 25267 6262 25281 6282
rect 25301 6262 25309 6282
rect 25267 6224 25309 6262
rect 25383 6282 25425 6324
rect 25383 6262 25391 6282
rect 25411 6262 25425 6282
rect 25383 6224 25425 6262
rect 25475 6282 25519 6324
rect 25475 6262 25487 6282
rect 25507 6262 25519 6282
rect 25475 6224 25519 6262
rect 25601 6282 25643 6324
rect 25601 6262 25609 6282
rect 25629 6262 25643 6282
rect 25601 6224 25643 6262
rect 25693 6282 25737 6324
rect 27294 6296 27338 6338
rect 27388 6358 27430 6396
rect 27388 6338 27402 6358
rect 27422 6338 27430 6358
rect 27388 6296 27430 6338
rect 27512 6358 27556 6396
rect 27512 6338 27524 6358
rect 27544 6338 27556 6358
rect 27512 6296 27556 6338
rect 27606 6358 27648 6396
rect 27606 6338 27620 6358
rect 27640 6338 27648 6358
rect 27606 6296 27648 6338
rect 27722 6358 27764 6396
rect 27722 6338 27730 6358
rect 27750 6338 27764 6358
rect 27722 6296 27764 6338
rect 27814 6365 27859 6396
rect 27814 6358 27858 6365
rect 27814 6338 27826 6358
rect 27846 6338 27858 6358
rect 27814 6296 27858 6338
rect 33116 6491 33160 6533
rect 33116 6471 33128 6491
rect 33148 6471 33160 6491
rect 33116 6464 33160 6471
rect 33115 6433 33160 6464
rect 33210 6491 33252 6533
rect 33210 6471 33224 6491
rect 33244 6471 33252 6491
rect 33210 6433 33252 6471
rect 33326 6491 33368 6533
rect 33326 6471 33334 6491
rect 33354 6471 33368 6491
rect 33326 6433 33368 6471
rect 33418 6491 33462 6533
rect 33418 6471 33430 6491
rect 33450 6471 33462 6491
rect 33418 6433 33462 6471
rect 33544 6491 33586 6533
rect 33544 6471 33552 6491
rect 33572 6471 33586 6491
rect 33544 6433 33586 6471
rect 33636 6491 33680 6533
rect 33636 6471 33648 6491
rect 33668 6471 33680 6491
rect 33636 6433 33680 6471
rect 31658 6371 31702 6409
rect 31658 6351 31670 6371
rect 31690 6351 31702 6371
rect 25693 6262 25705 6282
rect 25725 6262 25737 6282
rect 25693 6224 25737 6262
rect 14010 6069 14054 6111
rect 15646 6069 15690 6111
rect 11802 5998 11846 6036
rect 15646 6049 15658 6069
rect 15678 6049 15690 6069
rect 15646 6042 15690 6049
rect 15645 6011 15690 6042
rect 15740 6069 15782 6111
rect 15740 6049 15754 6069
rect 15774 6049 15782 6069
rect 15740 6011 15782 6049
rect 15856 6069 15898 6111
rect 15856 6049 15864 6069
rect 15884 6049 15898 6069
rect 15856 6011 15898 6049
rect 15948 6069 15992 6111
rect 15948 6049 15960 6069
rect 15980 6049 15992 6069
rect 15948 6011 15992 6049
rect 16074 6069 16116 6111
rect 16074 6049 16082 6069
rect 16102 6049 16116 6069
rect 16074 6011 16116 6049
rect 16166 6069 16210 6111
rect 16166 6049 16178 6069
rect 16198 6049 16210 6069
rect 17756 6105 17800 6143
rect 17756 6085 17768 6105
rect 17788 6085 17800 6105
rect 16166 6011 16210 6049
rect 17756 6043 17800 6085
rect 17850 6105 17892 6143
rect 17850 6085 17864 6105
rect 17884 6085 17892 6105
rect 17850 6043 17892 6085
rect 17974 6105 18018 6143
rect 17974 6085 17986 6105
rect 18006 6085 18018 6105
rect 17974 6043 18018 6085
rect 18068 6105 18110 6143
rect 18068 6085 18082 6105
rect 18102 6085 18110 6105
rect 18068 6043 18110 6085
rect 18184 6105 18226 6143
rect 18184 6085 18192 6105
rect 18212 6085 18226 6105
rect 18184 6043 18226 6085
rect 18276 6112 18321 6143
rect 18276 6105 18320 6112
rect 18276 6085 18288 6105
rect 18308 6085 18320 6105
rect 29550 6294 29594 6336
rect 29550 6274 29562 6294
rect 29582 6274 29594 6294
rect 29550 6267 29594 6274
rect 29549 6236 29594 6267
rect 29644 6294 29686 6336
rect 29644 6274 29658 6294
rect 29678 6274 29686 6294
rect 29644 6236 29686 6274
rect 29760 6294 29802 6336
rect 29760 6274 29768 6294
rect 29788 6274 29802 6294
rect 29760 6236 29802 6274
rect 29852 6294 29896 6336
rect 29852 6274 29864 6294
rect 29884 6274 29896 6294
rect 29852 6236 29896 6274
rect 29978 6294 30020 6336
rect 29978 6274 29986 6294
rect 30006 6274 30020 6294
rect 29978 6236 30020 6274
rect 30070 6294 30114 6336
rect 31658 6309 31702 6351
rect 31752 6371 31794 6409
rect 31752 6351 31766 6371
rect 31786 6351 31794 6371
rect 31752 6309 31794 6351
rect 31876 6371 31920 6409
rect 31876 6351 31888 6371
rect 31908 6351 31920 6371
rect 31876 6309 31920 6351
rect 31970 6371 32012 6409
rect 31970 6351 31984 6371
rect 32004 6351 32012 6371
rect 31970 6309 32012 6351
rect 32086 6371 32128 6409
rect 32086 6351 32094 6371
rect 32114 6351 32128 6371
rect 32086 6309 32128 6351
rect 32178 6378 32223 6409
rect 32178 6371 32222 6378
rect 32178 6351 32190 6371
rect 32210 6351 32222 6371
rect 32178 6309 32222 6351
rect 30070 6274 30082 6294
rect 30102 6274 30114 6294
rect 30070 6236 30114 6274
rect 22120 6118 22164 6156
rect 18276 6043 18320 6085
rect 19912 6043 19956 6085
rect 19912 6023 19924 6043
rect 19944 6023 19956 6043
rect 19912 6016 19956 6023
rect 19911 5985 19956 6016
rect 20006 6043 20048 6085
rect 20006 6023 20020 6043
rect 20040 6023 20048 6043
rect 20006 5985 20048 6023
rect 20122 6043 20164 6085
rect 20122 6023 20130 6043
rect 20150 6023 20164 6043
rect 20122 5985 20164 6023
rect 20214 6043 20258 6085
rect 20214 6023 20226 6043
rect 20246 6023 20258 6043
rect 20214 5985 20258 6023
rect 20340 6043 20382 6085
rect 20340 6023 20348 6043
rect 20368 6023 20382 6043
rect 20340 5985 20382 6023
rect 20432 6043 20476 6085
rect 22120 6098 22132 6118
rect 22152 6098 22164 6118
rect 20432 6023 20444 6043
rect 20464 6023 20476 6043
rect 22120 6056 22164 6098
rect 22214 6118 22256 6156
rect 22214 6098 22228 6118
rect 22248 6098 22256 6118
rect 22214 6056 22256 6098
rect 22338 6118 22382 6156
rect 22338 6098 22350 6118
rect 22370 6098 22382 6118
rect 22338 6056 22382 6098
rect 22432 6118 22474 6156
rect 22432 6098 22446 6118
rect 22466 6098 22474 6118
rect 22432 6056 22474 6098
rect 22548 6118 22590 6156
rect 22548 6098 22556 6118
rect 22576 6098 22590 6118
rect 22548 6056 22590 6098
rect 22640 6125 22685 6156
rect 22640 6118 22684 6125
rect 22640 6098 22652 6118
rect 22672 6098 22684 6118
rect 33914 6307 33958 6349
rect 33914 6287 33926 6307
rect 33946 6287 33958 6307
rect 33914 6280 33958 6287
rect 33913 6249 33958 6280
rect 34008 6307 34050 6349
rect 34008 6287 34022 6307
rect 34042 6287 34050 6307
rect 34008 6249 34050 6287
rect 34124 6307 34166 6349
rect 34124 6287 34132 6307
rect 34152 6287 34166 6307
rect 34124 6249 34166 6287
rect 34216 6307 34260 6349
rect 34216 6287 34228 6307
rect 34248 6287 34260 6307
rect 34216 6249 34260 6287
rect 34342 6307 34384 6349
rect 34342 6287 34350 6307
rect 34370 6287 34384 6307
rect 34342 6249 34384 6287
rect 34434 6307 34478 6349
rect 34434 6287 34446 6307
rect 34466 6287 34478 6307
rect 34434 6249 34478 6287
rect 26497 6130 26541 6168
rect 22640 6056 22684 6098
rect 24276 6056 24320 6098
rect 20432 5985 20476 6023
rect 24276 6036 24288 6056
rect 24308 6036 24320 6056
rect 24276 6029 24320 6036
rect 24275 5998 24320 6029
rect 24370 6056 24412 6098
rect 24370 6036 24384 6056
rect 24404 6036 24412 6056
rect 24370 5998 24412 6036
rect 24486 6056 24528 6098
rect 24486 6036 24494 6056
rect 24514 6036 24528 6056
rect 24486 5998 24528 6036
rect 24578 6056 24622 6098
rect 24578 6036 24590 6056
rect 24610 6036 24622 6056
rect 24578 5998 24622 6036
rect 24704 6056 24746 6098
rect 24704 6036 24712 6056
rect 24732 6036 24746 6056
rect 24704 5998 24746 6036
rect 24796 6056 24840 6098
rect 26497 6110 26509 6130
rect 26529 6110 26541 6130
rect 24796 6036 24808 6056
rect 24828 6036 24840 6056
rect 26497 6068 26541 6110
rect 26591 6130 26633 6168
rect 26591 6110 26605 6130
rect 26625 6110 26633 6130
rect 26591 6068 26633 6110
rect 26715 6130 26759 6168
rect 26715 6110 26727 6130
rect 26747 6110 26759 6130
rect 26715 6068 26759 6110
rect 26809 6130 26851 6168
rect 26809 6110 26823 6130
rect 26843 6110 26851 6130
rect 26809 6068 26851 6110
rect 26925 6130 26967 6168
rect 26925 6110 26933 6130
rect 26953 6110 26967 6130
rect 26925 6068 26967 6110
rect 27017 6137 27062 6168
rect 27017 6130 27061 6137
rect 27017 6110 27029 6130
rect 27049 6110 27061 6130
rect 30861 6143 30905 6181
rect 27017 6068 27061 6110
rect 28653 6068 28697 6110
rect 24796 5998 24840 6036
rect 28653 6048 28665 6068
rect 28685 6048 28697 6068
rect 28653 6041 28697 6048
rect 28652 6010 28697 6041
rect 28747 6068 28789 6110
rect 28747 6048 28761 6068
rect 28781 6048 28789 6068
rect 28747 6010 28789 6048
rect 28863 6068 28905 6110
rect 28863 6048 28871 6068
rect 28891 6048 28905 6068
rect 28863 6010 28905 6048
rect 28955 6068 28999 6110
rect 28955 6048 28967 6068
rect 28987 6048 28999 6068
rect 28955 6010 28999 6048
rect 29081 6068 29123 6110
rect 29081 6048 29089 6068
rect 29109 6048 29123 6068
rect 29081 6010 29123 6048
rect 29173 6068 29217 6110
rect 30861 6123 30873 6143
rect 30893 6123 30905 6143
rect 29173 6048 29185 6068
rect 29205 6048 29217 6068
rect 30861 6081 30905 6123
rect 30955 6143 30997 6181
rect 30955 6123 30969 6143
rect 30989 6123 30997 6143
rect 30955 6081 30997 6123
rect 31079 6143 31123 6181
rect 31079 6123 31091 6143
rect 31111 6123 31123 6143
rect 31079 6081 31123 6123
rect 31173 6143 31215 6181
rect 31173 6123 31187 6143
rect 31207 6123 31215 6143
rect 31173 6081 31215 6123
rect 31289 6143 31331 6181
rect 31289 6123 31297 6143
rect 31317 6123 31331 6143
rect 31289 6081 31331 6123
rect 31381 6150 31426 6181
rect 31381 6143 31425 6150
rect 31381 6123 31393 6143
rect 31413 6123 31425 6143
rect 31381 6081 31425 6123
rect 33017 6081 33061 6123
rect 29173 6010 29217 6048
rect 33017 6061 33029 6081
rect 33049 6061 33061 6081
rect 33017 6054 33061 6061
rect 33016 6023 33061 6054
rect 33111 6081 33153 6123
rect 33111 6061 33125 6081
rect 33145 6061 33153 6081
rect 33111 6023 33153 6061
rect 33227 6081 33269 6123
rect 33227 6061 33235 6081
rect 33255 6061 33269 6081
rect 33227 6023 33269 6061
rect 33319 6081 33363 6123
rect 33319 6061 33331 6081
rect 33351 6061 33363 6081
rect 33319 6023 33363 6061
rect 33445 6081 33487 6123
rect 33445 6061 33453 6081
rect 33473 6061 33487 6081
rect 33445 6023 33487 6061
rect 33537 6081 33581 6123
rect 33537 6061 33549 6081
rect 33569 6061 33581 6081
rect 33537 6023 33581 6061
rect 1264 5713 1308 5751
rect 1264 5693 1276 5713
rect 1296 5693 1308 5713
rect 1264 5651 1308 5693
rect 1358 5713 1400 5751
rect 1358 5693 1372 5713
rect 1392 5693 1400 5713
rect 1358 5651 1400 5693
rect 1482 5713 1526 5751
rect 1482 5693 1494 5713
rect 1514 5693 1526 5713
rect 1482 5651 1526 5693
rect 1576 5713 1618 5751
rect 1576 5693 1590 5713
rect 1610 5693 1618 5713
rect 1576 5651 1618 5693
rect 1692 5713 1734 5751
rect 1692 5693 1700 5713
rect 1720 5693 1734 5713
rect 1692 5651 1734 5693
rect 1784 5720 1829 5751
rect 1784 5713 1828 5720
rect 1784 5693 1796 5713
rect 1816 5693 1828 5713
rect 5628 5726 5672 5764
rect 1784 5651 1828 5693
rect 3420 5651 3464 5693
rect 3420 5631 3432 5651
rect 3452 5631 3464 5651
rect 3420 5624 3464 5631
rect 3419 5593 3464 5624
rect 3514 5651 3556 5693
rect 3514 5631 3528 5651
rect 3548 5631 3556 5651
rect 3514 5593 3556 5631
rect 3630 5651 3672 5693
rect 3630 5631 3638 5651
rect 3658 5631 3672 5651
rect 3630 5593 3672 5631
rect 3722 5651 3766 5693
rect 3722 5631 3734 5651
rect 3754 5631 3766 5651
rect 3722 5593 3766 5631
rect 3848 5651 3890 5693
rect 3848 5631 3856 5651
rect 3876 5631 3890 5651
rect 3848 5593 3890 5631
rect 3940 5651 3984 5693
rect 5628 5706 5640 5726
rect 5660 5706 5672 5726
rect 3940 5631 3952 5651
rect 3972 5631 3984 5651
rect 5628 5664 5672 5706
rect 5722 5726 5764 5764
rect 5722 5706 5736 5726
rect 5756 5706 5764 5726
rect 5722 5664 5764 5706
rect 5846 5726 5890 5764
rect 5846 5706 5858 5726
rect 5878 5706 5890 5726
rect 5846 5664 5890 5706
rect 5940 5726 5982 5764
rect 5940 5706 5954 5726
rect 5974 5706 5982 5726
rect 5940 5664 5982 5706
rect 6056 5726 6098 5764
rect 6056 5706 6064 5726
rect 6084 5706 6098 5726
rect 6056 5664 6098 5706
rect 6148 5733 6193 5764
rect 6148 5726 6192 5733
rect 6148 5706 6160 5726
rect 6180 5706 6192 5726
rect 10005 5738 10049 5776
rect 6148 5664 6192 5706
rect 7784 5664 7828 5706
rect 3940 5593 3984 5631
rect 7784 5644 7796 5664
rect 7816 5644 7828 5664
rect 7784 5637 7828 5644
rect 7783 5606 7828 5637
rect 7878 5664 7920 5706
rect 7878 5644 7892 5664
rect 7912 5644 7920 5664
rect 7878 5606 7920 5644
rect 7994 5664 8036 5706
rect 7994 5644 8002 5664
rect 8022 5644 8036 5664
rect 7994 5606 8036 5644
rect 8086 5664 8130 5706
rect 8086 5644 8098 5664
rect 8118 5644 8130 5664
rect 8086 5606 8130 5644
rect 8212 5664 8254 5706
rect 8212 5644 8220 5664
rect 8240 5644 8254 5664
rect 8212 5606 8254 5644
rect 8304 5664 8348 5706
rect 10005 5718 10017 5738
rect 10037 5718 10049 5738
rect 8304 5644 8316 5664
rect 8336 5644 8348 5664
rect 10005 5676 10049 5718
rect 10099 5738 10141 5776
rect 10099 5718 10113 5738
rect 10133 5718 10141 5738
rect 10099 5676 10141 5718
rect 10223 5738 10267 5776
rect 10223 5718 10235 5738
rect 10255 5718 10267 5738
rect 10223 5676 10267 5718
rect 10317 5738 10359 5776
rect 10317 5718 10331 5738
rect 10351 5718 10359 5738
rect 10317 5676 10359 5718
rect 10433 5738 10475 5776
rect 10433 5718 10441 5738
rect 10461 5718 10475 5738
rect 10433 5676 10475 5718
rect 10525 5745 10570 5776
rect 10525 5738 10569 5745
rect 10525 5718 10537 5738
rect 10557 5718 10569 5738
rect 14369 5751 14413 5789
rect 10525 5676 10569 5718
rect 12161 5676 12205 5718
rect 8304 5606 8348 5644
rect 367 5487 411 5525
rect 367 5467 379 5487
rect 399 5467 411 5487
rect 367 5425 411 5467
rect 461 5487 503 5525
rect 461 5467 475 5487
rect 495 5467 503 5487
rect 461 5425 503 5467
rect 585 5487 629 5525
rect 585 5467 597 5487
rect 617 5467 629 5487
rect 585 5425 629 5467
rect 679 5487 721 5525
rect 679 5467 693 5487
rect 713 5467 721 5487
rect 679 5425 721 5467
rect 795 5487 837 5525
rect 795 5467 803 5487
rect 823 5467 837 5487
rect 795 5425 837 5467
rect 887 5494 932 5525
rect 887 5487 931 5494
rect 887 5467 899 5487
rect 919 5467 931 5487
rect 887 5425 931 5467
rect 12161 5656 12173 5676
rect 12193 5656 12205 5676
rect 12161 5649 12205 5656
rect 12160 5618 12205 5649
rect 12255 5676 12297 5718
rect 12255 5656 12269 5676
rect 12289 5656 12297 5676
rect 12255 5618 12297 5656
rect 12371 5676 12413 5718
rect 12371 5656 12379 5676
rect 12399 5656 12413 5676
rect 12371 5618 12413 5656
rect 12463 5676 12507 5718
rect 12463 5656 12475 5676
rect 12495 5656 12507 5676
rect 12463 5618 12507 5656
rect 12589 5676 12631 5718
rect 12589 5656 12597 5676
rect 12617 5656 12631 5676
rect 12589 5618 12631 5656
rect 12681 5676 12725 5718
rect 14369 5731 14381 5751
rect 14401 5731 14413 5751
rect 12681 5656 12693 5676
rect 12713 5656 12725 5676
rect 14369 5689 14413 5731
rect 14463 5751 14505 5789
rect 14463 5731 14477 5751
rect 14497 5731 14505 5751
rect 14463 5689 14505 5731
rect 14587 5751 14631 5789
rect 14587 5731 14599 5751
rect 14619 5731 14631 5751
rect 14587 5689 14631 5731
rect 14681 5751 14723 5789
rect 14681 5731 14695 5751
rect 14715 5731 14723 5751
rect 14681 5689 14723 5731
rect 14797 5751 14839 5789
rect 14797 5731 14805 5751
rect 14825 5731 14839 5751
rect 14797 5689 14839 5731
rect 14889 5758 14934 5789
rect 14889 5751 14933 5758
rect 14889 5731 14901 5751
rect 14921 5731 14933 5751
rect 14889 5689 14933 5731
rect 16525 5689 16569 5731
rect 12681 5618 12725 5656
rect 4731 5500 4775 5538
rect 4731 5480 4743 5500
rect 4763 5480 4775 5500
rect 2623 5423 2667 5465
rect 2623 5403 2635 5423
rect 2655 5403 2667 5423
rect 2623 5396 2667 5403
rect 2622 5365 2667 5396
rect 2717 5423 2759 5465
rect 2717 5403 2731 5423
rect 2751 5403 2759 5423
rect 2717 5365 2759 5403
rect 2833 5423 2875 5465
rect 2833 5403 2841 5423
rect 2861 5403 2875 5423
rect 2833 5365 2875 5403
rect 2925 5423 2969 5465
rect 2925 5403 2937 5423
rect 2957 5403 2969 5423
rect 2925 5365 2969 5403
rect 3051 5423 3093 5465
rect 3051 5403 3059 5423
rect 3079 5403 3093 5423
rect 3051 5365 3093 5403
rect 3143 5423 3187 5465
rect 4731 5438 4775 5480
rect 4825 5500 4867 5538
rect 4825 5480 4839 5500
rect 4859 5480 4867 5500
rect 4825 5438 4867 5480
rect 4949 5500 4993 5538
rect 4949 5480 4961 5500
rect 4981 5480 4993 5500
rect 4949 5438 4993 5480
rect 5043 5500 5085 5538
rect 5043 5480 5057 5500
rect 5077 5480 5085 5500
rect 5043 5438 5085 5480
rect 5159 5500 5201 5538
rect 5159 5480 5167 5500
rect 5187 5480 5201 5500
rect 5159 5438 5201 5480
rect 5251 5507 5296 5538
rect 5251 5500 5295 5507
rect 5251 5480 5263 5500
rect 5283 5480 5295 5500
rect 5251 5438 5295 5480
rect 16525 5669 16537 5689
rect 16557 5669 16569 5689
rect 16525 5662 16569 5669
rect 16524 5631 16569 5662
rect 16619 5689 16661 5731
rect 16619 5669 16633 5689
rect 16653 5669 16661 5689
rect 16619 5631 16661 5669
rect 16735 5689 16777 5731
rect 16735 5669 16743 5689
rect 16763 5669 16777 5689
rect 16735 5631 16777 5669
rect 16827 5689 16871 5731
rect 16827 5669 16839 5689
rect 16859 5669 16871 5689
rect 16827 5631 16871 5669
rect 16953 5689 16995 5731
rect 16953 5669 16961 5689
rect 16981 5669 16995 5689
rect 16953 5631 16995 5669
rect 17045 5689 17089 5731
rect 18635 5725 18679 5763
rect 17045 5669 17057 5689
rect 17077 5669 17089 5689
rect 17045 5631 17089 5669
rect 18635 5705 18647 5725
rect 18667 5705 18679 5725
rect 18635 5663 18679 5705
rect 18729 5725 18771 5763
rect 18729 5705 18743 5725
rect 18763 5705 18771 5725
rect 18729 5663 18771 5705
rect 18853 5725 18897 5763
rect 18853 5705 18865 5725
rect 18885 5705 18897 5725
rect 18853 5663 18897 5705
rect 18947 5725 18989 5763
rect 18947 5705 18961 5725
rect 18981 5705 18989 5725
rect 18947 5663 18989 5705
rect 19063 5725 19105 5763
rect 19063 5705 19071 5725
rect 19091 5705 19105 5725
rect 19063 5663 19105 5705
rect 19155 5732 19200 5763
rect 19155 5725 19199 5732
rect 19155 5705 19167 5725
rect 19187 5705 19199 5725
rect 22999 5738 23043 5776
rect 19155 5663 19199 5705
rect 20791 5663 20835 5705
rect 9108 5512 9152 5550
rect 9108 5492 9120 5512
rect 9140 5492 9152 5512
rect 3143 5403 3155 5423
rect 3175 5403 3187 5423
rect 3143 5365 3187 5403
rect 1165 5303 1209 5341
rect 1165 5283 1177 5303
rect 1197 5283 1209 5303
rect 1165 5241 1209 5283
rect 1259 5303 1301 5341
rect 1259 5283 1273 5303
rect 1293 5283 1301 5303
rect 1259 5241 1301 5283
rect 1383 5303 1427 5341
rect 1383 5283 1395 5303
rect 1415 5283 1427 5303
rect 1383 5241 1427 5283
rect 1477 5303 1519 5341
rect 1477 5283 1491 5303
rect 1511 5283 1519 5303
rect 1477 5241 1519 5283
rect 1593 5303 1635 5341
rect 1593 5283 1601 5303
rect 1621 5283 1635 5303
rect 1593 5241 1635 5283
rect 1685 5310 1730 5341
rect 1685 5303 1729 5310
rect 1685 5283 1697 5303
rect 1717 5283 1729 5303
rect 1685 5241 1729 5283
rect 6987 5436 7031 5478
rect 6987 5416 6999 5436
rect 7019 5416 7031 5436
rect 6987 5409 7031 5416
rect 6986 5378 7031 5409
rect 7081 5436 7123 5478
rect 7081 5416 7095 5436
rect 7115 5416 7123 5436
rect 7081 5378 7123 5416
rect 7197 5436 7239 5478
rect 7197 5416 7205 5436
rect 7225 5416 7239 5436
rect 7197 5378 7239 5416
rect 7289 5436 7333 5478
rect 7289 5416 7301 5436
rect 7321 5416 7333 5436
rect 7289 5378 7333 5416
rect 7415 5436 7457 5478
rect 7415 5416 7423 5436
rect 7443 5416 7457 5436
rect 7415 5378 7457 5416
rect 7507 5436 7551 5478
rect 9108 5450 9152 5492
rect 9202 5512 9244 5550
rect 9202 5492 9216 5512
rect 9236 5492 9244 5512
rect 9202 5450 9244 5492
rect 9326 5512 9370 5550
rect 9326 5492 9338 5512
rect 9358 5492 9370 5512
rect 9326 5450 9370 5492
rect 9420 5512 9462 5550
rect 9420 5492 9434 5512
rect 9454 5492 9462 5512
rect 9420 5450 9462 5492
rect 9536 5512 9578 5550
rect 9536 5492 9544 5512
rect 9564 5492 9578 5512
rect 9536 5450 9578 5492
rect 9628 5519 9673 5550
rect 9628 5512 9672 5519
rect 9628 5492 9640 5512
rect 9660 5492 9672 5512
rect 9628 5450 9672 5492
rect 20791 5643 20803 5663
rect 20823 5643 20835 5663
rect 20791 5636 20835 5643
rect 20790 5605 20835 5636
rect 20885 5663 20927 5705
rect 20885 5643 20899 5663
rect 20919 5643 20927 5663
rect 20885 5605 20927 5643
rect 21001 5663 21043 5705
rect 21001 5643 21009 5663
rect 21029 5643 21043 5663
rect 21001 5605 21043 5643
rect 21093 5663 21137 5705
rect 21093 5643 21105 5663
rect 21125 5643 21137 5663
rect 21093 5605 21137 5643
rect 21219 5663 21261 5705
rect 21219 5643 21227 5663
rect 21247 5643 21261 5663
rect 21219 5605 21261 5643
rect 21311 5663 21355 5705
rect 22999 5718 23011 5738
rect 23031 5718 23043 5738
rect 21311 5643 21323 5663
rect 21343 5643 21355 5663
rect 22999 5676 23043 5718
rect 23093 5738 23135 5776
rect 23093 5718 23107 5738
rect 23127 5718 23135 5738
rect 23093 5676 23135 5718
rect 23217 5738 23261 5776
rect 23217 5718 23229 5738
rect 23249 5718 23261 5738
rect 23217 5676 23261 5718
rect 23311 5738 23353 5776
rect 23311 5718 23325 5738
rect 23345 5718 23353 5738
rect 23311 5676 23353 5718
rect 23427 5738 23469 5776
rect 23427 5718 23435 5738
rect 23455 5718 23469 5738
rect 23427 5676 23469 5718
rect 23519 5745 23564 5776
rect 23519 5738 23563 5745
rect 23519 5718 23531 5738
rect 23551 5718 23563 5738
rect 27376 5750 27420 5788
rect 23519 5676 23563 5718
rect 25155 5676 25199 5718
rect 21311 5605 21355 5643
rect 13472 5525 13516 5563
rect 13472 5505 13484 5525
rect 13504 5505 13516 5525
rect 7507 5416 7519 5436
rect 7539 5416 7551 5436
rect 7507 5378 7551 5416
rect 5529 5316 5573 5354
rect 5529 5296 5541 5316
rect 5561 5296 5573 5316
rect 3421 5239 3465 5281
rect 3421 5219 3433 5239
rect 3453 5219 3465 5239
rect 3421 5212 3465 5219
rect 3420 5181 3465 5212
rect 3515 5239 3557 5281
rect 3515 5219 3529 5239
rect 3549 5219 3557 5239
rect 3515 5181 3557 5219
rect 3631 5239 3673 5281
rect 3631 5219 3639 5239
rect 3659 5219 3673 5239
rect 3631 5181 3673 5219
rect 3723 5239 3767 5281
rect 3723 5219 3735 5239
rect 3755 5219 3767 5239
rect 3723 5181 3767 5219
rect 3849 5239 3891 5281
rect 3849 5219 3857 5239
rect 3877 5219 3891 5239
rect 3849 5181 3891 5219
rect 3941 5239 3985 5281
rect 5529 5254 5573 5296
rect 5623 5316 5665 5354
rect 5623 5296 5637 5316
rect 5657 5296 5665 5316
rect 5623 5254 5665 5296
rect 5747 5316 5791 5354
rect 5747 5296 5759 5316
rect 5779 5296 5791 5316
rect 5747 5254 5791 5296
rect 5841 5316 5883 5354
rect 5841 5296 5855 5316
rect 5875 5296 5883 5316
rect 5841 5254 5883 5296
rect 5957 5316 5999 5354
rect 5957 5296 5965 5316
rect 5985 5296 5999 5316
rect 5957 5254 5999 5296
rect 6049 5323 6094 5354
rect 6049 5316 6093 5323
rect 6049 5296 6061 5316
rect 6081 5296 6093 5316
rect 6049 5254 6093 5296
rect 11364 5448 11408 5490
rect 11364 5428 11376 5448
rect 11396 5428 11408 5448
rect 11364 5421 11408 5428
rect 11363 5390 11408 5421
rect 11458 5448 11500 5490
rect 11458 5428 11472 5448
rect 11492 5428 11500 5448
rect 11458 5390 11500 5428
rect 11574 5448 11616 5490
rect 11574 5428 11582 5448
rect 11602 5428 11616 5448
rect 11574 5390 11616 5428
rect 11666 5448 11710 5490
rect 11666 5428 11678 5448
rect 11698 5428 11710 5448
rect 11666 5390 11710 5428
rect 11792 5448 11834 5490
rect 11792 5428 11800 5448
rect 11820 5428 11834 5448
rect 11792 5390 11834 5428
rect 11884 5448 11928 5490
rect 13472 5463 13516 5505
rect 13566 5525 13608 5563
rect 13566 5505 13580 5525
rect 13600 5505 13608 5525
rect 13566 5463 13608 5505
rect 13690 5525 13734 5563
rect 13690 5505 13702 5525
rect 13722 5505 13734 5525
rect 13690 5463 13734 5505
rect 13784 5525 13826 5563
rect 13784 5505 13798 5525
rect 13818 5505 13826 5525
rect 13784 5463 13826 5505
rect 13900 5525 13942 5563
rect 13900 5505 13908 5525
rect 13928 5505 13942 5525
rect 13900 5463 13942 5505
rect 13992 5532 14037 5563
rect 13992 5525 14036 5532
rect 13992 5505 14004 5525
rect 14024 5505 14036 5525
rect 13992 5463 14036 5505
rect 25155 5656 25167 5676
rect 25187 5656 25199 5676
rect 25155 5649 25199 5656
rect 25154 5618 25199 5649
rect 25249 5676 25291 5718
rect 25249 5656 25263 5676
rect 25283 5656 25291 5676
rect 25249 5618 25291 5656
rect 25365 5676 25407 5718
rect 25365 5656 25373 5676
rect 25393 5656 25407 5676
rect 25365 5618 25407 5656
rect 25457 5676 25501 5718
rect 25457 5656 25469 5676
rect 25489 5656 25501 5676
rect 25457 5618 25501 5656
rect 25583 5676 25625 5718
rect 25583 5656 25591 5676
rect 25611 5656 25625 5676
rect 25583 5618 25625 5656
rect 25675 5676 25719 5718
rect 27376 5730 27388 5750
rect 27408 5730 27420 5750
rect 25675 5656 25687 5676
rect 25707 5656 25719 5676
rect 27376 5688 27420 5730
rect 27470 5750 27512 5788
rect 27470 5730 27484 5750
rect 27504 5730 27512 5750
rect 27470 5688 27512 5730
rect 27594 5750 27638 5788
rect 27594 5730 27606 5750
rect 27626 5730 27638 5750
rect 27594 5688 27638 5730
rect 27688 5750 27730 5788
rect 27688 5730 27702 5750
rect 27722 5730 27730 5750
rect 27688 5688 27730 5730
rect 27804 5750 27846 5788
rect 27804 5730 27812 5750
rect 27832 5730 27846 5750
rect 27804 5688 27846 5730
rect 27896 5757 27941 5788
rect 27896 5750 27940 5757
rect 27896 5730 27908 5750
rect 27928 5730 27940 5750
rect 31740 5763 31784 5801
rect 27896 5688 27940 5730
rect 29532 5688 29576 5730
rect 25675 5618 25719 5656
rect 11884 5428 11896 5448
rect 11916 5428 11928 5448
rect 11884 5390 11928 5428
rect 9906 5328 9950 5366
rect 9906 5308 9918 5328
rect 9938 5308 9950 5328
rect 3941 5219 3953 5239
rect 3973 5219 3985 5239
rect 3941 5181 3985 5219
rect 7785 5252 7829 5294
rect 7785 5232 7797 5252
rect 7817 5232 7829 5252
rect 7785 5225 7829 5232
rect 7784 5194 7829 5225
rect 7879 5252 7921 5294
rect 7879 5232 7893 5252
rect 7913 5232 7921 5252
rect 7879 5194 7921 5232
rect 7995 5252 8037 5294
rect 7995 5232 8003 5252
rect 8023 5232 8037 5252
rect 7995 5194 8037 5232
rect 8087 5252 8131 5294
rect 8087 5232 8099 5252
rect 8119 5232 8131 5252
rect 8087 5194 8131 5232
rect 8213 5252 8255 5294
rect 8213 5232 8221 5252
rect 8241 5232 8255 5252
rect 8213 5194 8255 5232
rect 8305 5252 8349 5294
rect 9906 5266 9950 5308
rect 10000 5328 10042 5366
rect 10000 5308 10014 5328
rect 10034 5308 10042 5328
rect 10000 5266 10042 5308
rect 10124 5328 10168 5366
rect 10124 5308 10136 5328
rect 10156 5308 10168 5328
rect 10124 5266 10168 5308
rect 10218 5328 10260 5366
rect 10218 5308 10232 5328
rect 10252 5308 10260 5328
rect 10218 5266 10260 5308
rect 10334 5328 10376 5366
rect 10334 5308 10342 5328
rect 10362 5308 10376 5328
rect 10334 5266 10376 5308
rect 10426 5335 10471 5366
rect 10426 5328 10470 5335
rect 10426 5308 10438 5328
rect 10458 5308 10470 5328
rect 10426 5266 10470 5308
rect 15728 5461 15772 5503
rect 15728 5441 15740 5461
rect 15760 5441 15772 5461
rect 15728 5434 15772 5441
rect 15727 5403 15772 5434
rect 15822 5461 15864 5503
rect 15822 5441 15836 5461
rect 15856 5441 15864 5461
rect 15822 5403 15864 5441
rect 15938 5461 15980 5503
rect 15938 5441 15946 5461
rect 15966 5441 15980 5461
rect 15938 5403 15980 5441
rect 16030 5461 16074 5503
rect 16030 5441 16042 5461
rect 16062 5441 16074 5461
rect 16030 5403 16074 5441
rect 16156 5461 16198 5503
rect 16156 5441 16164 5461
rect 16184 5441 16198 5461
rect 16156 5403 16198 5441
rect 16248 5461 16292 5503
rect 17738 5499 17782 5537
rect 17738 5479 17750 5499
rect 17770 5479 17782 5499
rect 16248 5441 16260 5461
rect 16280 5441 16292 5461
rect 16248 5403 16292 5441
rect 17738 5437 17782 5479
rect 17832 5499 17874 5537
rect 17832 5479 17846 5499
rect 17866 5479 17874 5499
rect 17832 5437 17874 5479
rect 17956 5499 18000 5537
rect 17956 5479 17968 5499
rect 17988 5479 18000 5499
rect 17956 5437 18000 5479
rect 18050 5499 18092 5537
rect 18050 5479 18064 5499
rect 18084 5479 18092 5499
rect 18050 5437 18092 5479
rect 18166 5499 18208 5537
rect 18166 5479 18174 5499
rect 18194 5479 18208 5499
rect 18166 5437 18208 5479
rect 18258 5506 18303 5537
rect 18258 5499 18302 5506
rect 18258 5479 18270 5499
rect 18290 5479 18302 5499
rect 18258 5437 18302 5479
rect 29532 5668 29544 5688
rect 29564 5668 29576 5688
rect 29532 5661 29576 5668
rect 29531 5630 29576 5661
rect 29626 5688 29668 5730
rect 29626 5668 29640 5688
rect 29660 5668 29668 5688
rect 29626 5630 29668 5668
rect 29742 5688 29784 5730
rect 29742 5668 29750 5688
rect 29770 5668 29784 5688
rect 29742 5630 29784 5668
rect 29834 5688 29878 5730
rect 29834 5668 29846 5688
rect 29866 5668 29878 5688
rect 29834 5630 29878 5668
rect 29960 5688 30002 5730
rect 29960 5668 29968 5688
rect 29988 5668 30002 5688
rect 29960 5630 30002 5668
rect 30052 5688 30096 5730
rect 31740 5743 31752 5763
rect 31772 5743 31784 5763
rect 30052 5668 30064 5688
rect 30084 5668 30096 5688
rect 31740 5701 31784 5743
rect 31834 5763 31876 5801
rect 31834 5743 31848 5763
rect 31868 5743 31876 5763
rect 31834 5701 31876 5743
rect 31958 5763 32002 5801
rect 31958 5743 31970 5763
rect 31990 5743 32002 5763
rect 31958 5701 32002 5743
rect 32052 5763 32094 5801
rect 32052 5743 32066 5763
rect 32086 5743 32094 5763
rect 32052 5701 32094 5743
rect 32168 5763 32210 5801
rect 32168 5743 32176 5763
rect 32196 5743 32210 5763
rect 32168 5701 32210 5743
rect 32260 5770 32305 5801
rect 32260 5763 32304 5770
rect 32260 5743 32272 5763
rect 32292 5743 32304 5763
rect 32260 5701 32304 5743
rect 33896 5701 33940 5743
rect 30052 5630 30096 5668
rect 22102 5512 22146 5550
rect 22102 5492 22114 5512
rect 22134 5492 22146 5512
rect 14270 5341 14314 5379
rect 14270 5321 14282 5341
rect 14302 5321 14314 5341
rect 8305 5232 8317 5252
rect 8337 5232 8349 5252
rect 8305 5194 8349 5232
rect 368 5075 412 5113
rect 368 5055 380 5075
rect 400 5055 412 5075
rect 368 5013 412 5055
rect 462 5075 504 5113
rect 462 5055 476 5075
rect 496 5055 504 5075
rect 462 5013 504 5055
rect 586 5075 630 5113
rect 586 5055 598 5075
rect 618 5055 630 5075
rect 586 5013 630 5055
rect 680 5075 722 5113
rect 680 5055 694 5075
rect 714 5055 722 5075
rect 680 5013 722 5055
rect 796 5075 838 5113
rect 796 5055 804 5075
rect 824 5055 838 5075
rect 796 5013 838 5055
rect 888 5082 933 5113
rect 888 5075 932 5082
rect 888 5055 900 5075
rect 920 5055 932 5075
rect 12162 5264 12206 5306
rect 12162 5244 12174 5264
rect 12194 5244 12206 5264
rect 12162 5237 12206 5244
rect 12161 5206 12206 5237
rect 12256 5264 12298 5306
rect 12256 5244 12270 5264
rect 12290 5244 12298 5264
rect 12256 5206 12298 5244
rect 12372 5264 12414 5306
rect 12372 5244 12380 5264
rect 12400 5244 12414 5264
rect 12372 5206 12414 5244
rect 12464 5264 12508 5306
rect 12464 5244 12476 5264
rect 12496 5244 12508 5264
rect 12464 5206 12508 5244
rect 12590 5264 12632 5306
rect 12590 5244 12598 5264
rect 12618 5244 12632 5264
rect 12590 5206 12632 5244
rect 12682 5264 12726 5306
rect 14270 5279 14314 5321
rect 14364 5341 14406 5379
rect 14364 5321 14378 5341
rect 14398 5321 14406 5341
rect 14364 5279 14406 5321
rect 14488 5341 14532 5379
rect 14488 5321 14500 5341
rect 14520 5321 14532 5341
rect 14488 5279 14532 5321
rect 14582 5341 14624 5379
rect 14582 5321 14596 5341
rect 14616 5321 14624 5341
rect 14582 5279 14624 5321
rect 14698 5341 14740 5379
rect 14698 5321 14706 5341
rect 14726 5321 14740 5341
rect 14698 5279 14740 5321
rect 14790 5348 14835 5379
rect 14790 5341 14834 5348
rect 14790 5321 14802 5341
rect 14822 5321 14834 5341
rect 14790 5279 14834 5321
rect 19994 5435 20038 5477
rect 19994 5415 20006 5435
rect 20026 5415 20038 5435
rect 19994 5408 20038 5415
rect 19993 5377 20038 5408
rect 20088 5435 20130 5477
rect 20088 5415 20102 5435
rect 20122 5415 20130 5435
rect 20088 5377 20130 5415
rect 20204 5435 20246 5477
rect 20204 5415 20212 5435
rect 20232 5415 20246 5435
rect 20204 5377 20246 5415
rect 20296 5435 20340 5477
rect 20296 5415 20308 5435
rect 20328 5415 20340 5435
rect 20296 5377 20340 5415
rect 20422 5435 20464 5477
rect 20422 5415 20430 5435
rect 20450 5415 20464 5435
rect 20422 5377 20464 5415
rect 20514 5435 20558 5477
rect 22102 5450 22146 5492
rect 22196 5512 22238 5550
rect 22196 5492 22210 5512
rect 22230 5492 22238 5512
rect 22196 5450 22238 5492
rect 22320 5512 22364 5550
rect 22320 5492 22332 5512
rect 22352 5492 22364 5512
rect 22320 5450 22364 5492
rect 22414 5512 22456 5550
rect 22414 5492 22428 5512
rect 22448 5492 22456 5512
rect 22414 5450 22456 5492
rect 22530 5512 22572 5550
rect 22530 5492 22538 5512
rect 22558 5492 22572 5512
rect 22530 5450 22572 5492
rect 22622 5519 22667 5550
rect 22622 5512 22666 5519
rect 22622 5492 22634 5512
rect 22654 5492 22666 5512
rect 22622 5450 22666 5492
rect 33896 5681 33908 5701
rect 33928 5681 33940 5701
rect 33896 5674 33940 5681
rect 33895 5643 33940 5674
rect 33990 5701 34032 5743
rect 33990 5681 34004 5701
rect 34024 5681 34032 5701
rect 33990 5643 34032 5681
rect 34106 5701 34148 5743
rect 34106 5681 34114 5701
rect 34134 5681 34148 5701
rect 34106 5643 34148 5681
rect 34198 5701 34242 5743
rect 34198 5681 34210 5701
rect 34230 5681 34242 5701
rect 34198 5643 34242 5681
rect 34324 5701 34366 5743
rect 34324 5681 34332 5701
rect 34352 5681 34366 5701
rect 34324 5643 34366 5681
rect 34416 5701 34460 5743
rect 34416 5681 34428 5701
rect 34448 5681 34460 5701
rect 34416 5643 34460 5681
rect 26479 5524 26523 5562
rect 26479 5504 26491 5524
rect 26511 5504 26523 5524
rect 20514 5415 20526 5435
rect 20546 5415 20558 5435
rect 20514 5377 20558 5415
rect 12682 5244 12694 5264
rect 12714 5244 12726 5264
rect 12682 5206 12726 5244
rect 4732 5088 4776 5126
rect 888 5013 932 5055
rect 2319 5017 2363 5059
rect 2319 4997 2331 5017
rect 2351 4997 2363 5017
rect 2319 4990 2363 4997
rect 2318 4959 2363 4990
rect 2413 5017 2455 5059
rect 2413 4997 2427 5017
rect 2447 4997 2455 5017
rect 2413 4959 2455 4997
rect 2529 5017 2571 5059
rect 2529 4997 2537 5017
rect 2557 4997 2571 5017
rect 2529 4959 2571 4997
rect 2621 5017 2665 5059
rect 2621 4997 2633 5017
rect 2653 4997 2665 5017
rect 2621 4959 2665 4997
rect 2747 5017 2789 5059
rect 2747 4997 2755 5017
rect 2775 4997 2789 5017
rect 2747 4959 2789 4997
rect 2839 5017 2883 5059
rect 4732 5068 4744 5088
rect 4764 5068 4776 5088
rect 2839 4997 2851 5017
rect 2871 4997 2883 5017
rect 4732 5026 4776 5068
rect 4826 5088 4868 5126
rect 4826 5068 4840 5088
rect 4860 5068 4868 5088
rect 4826 5026 4868 5068
rect 4950 5088 4994 5126
rect 4950 5068 4962 5088
rect 4982 5068 4994 5088
rect 4950 5026 4994 5068
rect 5044 5088 5086 5126
rect 5044 5068 5058 5088
rect 5078 5068 5086 5088
rect 5044 5026 5086 5068
rect 5160 5088 5202 5126
rect 5160 5068 5168 5088
rect 5188 5068 5202 5088
rect 5160 5026 5202 5068
rect 5252 5095 5297 5126
rect 5252 5088 5296 5095
rect 5252 5068 5264 5088
rect 5284 5068 5296 5088
rect 16526 5277 16570 5319
rect 16526 5257 16538 5277
rect 16558 5257 16570 5277
rect 16526 5250 16570 5257
rect 16525 5219 16570 5250
rect 16620 5277 16662 5319
rect 16620 5257 16634 5277
rect 16654 5257 16662 5277
rect 16620 5219 16662 5257
rect 16736 5277 16778 5319
rect 16736 5257 16744 5277
rect 16764 5257 16778 5277
rect 16736 5219 16778 5257
rect 16828 5277 16872 5319
rect 16828 5257 16840 5277
rect 16860 5257 16872 5277
rect 16828 5219 16872 5257
rect 16954 5277 16996 5319
rect 16954 5257 16962 5277
rect 16982 5257 16996 5277
rect 16954 5219 16996 5257
rect 17046 5277 17090 5319
rect 18536 5315 18580 5353
rect 18536 5295 18548 5315
rect 18568 5295 18580 5315
rect 17046 5257 17058 5277
rect 17078 5257 17090 5277
rect 17046 5219 17090 5257
rect 18536 5253 18580 5295
rect 18630 5315 18672 5353
rect 18630 5295 18644 5315
rect 18664 5295 18672 5315
rect 18630 5253 18672 5295
rect 18754 5315 18798 5353
rect 18754 5295 18766 5315
rect 18786 5295 18798 5315
rect 18754 5253 18798 5295
rect 18848 5315 18890 5353
rect 18848 5295 18862 5315
rect 18882 5295 18890 5315
rect 18848 5253 18890 5295
rect 18964 5315 19006 5353
rect 18964 5295 18972 5315
rect 18992 5295 19006 5315
rect 18964 5253 19006 5295
rect 19056 5322 19101 5353
rect 19056 5315 19100 5322
rect 19056 5295 19068 5315
rect 19088 5295 19100 5315
rect 19056 5253 19100 5295
rect 24358 5448 24402 5490
rect 24358 5428 24370 5448
rect 24390 5428 24402 5448
rect 24358 5421 24402 5428
rect 24357 5390 24402 5421
rect 24452 5448 24494 5490
rect 24452 5428 24466 5448
rect 24486 5428 24494 5448
rect 24452 5390 24494 5428
rect 24568 5448 24610 5490
rect 24568 5428 24576 5448
rect 24596 5428 24610 5448
rect 24568 5390 24610 5428
rect 24660 5448 24704 5490
rect 24660 5428 24672 5448
rect 24692 5428 24704 5448
rect 24660 5390 24704 5428
rect 24786 5448 24828 5490
rect 24786 5428 24794 5448
rect 24814 5428 24828 5448
rect 24786 5390 24828 5428
rect 24878 5448 24922 5490
rect 26479 5462 26523 5504
rect 26573 5524 26615 5562
rect 26573 5504 26587 5524
rect 26607 5504 26615 5524
rect 26573 5462 26615 5504
rect 26697 5524 26741 5562
rect 26697 5504 26709 5524
rect 26729 5504 26741 5524
rect 26697 5462 26741 5504
rect 26791 5524 26833 5562
rect 26791 5504 26805 5524
rect 26825 5504 26833 5524
rect 26791 5462 26833 5504
rect 26907 5524 26949 5562
rect 26907 5504 26915 5524
rect 26935 5504 26949 5524
rect 26907 5462 26949 5504
rect 26999 5531 27044 5562
rect 26999 5524 27043 5531
rect 26999 5504 27011 5524
rect 27031 5504 27043 5524
rect 26999 5462 27043 5504
rect 30843 5537 30887 5575
rect 30843 5517 30855 5537
rect 30875 5517 30887 5537
rect 24878 5428 24890 5448
rect 24910 5428 24922 5448
rect 24878 5390 24922 5428
rect 22900 5328 22944 5366
rect 22900 5308 22912 5328
rect 22932 5308 22944 5328
rect 9109 5100 9153 5138
rect 5252 5026 5296 5068
rect 6683 5030 6727 5072
rect 2839 4959 2883 4997
rect 6683 5010 6695 5030
rect 6715 5010 6727 5030
rect 6683 5003 6727 5010
rect 6682 4972 6727 5003
rect 6777 5030 6819 5072
rect 6777 5010 6791 5030
rect 6811 5010 6819 5030
rect 6777 4972 6819 5010
rect 6893 5030 6935 5072
rect 6893 5010 6901 5030
rect 6921 5010 6935 5030
rect 6893 4972 6935 5010
rect 6985 5030 7029 5072
rect 6985 5010 6997 5030
rect 7017 5010 7029 5030
rect 6985 4972 7029 5010
rect 7111 5030 7153 5072
rect 7111 5010 7119 5030
rect 7139 5010 7153 5030
rect 7111 4972 7153 5010
rect 7203 5030 7247 5072
rect 9109 5080 9121 5100
rect 9141 5080 9153 5100
rect 7203 5010 7215 5030
rect 7235 5010 7247 5030
rect 9109 5038 9153 5080
rect 9203 5100 9245 5138
rect 9203 5080 9217 5100
rect 9237 5080 9245 5100
rect 9203 5038 9245 5080
rect 9327 5100 9371 5138
rect 9327 5080 9339 5100
rect 9359 5080 9371 5100
rect 9327 5038 9371 5080
rect 9421 5100 9463 5138
rect 9421 5080 9435 5100
rect 9455 5080 9463 5100
rect 9421 5038 9463 5080
rect 9537 5100 9579 5138
rect 9537 5080 9545 5100
rect 9565 5080 9579 5100
rect 9537 5038 9579 5080
rect 9629 5107 9674 5138
rect 9629 5100 9673 5107
rect 9629 5080 9641 5100
rect 9661 5080 9673 5100
rect 13473 5113 13517 5151
rect 9629 5038 9673 5080
rect 11060 5042 11104 5084
rect 7203 4972 7247 5010
rect 11060 5022 11072 5042
rect 11092 5022 11104 5042
rect 11060 5015 11104 5022
rect 11059 4984 11104 5015
rect 11154 5042 11196 5084
rect 11154 5022 11168 5042
rect 11188 5022 11196 5042
rect 11154 4984 11196 5022
rect 11270 5042 11312 5084
rect 11270 5022 11278 5042
rect 11298 5022 11312 5042
rect 11270 4984 11312 5022
rect 11362 5042 11406 5084
rect 11362 5022 11374 5042
rect 11394 5022 11406 5042
rect 11362 4984 11406 5022
rect 11488 5042 11530 5084
rect 11488 5022 11496 5042
rect 11516 5022 11530 5042
rect 11488 4984 11530 5022
rect 11580 5042 11624 5084
rect 13473 5093 13485 5113
rect 13505 5093 13517 5113
rect 11580 5022 11592 5042
rect 11612 5022 11624 5042
rect 13473 5051 13517 5093
rect 13567 5113 13609 5151
rect 13567 5093 13581 5113
rect 13601 5093 13609 5113
rect 13567 5051 13609 5093
rect 13691 5113 13735 5151
rect 13691 5093 13703 5113
rect 13723 5093 13735 5113
rect 13691 5051 13735 5093
rect 13785 5113 13827 5151
rect 13785 5093 13799 5113
rect 13819 5093 13827 5113
rect 13785 5051 13827 5093
rect 13901 5113 13943 5151
rect 13901 5093 13909 5113
rect 13929 5093 13943 5113
rect 13901 5051 13943 5093
rect 13993 5120 14038 5151
rect 13993 5113 14037 5120
rect 13993 5093 14005 5113
rect 14025 5093 14037 5113
rect 20792 5251 20836 5293
rect 20792 5231 20804 5251
rect 20824 5231 20836 5251
rect 20792 5224 20836 5231
rect 20791 5193 20836 5224
rect 20886 5251 20928 5293
rect 20886 5231 20900 5251
rect 20920 5231 20928 5251
rect 20886 5193 20928 5231
rect 21002 5251 21044 5293
rect 21002 5231 21010 5251
rect 21030 5231 21044 5251
rect 21002 5193 21044 5231
rect 21094 5251 21138 5293
rect 21094 5231 21106 5251
rect 21126 5231 21138 5251
rect 21094 5193 21138 5231
rect 21220 5251 21262 5293
rect 21220 5231 21228 5251
rect 21248 5231 21262 5251
rect 21220 5193 21262 5231
rect 21312 5251 21356 5293
rect 22900 5266 22944 5308
rect 22994 5328 23036 5366
rect 22994 5308 23008 5328
rect 23028 5308 23036 5328
rect 22994 5266 23036 5308
rect 23118 5328 23162 5366
rect 23118 5308 23130 5328
rect 23150 5308 23162 5328
rect 23118 5266 23162 5308
rect 23212 5328 23254 5366
rect 23212 5308 23226 5328
rect 23246 5308 23254 5328
rect 23212 5266 23254 5308
rect 23328 5328 23370 5366
rect 23328 5308 23336 5328
rect 23356 5308 23370 5328
rect 23328 5266 23370 5308
rect 23420 5335 23465 5366
rect 23420 5328 23464 5335
rect 23420 5308 23432 5328
rect 23452 5308 23464 5328
rect 23420 5266 23464 5308
rect 28735 5460 28779 5502
rect 28735 5440 28747 5460
rect 28767 5440 28779 5460
rect 28735 5433 28779 5440
rect 28734 5402 28779 5433
rect 28829 5460 28871 5502
rect 28829 5440 28843 5460
rect 28863 5440 28871 5460
rect 28829 5402 28871 5440
rect 28945 5460 28987 5502
rect 28945 5440 28953 5460
rect 28973 5440 28987 5460
rect 28945 5402 28987 5440
rect 29037 5460 29081 5502
rect 29037 5440 29049 5460
rect 29069 5440 29081 5460
rect 29037 5402 29081 5440
rect 29163 5460 29205 5502
rect 29163 5440 29171 5460
rect 29191 5440 29205 5460
rect 29163 5402 29205 5440
rect 29255 5460 29299 5502
rect 30843 5475 30887 5517
rect 30937 5537 30979 5575
rect 30937 5517 30951 5537
rect 30971 5517 30979 5537
rect 30937 5475 30979 5517
rect 31061 5537 31105 5575
rect 31061 5517 31073 5537
rect 31093 5517 31105 5537
rect 31061 5475 31105 5517
rect 31155 5537 31197 5575
rect 31155 5517 31169 5537
rect 31189 5517 31197 5537
rect 31155 5475 31197 5517
rect 31271 5537 31313 5575
rect 31271 5517 31279 5537
rect 31299 5517 31313 5537
rect 31271 5475 31313 5517
rect 31363 5544 31408 5575
rect 31363 5537 31407 5544
rect 31363 5517 31375 5537
rect 31395 5517 31407 5537
rect 31363 5475 31407 5517
rect 29255 5440 29267 5460
rect 29287 5440 29299 5460
rect 29255 5402 29299 5440
rect 27277 5340 27321 5378
rect 27277 5320 27289 5340
rect 27309 5320 27321 5340
rect 21312 5231 21324 5251
rect 21344 5231 21356 5251
rect 21312 5193 21356 5231
rect 25156 5264 25200 5306
rect 25156 5244 25168 5264
rect 25188 5244 25200 5264
rect 25156 5237 25200 5244
rect 25155 5206 25200 5237
rect 25250 5264 25292 5306
rect 25250 5244 25264 5264
rect 25284 5244 25292 5264
rect 25250 5206 25292 5244
rect 25366 5264 25408 5306
rect 25366 5244 25374 5264
rect 25394 5244 25408 5264
rect 25366 5206 25408 5244
rect 25458 5264 25502 5306
rect 25458 5244 25470 5264
rect 25490 5244 25502 5264
rect 25458 5206 25502 5244
rect 25584 5264 25626 5306
rect 25584 5244 25592 5264
rect 25612 5244 25626 5264
rect 25584 5206 25626 5244
rect 25676 5264 25720 5306
rect 27277 5278 27321 5320
rect 27371 5340 27413 5378
rect 27371 5320 27385 5340
rect 27405 5320 27413 5340
rect 27371 5278 27413 5320
rect 27495 5340 27539 5378
rect 27495 5320 27507 5340
rect 27527 5320 27539 5340
rect 27495 5278 27539 5320
rect 27589 5340 27631 5378
rect 27589 5320 27603 5340
rect 27623 5320 27631 5340
rect 27589 5278 27631 5320
rect 27705 5340 27747 5378
rect 27705 5320 27713 5340
rect 27733 5320 27747 5340
rect 27705 5278 27747 5320
rect 27797 5347 27842 5378
rect 27797 5340 27841 5347
rect 27797 5320 27809 5340
rect 27829 5320 27841 5340
rect 27797 5278 27841 5320
rect 33099 5473 33143 5515
rect 33099 5453 33111 5473
rect 33131 5453 33143 5473
rect 33099 5446 33143 5453
rect 33098 5415 33143 5446
rect 33193 5473 33235 5515
rect 33193 5453 33207 5473
rect 33227 5453 33235 5473
rect 33193 5415 33235 5453
rect 33309 5473 33351 5515
rect 33309 5453 33317 5473
rect 33337 5453 33351 5473
rect 33309 5415 33351 5453
rect 33401 5473 33445 5515
rect 33401 5453 33413 5473
rect 33433 5453 33445 5473
rect 33401 5415 33445 5453
rect 33527 5473 33569 5515
rect 33527 5453 33535 5473
rect 33555 5453 33569 5473
rect 33527 5415 33569 5453
rect 33619 5473 33663 5515
rect 33619 5453 33631 5473
rect 33651 5453 33663 5473
rect 33619 5415 33663 5453
rect 31641 5353 31685 5391
rect 31641 5333 31653 5353
rect 31673 5333 31685 5353
rect 25676 5244 25688 5264
rect 25708 5244 25720 5264
rect 25676 5206 25720 5244
rect 13993 5051 14037 5093
rect 15424 5055 15468 5097
rect 11580 4984 11624 5022
rect 15424 5035 15436 5055
rect 15456 5035 15468 5055
rect 15424 5028 15468 5035
rect 15423 4997 15468 5028
rect 15518 5055 15560 5097
rect 15518 5035 15532 5055
rect 15552 5035 15560 5055
rect 15518 4997 15560 5035
rect 15634 5055 15676 5097
rect 15634 5035 15642 5055
rect 15662 5035 15676 5055
rect 15634 4997 15676 5035
rect 15726 5055 15770 5097
rect 15726 5035 15738 5055
rect 15758 5035 15770 5055
rect 15726 4997 15770 5035
rect 15852 5055 15894 5097
rect 15852 5035 15860 5055
rect 15880 5035 15894 5055
rect 15852 4997 15894 5035
rect 15944 5055 15988 5097
rect 15944 5035 15956 5055
rect 15976 5035 15988 5055
rect 17739 5087 17783 5125
rect 17739 5067 17751 5087
rect 17771 5067 17783 5087
rect 15944 4997 15988 5035
rect 17739 5025 17783 5067
rect 17833 5087 17875 5125
rect 17833 5067 17847 5087
rect 17867 5067 17875 5087
rect 17833 5025 17875 5067
rect 17957 5087 18001 5125
rect 17957 5067 17969 5087
rect 17989 5067 18001 5087
rect 17957 5025 18001 5067
rect 18051 5087 18093 5125
rect 18051 5067 18065 5087
rect 18085 5067 18093 5087
rect 18051 5025 18093 5067
rect 18167 5087 18209 5125
rect 18167 5067 18175 5087
rect 18195 5067 18209 5087
rect 18167 5025 18209 5067
rect 18259 5094 18304 5125
rect 18259 5087 18303 5094
rect 18259 5067 18271 5087
rect 18291 5067 18303 5087
rect 29533 5276 29577 5318
rect 29533 5256 29545 5276
rect 29565 5256 29577 5276
rect 29533 5249 29577 5256
rect 29532 5218 29577 5249
rect 29627 5276 29669 5318
rect 29627 5256 29641 5276
rect 29661 5256 29669 5276
rect 29627 5218 29669 5256
rect 29743 5276 29785 5318
rect 29743 5256 29751 5276
rect 29771 5256 29785 5276
rect 29743 5218 29785 5256
rect 29835 5276 29879 5318
rect 29835 5256 29847 5276
rect 29867 5256 29879 5276
rect 29835 5218 29879 5256
rect 29961 5276 30003 5318
rect 29961 5256 29969 5276
rect 29989 5256 30003 5276
rect 29961 5218 30003 5256
rect 30053 5276 30097 5318
rect 31641 5291 31685 5333
rect 31735 5353 31777 5391
rect 31735 5333 31749 5353
rect 31769 5333 31777 5353
rect 31735 5291 31777 5333
rect 31859 5353 31903 5391
rect 31859 5333 31871 5353
rect 31891 5333 31903 5353
rect 31859 5291 31903 5333
rect 31953 5353 31995 5391
rect 31953 5333 31967 5353
rect 31987 5333 31995 5353
rect 31953 5291 31995 5333
rect 32069 5353 32111 5391
rect 32069 5333 32077 5353
rect 32097 5333 32111 5353
rect 32069 5291 32111 5333
rect 32161 5360 32206 5391
rect 32161 5353 32205 5360
rect 32161 5333 32173 5353
rect 32193 5333 32205 5353
rect 32161 5291 32205 5333
rect 30053 5256 30065 5276
rect 30085 5256 30097 5276
rect 30053 5218 30097 5256
rect 22103 5100 22147 5138
rect 18259 5025 18303 5067
rect 19690 5029 19734 5071
rect 19690 5009 19702 5029
rect 19722 5009 19734 5029
rect 19690 5002 19734 5009
rect 19689 4971 19734 5002
rect 19784 5029 19826 5071
rect 19784 5009 19798 5029
rect 19818 5009 19826 5029
rect 19784 4971 19826 5009
rect 19900 5029 19942 5071
rect 19900 5009 19908 5029
rect 19928 5009 19942 5029
rect 19900 4971 19942 5009
rect 19992 5029 20036 5071
rect 19992 5009 20004 5029
rect 20024 5009 20036 5029
rect 19992 4971 20036 5009
rect 20118 5029 20160 5071
rect 20118 5009 20126 5029
rect 20146 5009 20160 5029
rect 20118 4971 20160 5009
rect 20210 5029 20254 5071
rect 22103 5080 22115 5100
rect 22135 5080 22147 5100
rect 20210 5009 20222 5029
rect 20242 5009 20254 5029
rect 22103 5038 22147 5080
rect 22197 5100 22239 5138
rect 22197 5080 22211 5100
rect 22231 5080 22239 5100
rect 22197 5038 22239 5080
rect 22321 5100 22365 5138
rect 22321 5080 22333 5100
rect 22353 5080 22365 5100
rect 22321 5038 22365 5080
rect 22415 5100 22457 5138
rect 22415 5080 22429 5100
rect 22449 5080 22457 5100
rect 22415 5038 22457 5080
rect 22531 5100 22573 5138
rect 22531 5080 22539 5100
rect 22559 5080 22573 5100
rect 22531 5038 22573 5080
rect 22623 5107 22668 5138
rect 22623 5100 22667 5107
rect 22623 5080 22635 5100
rect 22655 5080 22667 5100
rect 33897 5289 33941 5331
rect 33897 5269 33909 5289
rect 33929 5269 33941 5289
rect 33897 5262 33941 5269
rect 33896 5231 33941 5262
rect 33991 5289 34033 5331
rect 33991 5269 34005 5289
rect 34025 5269 34033 5289
rect 33991 5231 34033 5269
rect 34107 5289 34149 5331
rect 34107 5269 34115 5289
rect 34135 5269 34149 5289
rect 34107 5231 34149 5269
rect 34199 5289 34243 5331
rect 34199 5269 34211 5289
rect 34231 5269 34243 5289
rect 34199 5231 34243 5269
rect 34325 5289 34367 5331
rect 34325 5269 34333 5289
rect 34353 5269 34367 5289
rect 34325 5231 34367 5269
rect 34417 5289 34461 5331
rect 34417 5269 34429 5289
rect 34449 5269 34461 5289
rect 34417 5231 34461 5269
rect 26480 5112 26524 5150
rect 22623 5038 22667 5080
rect 24054 5042 24098 5084
rect 20210 4971 20254 5009
rect 24054 5022 24066 5042
rect 24086 5022 24098 5042
rect 24054 5015 24098 5022
rect 24053 4984 24098 5015
rect 24148 5042 24190 5084
rect 24148 5022 24162 5042
rect 24182 5022 24190 5042
rect 24148 4984 24190 5022
rect 24264 5042 24306 5084
rect 24264 5022 24272 5042
rect 24292 5022 24306 5042
rect 24264 4984 24306 5022
rect 24356 5042 24400 5084
rect 24356 5022 24368 5042
rect 24388 5022 24400 5042
rect 24356 4984 24400 5022
rect 24482 5042 24524 5084
rect 24482 5022 24490 5042
rect 24510 5022 24524 5042
rect 24482 4984 24524 5022
rect 24574 5042 24618 5084
rect 26480 5092 26492 5112
rect 26512 5092 26524 5112
rect 24574 5022 24586 5042
rect 24606 5022 24618 5042
rect 26480 5050 26524 5092
rect 26574 5112 26616 5150
rect 26574 5092 26588 5112
rect 26608 5092 26616 5112
rect 26574 5050 26616 5092
rect 26698 5112 26742 5150
rect 26698 5092 26710 5112
rect 26730 5092 26742 5112
rect 26698 5050 26742 5092
rect 26792 5112 26834 5150
rect 26792 5092 26806 5112
rect 26826 5092 26834 5112
rect 26792 5050 26834 5092
rect 26908 5112 26950 5150
rect 26908 5092 26916 5112
rect 26936 5092 26950 5112
rect 26908 5050 26950 5092
rect 27000 5119 27045 5150
rect 27000 5112 27044 5119
rect 27000 5092 27012 5112
rect 27032 5092 27044 5112
rect 30844 5125 30888 5163
rect 27000 5050 27044 5092
rect 28431 5054 28475 5096
rect 24574 4984 24618 5022
rect 28431 5034 28443 5054
rect 28463 5034 28475 5054
rect 28431 5027 28475 5034
rect 28430 4996 28475 5027
rect 28525 5054 28567 5096
rect 28525 5034 28539 5054
rect 28559 5034 28567 5054
rect 28525 4996 28567 5034
rect 28641 5054 28683 5096
rect 28641 5034 28649 5054
rect 28669 5034 28683 5054
rect 28641 4996 28683 5034
rect 28733 5054 28777 5096
rect 28733 5034 28745 5054
rect 28765 5034 28777 5054
rect 28733 4996 28777 5034
rect 28859 5054 28901 5096
rect 28859 5034 28867 5054
rect 28887 5034 28901 5054
rect 28859 4996 28901 5034
rect 28951 5054 28995 5096
rect 30844 5105 30856 5125
rect 30876 5105 30888 5125
rect 28951 5034 28963 5054
rect 28983 5034 28995 5054
rect 30844 5063 30888 5105
rect 30938 5125 30980 5163
rect 30938 5105 30952 5125
rect 30972 5105 30980 5125
rect 30938 5063 30980 5105
rect 31062 5125 31106 5163
rect 31062 5105 31074 5125
rect 31094 5105 31106 5125
rect 31062 5063 31106 5105
rect 31156 5125 31198 5163
rect 31156 5105 31170 5125
rect 31190 5105 31198 5125
rect 31156 5063 31198 5105
rect 31272 5125 31314 5163
rect 31272 5105 31280 5125
rect 31300 5105 31314 5125
rect 31272 5063 31314 5105
rect 31364 5132 31409 5163
rect 31364 5125 31408 5132
rect 31364 5105 31376 5125
rect 31396 5105 31408 5125
rect 31364 5063 31408 5105
rect 32795 5067 32839 5109
rect 28951 4996 28995 5034
rect 32795 5047 32807 5067
rect 32827 5047 32839 5067
rect 32795 5040 32839 5047
rect 32794 5009 32839 5040
rect 32889 5067 32931 5109
rect 32889 5047 32903 5067
rect 32923 5047 32931 5067
rect 32889 5009 32931 5047
rect 33005 5067 33047 5109
rect 33005 5047 33013 5067
rect 33033 5047 33047 5067
rect 33005 5009 33047 5047
rect 33097 5067 33141 5109
rect 33097 5047 33109 5067
rect 33129 5047 33141 5067
rect 33097 5009 33141 5047
rect 33223 5067 33265 5109
rect 33223 5047 33231 5067
rect 33251 5047 33265 5067
rect 33223 5009 33265 5047
rect 33315 5067 33359 5109
rect 33315 5047 33327 5067
rect 33347 5047 33359 5067
rect 33315 5009 33359 5047
rect 1450 4691 1494 4729
rect 1450 4671 1462 4691
rect 1482 4671 1494 4691
rect 1450 4629 1494 4671
rect 1544 4691 1586 4729
rect 1544 4671 1558 4691
rect 1578 4671 1586 4691
rect 1544 4629 1586 4671
rect 1668 4691 1712 4729
rect 1668 4671 1680 4691
rect 1700 4671 1712 4691
rect 1668 4629 1712 4671
rect 1762 4691 1804 4729
rect 1762 4671 1776 4691
rect 1796 4671 1804 4691
rect 1762 4629 1804 4671
rect 1878 4691 1920 4729
rect 1878 4671 1886 4691
rect 1906 4671 1920 4691
rect 1878 4629 1920 4671
rect 1970 4698 2015 4729
rect 1970 4691 2014 4698
rect 1970 4671 1982 4691
rect 2002 4671 2014 4691
rect 5814 4704 5858 4742
rect 1970 4629 2014 4671
rect 3401 4633 3445 4675
rect 3401 4613 3413 4633
rect 3433 4613 3445 4633
rect 3401 4606 3445 4613
rect 3400 4575 3445 4606
rect 3495 4633 3537 4675
rect 3495 4613 3509 4633
rect 3529 4613 3537 4633
rect 3495 4575 3537 4613
rect 3611 4633 3653 4675
rect 3611 4613 3619 4633
rect 3639 4613 3653 4633
rect 3611 4575 3653 4613
rect 3703 4633 3747 4675
rect 3703 4613 3715 4633
rect 3735 4613 3747 4633
rect 3703 4575 3747 4613
rect 3829 4633 3871 4675
rect 3829 4613 3837 4633
rect 3857 4613 3871 4633
rect 3829 4575 3871 4613
rect 3921 4633 3965 4675
rect 5814 4684 5826 4704
rect 5846 4684 5858 4704
rect 3921 4613 3933 4633
rect 3953 4613 3965 4633
rect 5814 4642 5858 4684
rect 5908 4704 5950 4742
rect 5908 4684 5922 4704
rect 5942 4684 5950 4704
rect 5908 4642 5950 4684
rect 6032 4704 6076 4742
rect 6032 4684 6044 4704
rect 6064 4684 6076 4704
rect 6032 4642 6076 4684
rect 6126 4704 6168 4742
rect 6126 4684 6140 4704
rect 6160 4684 6168 4704
rect 6126 4642 6168 4684
rect 6242 4704 6284 4742
rect 6242 4684 6250 4704
rect 6270 4684 6284 4704
rect 6242 4642 6284 4684
rect 6334 4711 6379 4742
rect 6334 4704 6378 4711
rect 6334 4684 6346 4704
rect 6366 4684 6378 4704
rect 10191 4716 10235 4754
rect 6334 4642 6378 4684
rect 7765 4646 7809 4688
rect 3921 4575 3965 4613
rect 7765 4626 7777 4646
rect 7797 4626 7809 4646
rect 7765 4619 7809 4626
rect 7764 4588 7809 4619
rect 7859 4646 7901 4688
rect 7859 4626 7873 4646
rect 7893 4626 7901 4646
rect 7859 4588 7901 4626
rect 7975 4646 8017 4688
rect 7975 4626 7983 4646
rect 8003 4626 8017 4646
rect 7975 4588 8017 4626
rect 8067 4646 8111 4688
rect 8067 4626 8079 4646
rect 8099 4626 8111 4646
rect 8067 4588 8111 4626
rect 8193 4646 8235 4688
rect 8193 4626 8201 4646
rect 8221 4626 8235 4646
rect 8193 4588 8235 4626
rect 8285 4646 8329 4688
rect 10191 4696 10203 4716
rect 10223 4696 10235 4716
rect 8285 4626 8297 4646
rect 8317 4626 8329 4646
rect 10191 4654 10235 4696
rect 10285 4716 10327 4754
rect 10285 4696 10299 4716
rect 10319 4696 10327 4716
rect 10285 4654 10327 4696
rect 10409 4716 10453 4754
rect 10409 4696 10421 4716
rect 10441 4696 10453 4716
rect 10409 4654 10453 4696
rect 10503 4716 10545 4754
rect 10503 4696 10517 4716
rect 10537 4696 10545 4716
rect 10503 4654 10545 4696
rect 10619 4716 10661 4754
rect 10619 4696 10627 4716
rect 10647 4696 10661 4716
rect 10619 4654 10661 4696
rect 10711 4723 10756 4754
rect 10711 4716 10755 4723
rect 10711 4696 10723 4716
rect 10743 4696 10755 4716
rect 14555 4729 14599 4767
rect 10711 4654 10755 4696
rect 12142 4658 12186 4700
rect 8285 4588 8329 4626
rect 348 4469 392 4507
rect 348 4449 360 4469
rect 380 4449 392 4469
rect 348 4407 392 4449
rect 442 4469 484 4507
rect 442 4449 456 4469
rect 476 4449 484 4469
rect 442 4407 484 4449
rect 566 4469 610 4507
rect 566 4449 578 4469
rect 598 4449 610 4469
rect 566 4407 610 4449
rect 660 4469 702 4507
rect 660 4449 674 4469
rect 694 4449 702 4469
rect 660 4407 702 4449
rect 776 4469 818 4507
rect 776 4449 784 4469
rect 804 4449 818 4469
rect 776 4407 818 4449
rect 868 4476 913 4507
rect 868 4469 912 4476
rect 868 4449 880 4469
rect 900 4449 912 4469
rect 868 4407 912 4449
rect 12142 4638 12154 4658
rect 12174 4638 12186 4658
rect 12142 4631 12186 4638
rect 12141 4600 12186 4631
rect 12236 4658 12278 4700
rect 12236 4638 12250 4658
rect 12270 4638 12278 4658
rect 12236 4600 12278 4638
rect 12352 4658 12394 4700
rect 12352 4638 12360 4658
rect 12380 4638 12394 4658
rect 12352 4600 12394 4638
rect 12444 4658 12488 4700
rect 12444 4638 12456 4658
rect 12476 4638 12488 4658
rect 12444 4600 12488 4638
rect 12570 4658 12612 4700
rect 12570 4638 12578 4658
rect 12598 4638 12612 4658
rect 12570 4600 12612 4638
rect 12662 4658 12706 4700
rect 14555 4709 14567 4729
rect 14587 4709 14599 4729
rect 12662 4638 12674 4658
rect 12694 4638 12706 4658
rect 14555 4667 14599 4709
rect 14649 4729 14691 4767
rect 14649 4709 14663 4729
rect 14683 4709 14691 4729
rect 14649 4667 14691 4709
rect 14773 4729 14817 4767
rect 14773 4709 14785 4729
rect 14805 4709 14817 4729
rect 14773 4667 14817 4709
rect 14867 4729 14909 4767
rect 14867 4709 14881 4729
rect 14901 4709 14909 4729
rect 14867 4667 14909 4709
rect 14983 4729 15025 4767
rect 14983 4709 14991 4729
rect 15011 4709 15025 4729
rect 14983 4667 15025 4709
rect 15075 4736 15120 4767
rect 15075 4729 15119 4736
rect 15075 4709 15087 4729
rect 15107 4709 15119 4729
rect 15075 4667 15119 4709
rect 16506 4671 16550 4713
rect 12662 4600 12706 4638
rect 4712 4482 4756 4520
rect 4712 4462 4724 4482
rect 4744 4462 4756 4482
rect 2604 4405 2648 4447
rect 2604 4385 2616 4405
rect 2636 4385 2648 4405
rect 2604 4378 2648 4385
rect 2603 4347 2648 4378
rect 2698 4405 2740 4447
rect 2698 4385 2712 4405
rect 2732 4385 2740 4405
rect 2698 4347 2740 4385
rect 2814 4405 2856 4447
rect 2814 4385 2822 4405
rect 2842 4385 2856 4405
rect 2814 4347 2856 4385
rect 2906 4405 2950 4447
rect 2906 4385 2918 4405
rect 2938 4385 2950 4405
rect 2906 4347 2950 4385
rect 3032 4405 3074 4447
rect 3032 4385 3040 4405
rect 3060 4385 3074 4405
rect 3032 4347 3074 4385
rect 3124 4405 3168 4447
rect 4712 4420 4756 4462
rect 4806 4482 4848 4520
rect 4806 4462 4820 4482
rect 4840 4462 4848 4482
rect 4806 4420 4848 4462
rect 4930 4482 4974 4520
rect 4930 4462 4942 4482
rect 4962 4462 4974 4482
rect 4930 4420 4974 4462
rect 5024 4482 5066 4520
rect 5024 4462 5038 4482
rect 5058 4462 5066 4482
rect 5024 4420 5066 4462
rect 5140 4482 5182 4520
rect 5140 4462 5148 4482
rect 5168 4462 5182 4482
rect 5140 4420 5182 4462
rect 5232 4489 5277 4520
rect 5232 4482 5276 4489
rect 5232 4462 5244 4482
rect 5264 4462 5276 4482
rect 5232 4420 5276 4462
rect 16506 4651 16518 4671
rect 16538 4651 16550 4671
rect 16506 4644 16550 4651
rect 16505 4613 16550 4644
rect 16600 4671 16642 4713
rect 16600 4651 16614 4671
rect 16634 4651 16642 4671
rect 16600 4613 16642 4651
rect 16716 4671 16758 4713
rect 16716 4651 16724 4671
rect 16744 4651 16758 4671
rect 16716 4613 16758 4651
rect 16808 4671 16852 4713
rect 16808 4651 16820 4671
rect 16840 4651 16852 4671
rect 16808 4613 16852 4651
rect 16934 4671 16976 4713
rect 16934 4651 16942 4671
rect 16962 4651 16976 4671
rect 16934 4613 16976 4651
rect 17026 4671 17070 4713
rect 18821 4703 18865 4741
rect 17026 4651 17038 4671
rect 17058 4651 17070 4671
rect 17026 4613 17070 4651
rect 18821 4683 18833 4703
rect 18853 4683 18865 4703
rect 18821 4641 18865 4683
rect 18915 4703 18957 4741
rect 18915 4683 18929 4703
rect 18949 4683 18957 4703
rect 18915 4641 18957 4683
rect 19039 4703 19083 4741
rect 19039 4683 19051 4703
rect 19071 4683 19083 4703
rect 19039 4641 19083 4683
rect 19133 4703 19175 4741
rect 19133 4683 19147 4703
rect 19167 4683 19175 4703
rect 19133 4641 19175 4683
rect 19249 4703 19291 4741
rect 19249 4683 19257 4703
rect 19277 4683 19291 4703
rect 19249 4641 19291 4683
rect 19341 4710 19386 4741
rect 19341 4703 19385 4710
rect 19341 4683 19353 4703
rect 19373 4683 19385 4703
rect 23185 4716 23229 4754
rect 19341 4641 19385 4683
rect 20772 4645 20816 4687
rect 9089 4494 9133 4532
rect 9089 4474 9101 4494
rect 9121 4474 9133 4494
rect 3124 4385 3136 4405
rect 3156 4385 3168 4405
rect 3124 4347 3168 4385
rect 1146 4285 1190 4323
rect 1146 4265 1158 4285
rect 1178 4265 1190 4285
rect 1146 4223 1190 4265
rect 1240 4285 1282 4323
rect 1240 4265 1254 4285
rect 1274 4265 1282 4285
rect 1240 4223 1282 4265
rect 1364 4285 1408 4323
rect 1364 4265 1376 4285
rect 1396 4265 1408 4285
rect 1364 4223 1408 4265
rect 1458 4285 1500 4323
rect 1458 4265 1472 4285
rect 1492 4265 1500 4285
rect 1458 4223 1500 4265
rect 1574 4285 1616 4323
rect 1574 4265 1582 4285
rect 1602 4265 1616 4285
rect 1574 4223 1616 4265
rect 1666 4292 1711 4323
rect 1666 4285 1710 4292
rect 1666 4265 1678 4285
rect 1698 4265 1710 4285
rect 1666 4223 1710 4265
rect 6968 4418 7012 4460
rect 6968 4398 6980 4418
rect 7000 4398 7012 4418
rect 6968 4391 7012 4398
rect 6967 4360 7012 4391
rect 7062 4418 7104 4460
rect 7062 4398 7076 4418
rect 7096 4398 7104 4418
rect 7062 4360 7104 4398
rect 7178 4418 7220 4460
rect 7178 4398 7186 4418
rect 7206 4398 7220 4418
rect 7178 4360 7220 4398
rect 7270 4418 7314 4460
rect 7270 4398 7282 4418
rect 7302 4398 7314 4418
rect 7270 4360 7314 4398
rect 7396 4418 7438 4460
rect 7396 4398 7404 4418
rect 7424 4398 7438 4418
rect 7396 4360 7438 4398
rect 7488 4418 7532 4460
rect 9089 4432 9133 4474
rect 9183 4494 9225 4532
rect 9183 4474 9197 4494
rect 9217 4474 9225 4494
rect 9183 4432 9225 4474
rect 9307 4494 9351 4532
rect 9307 4474 9319 4494
rect 9339 4474 9351 4494
rect 9307 4432 9351 4474
rect 9401 4494 9443 4532
rect 9401 4474 9415 4494
rect 9435 4474 9443 4494
rect 9401 4432 9443 4474
rect 9517 4494 9559 4532
rect 9517 4474 9525 4494
rect 9545 4474 9559 4494
rect 9517 4432 9559 4474
rect 9609 4501 9654 4532
rect 9609 4494 9653 4501
rect 9609 4474 9621 4494
rect 9641 4474 9653 4494
rect 9609 4432 9653 4474
rect 13453 4507 13497 4545
rect 13453 4487 13465 4507
rect 13485 4487 13497 4507
rect 7488 4398 7500 4418
rect 7520 4398 7532 4418
rect 7488 4360 7532 4398
rect 5510 4298 5554 4336
rect 5510 4278 5522 4298
rect 5542 4278 5554 4298
rect 3402 4221 3446 4263
rect 3402 4201 3414 4221
rect 3434 4201 3446 4221
rect 3402 4194 3446 4201
rect 3401 4163 3446 4194
rect 3496 4221 3538 4263
rect 3496 4201 3510 4221
rect 3530 4201 3538 4221
rect 3496 4163 3538 4201
rect 3612 4221 3654 4263
rect 3612 4201 3620 4221
rect 3640 4201 3654 4221
rect 3612 4163 3654 4201
rect 3704 4221 3748 4263
rect 3704 4201 3716 4221
rect 3736 4201 3748 4221
rect 3704 4163 3748 4201
rect 3830 4221 3872 4263
rect 3830 4201 3838 4221
rect 3858 4201 3872 4221
rect 3830 4163 3872 4201
rect 3922 4221 3966 4263
rect 5510 4236 5554 4278
rect 5604 4298 5646 4336
rect 5604 4278 5618 4298
rect 5638 4278 5646 4298
rect 5604 4236 5646 4278
rect 5728 4298 5772 4336
rect 5728 4278 5740 4298
rect 5760 4278 5772 4298
rect 5728 4236 5772 4278
rect 5822 4298 5864 4336
rect 5822 4278 5836 4298
rect 5856 4278 5864 4298
rect 5822 4236 5864 4278
rect 5938 4298 5980 4336
rect 5938 4278 5946 4298
rect 5966 4278 5980 4298
rect 5938 4236 5980 4278
rect 6030 4305 6075 4336
rect 6030 4298 6074 4305
rect 6030 4278 6042 4298
rect 6062 4278 6074 4298
rect 6030 4236 6074 4278
rect 11345 4430 11389 4472
rect 11345 4410 11357 4430
rect 11377 4410 11389 4430
rect 11345 4403 11389 4410
rect 11344 4372 11389 4403
rect 11439 4430 11481 4472
rect 11439 4410 11453 4430
rect 11473 4410 11481 4430
rect 11439 4372 11481 4410
rect 11555 4430 11597 4472
rect 11555 4410 11563 4430
rect 11583 4410 11597 4430
rect 11555 4372 11597 4410
rect 11647 4430 11691 4472
rect 11647 4410 11659 4430
rect 11679 4410 11691 4430
rect 11647 4372 11691 4410
rect 11773 4430 11815 4472
rect 11773 4410 11781 4430
rect 11801 4410 11815 4430
rect 11773 4372 11815 4410
rect 11865 4430 11909 4472
rect 13453 4445 13497 4487
rect 13547 4507 13589 4545
rect 13547 4487 13561 4507
rect 13581 4487 13589 4507
rect 13547 4445 13589 4487
rect 13671 4507 13715 4545
rect 13671 4487 13683 4507
rect 13703 4487 13715 4507
rect 13671 4445 13715 4487
rect 13765 4507 13807 4545
rect 13765 4487 13779 4507
rect 13799 4487 13807 4507
rect 13765 4445 13807 4487
rect 13881 4507 13923 4545
rect 13881 4487 13889 4507
rect 13909 4487 13923 4507
rect 13881 4445 13923 4487
rect 13973 4514 14018 4545
rect 13973 4507 14017 4514
rect 13973 4487 13985 4507
rect 14005 4487 14017 4507
rect 13973 4445 14017 4487
rect 20772 4625 20784 4645
rect 20804 4625 20816 4645
rect 20772 4618 20816 4625
rect 20771 4587 20816 4618
rect 20866 4645 20908 4687
rect 20866 4625 20880 4645
rect 20900 4625 20908 4645
rect 20866 4587 20908 4625
rect 20982 4645 21024 4687
rect 20982 4625 20990 4645
rect 21010 4625 21024 4645
rect 20982 4587 21024 4625
rect 21074 4645 21118 4687
rect 21074 4625 21086 4645
rect 21106 4625 21118 4645
rect 21074 4587 21118 4625
rect 21200 4645 21242 4687
rect 21200 4625 21208 4645
rect 21228 4625 21242 4645
rect 21200 4587 21242 4625
rect 21292 4645 21336 4687
rect 23185 4696 23197 4716
rect 23217 4696 23229 4716
rect 21292 4625 21304 4645
rect 21324 4625 21336 4645
rect 23185 4654 23229 4696
rect 23279 4716 23321 4754
rect 23279 4696 23293 4716
rect 23313 4696 23321 4716
rect 23279 4654 23321 4696
rect 23403 4716 23447 4754
rect 23403 4696 23415 4716
rect 23435 4696 23447 4716
rect 23403 4654 23447 4696
rect 23497 4716 23539 4754
rect 23497 4696 23511 4716
rect 23531 4696 23539 4716
rect 23497 4654 23539 4696
rect 23613 4716 23655 4754
rect 23613 4696 23621 4716
rect 23641 4696 23655 4716
rect 23613 4654 23655 4696
rect 23705 4723 23750 4754
rect 23705 4716 23749 4723
rect 23705 4696 23717 4716
rect 23737 4696 23749 4716
rect 27562 4728 27606 4766
rect 23705 4654 23749 4696
rect 25136 4658 25180 4700
rect 21292 4587 21336 4625
rect 25136 4638 25148 4658
rect 25168 4638 25180 4658
rect 25136 4631 25180 4638
rect 25135 4600 25180 4631
rect 25230 4658 25272 4700
rect 25230 4638 25244 4658
rect 25264 4638 25272 4658
rect 25230 4600 25272 4638
rect 25346 4658 25388 4700
rect 25346 4638 25354 4658
rect 25374 4638 25388 4658
rect 25346 4600 25388 4638
rect 25438 4658 25482 4700
rect 25438 4638 25450 4658
rect 25470 4638 25482 4658
rect 25438 4600 25482 4638
rect 25564 4658 25606 4700
rect 25564 4638 25572 4658
rect 25592 4638 25606 4658
rect 25564 4600 25606 4638
rect 25656 4658 25700 4700
rect 27562 4708 27574 4728
rect 27594 4708 27606 4728
rect 25656 4638 25668 4658
rect 25688 4638 25700 4658
rect 27562 4666 27606 4708
rect 27656 4728 27698 4766
rect 27656 4708 27670 4728
rect 27690 4708 27698 4728
rect 27656 4666 27698 4708
rect 27780 4728 27824 4766
rect 27780 4708 27792 4728
rect 27812 4708 27824 4728
rect 27780 4666 27824 4708
rect 27874 4728 27916 4766
rect 27874 4708 27888 4728
rect 27908 4708 27916 4728
rect 27874 4666 27916 4708
rect 27990 4728 28032 4766
rect 27990 4708 27998 4728
rect 28018 4708 28032 4728
rect 27990 4666 28032 4708
rect 28082 4735 28127 4766
rect 28082 4728 28126 4735
rect 28082 4708 28094 4728
rect 28114 4708 28126 4728
rect 31926 4741 31970 4779
rect 28082 4666 28126 4708
rect 29513 4670 29557 4712
rect 25656 4600 25700 4638
rect 11865 4410 11877 4430
rect 11897 4410 11909 4430
rect 11865 4372 11909 4410
rect 9887 4310 9931 4348
rect 9887 4290 9899 4310
rect 9919 4290 9931 4310
rect 3922 4201 3934 4221
rect 3954 4201 3966 4221
rect 3922 4163 3966 4201
rect 7766 4234 7810 4276
rect 7766 4214 7778 4234
rect 7798 4214 7810 4234
rect 7766 4207 7810 4214
rect 7765 4176 7810 4207
rect 7860 4234 7902 4276
rect 7860 4214 7874 4234
rect 7894 4214 7902 4234
rect 7860 4176 7902 4214
rect 7976 4234 8018 4276
rect 7976 4214 7984 4234
rect 8004 4214 8018 4234
rect 7976 4176 8018 4214
rect 8068 4234 8112 4276
rect 8068 4214 8080 4234
rect 8100 4214 8112 4234
rect 8068 4176 8112 4214
rect 8194 4234 8236 4276
rect 8194 4214 8202 4234
rect 8222 4214 8236 4234
rect 8194 4176 8236 4214
rect 8286 4234 8330 4276
rect 9887 4248 9931 4290
rect 9981 4310 10023 4348
rect 9981 4290 9995 4310
rect 10015 4290 10023 4310
rect 9981 4248 10023 4290
rect 10105 4310 10149 4348
rect 10105 4290 10117 4310
rect 10137 4290 10149 4310
rect 10105 4248 10149 4290
rect 10199 4310 10241 4348
rect 10199 4290 10213 4310
rect 10233 4290 10241 4310
rect 10199 4248 10241 4290
rect 10315 4310 10357 4348
rect 10315 4290 10323 4310
rect 10343 4290 10357 4310
rect 10315 4248 10357 4290
rect 10407 4317 10452 4348
rect 10407 4310 10451 4317
rect 10407 4290 10419 4310
rect 10439 4290 10451 4310
rect 10407 4248 10451 4290
rect 15709 4443 15753 4485
rect 15709 4423 15721 4443
rect 15741 4423 15753 4443
rect 15709 4416 15753 4423
rect 15708 4385 15753 4416
rect 15803 4443 15845 4485
rect 15803 4423 15817 4443
rect 15837 4423 15845 4443
rect 15803 4385 15845 4423
rect 15919 4443 15961 4485
rect 15919 4423 15927 4443
rect 15947 4423 15961 4443
rect 15919 4385 15961 4423
rect 16011 4443 16055 4485
rect 16011 4423 16023 4443
rect 16043 4423 16055 4443
rect 16011 4385 16055 4423
rect 16137 4443 16179 4485
rect 16137 4423 16145 4443
rect 16165 4423 16179 4443
rect 16137 4385 16179 4423
rect 16229 4443 16273 4485
rect 17719 4481 17763 4519
rect 17719 4461 17731 4481
rect 17751 4461 17763 4481
rect 16229 4423 16241 4443
rect 16261 4423 16273 4443
rect 16229 4385 16273 4423
rect 17719 4419 17763 4461
rect 17813 4481 17855 4519
rect 17813 4461 17827 4481
rect 17847 4461 17855 4481
rect 17813 4419 17855 4461
rect 17937 4481 17981 4519
rect 17937 4461 17949 4481
rect 17969 4461 17981 4481
rect 17937 4419 17981 4461
rect 18031 4481 18073 4519
rect 18031 4461 18045 4481
rect 18065 4461 18073 4481
rect 18031 4419 18073 4461
rect 18147 4481 18189 4519
rect 18147 4461 18155 4481
rect 18175 4461 18189 4481
rect 18147 4419 18189 4461
rect 18239 4488 18284 4519
rect 18239 4481 18283 4488
rect 18239 4461 18251 4481
rect 18271 4461 18283 4481
rect 18239 4419 18283 4461
rect 29513 4650 29525 4670
rect 29545 4650 29557 4670
rect 29513 4643 29557 4650
rect 29512 4612 29557 4643
rect 29607 4670 29649 4712
rect 29607 4650 29621 4670
rect 29641 4650 29649 4670
rect 29607 4612 29649 4650
rect 29723 4670 29765 4712
rect 29723 4650 29731 4670
rect 29751 4650 29765 4670
rect 29723 4612 29765 4650
rect 29815 4670 29859 4712
rect 29815 4650 29827 4670
rect 29847 4650 29859 4670
rect 29815 4612 29859 4650
rect 29941 4670 29983 4712
rect 29941 4650 29949 4670
rect 29969 4650 29983 4670
rect 29941 4612 29983 4650
rect 30033 4670 30077 4712
rect 31926 4721 31938 4741
rect 31958 4721 31970 4741
rect 30033 4650 30045 4670
rect 30065 4650 30077 4670
rect 31926 4679 31970 4721
rect 32020 4741 32062 4779
rect 32020 4721 32034 4741
rect 32054 4721 32062 4741
rect 32020 4679 32062 4721
rect 32144 4741 32188 4779
rect 32144 4721 32156 4741
rect 32176 4721 32188 4741
rect 32144 4679 32188 4721
rect 32238 4741 32280 4779
rect 32238 4721 32252 4741
rect 32272 4721 32280 4741
rect 32238 4679 32280 4721
rect 32354 4741 32396 4779
rect 32354 4721 32362 4741
rect 32382 4721 32396 4741
rect 32354 4679 32396 4721
rect 32446 4748 32491 4779
rect 32446 4741 32490 4748
rect 32446 4721 32458 4741
rect 32478 4721 32490 4741
rect 32446 4679 32490 4721
rect 33877 4683 33921 4725
rect 30033 4612 30077 4650
rect 22083 4494 22127 4532
rect 22083 4474 22095 4494
rect 22115 4474 22127 4494
rect 14251 4323 14295 4361
rect 14251 4303 14263 4323
rect 14283 4303 14295 4323
rect 8286 4214 8298 4234
rect 8318 4214 8330 4234
rect 8286 4176 8330 4214
rect 349 4057 393 4095
rect 349 4037 361 4057
rect 381 4037 393 4057
rect 349 3995 393 4037
rect 443 4057 485 4095
rect 443 4037 457 4057
rect 477 4037 485 4057
rect 443 3995 485 4037
rect 567 4057 611 4095
rect 567 4037 579 4057
rect 599 4037 611 4057
rect 567 3995 611 4037
rect 661 4057 703 4095
rect 661 4037 675 4057
rect 695 4037 703 4057
rect 661 3995 703 4037
rect 777 4057 819 4095
rect 777 4037 785 4057
rect 805 4037 819 4057
rect 777 3995 819 4037
rect 869 4064 914 4095
rect 869 4057 913 4064
rect 869 4037 881 4057
rect 901 4037 913 4057
rect 12143 4246 12187 4288
rect 12143 4226 12155 4246
rect 12175 4226 12187 4246
rect 12143 4219 12187 4226
rect 12142 4188 12187 4219
rect 12237 4246 12279 4288
rect 12237 4226 12251 4246
rect 12271 4226 12279 4246
rect 12237 4188 12279 4226
rect 12353 4246 12395 4288
rect 12353 4226 12361 4246
rect 12381 4226 12395 4246
rect 12353 4188 12395 4226
rect 12445 4246 12489 4288
rect 12445 4226 12457 4246
rect 12477 4226 12489 4246
rect 12445 4188 12489 4226
rect 12571 4246 12613 4288
rect 12571 4226 12579 4246
rect 12599 4226 12613 4246
rect 12571 4188 12613 4226
rect 12663 4246 12707 4288
rect 14251 4261 14295 4303
rect 14345 4323 14387 4361
rect 14345 4303 14359 4323
rect 14379 4303 14387 4323
rect 14345 4261 14387 4303
rect 14469 4323 14513 4361
rect 14469 4303 14481 4323
rect 14501 4303 14513 4323
rect 14469 4261 14513 4303
rect 14563 4323 14605 4361
rect 14563 4303 14577 4323
rect 14597 4303 14605 4323
rect 14563 4261 14605 4303
rect 14679 4323 14721 4361
rect 14679 4303 14687 4323
rect 14707 4303 14721 4323
rect 14679 4261 14721 4303
rect 14771 4330 14816 4361
rect 14771 4323 14815 4330
rect 14771 4303 14783 4323
rect 14803 4303 14815 4323
rect 14771 4261 14815 4303
rect 19975 4417 20019 4459
rect 19975 4397 19987 4417
rect 20007 4397 20019 4417
rect 19975 4390 20019 4397
rect 19974 4359 20019 4390
rect 20069 4417 20111 4459
rect 20069 4397 20083 4417
rect 20103 4397 20111 4417
rect 20069 4359 20111 4397
rect 20185 4417 20227 4459
rect 20185 4397 20193 4417
rect 20213 4397 20227 4417
rect 20185 4359 20227 4397
rect 20277 4417 20321 4459
rect 20277 4397 20289 4417
rect 20309 4397 20321 4417
rect 20277 4359 20321 4397
rect 20403 4417 20445 4459
rect 20403 4397 20411 4417
rect 20431 4397 20445 4417
rect 20403 4359 20445 4397
rect 20495 4417 20539 4459
rect 22083 4432 22127 4474
rect 22177 4494 22219 4532
rect 22177 4474 22191 4494
rect 22211 4474 22219 4494
rect 22177 4432 22219 4474
rect 22301 4494 22345 4532
rect 22301 4474 22313 4494
rect 22333 4474 22345 4494
rect 22301 4432 22345 4474
rect 22395 4494 22437 4532
rect 22395 4474 22409 4494
rect 22429 4474 22437 4494
rect 22395 4432 22437 4474
rect 22511 4494 22553 4532
rect 22511 4474 22519 4494
rect 22539 4474 22553 4494
rect 22511 4432 22553 4474
rect 22603 4501 22648 4532
rect 22603 4494 22647 4501
rect 22603 4474 22615 4494
rect 22635 4474 22647 4494
rect 22603 4432 22647 4474
rect 33877 4663 33889 4683
rect 33909 4663 33921 4683
rect 33877 4656 33921 4663
rect 33876 4625 33921 4656
rect 33971 4683 34013 4725
rect 33971 4663 33985 4683
rect 34005 4663 34013 4683
rect 33971 4625 34013 4663
rect 34087 4683 34129 4725
rect 34087 4663 34095 4683
rect 34115 4663 34129 4683
rect 34087 4625 34129 4663
rect 34179 4683 34223 4725
rect 34179 4663 34191 4683
rect 34211 4663 34223 4683
rect 34179 4625 34223 4663
rect 34305 4683 34347 4725
rect 34305 4663 34313 4683
rect 34333 4663 34347 4683
rect 34305 4625 34347 4663
rect 34397 4683 34441 4725
rect 34397 4663 34409 4683
rect 34429 4663 34441 4683
rect 34397 4625 34441 4663
rect 26460 4506 26504 4544
rect 26460 4486 26472 4506
rect 26492 4486 26504 4506
rect 20495 4397 20507 4417
rect 20527 4397 20539 4417
rect 20495 4359 20539 4397
rect 12663 4226 12675 4246
rect 12695 4226 12707 4246
rect 12663 4188 12707 4226
rect 4713 4070 4757 4108
rect 869 3995 913 4037
rect 2505 3995 2549 4037
rect 2505 3975 2517 3995
rect 2537 3975 2549 3995
rect 2505 3968 2549 3975
rect 2504 3937 2549 3968
rect 2599 3995 2641 4037
rect 2599 3975 2613 3995
rect 2633 3975 2641 3995
rect 2599 3937 2641 3975
rect 2715 3995 2757 4037
rect 2715 3975 2723 3995
rect 2743 3975 2757 3995
rect 2715 3937 2757 3975
rect 2807 3995 2851 4037
rect 2807 3975 2819 3995
rect 2839 3975 2851 3995
rect 2807 3937 2851 3975
rect 2933 3995 2975 4037
rect 2933 3975 2941 3995
rect 2961 3975 2975 3995
rect 2933 3937 2975 3975
rect 3025 3995 3069 4037
rect 4713 4050 4725 4070
rect 4745 4050 4757 4070
rect 3025 3975 3037 3995
rect 3057 3975 3069 3995
rect 4713 4008 4757 4050
rect 4807 4070 4849 4108
rect 4807 4050 4821 4070
rect 4841 4050 4849 4070
rect 4807 4008 4849 4050
rect 4931 4070 4975 4108
rect 4931 4050 4943 4070
rect 4963 4050 4975 4070
rect 4931 4008 4975 4050
rect 5025 4070 5067 4108
rect 5025 4050 5039 4070
rect 5059 4050 5067 4070
rect 5025 4008 5067 4050
rect 5141 4070 5183 4108
rect 5141 4050 5149 4070
rect 5169 4050 5183 4070
rect 5141 4008 5183 4050
rect 5233 4077 5278 4108
rect 5233 4070 5277 4077
rect 5233 4050 5245 4070
rect 5265 4050 5277 4070
rect 16507 4259 16551 4301
rect 16507 4239 16519 4259
rect 16539 4239 16551 4259
rect 16507 4232 16551 4239
rect 16506 4201 16551 4232
rect 16601 4259 16643 4301
rect 16601 4239 16615 4259
rect 16635 4239 16643 4259
rect 16601 4201 16643 4239
rect 16717 4259 16759 4301
rect 16717 4239 16725 4259
rect 16745 4239 16759 4259
rect 16717 4201 16759 4239
rect 16809 4259 16853 4301
rect 16809 4239 16821 4259
rect 16841 4239 16853 4259
rect 16809 4201 16853 4239
rect 16935 4259 16977 4301
rect 16935 4239 16943 4259
rect 16963 4239 16977 4259
rect 16935 4201 16977 4239
rect 17027 4259 17071 4301
rect 18517 4297 18561 4335
rect 18517 4277 18529 4297
rect 18549 4277 18561 4297
rect 17027 4239 17039 4259
rect 17059 4239 17071 4259
rect 17027 4201 17071 4239
rect 18517 4235 18561 4277
rect 18611 4297 18653 4335
rect 18611 4277 18625 4297
rect 18645 4277 18653 4297
rect 18611 4235 18653 4277
rect 18735 4297 18779 4335
rect 18735 4277 18747 4297
rect 18767 4277 18779 4297
rect 18735 4235 18779 4277
rect 18829 4297 18871 4335
rect 18829 4277 18843 4297
rect 18863 4277 18871 4297
rect 18829 4235 18871 4277
rect 18945 4297 18987 4335
rect 18945 4277 18953 4297
rect 18973 4277 18987 4297
rect 18945 4235 18987 4277
rect 19037 4304 19082 4335
rect 19037 4297 19081 4304
rect 19037 4277 19049 4297
rect 19069 4277 19081 4297
rect 19037 4235 19081 4277
rect 24339 4430 24383 4472
rect 24339 4410 24351 4430
rect 24371 4410 24383 4430
rect 24339 4403 24383 4410
rect 24338 4372 24383 4403
rect 24433 4430 24475 4472
rect 24433 4410 24447 4430
rect 24467 4410 24475 4430
rect 24433 4372 24475 4410
rect 24549 4430 24591 4472
rect 24549 4410 24557 4430
rect 24577 4410 24591 4430
rect 24549 4372 24591 4410
rect 24641 4430 24685 4472
rect 24641 4410 24653 4430
rect 24673 4410 24685 4430
rect 24641 4372 24685 4410
rect 24767 4430 24809 4472
rect 24767 4410 24775 4430
rect 24795 4410 24809 4430
rect 24767 4372 24809 4410
rect 24859 4430 24903 4472
rect 26460 4444 26504 4486
rect 26554 4506 26596 4544
rect 26554 4486 26568 4506
rect 26588 4486 26596 4506
rect 26554 4444 26596 4486
rect 26678 4506 26722 4544
rect 26678 4486 26690 4506
rect 26710 4486 26722 4506
rect 26678 4444 26722 4486
rect 26772 4506 26814 4544
rect 26772 4486 26786 4506
rect 26806 4486 26814 4506
rect 26772 4444 26814 4486
rect 26888 4506 26930 4544
rect 26888 4486 26896 4506
rect 26916 4486 26930 4506
rect 26888 4444 26930 4486
rect 26980 4513 27025 4544
rect 26980 4506 27024 4513
rect 26980 4486 26992 4506
rect 27012 4486 27024 4506
rect 26980 4444 27024 4486
rect 30824 4519 30868 4557
rect 30824 4499 30836 4519
rect 30856 4499 30868 4519
rect 24859 4410 24871 4430
rect 24891 4410 24903 4430
rect 24859 4372 24903 4410
rect 22881 4310 22925 4348
rect 22881 4290 22893 4310
rect 22913 4290 22925 4310
rect 9090 4082 9134 4120
rect 5233 4008 5277 4050
rect 6869 4008 6913 4050
rect 3025 3937 3069 3975
rect 6869 3988 6881 4008
rect 6901 3988 6913 4008
rect 6869 3981 6913 3988
rect 6868 3950 6913 3981
rect 6963 4008 7005 4050
rect 6963 3988 6977 4008
rect 6997 3988 7005 4008
rect 6963 3950 7005 3988
rect 7079 4008 7121 4050
rect 7079 3988 7087 4008
rect 7107 3988 7121 4008
rect 7079 3950 7121 3988
rect 7171 4008 7215 4050
rect 7171 3988 7183 4008
rect 7203 3988 7215 4008
rect 7171 3950 7215 3988
rect 7297 4008 7339 4050
rect 7297 3988 7305 4008
rect 7325 3988 7339 4008
rect 7297 3950 7339 3988
rect 7389 4008 7433 4050
rect 9090 4062 9102 4082
rect 9122 4062 9134 4082
rect 7389 3988 7401 4008
rect 7421 3988 7433 4008
rect 9090 4020 9134 4062
rect 9184 4082 9226 4120
rect 9184 4062 9198 4082
rect 9218 4062 9226 4082
rect 9184 4020 9226 4062
rect 9308 4082 9352 4120
rect 9308 4062 9320 4082
rect 9340 4062 9352 4082
rect 9308 4020 9352 4062
rect 9402 4082 9444 4120
rect 9402 4062 9416 4082
rect 9436 4062 9444 4082
rect 9402 4020 9444 4062
rect 9518 4082 9560 4120
rect 9518 4062 9526 4082
rect 9546 4062 9560 4082
rect 9518 4020 9560 4062
rect 9610 4089 9655 4120
rect 9610 4082 9654 4089
rect 9610 4062 9622 4082
rect 9642 4062 9654 4082
rect 20773 4233 20817 4275
rect 20773 4213 20785 4233
rect 20805 4213 20817 4233
rect 20773 4206 20817 4213
rect 20772 4175 20817 4206
rect 20867 4233 20909 4275
rect 20867 4213 20881 4233
rect 20901 4213 20909 4233
rect 20867 4175 20909 4213
rect 20983 4233 21025 4275
rect 20983 4213 20991 4233
rect 21011 4213 21025 4233
rect 20983 4175 21025 4213
rect 21075 4233 21119 4275
rect 21075 4213 21087 4233
rect 21107 4213 21119 4233
rect 21075 4175 21119 4213
rect 21201 4233 21243 4275
rect 21201 4213 21209 4233
rect 21229 4213 21243 4233
rect 21201 4175 21243 4213
rect 21293 4233 21337 4275
rect 22881 4248 22925 4290
rect 22975 4310 23017 4348
rect 22975 4290 22989 4310
rect 23009 4290 23017 4310
rect 22975 4248 23017 4290
rect 23099 4310 23143 4348
rect 23099 4290 23111 4310
rect 23131 4290 23143 4310
rect 23099 4248 23143 4290
rect 23193 4310 23235 4348
rect 23193 4290 23207 4310
rect 23227 4290 23235 4310
rect 23193 4248 23235 4290
rect 23309 4310 23351 4348
rect 23309 4290 23317 4310
rect 23337 4290 23351 4310
rect 23309 4248 23351 4290
rect 23401 4317 23446 4348
rect 23401 4310 23445 4317
rect 23401 4290 23413 4310
rect 23433 4290 23445 4310
rect 23401 4248 23445 4290
rect 28716 4442 28760 4484
rect 28716 4422 28728 4442
rect 28748 4422 28760 4442
rect 28716 4415 28760 4422
rect 28715 4384 28760 4415
rect 28810 4442 28852 4484
rect 28810 4422 28824 4442
rect 28844 4422 28852 4442
rect 28810 4384 28852 4422
rect 28926 4442 28968 4484
rect 28926 4422 28934 4442
rect 28954 4422 28968 4442
rect 28926 4384 28968 4422
rect 29018 4442 29062 4484
rect 29018 4422 29030 4442
rect 29050 4422 29062 4442
rect 29018 4384 29062 4422
rect 29144 4442 29186 4484
rect 29144 4422 29152 4442
rect 29172 4422 29186 4442
rect 29144 4384 29186 4422
rect 29236 4442 29280 4484
rect 30824 4457 30868 4499
rect 30918 4519 30960 4557
rect 30918 4499 30932 4519
rect 30952 4499 30960 4519
rect 30918 4457 30960 4499
rect 31042 4519 31086 4557
rect 31042 4499 31054 4519
rect 31074 4499 31086 4519
rect 31042 4457 31086 4499
rect 31136 4519 31178 4557
rect 31136 4499 31150 4519
rect 31170 4499 31178 4519
rect 31136 4457 31178 4499
rect 31252 4519 31294 4557
rect 31252 4499 31260 4519
rect 31280 4499 31294 4519
rect 31252 4457 31294 4499
rect 31344 4526 31389 4557
rect 31344 4519 31388 4526
rect 31344 4499 31356 4519
rect 31376 4499 31388 4519
rect 31344 4457 31388 4499
rect 29236 4422 29248 4442
rect 29268 4422 29280 4442
rect 29236 4384 29280 4422
rect 27258 4322 27302 4360
rect 27258 4302 27270 4322
rect 27290 4302 27302 4322
rect 21293 4213 21305 4233
rect 21325 4213 21337 4233
rect 21293 4175 21337 4213
rect 13454 4095 13498 4133
rect 9610 4020 9654 4062
rect 11246 4020 11290 4062
rect 7389 3950 7433 3988
rect 11246 4000 11258 4020
rect 11278 4000 11290 4020
rect 11246 3993 11290 4000
rect 11245 3962 11290 3993
rect 11340 4020 11382 4062
rect 11340 4000 11354 4020
rect 11374 4000 11382 4020
rect 11340 3962 11382 4000
rect 11456 4020 11498 4062
rect 11456 4000 11464 4020
rect 11484 4000 11498 4020
rect 11456 3962 11498 4000
rect 11548 4020 11592 4062
rect 11548 4000 11560 4020
rect 11580 4000 11592 4020
rect 11548 3962 11592 4000
rect 11674 4020 11716 4062
rect 11674 4000 11682 4020
rect 11702 4000 11716 4020
rect 11674 3962 11716 4000
rect 11766 4020 11810 4062
rect 13454 4075 13466 4095
rect 13486 4075 13498 4095
rect 11766 4000 11778 4020
rect 11798 4000 11810 4020
rect 13454 4033 13498 4075
rect 13548 4095 13590 4133
rect 13548 4075 13562 4095
rect 13582 4075 13590 4095
rect 13548 4033 13590 4075
rect 13672 4095 13716 4133
rect 13672 4075 13684 4095
rect 13704 4075 13716 4095
rect 13672 4033 13716 4075
rect 13766 4095 13808 4133
rect 13766 4075 13780 4095
rect 13800 4075 13808 4095
rect 13766 4033 13808 4075
rect 13882 4095 13924 4133
rect 13882 4075 13890 4095
rect 13910 4075 13924 4095
rect 13882 4033 13924 4075
rect 13974 4102 14019 4133
rect 13974 4095 14018 4102
rect 13974 4075 13986 4095
rect 14006 4075 14018 4095
rect 25137 4246 25181 4288
rect 25137 4226 25149 4246
rect 25169 4226 25181 4246
rect 25137 4219 25181 4226
rect 25136 4188 25181 4219
rect 25231 4246 25273 4288
rect 25231 4226 25245 4246
rect 25265 4226 25273 4246
rect 25231 4188 25273 4226
rect 25347 4246 25389 4288
rect 25347 4226 25355 4246
rect 25375 4226 25389 4246
rect 25347 4188 25389 4226
rect 25439 4246 25483 4288
rect 25439 4226 25451 4246
rect 25471 4226 25483 4246
rect 25439 4188 25483 4226
rect 25565 4246 25607 4288
rect 25565 4226 25573 4246
rect 25593 4226 25607 4246
rect 25565 4188 25607 4226
rect 25657 4246 25701 4288
rect 27258 4260 27302 4302
rect 27352 4322 27394 4360
rect 27352 4302 27366 4322
rect 27386 4302 27394 4322
rect 27352 4260 27394 4302
rect 27476 4322 27520 4360
rect 27476 4302 27488 4322
rect 27508 4302 27520 4322
rect 27476 4260 27520 4302
rect 27570 4322 27612 4360
rect 27570 4302 27584 4322
rect 27604 4302 27612 4322
rect 27570 4260 27612 4302
rect 27686 4322 27728 4360
rect 27686 4302 27694 4322
rect 27714 4302 27728 4322
rect 27686 4260 27728 4302
rect 27778 4329 27823 4360
rect 27778 4322 27822 4329
rect 27778 4302 27790 4322
rect 27810 4302 27822 4322
rect 27778 4260 27822 4302
rect 33080 4455 33124 4497
rect 33080 4435 33092 4455
rect 33112 4435 33124 4455
rect 33080 4428 33124 4435
rect 33079 4397 33124 4428
rect 33174 4455 33216 4497
rect 33174 4435 33188 4455
rect 33208 4435 33216 4455
rect 33174 4397 33216 4435
rect 33290 4455 33332 4497
rect 33290 4435 33298 4455
rect 33318 4435 33332 4455
rect 33290 4397 33332 4435
rect 33382 4455 33426 4497
rect 33382 4435 33394 4455
rect 33414 4435 33426 4455
rect 33382 4397 33426 4435
rect 33508 4455 33550 4497
rect 33508 4435 33516 4455
rect 33536 4435 33550 4455
rect 33508 4397 33550 4435
rect 33600 4455 33644 4497
rect 33600 4435 33612 4455
rect 33632 4435 33644 4455
rect 33600 4397 33644 4435
rect 31622 4335 31666 4373
rect 31622 4315 31634 4335
rect 31654 4315 31666 4335
rect 25657 4226 25669 4246
rect 25689 4226 25701 4246
rect 25657 4188 25701 4226
rect 13974 4033 14018 4075
rect 15610 4033 15654 4075
rect 11766 3962 11810 4000
rect 15610 4013 15622 4033
rect 15642 4013 15654 4033
rect 15610 4006 15654 4013
rect 15609 3975 15654 4006
rect 15704 4033 15746 4075
rect 15704 4013 15718 4033
rect 15738 4013 15746 4033
rect 15704 3975 15746 4013
rect 15820 4033 15862 4075
rect 15820 4013 15828 4033
rect 15848 4013 15862 4033
rect 15820 3975 15862 4013
rect 15912 4033 15956 4075
rect 15912 4013 15924 4033
rect 15944 4013 15956 4033
rect 15912 3975 15956 4013
rect 16038 4033 16080 4075
rect 16038 4013 16046 4033
rect 16066 4013 16080 4033
rect 16038 3975 16080 4013
rect 16130 4033 16174 4075
rect 16130 4013 16142 4033
rect 16162 4013 16174 4033
rect 17720 4069 17764 4107
rect 17720 4049 17732 4069
rect 17752 4049 17764 4069
rect 16130 3975 16174 4013
rect 17720 4007 17764 4049
rect 17814 4069 17856 4107
rect 17814 4049 17828 4069
rect 17848 4049 17856 4069
rect 17814 4007 17856 4049
rect 17938 4069 17982 4107
rect 17938 4049 17950 4069
rect 17970 4049 17982 4069
rect 17938 4007 17982 4049
rect 18032 4069 18074 4107
rect 18032 4049 18046 4069
rect 18066 4049 18074 4069
rect 18032 4007 18074 4049
rect 18148 4069 18190 4107
rect 18148 4049 18156 4069
rect 18176 4049 18190 4069
rect 18148 4007 18190 4049
rect 18240 4076 18285 4107
rect 18240 4069 18284 4076
rect 18240 4049 18252 4069
rect 18272 4049 18284 4069
rect 29514 4258 29558 4300
rect 29514 4238 29526 4258
rect 29546 4238 29558 4258
rect 29514 4231 29558 4238
rect 29513 4200 29558 4231
rect 29608 4258 29650 4300
rect 29608 4238 29622 4258
rect 29642 4238 29650 4258
rect 29608 4200 29650 4238
rect 29724 4258 29766 4300
rect 29724 4238 29732 4258
rect 29752 4238 29766 4258
rect 29724 4200 29766 4238
rect 29816 4258 29860 4300
rect 29816 4238 29828 4258
rect 29848 4238 29860 4258
rect 29816 4200 29860 4238
rect 29942 4258 29984 4300
rect 29942 4238 29950 4258
rect 29970 4238 29984 4258
rect 29942 4200 29984 4238
rect 30034 4258 30078 4300
rect 31622 4273 31666 4315
rect 31716 4335 31758 4373
rect 31716 4315 31730 4335
rect 31750 4315 31758 4335
rect 31716 4273 31758 4315
rect 31840 4335 31884 4373
rect 31840 4315 31852 4335
rect 31872 4315 31884 4335
rect 31840 4273 31884 4315
rect 31934 4335 31976 4373
rect 31934 4315 31948 4335
rect 31968 4315 31976 4335
rect 31934 4273 31976 4315
rect 32050 4335 32092 4373
rect 32050 4315 32058 4335
rect 32078 4315 32092 4335
rect 32050 4273 32092 4315
rect 32142 4342 32187 4373
rect 32142 4335 32186 4342
rect 32142 4315 32154 4335
rect 32174 4315 32186 4335
rect 32142 4273 32186 4315
rect 30034 4238 30046 4258
rect 30066 4238 30078 4258
rect 30034 4200 30078 4238
rect 22084 4082 22128 4120
rect 18240 4007 18284 4049
rect 19876 4007 19920 4049
rect 19876 3987 19888 4007
rect 19908 3987 19920 4007
rect 19876 3980 19920 3987
rect 19875 3949 19920 3980
rect 19970 4007 20012 4049
rect 19970 3987 19984 4007
rect 20004 3987 20012 4007
rect 19970 3949 20012 3987
rect 20086 4007 20128 4049
rect 20086 3987 20094 4007
rect 20114 3987 20128 4007
rect 20086 3949 20128 3987
rect 20178 4007 20222 4049
rect 20178 3987 20190 4007
rect 20210 3987 20222 4007
rect 20178 3949 20222 3987
rect 20304 4007 20346 4049
rect 20304 3987 20312 4007
rect 20332 3987 20346 4007
rect 20304 3949 20346 3987
rect 20396 4007 20440 4049
rect 22084 4062 22096 4082
rect 22116 4062 22128 4082
rect 20396 3987 20408 4007
rect 20428 3987 20440 4007
rect 22084 4020 22128 4062
rect 22178 4082 22220 4120
rect 22178 4062 22192 4082
rect 22212 4062 22220 4082
rect 22178 4020 22220 4062
rect 22302 4082 22346 4120
rect 22302 4062 22314 4082
rect 22334 4062 22346 4082
rect 22302 4020 22346 4062
rect 22396 4082 22438 4120
rect 22396 4062 22410 4082
rect 22430 4062 22438 4082
rect 22396 4020 22438 4062
rect 22512 4082 22554 4120
rect 22512 4062 22520 4082
rect 22540 4062 22554 4082
rect 22512 4020 22554 4062
rect 22604 4089 22649 4120
rect 22604 4082 22648 4089
rect 22604 4062 22616 4082
rect 22636 4062 22648 4082
rect 33878 4271 33922 4313
rect 33878 4251 33890 4271
rect 33910 4251 33922 4271
rect 33878 4244 33922 4251
rect 33877 4213 33922 4244
rect 33972 4271 34014 4313
rect 33972 4251 33986 4271
rect 34006 4251 34014 4271
rect 33972 4213 34014 4251
rect 34088 4271 34130 4313
rect 34088 4251 34096 4271
rect 34116 4251 34130 4271
rect 34088 4213 34130 4251
rect 34180 4271 34224 4313
rect 34180 4251 34192 4271
rect 34212 4251 34224 4271
rect 34180 4213 34224 4251
rect 34306 4271 34348 4313
rect 34306 4251 34314 4271
rect 34334 4251 34348 4271
rect 34306 4213 34348 4251
rect 34398 4271 34442 4313
rect 34398 4251 34410 4271
rect 34430 4251 34442 4271
rect 34398 4213 34442 4251
rect 26461 4094 26505 4132
rect 22604 4020 22648 4062
rect 24240 4020 24284 4062
rect 20396 3949 20440 3987
rect 24240 4000 24252 4020
rect 24272 4000 24284 4020
rect 24240 3993 24284 4000
rect 24239 3962 24284 3993
rect 24334 4020 24376 4062
rect 24334 4000 24348 4020
rect 24368 4000 24376 4020
rect 24334 3962 24376 4000
rect 24450 4020 24492 4062
rect 24450 4000 24458 4020
rect 24478 4000 24492 4020
rect 24450 3962 24492 4000
rect 24542 4020 24586 4062
rect 24542 4000 24554 4020
rect 24574 4000 24586 4020
rect 24542 3962 24586 4000
rect 24668 4020 24710 4062
rect 24668 4000 24676 4020
rect 24696 4000 24710 4020
rect 24668 3962 24710 4000
rect 24760 4020 24804 4062
rect 26461 4074 26473 4094
rect 26493 4074 26505 4094
rect 24760 4000 24772 4020
rect 24792 4000 24804 4020
rect 26461 4032 26505 4074
rect 26555 4094 26597 4132
rect 26555 4074 26569 4094
rect 26589 4074 26597 4094
rect 26555 4032 26597 4074
rect 26679 4094 26723 4132
rect 26679 4074 26691 4094
rect 26711 4074 26723 4094
rect 26679 4032 26723 4074
rect 26773 4094 26815 4132
rect 26773 4074 26787 4094
rect 26807 4074 26815 4094
rect 26773 4032 26815 4074
rect 26889 4094 26931 4132
rect 26889 4074 26897 4094
rect 26917 4074 26931 4094
rect 26889 4032 26931 4074
rect 26981 4101 27026 4132
rect 26981 4094 27025 4101
rect 26981 4074 26993 4094
rect 27013 4074 27025 4094
rect 30825 4107 30869 4145
rect 26981 4032 27025 4074
rect 28617 4032 28661 4074
rect 24760 3962 24804 4000
rect 28617 4012 28629 4032
rect 28649 4012 28661 4032
rect 28617 4005 28661 4012
rect 28616 3974 28661 4005
rect 28711 4032 28753 4074
rect 28711 4012 28725 4032
rect 28745 4012 28753 4032
rect 28711 3974 28753 4012
rect 28827 4032 28869 4074
rect 28827 4012 28835 4032
rect 28855 4012 28869 4032
rect 28827 3974 28869 4012
rect 28919 4032 28963 4074
rect 28919 4012 28931 4032
rect 28951 4012 28963 4032
rect 28919 3974 28963 4012
rect 29045 4032 29087 4074
rect 29045 4012 29053 4032
rect 29073 4012 29087 4032
rect 29045 3974 29087 4012
rect 29137 4032 29181 4074
rect 30825 4087 30837 4107
rect 30857 4087 30869 4107
rect 29137 4012 29149 4032
rect 29169 4012 29181 4032
rect 30825 4045 30869 4087
rect 30919 4107 30961 4145
rect 30919 4087 30933 4107
rect 30953 4087 30961 4107
rect 30919 4045 30961 4087
rect 31043 4107 31087 4145
rect 31043 4087 31055 4107
rect 31075 4087 31087 4107
rect 31043 4045 31087 4087
rect 31137 4107 31179 4145
rect 31137 4087 31151 4107
rect 31171 4087 31179 4107
rect 31137 4045 31179 4087
rect 31253 4107 31295 4145
rect 31253 4087 31261 4107
rect 31281 4087 31295 4107
rect 31253 4045 31295 4087
rect 31345 4114 31390 4145
rect 31345 4107 31389 4114
rect 31345 4087 31357 4107
rect 31377 4087 31389 4107
rect 31345 4045 31389 4087
rect 32981 4045 33025 4087
rect 29137 3974 29181 4012
rect 32981 4025 32993 4045
rect 33013 4025 33025 4045
rect 32981 4018 33025 4025
rect 32980 3987 33025 4018
rect 33075 4045 33117 4087
rect 33075 4025 33089 4045
rect 33109 4025 33117 4045
rect 33075 3987 33117 4025
rect 33191 4045 33233 4087
rect 33191 4025 33199 4045
rect 33219 4025 33233 4045
rect 33191 3987 33233 4025
rect 33283 4045 33327 4087
rect 33283 4025 33295 4045
rect 33315 4025 33327 4045
rect 33283 3987 33327 4025
rect 33409 4045 33451 4087
rect 33409 4025 33417 4045
rect 33437 4025 33451 4045
rect 33409 3987 33451 4025
rect 33501 4045 33545 4087
rect 33501 4025 33513 4045
rect 33533 4025 33545 4045
rect 33501 3987 33545 4025
rect 1228 3677 1272 3715
rect 1228 3657 1240 3677
rect 1260 3657 1272 3677
rect 1228 3615 1272 3657
rect 1322 3677 1364 3715
rect 1322 3657 1336 3677
rect 1356 3657 1364 3677
rect 1322 3615 1364 3657
rect 1446 3677 1490 3715
rect 1446 3657 1458 3677
rect 1478 3657 1490 3677
rect 1446 3615 1490 3657
rect 1540 3677 1582 3715
rect 1540 3657 1554 3677
rect 1574 3657 1582 3677
rect 1540 3615 1582 3657
rect 1656 3677 1698 3715
rect 1656 3657 1664 3677
rect 1684 3657 1698 3677
rect 1656 3615 1698 3657
rect 1748 3684 1793 3715
rect 1748 3677 1792 3684
rect 1748 3657 1760 3677
rect 1780 3657 1792 3677
rect 5592 3690 5636 3728
rect 1748 3615 1792 3657
rect 3384 3615 3428 3657
rect 3384 3595 3396 3615
rect 3416 3595 3428 3615
rect 3384 3588 3428 3595
rect 3383 3557 3428 3588
rect 3478 3615 3520 3657
rect 3478 3595 3492 3615
rect 3512 3595 3520 3615
rect 3478 3557 3520 3595
rect 3594 3615 3636 3657
rect 3594 3595 3602 3615
rect 3622 3595 3636 3615
rect 3594 3557 3636 3595
rect 3686 3615 3730 3657
rect 3686 3595 3698 3615
rect 3718 3595 3730 3615
rect 3686 3557 3730 3595
rect 3812 3615 3854 3657
rect 3812 3595 3820 3615
rect 3840 3595 3854 3615
rect 3812 3557 3854 3595
rect 3904 3615 3948 3657
rect 5592 3670 5604 3690
rect 5624 3670 5636 3690
rect 3904 3595 3916 3615
rect 3936 3595 3948 3615
rect 5592 3628 5636 3670
rect 5686 3690 5728 3728
rect 5686 3670 5700 3690
rect 5720 3670 5728 3690
rect 5686 3628 5728 3670
rect 5810 3690 5854 3728
rect 5810 3670 5822 3690
rect 5842 3670 5854 3690
rect 5810 3628 5854 3670
rect 5904 3690 5946 3728
rect 5904 3670 5918 3690
rect 5938 3670 5946 3690
rect 5904 3628 5946 3670
rect 6020 3690 6062 3728
rect 6020 3670 6028 3690
rect 6048 3670 6062 3690
rect 6020 3628 6062 3670
rect 6112 3697 6157 3728
rect 6112 3690 6156 3697
rect 6112 3670 6124 3690
rect 6144 3670 6156 3690
rect 9969 3702 10013 3740
rect 6112 3628 6156 3670
rect 7748 3628 7792 3670
rect 3904 3557 3948 3595
rect 7748 3608 7760 3628
rect 7780 3608 7792 3628
rect 7748 3601 7792 3608
rect 7747 3570 7792 3601
rect 7842 3628 7884 3670
rect 7842 3608 7856 3628
rect 7876 3608 7884 3628
rect 7842 3570 7884 3608
rect 7958 3628 8000 3670
rect 7958 3608 7966 3628
rect 7986 3608 8000 3628
rect 7958 3570 8000 3608
rect 8050 3628 8094 3670
rect 8050 3608 8062 3628
rect 8082 3608 8094 3628
rect 8050 3570 8094 3608
rect 8176 3628 8218 3670
rect 8176 3608 8184 3628
rect 8204 3608 8218 3628
rect 8176 3570 8218 3608
rect 8268 3628 8312 3670
rect 9969 3682 9981 3702
rect 10001 3682 10013 3702
rect 8268 3608 8280 3628
rect 8300 3608 8312 3628
rect 9969 3640 10013 3682
rect 10063 3702 10105 3740
rect 10063 3682 10077 3702
rect 10097 3682 10105 3702
rect 10063 3640 10105 3682
rect 10187 3702 10231 3740
rect 10187 3682 10199 3702
rect 10219 3682 10231 3702
rect 10187 3640 10231 3682
rect 10281 3702 10323 3740
rect 10281 3682 10295 3702
rect 10315 3682 10323 3702
rect 10281 3640 10323 3682
rect 10397 3702 10439 3740
rect 10397 3682 10405 3702
rect 10425 3682 10439 3702
rect 10397 3640 10439 3682
rect 10489 3709 10534 3740
rect 10489 3702 10533 3709
rect 10489 3682 10501 3702
rect 10521 3682 10533 3702
rect 14333 3715 14377 3753
rect 10489 3640 10533 3682
rect 12125 3640 12169 3682
rect 8268 3570 8312 3608
rect 331 3451 375 3489
rect 331 3431 343 3451
rect 363 3431 375 3451
rect 331 3389 375 3431
rect 425 3451 467 3489
rect 425 3431 439 3451
rect 459 3431 467 3451
rect 425 3389 467 3431
rect 549 3451 593 3489
rect 549 3431 561 3451
rect 581 3431 593 3451
rect 549 3389 593 3431
rect 643 3451 685 3489
rect 643 3431 657 3451
rect 677 3431 685 3451
rect 643 3389 685 3431
rect 759 3451 801 3489
rect 759 3431 767 3451
rect 787 3431 801 3451
rect 759 3389 801 3431
rect 851 3458 896 3489
rect 851 3451 895 3458
rect 851 3431 863 3451
rect 883 3431 895 3451
rect 851 3389 895 3431
rect 12125 3620 12137 3640
rect 12157 3620 12169 3640
rect 12125 3613 12169 3620
rect 12124 3582 12169 3613
rect 12219 3640 12261 3682
rect 12219 3620 12233 3640
rect 12253 3620 12261 3640
rect 12219 3582 12261 3620
rect 12335 3640 12377 3682
rect 12335 3620 12343 3640
rect 12363 3620 12377 3640
rect 12335 3582 12377 3620
rect 12427 3640 12471 3682
rect 12427 3620 12439 3640
rect 12459 3620 12471 3640
rect 12427 3582 12471 3620
rect 12553 3640 12595 3682
rect 12553 3620 12561 3640
rect 12581 3620 12595 3640
rect 12553 3582 12595 3620
rect 12645 3640 12689 3682
rect 14333 3695 14345 3715
rect 14365 3695 14377 3715
rect 12645 3620 12657 3640
rect 12677 3620 12689 3640
rect 14333 3653 14377 3695
rect 14427 3715 14469 3753
rect 14427 3695 14441 3715
rect 14461 3695 14469 3715
rect 14427 3653 14469 3695
rect 14551 3715 14595 3753
rect 14551 3695 14563 3715
rect 14583 3695 14595 3715
rect 14551 3653 14595 3695
rect 14645 3715 14687 3753
rect 14645 3695 14659 3715
rect 14679 3695 14687 3715
rect 14645 3653 14687 3695
rect 14761 3715 14803 3753
rect 14761 3695 14769 3715
rect 14789 3695 14803 3715
rect 14761 3653 14803 3695
rect 14853 3722 14898 3753
rect 14853 3715 14897 3722
rect 14853 3695 14865 3715
rect 14885 3695 14897 3715
rect 14853 3653 14897 3695
rect 16489 3653 16533 3695
rect 12645 3582 12689 3620
rect 4695 3464 4739 3502
rect 4695 3444 4707 3464
rect 4727 3444 4739 3464
rect 2587 3387 2631 3429
rect 2587 3367 2599 3387
rect 2619 3367 2631 3387
rect 2587 3360 2631 3367
rect 2586 3329 2631 3360
rect 2681 3387 2723 3429
rect 2681 3367 2695 3387
rect 2715 3367 2723 3387
rect 2681 3329 2723 3367
rect 2797 3387 2839 3429
rect 2797 3367 2805 3387
rect 2825 3367 2839 3387
rect 2797 3329 2839 3367
rect 2889 3387 2933 3429
rect 2889 3367 2901 3387
rect 2921 3367 2933 3387
rect 2889 3329 2933 3367
rect 3015 3387 3057 3429
rect 3015 3367 3023 3387
rect 3043 3367 3057 3387
rect 3015 3329 3057 3367
rect 3107 3387 3151 3429
rect 4695 3402 4739 3444
rect 4789 3464 4831 3502
rect 4789 3444 4803 3464
rect 4823 3444 4831 3464
rect 4789 3402 4831 3444
rect 4913 3464 4957 3502
rect 4913 3444 4925 3464
rect 4945 3444 4957 3464
rect 4913 3402 4957 3444
rect 5007 3464 5049 3502
rect 5007 3444 5021 3464
rect 5041 3444 5049 3464
rect 5007 3402 5049 3444
rect 5123 3464 5165 3502
rect 5123 3444 5131 3464
rect 5151 3444 5165 3464
rect 5123 3402 5165 3444
rect 5215 3471 5260 3502
rect 5215 3464 5259 3471
rect 5215 3444 5227 3464
rect 5247 3444 5259 3464
rect 5215 3402 5259 3444
rect 16489 3633 16501 3653
rect 16521 3633 16533 3653
rect 16489 3626 16533 3633
rect 16488 3595 16533 3626
rect 16583 3653 16625 3695
rect 16583 3633 16597 3653
rect 16617 3633 16625 3653
rect 16583 3595 16625 3633
rect 16699 3653 16741 3695
rect 16699 3633 16707 3653
rect 16727 3633 16741 3653
rect 16699 3595 16741 3633
rect 16791 3653 16835 3695
rect 16791 3633 16803 3653
rect 16823 3633 16835 3653
rect 16791 3595 16835 3633
rect 16917 3653 16959 3695
rect 16917 3633 16925 3653
rect 16945 3633 16959 3653
rect 16917 3595 16959 3633
rect 17009 3653 17053 3695
rect 18599 3689 18643 3727
rect 17009 3633 17021 3653
rect 17041 3633 17053 3653
rect 17009 3595 17053 3633
rect 18599 3669 18611 3689
rect 18631 3669 18643 3689
rect 18599 3627 18643 3669
rect 18693 3689 18735 3727
rect 18693 3669 18707 3689
rect 18727 3669 18735 3689
rect 18693 3627 18735 3669
rect 18817 3689 18861 3727
rect 18817 3669 18829 3689
rect 18849 3669 18861 3689
rect 18817 3627 18861 3669
rect 18911 3689 18953 3727
rect 18911 3669 18925 3689
rect 18945 3669 18953 3689
rect 18911 3627 18953 3669
rect 19027 3689 19069 3727
rect 19027 3669 19035 3689
rect 19055 3669 19069 3689
rect 19027 3627 19069 3669
rect 19119 3696 19164 3727
rect 19119 3689 19163 3696
rect 19119 3669 19131 3689
rect 19151 3669 19163 3689
rect 22963 3702 23007 3740
rect 19119 3627 19163 3669
rect 20755 3627 20799 3669
rect 9072 3476 9116 3514
rect 9072 3456 9084 3476
rect 9104 3456 9116 3476
rect 3107 3367 3119 3387
rect 3139 3367 3151 3387
rect 3107 3329 3151 3367
rect 1129 3267 1173 3305
rect 1129 3247 1141 3267
rect 1161 3247 1173 3267
rect 1129 3205 1173 3247
rect 1223 3267 1265 3305
rect 1223 3247 1237 3267
rect 1257 3247 1265 3267
rect 1223 3205 1265 3247
rect 1347 3267 1391 3305
rect 1347 3247 1359 3267
rect 1379 3247 1391 3267
rect 1347 3205 1391 3247
rect 1441 3267 1483 3305
rect 1441 3247 1455 3267
rect 1475 3247 1483 3267
rect 1441 3205 1483 3247
rect 1557 3267 1599 3305
rect 1557 3247 1565 3267
rect 1585 3247 1599 3267
rect 1557 3205 1599 3247
rect 1649 3274 1694 3305
rect 1649 3267 1693 3274
rect 1649 3247 1661 3267
rect 1681 3247 1693 3267
rect 1649 3205 1693 3247
rect 6951 3400 6995 3442
rect 6951 3380 6963 3400
rect 6983 3380 6995 3400
rect 6951 3373 6995 3380
rect 6950 3342 6995 3373
rect 7045 3400 7087 3442
rect 7045 3380 7059 3400
rect 7079 3380 7087 3400
rect 7045 3342 7087 3380
rect 7161 3400 7203 3442
rect 7161 3380 7169 3400
rect 7189 3380 7203 3400
rect 7161 3342 7203 3380
rect 7253 3400 7297 3442
rect 7253 3380 7265 3400
rect 7285 3380 7297 3400
rect 7253 3342 7297 3380
rect 7379 3400 7421 3442
rect 7379 3380 7387 3400
rect 7407 3380 7421 3400
rect 7379 3342 7421 3380
rect 7471 3400 7515 3442
rect 9072 3414 9116 3456
rect 9166 3476 9208 3514
rect 9166 3456 9180 3476
rect 9200 3456 9208 3476
rect 9166 3414 9208 3456
rect 9290 3476 9334 3514
rect 9290 3456 9302 3476
rect 9322 3456 9334 3476
rect 9290 3414 9334 3456
rect 9384 3476 9426 3514
rect 9384 3456 9398 3476
rect 9418 3456 9426 3476
rect 9384 3414 9426 3456
rect 9500 3476 9542 3514
rect 9500 3456 9508 3476
rect 9528 3456 9542 3476
rect 9500 3414 9542 3456
rect 9592 3483 9637 3514
rect 9592 3476 9636 3483
rect 9592 3456 9604 3476
rect 9624 3456 9636 3476
rect 9592 3414 9636 3456
rect 20755 3607 20767 3627
rect 20787 3607 20799 3627
rect 20755 3600 20799 3607
rect 20754 3569 20799 3600
rect 20849 3627 20891 3669
rect 20849 3607 20863 3627
rect 20883 3607 20891 3627
rect 20849 3569 20891 3607
rect 20965 3627 21007 3669
rect 20965 3607 20973 3627
rect 20993 3607 21007 3627
rect 20965 3569 21007 3607
rect 21057 3627 21101 3669
rect 21057 3607 21069 3627
rect 21089 3607 21101 3627
rect 21057 3569 21101 3607
rect 21183 3627 21225 3669
rect 21183 3607 21191 3627
rect 21211 3607 21225 3627
rect 21183 3569 21225 3607
rect 21275 3627 21319 3669
rect 22963 3682 22975 3702
rect 22995 3682 23007 3702
rect 21275 3607 21287 3627
rect 21307 3607 21319 3627
rect 22963 3640 23007 3682
rect 23057 3702 23099 3740
rect 23057 3682 23071 3702
rect 23091 3682 23099 3702
rect 23057 3640 23099 3682
rect 23181 3702 23225 3740
rect 23181 3682 23193 3702
rect 23213 3682 23225 3702
rect 23181 3640 23225 3682
rect 23275 3702 23317 3740
rect 23275 3682 23289 3702
rect 23309 3682 23317 3702
rect 23275 3640 23317 3682
rect 23391 3702 23433 3740
rect 23391 3682 23399 3702
rect 23419 3682 23433 3702
rect 23391 3640 23433 3682
rect 23483 3709 23528 3740
rect 23483 3702 23527 3709
rect 23483 3682 23495 3702
rect 23515 3682 23527 3702
rect 27340 3714 27384 3752
rect 23483 3640 23527 3682
rect 25119 3640 25163 3682
rect 21275 3569 21319 3607
rect 13436 3489 13480 3527
rect 13436 3469 13448 3489
rect 13468 3469 13480 3489
rect 7471 3380 7483 3400
rect 7503 3380 7515 3400
rect 7471 3342 7515 3380
rect 5493 3280 5537 3318
rect 5493 3260 5505 3280
rect 5525 3260 5537 3280
rect 3385 3203 3429 3245
rect 3385 3183 3397 3203
rect 3417 3183 3429 3203
rect 3385 3176 3429 3183
rect 3384 3145 3429 3176
rect 3479 3203 3521 3245
rect 3479 3183 3493 3203
rect 3513 3183 3521 3203
rect 3479 3145 3521 3183
rect 3595 3203 3637 3245
rect 3595 3183 3603 3203
rect 3623 3183 3637 3203
rect 3595 3145 3637 3183
rect 3687 3203 3731 3245
rect 3687 3183 3699 3203
rect 3719 3183 3731 3203
rect 3687 3145 3731 3183
rect 3813 3203 3855 3245
rect 3813 3183 3821 3203
rect 3841 3183 3855 3203
rect 3813 3145 3855 3183
rect 3905 3203 3949 3245
rect 5493 3218 5537 3260
rect 5587 3280 5629 3318
rect 5587 3260 5601 3280
rect 5621 3260 5629 3280
rect 5587 3218 5629 3260
rect 5711 3280 5755 3318
rect 5711 3260 5723 3280
rect 5743 3260 5755 3280
rect 5711 3218 5755 3260
rect 5805 3280 5847 3318
rect 5805 3260 5819 3280
rect 5839 3260 5847 3280
rect 5805 3218 5847 3260
rect 5921 3280 5963 3318
rect 5921 3260 5929 3280
rect 5949 3260 5963 3280
rect 5921 3218 5963 3260
rect 6013 3287 6058 3318
rect 6013 3280 6057 3287
rect 6013 3260 6025 3280
rect 6045 3260 6057 3280
rect 6013 3218 6057 3260
rect 11328 3412 11372 3454
rect 11328 3392 11340 3412
rect 11360 3392 11372 3412
rect 11328 3385 11372 3392
rect 11327 3354 11372 3385
rect 11422 3412 11464 3454
rect 11422 3392 11436 3412
rect 11456 3392 11464 3412
rect 11422 3354 11464 3392
rect 11538 3412 11580 3454
rect 11538 3392 11546 3412
rect 11566 3392 11580 3412
rect 11538 3354 11580 3392
rect 11630 3412 11674 3454
rect 11630 3392 11642 3412
rect 11662 3392 11674 3412
rect 11630 3354 11674 3392
rect 11756 3412 11798 3454
rect 11756 3392 11764 3412
rect 11784 3392 11798 3412
rect 11756 3354 11798 3392
rect 11848 3412 11892 3454
rect 13436 3427 13480 3469
rect 13530 3489 13572 3527
rect 13530 3469 13544 3489
rect 13564 3469 13572 3489
rect 13530 3427 13572 3469
rect 13654 3489 13698 3527
rect 13654 3469 13666 3489
rect 13686 3469 13698 3489
rect 13654 3427 13698 3469
rect 13748 3489 13790 3527
rect 13748 3469 13762 3489
rect 13782 3469 13790 3489
rect 13748 3427 13790 3469
rect 13864 3489 13906 3527
rect 13864 3469 13872 3489
rect 13892 3469 13906 3489
rect 13864 3427 13906 3469
rect 13956 3496 14001 3527
rect 13956 3489 14000 3496
rect 13956 3469 13968 3489
rect 13988 3469 14000 3489
rect 13956 3427 14000 3469
rect 25119 3620 25131 3640
rect 25151 3620 25163 3640
rect 25119 3613 25163 3620
rect 25118 3582 25163 3613
rect 25213 3640 25255 3682
rect 25213 3620 25227 3640
rect 25247 3620 25255 3640
rect 25213 3582 25255 3620
rect 25329 3640 25371 3682
rect 25329 3620 25337 3640
rect 25357 3620 25371 3640
rect 25329 3582 25371 3620
rect 25421 3640 25465 3682
rect 25421 3620 25433 3640
rect 25453 3620 25465 3640
rect 25421 3582 25465 3620
rect 25547 3640 25589 3682
rect 25547 3620 25555 3640
rect 25575 3620 25589 3640
rect 25547 3582 25589 3620
rect 25639 3640 25683 3682
rect 27340 3694 27352 3714
rect 27372 3694 27384 3714
rect 25639 3620 25651 3640
rect 25671 3620 25683 3640
rect 27340 3652 27384 3694
rect 27434 3714 27476 3752
rect 27434 3694 27448 3714
rect 27468 3694 27476 3714
rect 27434 3652 27476 3694
rect 27558 3714 27602 3752
rect 27558 3694 27570 3714
rect 27590 3694 27602 3714
rect 27558 3652 27602 3694
rect 27652 3714 27694 3752
rect 27652 3694 27666 3714
rect 27686 3694 27694 3714
rect 27652 3652 27694 3694
rect 27768 3714 27810 3752
rect 27768 3694 27776 3714
rect 27796 3694 27810 3714
rect 27768 3652 27810 3694
rect 27860 3721 27905 3752
rect 27860 3714 27904 3721
rect 27860 3694 27872 3714
rect 27892 3694 27904 3714
rect 31704 3727 31748 3765
rect 27860 3652 27904 3694
rect 29496 3652 29540 3694
rect 25639 3582 25683 3620
rect 11848 3392 11860 3412
rect 11880 3392 11892 3412
rect 11848 3354 11892 3392
rect 9870 3292 9914 3330
rect 9870 3272 9882 3292
rect 9902 3272 9914 3292
rect 3905 3183 3917 3203
rect 3937 3183 3949 3203
rect 3905 3145 3949 3183
rect 7749 3216 7793 3258
rect 7749 3196 7761 3216
rect 7781 3196 7793 3216
rect 7749 3189 7793 3196
rect 7748 3158 7793 3189
rect 7843 3216 7885 3258
rect 7843 3196 7857 3216
rect 7877 3196 7885 3216
rect 7843 3158 7885 3196
rect 7959 3216 8001 3258
rect 7959 3196 7967 3216
rect 7987 3196 8001 3216
rect 7959 3158 8001 3196
rect 8051 3216 8095 3258
rect 8051 3196 8063 3216
rect 8083 3196 8095 3216
rect 8051 3158 8095 3196
rect 8177 3216 8219 3258
rect 8177 3196 8185 3216
rect 8205 3196 8219 3216
rect 8177 3158 8219 3196
rect 8269 3216 8313 3258
rect 9870 3230 9914 3272
rect 9964 3292 10006 3330
rect 9964 3272 9978 3292
rect 9998 3272 10006 3292
rect 9964 3230 10006 3272
rect 10088 3292 10132 3330
rect 10088 3272 10100 3292
rect 10120 3272 10132 3292
rect 10088 3230 10132 3272
rect 10182 3292 10224 3330
rect 10182 3272 10196 3292
rect 10216 3272 10224 3292
rect 10182 3230 10224 3272
rect 10298 3292 10340 3330
rect 10298 3272 10306 3292
rect 10326 3272 10340 3292
rect 10298 3230 10340 3272
rect 10390 3299 10435 3330
rect 10390 3292 10434 3299
rect 10390 3272 10402 3292
rect 10422 3272 10434 3292
rect 10390 3230 10434 3272
rect 15692 3425 15736 3467
rect 15692 3405 15704 3425
rect 15724 3405 15736 3425
rect 15692 3398 15736 3405
rect 15691 3367 15736 3398
rect 15786 3425 15828 3467
rect 15786 3405 15800 3425
rect 15820 3405 15828 3425
rect 15786 3367 15828 3405
rect 15902 3425 15944 3467
rect 15902 3405 15910 3425
rect 15930 3405 15944 3425
rect 15902 3367 15944 3405
rect 15994 3425 16038 3467
rect 15994 3405 16006 3425
rect 16026 3405 16038 3425
rect 15994 3367 16038 3405
rect 16120 3425 16162 3467
rect 16120 3405 16128 3425
rect 16148 3405 16162 3425
rect 16120 3367 16162 3405
rect 16212 3425 16256 3467
rect 17702 3463 17746 3501
rect 17702 3443 17714 3463
rect 17734 3443 17746 3463
rect 16212 3405 16224 3425
rect 16244 3405 16256 3425
rect 16212 3367 16256 3405
rect 17702 3401 17746 3443
rect 17796 3463 17838 3501
rect 17796 3443 17810 3463
rect 17830 3443 17838 3463
rect 17796 3401 17838 3443
rect 17920 3463 17964 3501
rect 17920 3443 17932 3463
rect 17952 3443 17964 3463
rect 17920 3401 17964 3443
rect 18014 3463 18056 3501
rect 18014 3443 18028 3463
rect 18048 3443 18056 3463
rect 18014 3401 18056 3443
rect 18130 3463 18172 3501
rect 18130 3443 18138 3463
rect 18158 3443 18172 3463
rect 18130 3401 18172 3443
rect 18222 3470 18267 3501
rect 18222 3463 18266 3470
rect 18222 3443 18234 3463
rect 18254 3443 18266 3463
rect 18222 3401 18266 3443
rect 29496 3632 29508 3652
rect 29528 3632 29540 3652
rect 29496 3625 29540 3632
rect 29495 3594 29540 3625
rect 29590 3652 29632 3694
rect 29590 3632 29604 3652
rect 29624 3632 29632 3652
rect 29590 3594 29632 3632
rect 29706 3652 29748 3694
rect 29706 3632 29714 3652
rect 29734 3632 29748 3652
rect 29706 3594 29748 3632
rect 29798 3652 29842 3694
rect 29798 3632 29810 3652
rect 29830 3632 29842 3652
rect 29798 3594 29842 3632
rect 29924 3652 29966 3694
rect 29924 3632 29932 3652
rect 29952 3632 29966 3652
rect 29924 3594 29966 3632
rect 30016 3652 30060 3694
rect 31704 3707 31716 3727
rect 31736 3707 31748 3727
rect 30016 3632 30028 3652
rect 30048 3632 30060 3652
rect 31704 3665 31748 3707
rect 31798 3727 31840 3765
rect 31798 3707 31812 3727
rect 31832 3707 31840 3727
rect 31798 3665 31840 3707
rect 31922 3727 31966 3765
rect 31922 3707 31934 3727
rect 31954 3707 31966 3727
rect 31922 3665 31966 3707
rect 32016 3727 32058 3765
rect 32016 3707 32030 3727
rect 32050 3707 32058 3727
rect 32016 3665 32058 3707
rect 32132 3727 32174 3765
rect 32132 3707 32140 3727
rect 32160 3707 32174 3727
rect 32132 3665 32174 3707
rect 32224 3734 32269 3765
rect 32224 3727 32268 3734
rect 32224 3707 32236 3727
rect 32256 3707 32268 3727
rect 32224 3665 32268 3707
rect 33860 3665 33904 3707
rect 30016 3594 30060 3632
rect 22066 3476 22110 3514
rect 22066 3456 22078 3476
rect 22098 3456 22110 3476
rect 14234 3305 14278 3343
rect 14234 3285 14246 3305
rect 14266 3285 14278 3305
rect 8269 3196 8281 3216
rect 8301 3196 8313 3216
rect 8269 3158 8313 3196
rect 332 3039 376 3077
rect 332 3019 344 3039
rect 364 3019 376 3039
rect 332 2977 376 3019
rect 426 3039 468 3077
rect 426 3019 440 3039
rect 460 3019 468 3039
rect 426 2977 468 3019
rect 550 3039 594 3077
rect 550 3019 562 3039
rect 582 3019 594 3039
rect 550 2977 594 3019
rect 644 3039 686 3077
rect 644 3019 658 3039
rect 678 3019 686 3039
rect 644 2977 686 3019
rect 760 3039 802 3077
rect 760 3019 768 3039
rect 788 3019 802 3039
rect 760 2977 802 3019
rect 852 3046 897 3077
rect 852 3039 896 3046
rect 852 3019 864 3039
rect 884 3019 896 3039
rect 12126 3228 12170 3270
rect 12126 3208 12138 3228
rect 12158 3208 12170 3228
rect 12126 3201 12170 3208
rect 12125 3170 12170 3201
rect 12220 3228 12262 3270
rect 12220 3208 12234 3228
rect 12254 3208 12262 3228
rect 12220 3170 12262 3208
rect 12336 3228 12378 3270
rect 12336 3208 12344 3228
rect 12364 3208 12378 3228
rect 12336 3170 12378 3208
rect 12428 3228 12472 3270
rect 12428 3208 12440 3228
rect 12460 3208 12472 3228
rect 12428 3170 12472 3208
rect 12554 3228 12596 3270
rect 12554 3208 12562 3228
rect 12582 3208 12596 3228
rect 12554 3170 12596 3208
rect 12646 3228 12690 3270
rect 14234 3243 14278 3285
rect 14328 3305 14370 3343
rect 14328 3285 14342 3305
rect 14362 3285 14370 3305
rect 14328 3243 14370 3285
rect 14452 3305 14496 3343
rect 14452 3285 14464 3305
rect 14484 3285 14496 3305
rect 14452 3243 14496 3285
rect 14546 3305 14588 3343
rect 14546 3285 14560 3305
rect 14580 3285 14588 3305
rect 14546 3243 14588 3285
rect 14662 3305 14704 3343
rect 14662 3285 14670 3305
rect 14690 3285 14704 3305
rect 14662 3243 14704 3285
rect 14754 3312 14799 3343
rect 14754 3305 14798 3312
rect 14754 3285 14766 3305
rect 14786 3285 14798 3305
rect 14754 3243 14798 3285
rect 19958 3399 20002 3441
rect 19958 3379 19970 3399
rect 19990 3379 20002 3399
rect 19958 3372 20002 3379
rect 19957 3341 20002 3372
rect 20052 3399 20094 3441
rect 20052 3379 20066 3399
rect 20086 3379 20094 3399
rect 20052 3341 20094 3379
rect 20168 3399 20210 3441
rect 20168 3379 20176 3399
rect 20196 3379 20210 3399
rect 20168 3341 20210 3379
rect 20260 3399 20304 3441
rect 20260 3379 20272 3399
rect 20292 3379 20304 3399
rect 20260 3341 20304 3379
rect 20386 3399 20428 3441
rect 20386 3379 20394 3399
rect 20414 3379 20428 3399
rect 20386 3341 20428 3379
rect 20478 3399 20522 3441
rect 22066 3414 22110 3456
rect 22160 3476 22202 3514
rect 22160 3456 22174 3476
rect 22194 3456 22202 3476
rect 22160 3414 22202 3456
rect 22284 3476 22328 3514
rect 22284 3456 22296 3476
rect 22316 3456 22328 3476
rect 22284 3414 22328 3456
rect 22378 3476 22420 3514
rect 22378 3456 22392 3476
rect 22412 3456 22420 3476
rect 22378 3414 22420 3456
rect 22494 3476 22536 3514
rect 22494 3456 22502 3476
rect 22522 3456 22536 3476
rect 22494 3414 22536 3456
rect 22586 3483 22631 3514
rect 22586 3476 22630 3483
rect 22586 3456 22598 3476
rect 22618 3456 22630 3476
rect 22586 3414 22630 3456
rect 33860 3645 33872 3665
rect 33892 3645 33904 3665
rect 33860 3638 33904 3645
rect 33859 3607 33904 3638
rect 33954 3665 33996 3707
rect 33954 3645 33968 3665
rect 33988 3645 33996 3665
rect 33954 3607 33996 3645
rect 34070 3665 34112 3707
rect 34070 3645 34078 3665
rect 34098 3645 34112 3665
rect 34070 3607 34112 3645
rect 34162 3665 34206 3707
rect 34162 3645 34174 3665
rect 34194 3645 34206 3665
rect 34162 3607 34206 3645
rect 34288 3665 34330 3707
rect 34288 3645 34296 3665
rect 34316 3645 34330 3665
rect 34288 3607 34330 3645
rect 34380 3665 34424 3707
rect 34380 3645 34392 3665
rect 34412 3645 34424 3665
rect 34380 3607 34424 3645
rect 26443 3488 26487 3526
rect 26443 3468 26455 3488
rect 26475 3468 26487 3488
rect 20478 3379 20490 3399
rect 20510 3379 20522 3399
rect 20478 3341 20522 3379
rect 12646 3208 12658 3228
rect 12678 3208 12690 3228
rect 12646 3170 12690 3208
rect 4696 3052 4740 3090
rect 852 2977 896 3019
rect 2422 2979 2466 3021
rect 2422 2959 2434 2979
rect 2454 2959 2466 2979
rect 2422 2952 2466 2959
rect 2421 2921 2466 2952
rect 2516 2979 2558 3021
rect 2516 2959 2530 2979
rect 2550 2959 2558 2979
rect 2516 2921 2558 2959
rect 2632 2979 2674 3021
rect 2632 2959 2640 2979
rect 2660 2959 2674 2979
rect 2632 2921 2674 2959
rect 2724 2979 2768 3021
rect 2724 2959 2736 2979
rect 2756 2959 2768 2979
rect 2724 2921 2768 2959
rect 2850 2979 2892 3021
rect 2850 2959 2858 2979
rect 2878 2959 2892 2979
rect 2850 2921 2892 2959
rect 2942 2979 2986 3021
rect 4696 3032 4708 3052
rect 4728 3032 4740 3052
rect 2942 2959 2954 2979
rect 2974 2959 2986 2979
rect 4696 2990 4740 3032
rect 4790 3052 4832 3090
rect 4790 3032 4804 3052
rect 4824 3032 4832 3052
rect 4790 2990 4832 3032
rect 4914 3052 4958 3090
rect 4914 3032 4926 3052
rect 4946 3032 4958 3052
rect 4914 2990 4958 3032
rect 5008 3052 5050 3090
rect 5008 3032 5022 3052
rect 5042 3032 5050 3052
rect 5008 2990 5050 3032
rect 5124 3052 5166 3090
rect 5124 3032 5132 3052
rect 5152 3032 5166 3052
rect 5124 2990 5166 3032
rect 5216 3059 5261 3090
rect 5216 3052 5260 3059
rect 5216 3032 5228 3052
rect 5248 3032 5260 3052
rect 16490 3241 16534 3283
rect 16490 3221 16502 3241
rect 16522 3221 16534 3241
rect 16490 3214 16534 3221
rect 16489 3183 16534 3214
rect 16584 3241 16626 3283
rect 16584 3221 16598 3241
rect 16618 3221 16626 3241
rect 16584 3183 16626 3221
rect 16700 3241 16742 3283
rect 16700 3221 16708 3241
rect 16728 3221 16742 3241
rect 16700 3183 16742 3221
rect 16792 3241 16836 3283
rect 16792 3221 16804 3241
rect 16824 3221 16836 3241
rect 16792 3183 16836 3221
rect 16918 3241 16960 3283
rect 16918 3221 16926 3241
rect 16946 3221 16960 3241
rect 16918 3183 16960 3221
rect 17010 3241 17054 3283
rect 18500 3279 18544 3317
rect 18500 3259 18512 3279
rect 18532 3259 18544 3279
rect 17010 3221 17022 3241
rect 17042 3221 17054 3241
rect 17010 3183 17054 3221
rect 18500 3217 18544 3259
rect 18594 3279 18636 3317
rect 18594 3259 18608 3279
rect 18628 3259 18636 3279
rect 18594 3217 18636 3259
rect 18718 3279 18762 3317
rect 18718 3259 18730 3279
rect 18750 3259 18762 3279
rect 18718 3217 18762 3259
rect 18812 3279 18854 3317
rect 18812 3259 18826 3279
rect 18846 3259 18854 3279
rect 18812 3217 18854 3259
rect 18928 3279 18970 3317
rect 18928 3259 18936 3279
rect 18956 3259 18970 3279
rect 18928 3217 18970 3259
rect 19020 3286 19065 3317
rect 19020 3279 19064 3286
rect 19020 3259 19032 3279
rect 19052 3259 19064 3279
rect 19020 3217 19064 3259
rect 24322 3412 24366 3454
rect 24322 3392 24334 3412
rect 24354 3392 24366 3412
rect 24322 3385 24366 3392
rect 24321 3354 24366 3385
rect 24416 3412 24458 3454
rect 24416 3392 24430 3412
rect 24450 3392 24458 3412
rect 24416 3354 24458 3392
rect 24532 3412 24574 3454
rect 24532 3392 24540 3412
rect 24560 3392 24574 3412
rect 24532 3354 24574 3392
rect 24624 3412 24668 3454
rect 24624 3392 24636 3412
rect 24656 3392 24668 3412
rect 24624 3354 24668 3392
rect 24750 3412 24792 3454
rect 24750 3392 24758 3412
rect 24778 3392 24792 3412
rect 24750 3354 24792 3392
rect 24842 3412 24886 3454
rect 26443 3426 26487 3468
rect 26537 3488 26579 3526
rect 26537 3468 26551 3488
rect 26571 3468 26579 3488
rect 26537 3426 26579 3468
rect 26661 3488 26705 3526
rect 26661 3468 26673 3488
rect 26693 3468 26705 3488
rect 26661 3426 26705 3468
rect 26755 3488 26797 3526
rect 26755 3468 26769 3488
rect 26789 3468 26797 3488
rect 26755 3426 26797 3468
rect 26871 3488 26913 3526
rect 26871 3468 26879 3488
rect 26899 3468 26913 3488
rect 26871 3426 26913 3468
rect 26963 3495 27008 3526
rect 26963 3488 27007 3495
rect 26963 3468 26975 3488
rect 26995 3468 27007 3488
rect 26963 3426 27007 3468
rect 30807 3501 30851 3539
rect 30807 3481 30819 3501
rect 30839 3481 30851 3501
rect 24842 3392 24854 3412
rect 24874 3392 24886 3412
rect 24842 3354 24886 3392
rect 22864 3292 22908 3330
rect 22864 3272 22876 3292
rect 22896 3272 22908 3292
rect 9073 3064 9117 3102
rect 5216 2990 5260 3032
rect 6786 2992 6830 3034
rect 2942 2921 2986 2959
rect 6786 2972 6798 2992
rect 6818 2972 6830 2992
rect 6786 2965 6830 2972
rect 6785 2934 6830 2965
rect 6880 2992 6922 3034
rect 6880 2972 6894 2992
rect 6914 2972 6922 2992
rect 6880 2934 6922 2972
rect 6996 2992 7038 3034
rect 6996 2972 7004 2992
rect 7024 2972 7038 2992
rect 6996 2934 7038 2972
rect 7088 2992 7132 3034
rect 7088 2972 7100 2992
rect 7120 2972 7132 2992
rect 7088 2934 7132 2972
rect 7214 2992 7256 3034
rect 7214 2972 7222 2992
rect 7242 2972 7256 2992
rect 7214 2934 7256 2972
rect 7306 2992 7350 3034
rect 9073 3044 9085 3064
rect 9105 3044 9117 3064
rect 7306 2972 7318 2992
rect 7338 2972 7350 2992
rect 9073 3002 9117 3044
rect 9167 3064 9209 3102
rect 9167 3044 9181 3064
rect 9201 3044 9209 3064
rect 9167 3002 9209 3044
rect 9291 3064 9335 3102
rect 9291 3044 9303 3064
rect 9323 3044 9335 3064
rect 9291 3002 9335 3044
rect 9385 3064 9427 3102
rect 9385 3044 9399 3064
rect 9419 3044 9427 3064
rect 9385 3002 9427 3044
rect 9501 3064 9543 3102
rect 9501 3044 9509 3064
rect 9529 3044 9543 3064
rect 9501 3002 9543 3044
rect 9593 3071 9638 3102
rect 9593 3064 9637 3071
rect 9593 3044 9605 3064
rect 9625 3044 9637 3064
rect 20756 3215 20800 3257
rect 20756 3195 20768 3215
rect 20788 3195 20800 3215
rect 20756 3188 20800 3195
rect 20755 3157 20800 3188
rect 20850 3215 20892 3257
rect 20850 3195 20864 3215
rect 20884 3195 20892 3215
rect 20850 3157 20892 3195
rect 20966 3215 21008 3257
rect 20966 3195 20974 3215
rect 20994 3195 21008 3215
rect 20966 3157 21008 3195
rect 21058 3215 21102 3257
rect 21058 3195 21070 3215
rect 21090 3195 21102 3215
rect 21058 3157 21102 3195
rect 21184 3215 21226 3257
rect 21184 3195 21192 3215
rect 21212 3195 21226 3215
rect 21184 3157 21226 3195
rect 21276 3215 21320 3257
rect 22864 3230 22908 3272
rect 22958 3292 23000 3330
rect 22958 3272 22972 3292
rect 22992 3272 23000 3292
rect 22958 3230 23000 3272
rect 23082 3292 23126 3330
rect 23082 3272 23094 3292
rect 23114 3272 23126 3292
rect 23082 3230 23126 3272
rect 23176 3292 23218 3330
rect 23176 3272 23190 3292
rect 23210 3272 23218 3292
rect 23176 3230 23218 3272
rect 23292 3292 23334 3330
rect 23292 3272 23300 3292
rect 23320 3272 23334 3292
rect 23292 3230 23334 3272
rect 23384 3299 23429 3330
rect 23384 3292 23428 3299
rect 23384 3272 23396 3292
rect 23416 3272 23428 3292
rect 23384 3230 23428 3272
rect 28699 3424 28743 3466
rect 28699 3404 28711 3424
rect 28731 3404 28743 3424
rect 28699 3397 28743 3404
rect 28698 3366 28743 3397
rect 28793 3424 28835 3466
rect 28793 3404 28807 3424
rect 28827 3404 28835 3424
rect 28793 3366 28835 3404
rect 28909 3424 28951 3466
rect 28909 3404 28917 3424
rect 28937 3404 28951 3424
rect 28909 3366 28951 3404
rect 29001 3424 29045 3466
rect 29001 3404 29013 3424
rect 29033 3404 29045 3424
rect 29001 3366 29045 3404
rect 29127 3424 29169 3466
rect 29127 3404 29135 3424
rect 29155 3404 29169 3424
rect 29127 3366 29169 3404
rect 29219 3424 29263 3466
rect 30807 3439 30851 3481
rect 30901 3501 30943 3539
rect 30901 3481 30915 3501
rect 30935 3481 30943 3501
rect 30901 3439 30943 3481
rect 31025 3501 31069 3539
rect 31025 3481 31037 3501
rect 31057 3481 31069 3501
rect 31025 3439 31069 3481
rect 31119 3501 31161 3539
rect 31119 3481 31133 3501
rect 31153 3481 31161 3501
rect 31119 3439 31161 3481
rect 31235 3501 31277 3539
rect 31235 3481 31243 3501
rect 31263 3481 31277 3501
rect 31235 3439 31277 3481
rect 31327 3508 31372 3539
rect 31327 3501 31371 3508
rect 31327 3481 31339 3501
rect 31359 3481 31371 3501
rect 31327 3439 31371 3481
rect 29219 3404 29231 3424
rect 29251 3404 29263 3424
rect 29219 3366 29263 3404
rect 27241 3304 27285 3342
rect 27241 3284 27253 3304
rect 27273 3284 27285 3304
rect 21276 3195 21288 3215
rect 21308 3195 21320 3215
rect 21276 3157 21320 3195
rect 13437 3077 13481 3115
rect 9593 3002 9637 3044
rect 11163 3004 11207 3046
rect 7306 2934 7350 2972
rect 11163 2984 11175 3004
rect 11195 2984 11207 3004
rect 11163 2977 11207 2984
rect 11162 2946 11207 2977
rect 11257 3004 11299 3046
rect 11257 2984 11271 3004
rect 11291 2984 11299 3004
rect 11257 2946 11299 2984
rect 11373 3004 11415 3046
rect 11373 2984 11381 3004
rect 11401 2984 11415 3004
rect 11373 2946 11415 2984
rect 11465 3004 11509 3046
rect 11465 2984 11477 3004
rect 11497 2984 11509 3004
rect 11465 2946 11509 2984
rect 11591 3004 11633 3046
rect 11591 2984 11599 3004
rect 11619 2984 11633 3004
rect 11591 2946 11633 2984
rect 11683 3004 11727 3046
rect 13437 3057 13449 3077
rect 13469 3057 13481 3077
rect 11683 2984 11695 3004
rect 11715 2984 11727 3004
rect 13437 3015 13481 3057
rect 13531 3077 13573 3115
rect 13531 3057 13545 3077
rect 13565 3057 13573 3077
rect 13531 3015 13573 3057
rect 13655 3077 13699 3115
rect 13655 3057 13667 3077
rect 13687 3057 13699 3077
rect 13655 3015 13699 3057
rect 13749 3077 13791 3115
rect 13749 3057 13763 3077
rect 13783 3057 13791 3077
rect 13749 3015 13791 3057
rect 13865 3077 13907 3115
rect 13865 3057 13873 3077
rect 13893 3057 13907 3077
rect 13865 3015 13907 3057
rect 13957 3084 14002 3115
rect 13957 3077 14001 3084
rect 13957 3057 13969 3077
rect 13989 3057 14001 3077
rect 25120 3228 25164 3270
rect 25120 3208 25132 3228
rect 25152 3208 25164 3228
rect 25120 3201 25164 3208
rect 25119 3170 25164 3201
rect 25214 3228 25256 3270
rect 25214 3208 25228 3228
rect 25248 3208 25256 3228
rect 25214 3170 25256 3208
rect 25330 3228 25372 3270
rect 25330 3208 25338 3228
rect 25358 3208 25372 3228
rect 25330 3170 25372 3208
rect 25422 3228 25466 3270
rect 25422 3208 25434 3228
rect 25454 3208 25466 3228
rect 25422 3170 25466 3208
rect 25548 3228 25590 3270
rect 25548 3208 25556 3228
rect 25576 3208 25590 3228
rect 25548 3170 25590 3208
rect 25640 3228 25684 3270
rect 27241 3242 27285 3284
rect 27335 3304 27377 3342
rect 27335 3284 27349 3304
rect 27369 3284 27377 3304
rect 27335 3242 27377 3284
rect 27459 3304 27503 3342
rect 27459 3284 27471 3304
rect 27491 3284 27503 3304
rect 27459 3242 27503 3284
rect 27553 3304 27595 3342
rect 27553 3284 27567 3304
rect 27587 3284 27595 3304
rect 27553 3242 27595 3284
rect 27669 3304 27711 3342
rect 27669 3284 27677 3304
rect 27697 3284 27711 3304
rect 27669 3242 27711 3284
rect 27761 3311 27806 3342
rect 27761 3304 27805 3311
rect 27761 3284 27773 3304
rect 27793 3284 27805 3304
rect 27761 3242 27805 3284
rect 33063 3437 33107 3479
rect 33063 3417 33075 3437
rect 33095 3417 33107 3437
rect 33063 3410 33107 3417
rect 33062 3379 33107 3410
rect 33157 3437 33199 3479
rect 33157 3417 33171 3437
rect 33191 3417 33199 3437
rect 33157 3379 33199 3417
rect 33273 3437 33315 3479
rect 33273 3417 33281 3437
rect 33301 3417 33315 3437
rect 33273 3379 33315 3417
rect 33365 3437 33409 3479
rect 33365 3417 33377 3437
rect 33397 3417 33409 3437
rect 33365 3379 33409 3417
rect 33491 3437 33533 3479
rect 33491 3417 33499 3437
rect 33519 3417 33533 3437
rect 33491 3379 33533 3417
rect 33583 3437 33627 3479
rect 33583 3417 33595 3437
rect 33615 3417 33627 3437
rect 33583 3379 33627 3417
rect 31605 3317 31649 3355
rect 31605 3297 31617 3317
rect 31637 3297 31649 3317
rect 25640 3208 25652 3228
rect 25672 3208 25684 3228
rect 25640 3170 25684 3208
rect 13957 3015 14001 3057
rect 15527 3017 15571 3059
rect 11683 2946 11727 2984
rect 15527 2997 15539 3017
rect 15559 2997 15571 3017
rect 15527 2990 15571 2997
rect 15526 2959 15571 2990
rect 15621 3017 15663 3059
rect 15621 2997 15635 3017
rect 15655 2997 15663 3017
rect 15621 2959 15663 2997
rect 15737 3017 15779 3059
rect 15737 2997 15745 3017
rect 15765 2997 15779 3017
rect 15737 2959 15779 2997
rect 15829 3017 15873 3059
rect 15829 2997 15841 3017
rect 15861 2997 15873 3017
rect 15829 2959 15873 2997
rect 15955 3017 15997 3059
rect 15955 2997 15963 3017
rect 15983 2997 15997 3017
rect 15955 2959 15997 2997
rect 16047 3017 16091 3059
rect 16047 2997 16059 3017
rect 16079 2997 16091 3017
rect 17703 3051 17747 3089
rect 17703 3031 17715 3051
rect 17735 3031 17747 3051
rect 16047 2959 16091 2997
rect 17703 2989 17747 3031
rect 17797 3051 17839 3089
rect 17797 3031 17811 3051
rect 17831 3031 17839 3051
rect 17797 2989 17839 3031
rect 17921 3051 17965 3089
rect 17921 3031 17933 3051
rect 17953 3031 17965 3051
rect 17921 2989 17965 3031
rect 18015 3051 18057 3089
rect 18015 3031 18029 3051
rect 18049 3031 18057 3051
rect 18015 2989 18057 3031
rect 18131 3051 18173 3089
rect 18131 3031 18139 3051
rect 18159 3031 18173 3051
rect 18131 2989 18173 3031
rect 18223 3058 18268 3089
rect 18223 3051 18267 3058
rect 18223 3031 18235 3051
rect 18255 3031 18267 3051
rect 29497 3240 29541 3282
rect 29497 3220 29509 3240
rect 29529 3220 29541 3240
rect 29497 3213 29541 3220
rect 29496 3182 29541 3213
rect 29591 3240 29633 3282
rect 29591 3220 29605 3240
rect 29625 3220 29633 3240
rect 29591 3182 29633 3220
rect 29707 3240 29749 3282
rect 29707 3220 29715 3240
rect 29735 3220 29749 3240
rect 29707 3182 29749 3220
rect 29799 3240 29843 3282
rect 29799 3220 29811 3240
rect 29831 3220 29843 3240
rect 29799 3182 29843 3220
rect 29925 3240 29967 3282
rect 29925 3220 29933 3240
rect 29953 3220 29967 3240
rect 29925 3182 29967 3220
rect 30017 3240 30061 3282
rect 31605 3255 31649 3297
rect 31699 3317 31741 3355
rect 31699 3297 31713 3317
rect 31733 3297 31741 3317
rect 31699 3255 31741 3297
rect 31823 3317 31867 3355
rect 31823 3297 31835 3317
rect 31855 3297 31867 3317
rect 31823 3255 31867 3297
rect 31917 3317 31959 3355
rect 31917 3297 31931 3317
rect 31951 3297 31959 3317
rect 31917 3255 31959 3297
rect 32033 3317 32075 3355
rect 32033 3297 32041 3317
rect 32061 3297 32075 3317
rect 32033 3255 32075 3297
rect 32125 3324 32170 3355
rect 32125 3317 32169 3324
rect 32125 3297 32137 3317
rect 32157 3297 32169 3317
rect 32125 3255 32169 3297
rect 30017 3220 30029 3240
rect 30049 3220 30061 3240
rect 30017 3182 30061 3220
rect 22067 3064 22111 3102
rect 18223 2989 18267 3031
rect 19793 2991 19837 3033
rect 19793 2971 19805 2991
rect 19825 2971 19837 2991
rect 19793 2964 19837 2971
rect 19792 2933 19837 2964
rect 19887 2991 19929 3033
rect 19887 2971 19901 2991
rect 19921 2971 19929 2991
rect 19887 2933 19929 2971
rect 20003 2991 20045 3033
rect 20003 2971 20011 2991
rect 20031 2971 20045 2991
rect 20003 2933 20045 2971
rect 20095 2991 20139 3033
rect 20095 2971 20107 2991
rect 20127 2971 20139 2991
rect 20095 2933 20139 2971
rect 20221 2991 20263 3033
rect 20221 2971 20229 2991
rect 20249 2971 20263 2991
rect 20221 2933 20263 2971
rect 20313 2991 20357 3033
rect 22067 3044 22079 3064
rect 22099 3044 22111 3064
rect 20313 2971 20325 2991
rect 20345 2971 20357 2991
rect 22067 3002 22111 3044
rect 22161 3064 22203 3102
rect 22161 3044 22175 3064
rect 22195 3044 22203 3064
rect 22161 3002 22203 3044
rect 22285 3064 22329 3102
rect 22285 3044 22297 3064
rect 22317 3044 22329 3064
rect 22285 3002 22329 3044
rect 22379 3064 22421 3102
rect 22379 3044 22393 3064
rect 22413 3044 22421 3064
rect 22379 3002 22421 3044
rect 22495 3064 22537 3102
rect 22495 3044 22503 3064
rect 22523 3044 22537 3064
rect 22495 3002 22537 3044
rect 22587 3071 22632 3102
rect 22587 3064 22631 3071
rect 22587 3044 22599 3064
rect 22619 3044 22631 3064
rect 33861 3253 33905 3295
rect 33861 3233 33873 3253
rect 33893 3233 33905 3253
rect 33861 3226 33905 3233
rect 33860 3195 33905 3226
rect 33955 3253 33997 3295
rect 33955 3233 33969 3253
rect 33989 3233 33997 3253
rect 33955 3195 33997 3233
rect 34071 3253 34113 3295
rect 34071 3233 34079 3253
rect 34099 3233 34113 3253
rect 34071 3195 34113 3233
rect 34163 3253 34207 3295
rect 34163 3233 34175 3253
rect 34195 3233 34207 3253
rect 34163 3195 34207 3233
rect 34289 3253 34331 3295
rect 34289 3233 34297 3253
rect 34317 3233 34331 3253
rect 34289 3195 34331 3233
rect 34381 3253 34425 3295
rect 34381 3233 34393 3253
rect 34413 3233 34425 3253
rect 34381 3195 34425 3233
rect 26444 3076 26488 3114
rect 22587 3002 22631 3044
rect 24157 3004 24201 3046
rect 20313 2933 20357 2971
rect 24157 2984 24169 3004
rect 24189 2984 24201 3004
rect 24157 2977 24201 2984
rect 24156 2946 24201 2977
rect 24251 3004 24293 3046
rect 24251 2984 24265 3004
rect 24285 2984 24293 3004
rect 24251 2946 24293 2984
rect 24367 3004 24409 3046
rect 24367 2984 24375 3004
rect 24395 2984 24409 3004
rect 24367 2946 24409 2984
rect 24459 3004 24503 3046
rect 24459 2984 24471 3004
rect 24491 2984 24503 3004
rect 24459 2946 24503 2984
rect 24585 3004 24627 3046
rect 24585 2984 24593 3004
rect 24613 2984 24627 3004
rect 24585 2946 24627 2984
rect 24677 3004 24721 3046
rect 26444 3056 26456 3076
rect 26476 3056 26488 3076
rect 24677 2984 24689 3004
rect 24709 2984 24721 3004
rect 26444 3014 26488 3056
rect 26538 3076 26580 3114
rect 26538 3056 26552 3076
rect 26572 3056 26580 3076
rect 26538 3014 26580 3056
rect 26662 3076 26706 3114
rect 26662 3056 26674 3076
rect 26694 3056 26706 3076
rect 26662 3014 26706 3056
rect 26756 3076 26798 3114
rect 26756 3056 26770 3076
rect 26790 3056 26798 3076
rect 26756 3014 26798 3056
rect 26872 3076 26914 3114
rect 26872 3056 26880 3076
rect 26900 3056 26914 3076
rect 26872 3014 26914 3056
rect 26964 3083 27009 3114
rect 26964 3076 27008 3083
rect 26964 3056 26976 3076
rect 26996 3056 27008 3076
rect 30808 3089 30852 3127
rect 26964 3014 27008 3056
rect 28534 3016 28578 3058
rect 24677 2946 24721 2984
rect 28534 2996 28546 3016
rect 28566 2996 28578 3016
rect 28534 2989 28578 2996
rect 28533 2958 28578 2989
rect 28628 3016 28670 3058
rect 28628 2996 28642 3016
rect 28662 2996 28670 3016
rect 28628 2958 28670 2996
rect 28744 3016 28786 3058
rect 28744 2996 28752 3016
rect 28772 2996 28786 3016
rect 28744 2958 28786 2996
rect 28836 3016 28880 3058
rect 28836 2996 28848 3016
rect 28868 2996 28880 3016
rect 28836 2958 28880 2996
rect 28962 3016 29004 3058
rect 28962 2996 28970 3016
rect 28990 2996 29004 3016
rect 28962 2958 29004 2996
rect 29054 3016 29098 3058
rect 30808 3069 30820 3089
rect 30840 3069 30852 3089
rect 29054 2996 29066 3016
rect 29086 2996 29098 3016
rect 30808 3027 30852 3069
rect 30902 3089 30944 3127
rect 30902 3069 30916 3089
rect 30936 3069 30944 3089
rect 30902 3027 30944 3069
rect 31026 3089 31070 3127
rect 31026 3069 31038 3089
rect 31058 3069 31070 3089
rect 31026 3027 31070 3069
rect 31120 3089 31162 3127
rect 31120 3069 31134 3089
rect 31154 3069 31162 3089
rect 31120 3027 31162 3069
rect 31236 3089 31278 3127
rect 31236 3069 31244 3089
rect 31264 3069 31278 3089
rect 31236 3027 31278 3069
rect 31328 3096 31373 3127
rect 31328 3089 31372 3096
rect 31328 3069 31340 3089
rect 31360 3069 31372 3089
rect 31328 3027 31372 3069
rect 32898 3029 32942 3071
rect 29054 2958 29098 2996
rect 32898 3009 32910 3029
rect 32930 3009 32942 3029
rect 32898 3002 32942 3009
rect 32897 2971 32942 3002
rect 32992 3029 33034 3071
rect 32992 3009 33006 3029
rect 33026 3009 33034 3029
rect 32992 2971 33034 3009
rect 33108 3029 33150 3071
rect 33108 3009 33116 3029
rect 33136 3009 33150 3029
rect 33108 2971 33150 3009
rect 33200 3029 33244 3071
rect 33200 3009 33212 3029
rect 33232 3009 33244 3029
rect 33200 2971 33244 3009
rect 33326 3029 33368 3071
rect 33326 3009 33334 3029
rect 33354 3009 33368 3029
rect 33326 2971 33368 3009
rect 33418 3029 33462 3071
rect 33418 3009 33430 3029
rect 33450 3009 33462 3029
rect 33418 2971 33462 3009
rect 1274 2657 1318 2695
rect 1274 2637 1286 2657
rect 1306 2637 1318 2657
rect 1274 2595 1318 2637
rect 1368 2657 1410 2695
rect 1368 2637 1382 2657
rect 1402 2637 1410 2657
rect 1368 2595 1410 2637
rect 1492 2657 1536 2695
rect 1492 2637 1504 2657
rect 1524 2637 1536 2657
rect 1492 2595 1536 2637
rect 1586 2657 1628 2695
rect 1586 2637 1600 2657
rect 1620 2637 1628 2657
rect 1586 2595 1628 2637
rect 1702 2657 1744 2695
rect 1702 2637 1710 2657
rect 1730 2637 1744 2657
rect 1702 2595 1744 2637
rect 1794 2664 1839 2695
rect 1794 2657 1838 2664
rect 1794 2637 1806 2657
rect 1826 2637 1838 2657
rect 5638 2670 5682 2708
rect 1794 2595 1838 2637
rect 3364 2597 3408 2639
rect 3364 2577 3376 2597
rect 3396 2577 3408 2597
rect 3364 2570 3408 2577
rect 3363 2539 3408 2570
rect 3458 2597 3500 2639
rect 3458 2577 3472 2597
rect 3492 2577 3500 2597
rect 3458 2539 3500 2577
rect 3574 2597 3616 2639
rect 3574 2577 3582 2597
rect 3602 2577 3616 2597
rect 3574 2539 3616 2577
rect 3666 2597 3710 2639
rect 3666 2577 3678 2597
rect 3698 2577 3710 2597
rect 3666 2539 3710 2577
rect 3792 2597 3834 2639
rect 3792 2577 3800 2597
rect 3820 2577 3834 2597
rect 3792 2539 3834 2577
rect 3884 2597 3928 2639
rect 5638 2650 5650 2670
rect 5670 2650 5682 2670
rect 3884 2577 3896 2597
rect 3916 2577 3928 2597
rect 5638 2608 5682 2650
rect 5732 2670 5774 2708
rect 5732 2650 5746 2670
rect 5766 2650 5774 2670
rect 5732 2608 5774 2650
rect 5856 2670 5900 2708
rect 5856 2650 5868 2670
rect 5888 2650 5900 2670
rect 5856 2608 5900 2650
rect 5950 2670 5992 2708
rect 5950 2650 5964 2670
rect 5984 2650 5992 2670
rect 5950 2608 5992 2650
rect 6066 2670 6108 2708
rect 6066 2650 6074 2670
rect 6094 2650 6108 2670
rect 6066 2608 6108 2650
rect 6158 2677 6203 2708
rect 6158 2670 6202 2677
rect 6158 2650 6170 2670
rect 6190 2650 6202 2670
rect 10015 2682 10059 2720
rect 6158 2608 6202 2650
rect 7728 2610 7772 2652
rect 3884 2539 3928 2577
rect 7728 2590 7740 2610
rect 7760 2590 7772 2610
rect 7728 2583 7772 2590
rect 7727 2552 7772 2583
rect 7822 2610 7864 2652
rect 7822 2590 7836 2610
rect 7856 2590 7864 2610
rect 7822 2552 7864 2590
rect 7938 2610 7980 2652
rect 7938 2590 7946 2610
rect 7966 2590 7980 2610
rect 7938 2552 7980 2590
rect 8030 2610 8074 2652
rect 8030 2590 8042 2610
rect 8062 2590 8074 2610
rect 8030 2552 8074 2590
rect 8156 2610 8198 2652
rect 8156 2590 8164 2610
rect 8184 2590 8198 2610
rect 8156 2552 8198 2590
rect 8248 2610 8292 2652
rect 10015 2662 10027 2682
rect 10047 2662 10059 2682
rect 8248 2590 8260 2610
rect 8280 2590 8292 2610
rect 10015 2620 10059 2662
rect 10109 2682 10151 2720
rect 10109 2662 10123 2682
rect 10143 2662 10151 2682
rect 10109 2620 10151 2662
rect 10233 2682 10277 2720
rect 10233 2662 10245 2682
rect 10265 2662 10277 2682
rect 10233 2620 10277 2662
rect 10327 2682 10369 2720
rect 10327 2662 10341 2682
rect 10361 2662 10369 2682
rect 10327 2620 10369 2662
rect 10443 2682 10485 2720
rect 10443 2662 10451 2682
rect 10471 2662 10485 2682
rect 10443 2620 10485 2662
rect 10535 2689 10580 2720
rect 10535 2682 10579 2689
rect 10535 2662 10547 2682
rect 10567 2662 10579 2682
rect 14379 2695 14423 2733
rect 10535 2620 10579 2662
rect 12105 2622 12149 2664
rect 8248 2552 8292 2590
rect 311 2433 355 2471
rect 311 2413 323 2433
rect 343 2413 355 2433
rect 311 2371 355 2413
rect 405 2433 447 2471
rect 405 2413 419 2433
rect 439 2413 447 2433
rect 405 2371 447 2413
rect 529 2433 573 2471
rect 529 2413 541 2433
rect 561 2413 573 2433
rect 529 2371 573 2413
rect 623 2433 665 2471
rect 623 2413 637 2433
rect 657 2413 665 2433
rect 623 2371 665 2413
rect 739 2433 781 2471
rect 739 2413 747 2433
rect 767 2413 781 2433
rect 739 2371 781 2413
rect 831 2440 876 2471
rect 831 2433 875 2440
rect 831 2413 843 2433
rect 863 2413 875 2433
rect 831 2371 875 2413
rect 12105 2602 12117 2622
rect 12137 2602 12149 2622
rect 12105 2595 12149 2602
rect 12104 2564 12149 2595
rect 12199 2622 12241 2664
rect 12199 2602 12213 2622
rect 12233 2602 12241 2622
rect 12199 2564 12241 2602
rect 12315 2622 12357 2664
rect 12315 2602 12323 2622
rect 12343 2602 12357 2622
rect 12315 2564 12357 2602
rect 12407 2622 12451 2664
rect 12407 2602 12419 2622
rect 12439 2602 12451 2622
rect 12407 2564 12451 2602
rect 12533 2622 12575 2664
rect 12533 2602 12541 2622
rect 12561 2602 12575 2622
rect 12533 2564 12575 2602
rect 12625 2622 12669 2664
rect 14379 2675 14391 2695
rect 14411 2675 14423 2695
rect 12625 2602 12637 2622
rect 12657 2602 12669 2622
rect 14379 2633 14423 2675
rect 14473 2695 14515 2733
rect 14473 2675 14487 2695
rect 14507 2675 14515 2695
rect 14473 2633 14515 2675
rect 14597 2695 14641 2733
rect 14597 2675 14609 2695
rect 14629 2675 14641 2695
rect 14597 2633 14641 2675
rect 14691 2695 14733 2733
rect 14691 2675 14705 2695
rect 14725 2675 14733 2695
rect 14691 2633 14733 2675
rect 14807 2695 14849 2733
rect 14807 2675 14815 2695
rect 14835 2675 14849 2695
rect 14807 2633 14849 2675
rect 14899 2702 14944 2733
rect 14899 2695 14943 2702
rect 14899 2675 14911 2695
rect 14931 2675 14943 2695
rect 14899 2633 14943 2675
rect 16469 2635 16513 2677
rect 12625 2564 12669 2602
rect 4675 2446 4719 2484
rect 4675 2426 4687 2446
rect 4707 2426 4719 2446
rect 2567 2369 2611 2411
rect 2567 2349 2579 2369
rect 2599 2349 2611 2369
rect 2567 2342 2611 2349
rect 2566 2311 2611 2342
rect 2661 2369 2703 2411
rect 2661 2349 2675 2369
rect 2695 2349 2703 2369
rect 2661 2311 2703 2349
rect 2777 2369 2819 2411
rect 2777 2349 2785 2369
rect 2805 2349 2819 2369
rect 2777 2311 2819 2349
rect 2869 2369 2913 2411
rect 2869 2349 2881 2369
rect 2901 2349 2913 2369
rect 2869 2311 2913 2349
rect 2995 2369 3037 2411
rect 2995 2349 3003 2369
rect 3023 2349 3037 2369
rect 2995 2311 3037 2349
rect 3087 2369 3131 2411
rect 4675 2384 4719 2426
rect 4769 2446 4811 2484
rect 4769 2426 4783 2446
rect 4803 2426 4811 2446
rect 4769 2384 4811 2426
rect 4893 2446 4937 2484
rect 4893 2426 4905 2446
rect 4925 2426 4937 2446
rect 4893 2384 4937 2426
rect 4987 2446 5029 2484
rect 4987 2426 5001 2446
rect 5021 2426 5029 2446
rect 4987 2384 5029 2426
rect 5103 2446 5145 2484
rect 5103 2426 5111 2446
rect 5131 2426 5145 2446
rect 5103 2384 5145 2426
rect 5195 2453 5240 2484
rect 5195 2446 5239 2453
rect 5195 2426 5207 2446
rect 5227 2426 5239 2446
rect 5195 2384 5239 2426
rect 16469 2615 16481 2635
rect 16501 2615 16513 2635
rect 16469 2608 16513 2615
rect 16468 2577 16513 2608
rect 16563 2635 16605 2677
rect 16563 2615 16577 2635
rect 16597 2615 16605 2635
rect 16563 2577 16605 2615
rect 16679 2635 16721 2677
rect 16679 2615 16687 2635
rect 16707 2615 16721 2635
rect 16679 2577 16721 2615
rect 16771 2635 16815 2677
rect 16771 2615 16783 2635
rect 16803 2615 16815 2635
rect 16771 2577 16815 2615
rect 16897 2635 16939 2677
rect 16897 2615 16905 2635
rect 16925 2615 16939 2635
rect 16897 2577 16939 2615
rect 16989 2635 17033 2677
rect 18645 2669 18689 2707
rect 16989 2615 17001 2635
rect 17021 2615 17033 2635
rect 16989 2577 17033 2615
rect 18645 2649 18657 2669
rect 18677 2649 18689 2669
rect 18645 2607 18689 2649
rect 18739 2669 18781 2707
rect 18739 2649 18753 2669
rect 18773 2649 18781 2669
rect 18739 2607 18781 2649
rect 18863 2669 18907 2707
rect 18863 2649 18875 2669
rect 18895 2649 18907 2669
rect 18863 2607 18907 2649
rect 18957 2669 18999 2707
rect 18957 2649 18971 2669
rect 18991 2649 18999 2669
rect 18957 2607 18999 2649
rect 19073 2669 19115 2707
rect 19073 2649 19081 2669
rect 19101 2649 19115 2669
rect 19073 2607 19115 2649
rect 19165 2676 19210 2707
rect 19165 2669 19209 2676
rect 19165 2649 19177 2669
rect 19197 2649 19209 2669
rect 23009 2682 23053 2720
rect 19165 2607 19209 2649
rect 20735 2609 20779 2651
rect 9052 2458 9096 2496
rect 9052 2438 9064 2458
rect 9084 2438 9096 2458
rect 3087 2349 3099 2369
rect 3119 2349 3131 2369
rect 3087 2311 3131 2349
rect 1109 2249 1153 2287
rect 1109 2229 1121 2249
rect 1141 2229 1153 2249
rect 1109 2187 1153 2229
rect 1203 2249 1245 2287
rect 1203 2229 1217 2249
rect 1237 2229 1245 2249
rect 1203 2187 1245 2229
rect 1327 2249 1371 2287
rect 1327 2229 1339 2249
rect 1359 2229 1371 2249
rect 1327 2187 1371 2229
rect 1421 2249 1463 2287
rect 1421 2229 1435 2249
rect 1455 2229 1463 2249
rect 1421 2187 1463 2229
rect 1537 2249 1579 2287
rect 1537 2229 1545 2249
rect 1565 2229 1579 2249
rect 1537 2187 1579 2229
rect 1629 2256 1674 2287
rect 1629 2249 1673 2256
rect 1629 2229 1641 2249
rect 1661 2229 1673 2249
rect 1629 2187 1673 2229
rect 6931 2382 6975 2424
rect 6931 2362 6943 2382
rect 6963 2362 6975 2382
rect 6931 2355 6975 2362
rect 6930 2324 6975 2355
rect 7025 2382 7067 2424
rect 7025 2362 7039 2382
rect 7059 2362 7067 2382
rect 7025 2324 7067 2362
rect 7141 2382 7183 2424
rect 7141 2362 7149 2382
rect 7169 2362 7183 2382
rect 7141 2324 7183 2362
rect 7233 2382 7277 2424
rect 7233 2362 7245 2382
rect 7265 2362 7277 2382
rect 7233 2324 7277 2362
rect 7359 2382 7401 2424
rect 7359 2362 7367 2382
rect 7387 2362 7401 2382
rect 7359 2324 7401 2362
rect 7451 2382 7495 2424
rect 9052 2396 9096 2438
rect 9146 2458 9188 2496
rect 9146 2438 9160 2458
rect 9180 2438 9188 2458
rect 9146 2396 9188 2438
rect 9270 2458 9314 2496
rect 9270 2438 9282 2458
rect 9302 2438 9314 2458
rect 9270 2396 9314 2438
rect 9364 2458 9406 2496
rect 9364 2438 9378 2458
rect 9398 2438 9406 2458
rect 9364 2396 9406 2438
rect 9480 2458 9522 2496
rect 9480 2438 9488 2458
rect 9508 2438 9522 2458
rect 9480 2396 9522 2438
rect 9572 2465 9617 2496
rect 9572 2458 9616 2465
rect 9572 2438 9584 2458
rect 9604 2438 9616 2458
rect 9572 2396 9616 2438
rect 20735 2589 20747 2609
rect 20767 2589 20779 2609
rect 20735 2582 20779 2589
rect 20734 2551 20779 2582
rect 20829 2609 20871 2651
rect 20829 2589 20843 2609
rect 20863 2589 20871 2609
rect 20829 2551 20871 2589
rect 20945 2609 20987 2651
rect 20945 2589 20953 2609
rect 20973 2589 20987 2609
rect 20945 2551 20987 2589
rect 21037 2609 21081 2651
rect 21037 2589 21049 2609
rect 21069 2589 21081 2609
rect 21037 2551 21081 2589
rect 21163 2609 21205 2651
rect 21163 2589 21171 2609
rect 21191 2589 21205 2609
rect 21163 2551 21205 2589
rect 21255 2609 21299 2651
rect 23009 2662 23021 2682
rect 23041 2662 23053 2682
rect 21255 2589 21267 2609
rect 21287 2589 21299 2609
rect 23009 2620 23053 2662
rect 23103 2682 23145 2720
rect 23103 2662 23117 2682
rect 23137 2662 23145 2682
rect 23103 2620 23145 2662
rect 23227 2682 23271 2720
rect 23227 2662 23239 2682
rect 23259 2662 23271 2682
rect 23227 2620 23271 2662
rect 23321 2682 23363 2720
rect 23321 2662 23335 2682
rect 23355 2662 23363 2682
rect 23321 2620 23363 2662
rect 23437 2682 23479 2720
rect 23437 2662 23445 2682
rect 23465 2662 23479 2682
rect 23437 2620 23479 2662
rect 23529 2689 23574 2720
rect 23529 2682 23573 2689
rect 23529 2662 23541 2682
rect 23561 2662 23573 2682
rect 27386 2694 27430 2732
rect 23529 2620 23573 2662
rect 25099 2622 25143 2664
rect 21255 2551 21299 2589
rect 13416 2471 13460 2509
rect 13416 2451 13428 2471
rect 13448 2451 13460 2471
rect 7451 2362 7463 2382
rect 7483 2362 7495 2382
rect 7451 2324 7495 2362
rect 5473 2262 5517 2300
rect 5473 2242 5485 2262
rect 5505 2242 5517 2262
rect 3365 2185 3409 2227
rect 3365 2165 3377 2185
rect 3397 2165 3409 2185
rect 3365 2158 3409 2165
rect 3364 2127 3409 2158
rect 3459 2185 3501 2227
rect 3459 2165 3473 2185
rect 3493 2165 3501 2185
rect 3459 2127 3501 2165
rect 3575 2185 3617 2227
rect 3575 2165 3583 2185
rect 3603 2165 3617 2185
rect 3575 2127 3617 2165
rect 3667 2185 3711 2227
rect 3667 2165 3679 2185
rect 3699 2165 3711 2185
rect 3667 2127 3711 2165
rect 3793 2185 3835 2227
rect 3793 2165 3801 2185
rect 3821 2165 3835 2185
rect 3793 2127 3835 2165
rect 3885 2185 3929 2227
rect 5473 2200 5517 2242
rect 5567 2262 5609 2300
rect 5567 2242 5581 2262
rect 5601 2242 5609 2262
rect 5567 2200 5609 2242
rect 5691 2262 5735 2300
rect 5691 2242 5703 2262
rect 5723 2242 5735 2262
rect 5691 2200 5735 2242
rect 5785 2262 5827 2300
rect 5785 2242 5799 2262
rect 5819 2242 5827 2262
rect 5785 2200 5827 2242
rect 5901 2262 5943 2300
rect 5901 2242 5909 2262
rect 5929 2242 5943 2262
rect 5901 2200 5943 2242
rect 5993 2269 6038 2300
rect 5993 2262 6037 2269
rect 5993 2242 6005 2262
rect 6025 2242 6037 2262
rect 5993 2200 6037 2242
rect 11308 2394 11352 2436
rect 11308 2374 11320 2394
rect 11340 2374 11352 2394
rect 11308 2367 11352 2374
rect 11307 2336 11352 2367
rect 11402 2394 11444 2436
rect 11402 2374 11416 2394
rect 11436 2374 11444 2394
rect 11402 2336 11444 2374
rect 11518 2394 11560 2436
rect 11518 2374 11526 2394
rect 11546 2374 11560 2394
rect 11518 2336 11560 2374
rect 11610 2394 11654 2436
rect 11610 2374 11622 2394
rect 11642 2374 11654 2394
rect 11610 2336 11654 2374
rect 11736 2394 11778 2436
rect 11736 2374 11744 2394
rect 11764 2374 11778 2394
rect 11736 2336 11778 2374
rect 11828 2394 11872 2436
rect 13416 2409 13460 2451
rect 13510 2471 13552 2509
rect 13510 2451 13524 2471
rect 13544 2451 13552 2471
rect 13510 2409 13552 2451
rect 13634 2471 13678 2509
rect 13634 2451 13646 2471
rect 13666 2451 13678 2471
rect 13634 2409 13678 2451
rect 13728 2471 13770 2509
rect 13728 2451 13742 2471
rect 13762 2451 13770 2471
rect 13728 2409 13770 2451
rect 13844 2471 13886 2509
rect 13844 2451 13852 2471
rect 13872 2451 13886 2471
rect 13844 2409 13886 2451
rect 13936 2478 13981 2509
rect 13936 2471 13980 2478
rect 13936 2451 13948 2471
rect 13968 2451 13980 2471
rect 13936 2409 13980 2451
rect 25099 2602 25111 2622
rect 25131 2602 25143 2622
rect 25099 2595 25143 2602
rect 25098 2564 25143 2595
rect 25193 2622 25235 2664
rect 25193 2602 25207 2622
rect 25227 2602 25235 2622
rect 25193 2564 25235 2602
rect 25309 2622 25351 2664
rect 25309 2602 25317 2622
rect 25337 2602 25351 2622
rect 25309 2564 25351 2602
rect 25401 2622 25445 2664
rect 25401 2602 25413 2622
rect 25433 2602 25445 2622
rect 25401 2564 25445 2602
rect 25527 2622 25569 2664
rect 25527 2602 25535 2622
rect 25555 2602 25569 2622
rect 25527 2564 25569 2602
rect 25619 2622 25663 2664
rect 27386 2674 27398 2694
rect 27418 2674 27430 2694
rect 25619 2602 25631 2622
rect 25651 2602 25663 2622
rect 27386 2632 27430 2674
rect 27480 2694 27522 2732
rect 27480 2674 27494 2694
rect 27514 2674 27522 2694
rect 27480 2632 27522 2674
rect 27604 2694 27648 2732
rect 27604 2674 27616 2694
rect 27636 2674 27648 2694
rect 27604 2632 27648 2674
rect 27698 2694 27740 2732
rect 27698 2674 27712 2694
rect 27732 2674 27740 2694
rect 27698 2632 27740 2674
rect 27814 2694 27856 2732
rect 27814 2674 27822 2694
rect 27842 2674 27856 2694
rect 27814 2632 27856 2674
rect 27906 2701 27951 2732
rect 27906 2694 27950 2701
rect 27906 2674 27918 2694
rect 27938 2674 27950 2694
rect 31750 2707 31794 2745
rect 27906 2632 27950 2674
rect 29476 2634 29520 2676
rect 25619 2564 25663 2602
rect 11828 2374 11840 2394
rect 11860 2374 11872 2394
rect 11828 2336 11872 2374
rect 9850 2274 9894 2312
rect 9850 2254 9862 2274
rect 9882 2254 9894 2274
rect 3885 2165 3897 2185
rect 3917 2165 3929 2185
rect 3885 2127 3929 2165
rect 7729 2198 7773 2240
rect 7729 2178 7741 2198
rect 7761 2178 7773 2198
rect 7729 2171 7773 2178
rect 7728 2140 7773 2171
rect 7823 2198 7865 2240
rect 7823 2178 7837 2198
rect 7857 2178 7865 2198
rect 7823 2140 7865 2178
rect 7939 2198 7981 2240
rect 7939 2178 7947 2198
rect 7967 2178 7981 2198
rect 7939 2140 7981 2178
rect 8031 2198 8075 2240
rect 8031 2178 8043 2198
rect 8063 2178 8075 2198
rect 8031 2140 8075 2178
rect 8157 2198 8199 2240
rect 8157 2178 8165 2198
rect 8185 2178 8199 2198
rect 8157 2140 8199 2178
rect 8249 2198 8293 2240
rect 9850 2212 9894 2254
rect 9944 2274 9986 2312
rect 9944 2254 9958 2274
rect 9978 2254 9986 2274
rect 9944 2212 9986 2254
rect 10068 2274 10112 2312
rect 10068 2254 10080 2274
rect 10100 2254 10112 2274
rect 10068 2212 10112 2254
rect 10162 2274 10204 2312
rect 10162 2254 10176 2274
rect 10196 2254 10204 2274
rect 10162 2212 10204 2254
rect 10278 2274 10320 2312
rect 10278 2254 10286 2274
rect 10306 2254 10320 2274
rect 10278 2212 10320 2254
rect 10370 2281 10415 2312
rect 10370 2274 10414 2281
rect 10370 2254 10382 2274
rect 10402 2254 10414 2274
rect 10370 2212 10414 2254
rect 15672 2407 15716 2449
rect 15672 2387 15684 2407
rect 15704 2387 15716 2407
rect 15672 2380 15716 2387
rect 15671 2349 15716 2380
rect 15766 2407 15808 2449
rect 15766 2387 15780 2407
rect 15800 2387 15808 2407
rect 15766 2349 15808 2387
rect 15882 2407 15924 2449
rect 15882 2387 15890 2407
rect 15910 2387 15924 2407
rect 15882 2349 15924 2387
rect 15974 2407 16018 2449
rect 15974 2387 15986 2407
rect 16006 2387 16018 2407
rect 15974 2349 16018 2387
rect 16100 2407 16142 2449
rect 16100 2387 16108 2407
rect 16128 2387 16142 2407
rect 16100 2349 16142 2387
rect 16192 2407 16236 2449
rect 17682 2445 17726 2483
rect 17682 2425 17694 2445
rect 17714 2425 17726 2445
rect 16192 2387 16204 2407
rect 16224 2387 16236 2407
rect 16192 2349 16236 2387
rect 17682 2383 17726 2425
rect 17776 2445 17818 2483
rect 17776 2425 17790 2445
rect 17810 2425 17818 2445
rect 17776 2383 17818 2425
rect 17900 2445 17944 2483
rect 17900 2425 17912 2445
rect 17932 2425 17944 2445
rect 17900 2383 17944 2425
rect 17994 2445 18036 2483
rect 17994 2425 18008 2445
rect 18028 2425 18036 2445
rect 17994 2383 18036 2425
rect 18110 2445 18152 2483
rect 18110 2425 18118 2445
rect 18138 2425 18152 2445
rect 18110 2383 18152 2425
rect 18202 2452 18247 2483
rect 18202 2445 18246 2452
rect 18202 2425 18214 2445
rect 18234 2425 18246 2445
rect 18202 2383 18246 2425
rect 29476 2614 29488 2634
rect 29508 2614 29520 2634
rect 29476 2607 29520 2614
rect 29475 2576 29520 2607
rect 29570 2634 29612 2676
rect 29570 2614 29584 2634
rect 29604 2614 29612 2634
rect 29570 2576 29612 2614
rect 29686 2634 29728 2676
rect 29686 2614 29694 2634
rect 29714 2614 29728 2634
rect 29686 2576 29728 2614
rect 29778 2634 29822 2676
rect 29778 2614 29790 2634
rect 29810 2614 29822 2634
rect 29778 2576 29822 2614
rect 29904 2634 29946 2676
rect 29904 2614 29912 2634
rect 29932 2614 29946 2634
rect 29904 2576 29946 2614
rect 29996 2634 30040 2676
rect 31750 2687 31762 2707
rect 31782 2687 31794 2707
rect 29996 2614 30008 2634
rect 30028 2614 30040 2634
rect 31750 2645 31794 2687
rect 31844 2707 31886 2745
rect 31844 2687 31858 2707
rect 31878 2687 31886 2707
rect 31844 2645 31886 2687
rect 31968 2707 32012 2745
rect 31968 2687 31980 2707
rect 32000 2687 32012 2707
rect 31968 2645 32012 2687
rect 32062 2707 32104 2745
rect 32062 2687 32076 2707
rect 32096 2687 32104 2707
rect 32062 2645 32104 2687
rect 32178 2707 32220 2745
rect 32178 2687 32186 2707
rect 32206 2687 32220 2707
rect 32178 2645 32220 2687
rect 32270 2714 32315 2745
rect 32270 2707 32314 2714
rect 32270 2687 32282 2707
rect 32302 2687 32314 2707
rect 32270 2645 32314 2687
rect 33840 2647 33884 2689
rect 29996 2576 30040 2614
rect 22046 2458 22090 2496
rect 22046 2438 22058 2458
rect 22078 2438 22090 2458
rect 14214 2287 14258 2325
rect 14214 2267 14226 2287
rect 14246 2267 14258 2287
rect 8249 2178 8261 2198
rect 8281 2178 8293 2198
rect 8249 2140 8293 2178
rect 312 2021 356 2059
rect 312 2001 324 2021
rect 344 2001 356 2021
rect 312 1959 356 2001
rect 406 2021 448 2059
rect 406 2001 420 2021
rect 440 2001 448 2021
rect 406 1959 448 2001
rect 530 2021 574 2059
rect 530 2001 542 2021
rect 562 2001 574 2021
rect 530 1959 574 2001
rect 624 2021 666 2059
rect 624 2001 638 2021
rect 658 2001 666 2021
rect 624 1959 666 2001
rect 740 2021 782 2059
rect 740 2001 748 2021
rect 768 2001 782 2021
rect 740 1959 782 2001
rect 832 2028 877 2059
rect 832 2021 876 2028
rect 832 2001 844 2021
rect 864 2001 876 2021
rect 12106 2210 12150 2252
rect 12106 2190 12118 2210
rect 12138 2190 12150 2210
rect 12106 2183 12150 2190
rect 12105 2152 12150 2183
rect 12200 2210 12242 2252
rect 12200 2190 12214 2210
rect 12234 2190 12242 2210
rect 12200 2152 12242 2190
rect 12316 2210 12358 2252
rect 12316 2190 12324 2210
rect 12344 2190 12358 2210
rect 12316 2152 12358 2190
rect 12408 2210 12452 2252
rect 12408 2190 12420 2210
rect 12440 2190 12452 2210
rect 12408 2152 12452 2190
rect 12534 2210 12576 2252
rect 12534 2190 12542 2210
rect 12562 2190 12576 2210
rect 12534 2152 12576 2190
rect 12626 2210 12670 2252
rect 14214 2225 14258 2267
rect 14308 2287 14350 2325
rect 14308 2267 14322 2287
rect 14342 2267 14350 2287
rect 14308 2225 14350 2267
rect 14432 2287 14476 2325
rect 14432 2267 14444 2287
rect 14464 2267 14476 2287
rect 14432 2225 14476 2267
rect 14526 2287 14568 2325
rect 14526 2267 14540 2287
rect 14560 2267 14568 2287
rect 14526 2225 14568 2267
rect 14642 2287 14684 2325
rect 14642 2267 14650 2287
rect 14670 2267 14684 2287
rect 14642 2225 14684 2267
rect 14734 2294 14779 2325
rect 14734 2287 14778 2294
rect 14734 2267 14746 2287
rect 14766 2267 14778 2287
rect 14734 2225 14778 2267
rect 19938 2381 19982 2423
rect 19938 2361 19950 2381
rect 19970 2361 19982 2381
rect 19938 2354 19982 2361
rect 19937 2323 19982 2354
rect 20032 2381 20074 2423
rect 20032 2361 20046 2381
rect 20066 2361 20074 2381
rect 20032 2323 20074 2361
rect 20148 2381 20190 2423
rect 20148 2361 20156 2381
rect 20176 2361 20190 2381
rect 20148 2323 20190 2361
rect 20240 2381 20284 2423
rect 20240 2361 20252 2381
rect 20272 2361 20284 2381
rect 20240 2323 20284 2361
rect 20366 2381 20408 2423
rect 20366 2361 20374 2381
rect 20394 2361 20408 2381
rect 20366 2323 20408 2361
rect 20458 2381 20502 2423
rect 22046 2396 22090 2438
rect 22140 2458 22182 2496
rect 22140 2438 22154 2458
rect 22174 2438 22182 2458
rect 22140 2396 22182 2438
rect 22264 2458 22308 2496
rect 22264 2438 22276 2458
rect 22296 2438 22308 2458
rect 22264 2396 22308 2438
rect 22358 2458 22400 2496
rect 22358 2438 22372 2458
rect 22392 2438 22400 2458
rect 22358 2396 22400 2438
rect 22474 2458 22516 2496
rect 22474 2438 22482 2458
rect 22502 2438 22516 2458
rect 22474 2396 22516 2438
rect 22566 2465 22611 2496
rect 22566 2458 22610 2465
rect 22566 2438 22578 2458
rect 22598 2438 22610 2458
rect 22566 2396 22610 2438
rect 33840 2627 33852 2647
rect 33872 2627 33884 2647
rect 33840 2620 33884 2627
rect 33839 2589 33884 2620
rect 33934 2647 33976 2689
rect 33934 2627 33948 2647
rect 33968 2627 33976 2647
rect 33934 2589 33976 2627
rect 34050 2647 34092 2689
rect 34050 2627 34058 2647
rect 34078 2627 34092 2647
rect 34050 2589 34092 2627
rect 34142 2647 34186 2689
rect 34142 2627 34154 2647
rect 34174 2627 34186 2647
rect 34142 2589 34186 2627
rect 34268 2647 34310 2689
rect 34268 2627 34276 2647
rect 34296 2627 34310 2647
rect 34268 2589 34310 2627
rect 34360 2647 34404 2689
rect 34360 2627 34372 2647
rect 34392 2627 34404 2647
rect 34360 2589 34404 2627
rect 26423 2470 26467 2508
rect 26423 2450 26435 2470
rect 26455 2450 26467 2470
rect 20458 2361 20470 2381
rect 20490 2361 20502 2381
rect 20458 2323 20502 2361
rect 12626 2190 12638 2210
rect 12658 2190 12670 2210
rect 12626 2152 12670 2190
rect 4676 2034 4720 2072
rect 832 1959 876 2001
rect 2468 1959 2512 2001
rect 2468 1939 2480 1959
rect 2500 1939 2512 1959
rect 2468 1932 2512 1939
rect 2467 1901 2512 1932
rect 2562 1959 2604 2001
rect 2562 1939 2576 1959
rect 2596 1939 2604 1959
rect 2562 1901 2604 1939
rect 2678 1959 2720 2001
rect 2678 1939 2686 1959
rect 2706 1939 2720 1959
rect 2678 1901 2720 1939
rect 2770 1959 2814 2001
rect 2770 1939 2782 1959
rect 2802 1939 2814 1959
rect 2770 1901 2814 1939
rect 2896 1959 2938 2001
rect 2896 1939 2904 1959
rect 2924 1939 2938 1959
rect 2896 1901 2938 1939
rect 2988 1959 3032 2001
rect 4676 2014 4688 2034
rect 4708 2014 4720 2034
rect 2988 1939 3000 1959
rect 3020 1939 3032 1959
rect 4676 1972 4720 2014
rect 4770 2034 4812 2072
rect 4770 2014 4784 2034
rect 4804 2014 4812 2034
rect 4770 1972 4812 2014
rect 4894 2034 4938 2072
rect 4894 2014 4906 2034
rect 4926 2014 4938 2034
rect 4894 1972 4938 2014
rect 4988 2034 5030 2072
rect 4988 2014 5002 2034
rect 5022 2014 5030 2034
rect 4988 1972 5030 2014
rect 5104 2034 5146 2072
rect 5104 2014 5112 2034
rect 5132 2014 5146 2034
rect 5104 1972 5146 2014
rect 5196 2041 5241 2072
rect 5196 2034 5240 2041
rect 5196 2014 5208 2034
rect 5228 2014 5240 2034
rect 16470 2223 16514 2265
rect 16470 2203 16482 2223
rect 16502 2203 16514 2223
rect 16470 2196 16514 2203
rect 16469 2165 16514 2196
rect 16564 2223 16606 2265
rect 16564 2203 16578 2223
rect 16598 2203 16606 2223
rect 16564 2165 16606 2203
rect 16680 2223 16722 2265
rect 16680 2203 16688 2223
rect 16708 2203 16722 2223
rect 16680 2165 16722 2203
rect 16772 2223 16816 2265
rect 16772 2203 16784 2223
rect 16804 2203 16816 2223
rect 16772 2165 16816 2203
rect 16898 2223 16940 2265
rect 16898 2203 16906 2223
rect 16926 2203 16940 2223
rect 16898 2165 16940 2203
rect 16990 2223 17034 2265
rect 18480 2261 18524 2299
rect 18480 2241 18492 2261
rect 18512 2241 18524 2261
rect 16990 2203 17002 2223
rect 17022 2203 17034 2223
rect 16990 2165 17034 2203
rect 18480 2199 18524 2241
rect 18574 2261 18616 2299
rect 18574 2241 18588 2261
rect 18608 2241 18616 2261
rect 18574 2199 18616 2241
rect 18698 2261 18742 2299
rect 18698 2241 18710 2261
rect 18730 2241 18742 2261
rect 18698 2199 18742 2241
rect 18792 2261 18834 2299
rect 18792 2241 18806 2261
rect 18826 2241 18834 2261
rect 18792 2199 18834 2241
rect 18908 2261 18950 2299
rect 18908 2241 18916 2261
rect 18936 2241 18950 2261
rect 18908 2199 18950 2241
rect 19000 2268 19045 2299
rect 19000 2261 19044 2268
rect 19000 2241 19012 2261
rect 19032 2241 19044 2261
rect 19000 2199 19044 2241
rect 24302 2394 24346 2436
rect 24302 2374 24314 2394
rect 24334 2374 24346 2394
rect 24302 2367 24346 2374
rect 24301 2336 24346 2367
rect 24396 2394 24438 2436
rect 24396 2374 24410 2394
rect 24430 2374 24438 2394
rect 24396 2336 24438 2374
rect 24512 2394 24554 2436
rect 24512 2374 24520 2394
rect 24540 2374 24554 2394
rect 24512 2336 24554 2374
rect 24604 2394 24648 2436
rect 24604 2374 24616 2394
rect 24636 2374 24648 2394
rect 24604 2336 24648 2374
rect 24730 2394 24772 2436
rect 24730 2374 24738 2394
rect 24758 2374 24772 2394
rect 24730 2336 24772 2374
rect 24822 2394 24866 2436
rect 26423 2408 26467 2450
rect 26517 2470 26559 2508
rect 26517 2450 26531 2470
rect 26551 2450 26559 2470
rect 26517 2408 26559 2450
rect 26641 2470 26685 2508
rect 26641 2450 26653 2470
rect 26673 2450 26685 2470
rect 26641 2408 26685 2450
rect 26735 2470 26777 2508
rect 26735 2450 26749 2470
rect 26769 2450 26777 2470
rect 26735 2408 26777 2450
rect 26851 2470 26893 2508
rect 26851 2450 26859 2470
rect 26879 2450 26893 2470
rect 26851 2408 26893 2450
rect 26943 2477 26988 2508
rect 26943 2470 26987 2477
rect 26943 2450 26955 2470
rect 26975 2450 26987 2470
rect 26943 2408 26987 2450
rect 30787 2483 30831 2521
rect 30787 2463 30799 2483
rect 30819 2463 30831 2483
rect 24822 2374 24834 2394
rect 24854 2374 24866 2394
rect 24822 2336 24866 2374
rect 22844 2274 22888 2312
rect 22844 2254 22856 2274
rect 22876 2254 22888 2274
rect 9053 2046 9097 2084
rect 5196 1972 5240 2014
rect 6832 1972 6876 2014
rect 2988 1901 3032 1939
rect 6832 1952 6844 1972
rect 6864 1952 6876 1972
rect 6832 1945 6876 1952
rect 6831 1914 6876 1945
rect 6926 1972 6968 2014
rect 6926 1952 6940 1972
rect 6960 1952 6968 1972
rect 6926 1914 6968 1952
rect 7042 1972 7084 2014
rect 7042 1952 7050 1972
rect 7070 1952 7084 1972
rect 7042 1914 7084 1952
rect 7134 1972 7178 2014
rect 7134 1952 7146 1972
rect 7166 1952 7178 1972
rect 7134 1914 7178 1952
rect 7260 1972 7302 2014
rect 7260 1952 7268 1972
rect 7288 1952 7302 1972
rect 7260 1914 7302 1952
rect 7352 1972 7396 2014
rect 9053 2026 9065 2046
rect 9085 2026 9097 2046
rect 7352 1952 7364 1972
rect 7384 1952 7396 1972
rect 9053 1984 9097 2026
rect 9147 2046 9189 2084
rect 9147 2026 9161 2046
rect 9181 2026 9189 2046
rect 9147 1984 9189 2026
rect 9271 2046 9315 2084
rect 9271 2026 9283 2046
rect 9303 2026 9315 2046
rect 9271 1984 9315 2026
rect 9365 2046 9407 2084
rect 9365 2026 9379 2046
rect 9399 2026 9407 2046
rect 9365 1984 9407 2026
rect 9481 2046 9523 2084
rect 9481 2026 9489 2046
rect 9509 2026 9523 2046
rect 9481 1984 9523 2026
rect 9573 2053 9618 2084
rect 9573 2046 9617 2053
rect 9573 2026 9585 2046
rect 9605 2026 9617 2046
rect 20736 2197 20780 2239
rect 20736 2177 20748 2197
rect 20768 2177 20780 2197
rect 20736 2170 20780 2177
rect 20735 2139 20780 2170
rect 20830 2197 20872 2239
rect 20830 2177 20844 2197
rect 20864 2177 20872 2197
rect 20830 2139 20872 2177
rect 20946 2197 20988 2239
rect 20946 2177 20954 2197
rect 20974 2177 20988 2197
rect 20946 2139 20988 2177
rect 21038 2197 21082 2239
rect 21038 2177 21050 2197
rect 21070 2177 21082 2197
rect 21038 2139 21082 2177
rect 21164 2197 21206 2239
rect 21164 2177 21172 2197
rect 21192 2177 21206 2197
rect 21164 2139 21206 2177
rect 21256 2197 21300 2239
rect 22844 2212 22888 2254
rect 22938 2274 22980 2312
rect 22938 2254 22952 2274
rect 22972 2254 22980 2274
rect 22938 2212 22980 2254
rect 23062 2274 23106 2312
rect 23062 2254 23074 2274
rect 23094 2254 23106 2274
rect 23062 2212 23106 2254
rect 23156 2274 23198 2312
rect 23156 2254 23170 2274
rect 23190 2254 23198 2274
rect 23156 2212 23198 2254
rect 23272 2274 23314 2312
rect 23272 2254 23280 2274
rect 23300 2254 23314 2274
rect 23272 2212 23314 2254
rect 23364 2281 23409 2312
rect 23364 2274 23408 2281
rect 23364 2254 23376 2274
rect 23396 2254 23408 2274
rect 23364 2212 23408 2254
rect 28679 2406 28723 2448
rect 28679 2386 28691 2406
rect 28711 2386 28723 2406
rect 28679 2379 28723 2386
rect 28678 2348 28723 2379
rect 28773 2406 28815 2448
rect 28773 2386 28787 2406
rect 28807 2386 28815 2406
rect 28773 2348 28815 2386
rect 28889 2406 28931 2448
rect 28889 2386 28897 2406
rect 28917 2386 28931 2406
rect 28889 2348 28931 2386
rect 28981 2406 29025 2448
rect 28981 2386 28993 2406
rect 29013 2386 29025 2406
rect 28981 2348 29025 2386
rect 29107 2406 29149 2448
rect 29107 2386 29115 2406
rect 29135 2386 29149 2406
rect 29107 2348 29149 2386
rect 29199 2406 29243 2448
rect 30787 2421 30831 2463
rect 30881 2483 30923 2521
rect 30881 2463 30895 2483
rect 30915 2463 30923 2483
rect 30881 2421 30923 2463
rect 31005 2483 31049 2521
rect 31005 2463 31017 2483
rect 31037 2463 31049 2483
rect 31005 2421 31049 2463
rect 31099 2483 31141 2521
rect 31099 2463 31113 2483
rect 31133 2463 31141 2483
rect 31099 2421 31141 2463
rect 31215 2483 31257 2521
rect 31215 2463 31223 2483
rect 31243 2463 31257 2483
rect 31215 2421 31257 2463
rect 31307 2490 31352 2521
rect 31307 2483 31351 2490
rect 31307 2463 31319 2483
rect 31339 2463 31351 2483
rect 31307 2421 31351 2463
rect 29199 2386 29211 2406
rect 29231 2386 29243 2406
rect 29199 2348 29243 2386
rect 27221 2286 27265 2324
rect 27221 2266 27233 2286
rect 27253 2266 27265 2286
rect 21256 2177 21268 2197
rect 21288 2177 21300 2197
rect 21256 2139 21300 2177
rect 13417 2059 13461 2097
rect 9573 1984 9617 2026
rect 11209 1984 11253 2026
rect 7352 1914 7396 1952
rect 11209 1964 11221 1984
rect 11241 1964 11253 1984
rect 11209 1957 11253 1964
rect 11208 1926 11253 1957
rect 11303 1984 11345 2026
rect 11303 1964 11317 1984
rect 11337 1964 11345 1984
rect 11303 1926 11345 1964
rect 11419 1984 11461 2026
rect 11419 1964 11427 1984
rect 11447 1964 11461 1984
rect 11419 1926 11461 1964
rect 11511 1984 11555 2026
rect 11511 1964 11523 1984
rect 11543 1964 11555 1984
rect 11511 1926 11555 1964
rect 11637 1984 11679 2026
rect 11637 1964 11645 1984
rect 11665 1964 11679 1984
rect 11637 1926 11679 1964
rect 11729 1984 11773 2026
rect 13417 2039 13429 2059
rect 13449 2039 13461 2059
rect 11729 1964 11741 1984
rect 11761 1964 11773 1984
rect 13417 1997 13461 2039
rect 13511 2059 13553 2097
rect 13511 2039 13525 2059
rect 13545 2039 13553 2059
rect 13511 1997 13553 2039
rect 13635 2059 13679 2097
rect 13635 2039 13647 2059
rect 13667 2039 13679 2059
rect 13635 1997 13679 2039
rect 13729 2059 13771 2097
rect 13729 2039 13743 2059
rect 13763 2039 13771 2059
rect 13729 1997 13771 2039
rect 13845 2059 13887 2097
rect 13845 2039 13853 2059
rect 13873 2039 13887 2059
rect 13845 1997 13887 2039
rect 13937 2066 13982 2097
rect 13937 2059 13981 2066
rect 13937 2039 13949 2059
rect 13969 2039 13981 2059
rect 25100 2210 25144 2252
rect 25100 2190 25112 2210
rect 25132 2190 25144 2210
rect 25100 2183 25144 2190
rect 25099 2152 25144 2183
rect 25194 2210 25236 2252
rect 25194 2190 25208 2210
rect 25228 2190 25236 2210
rect 25194 2152 25236 2190
rect 25310 2210 25352 2252
rect 25310 2190 25318 2210
rect 25338 2190 25352 2210
rect 25310 2152 25352 2190
rect 25402 2210 25446 2252
rect 25402 2190 25414 2210
rect 25434 2190 25446 2210
rect 25402 2152 25446 2190
rect 25528 2210 25570 2252
rect 25528 2190 25536 2210
rect 25556 2190 25570 2210
rect 25528 2152 25570 2190
rect 25620 2210 25664 2252
rect 27221 2224 27265 2266
rect 27315 2286 27357 2324
rect 27315 2266 27329 2286
rect 27349 2266 27357 2286
rect 27315 2224 27357 2266
rect 27439 2286 27483 2324
rect 27439 2266 27451 2286
rect 27471 2266 27483 2286
rect 27439 2224 27483 2266
rect 27533 2286 27575 2324
rect 27533 2266 27547 2286
rect 27567 2266 27575 2286
rect 27533 2224 27575 2266
rect 27649 2286 27691 2324
rect 27649 2266 27657 2286
rect 27677 2266 27691 2286
rect 27649 2224 27691 2266
rect 27741 2293 27786 2324
rect 27741 2286 27785 2293
rect 27741 2266 27753 2286
rect 27773 2266 27785 2286
rect 27741 2224 27785 2266
rect 33043 2419 33087 2461
rect 33043 2399 33055 2419
rect 33075 2399 33087 2419
rect 33043 2392 33087 2399
rect 33042 2361 33087 2392
rect 33137 2419 33179 2461
rect 33137 2399 33151 2419
rect 33171 2399 33179 2419
rect 33137 2361 33179 2399
rect 33253 2419 33295 2461
rect 33253 2399 33261 2419
rect 33281 2399 33295 2419
rect 33253 2361 33295 2399
rect 33345 2419 33389 2461
rect 33345 2399 33357 2419
rect 33377 2399 33389 2419
rect 33345 2361 33389 2399
rect 33471 2419 33513 2461
rect 33471 2399 33479 2419
rect 33499 2399 33513 2419
rect 33471 2361 33513 2399
rect 33563 2419 33607 2461
rect 33563 2399 33575 2419
rect 33595 2399 33607 2419
rect 33563 2361 33607 2399
rect 31585 2299 31629 2337
rect 31585 2279 31597 2299
rect 31617 2279 31629 2299
rect 25620 2190 25632 2210
rect 25652 2190 25664 2210
rect 25620 2152 25664 2190
rect 13937 1997 13981 2039
rect 15573 1997 15617 2039
rect 11729 1926 11773 1964
rect 15573 1977 15585 1997
rect 15605 1977 15617 1997
rect 15573 1970 15617 1977
rect 15572 1939 15617 1970
rect 15667 1997 15709 2039
rect 15667 1977 15681 1997
rect 15701 1977 15709 1997
rect 15667 1939 15709 1977
rect 15783 1997 15825 2039
rect 15783 1977 15791 1997
rect 15811 1977 15825 1997
rect 15783 1939 15825 1977
rect 15875 1997 15919 2039
rect 15875 1977 15887 1997
rect 15907 1977 15919 1997
rect 15875 1939 15919 1977
rect 16001 1997 16043 2039
rect 16001 1977 16009 1997
rect 16029 1977 16043 1997
rect 16001 1939 16043 1977
rect 16093 1997 16137 2039
rect 16093 1977 16105 1997
rect 16125 1977 16137 1997
rect 17683 2033 17727 2071
rect 17683 2013 17695 2033
rect 17715 2013 17727 2033
rect 16093 1939 16137 1977
rect 17683 1971 17727 2013
rect 17777 2033 17819 2071
rect 17777 2013 17791 2033
rect 17811 2013 17819 2033
rect 17777 1971 17819 2013
rect 17901 2033 17945 2071
rect 17901 2013 17913 2033
rect 17933 2013 17945 2033
rect 17901 1971 17945 2013
rect 17995 2033 18037 2071
rect 17995 2013 18009 2033
rect 18029 2013 18037 2033
rect 17995 1971 18037 2013
rect 18111 2033 18153 2071
rect 18111 2013 18119 2033
rect 18139 2013 18153 2033
rect 18111 1971 18153 2013
rect 18203 2040 18248 2071
rect 18203 2033 18247 2040
rect 18203 2013 18215 2033
rect 18235 2013 18247 2033
rect 29477 2222 29521 2264
rect 29477 2202 29489 2222
rect 29509 2202 29521 2222
rect 29477 2195 29521 2202
rect 29476 2164 29521 2195
rect 29571 2222 29613 2264
rect 29571 2202 29585 2222
rect 29605 2202 29613 2222
rect 29571 2164 29613 2202
rect 29687 2222 29729 2264
rect 29687 2202 29695 2222
rect 29715 2202 29729 2222
rect 29687 2164 29729 2202
rect 29779 2222 29823 2264
rect 29779 2202 29791 2222
rect 29811 2202 29823 2222
rect 29779 2164 29823 2202
rect 29905 2222 29947 2264
rect 29905 2202 29913 2222
rect 29933 2202 29947 2222
rect 29905 2164 29947 2202
rect 29997 2222 30041 2264
rect 31585 2237 31629 2279
rect 31679 2299 31721 2337
rect 31679 2279 31693 2299
rect 31713 2279 31721 2299
rect 31679 2237 31721 2279
rect 31803 2299 31847 2337
rect 31803 2279 31815 2299
rect 31835 2279 31847 2299
rect 31803 2237 31847 2279
rect 31897 2299 31939 2337
rect 31897 2279 31911 2299
rect 31931 2279 31939 2299
rect 31897 2237 31939 2279
rect 32013 2299 32055 2337
rect 32013 2279 32021 2299
rect 32041 2279 32055 2299
rect 32013 2237 32055 2279
rect 32105 2306 32150 2337
rect 32105 2299 32149 2306
rect 32105 2279 32117 2299
rect 32137 2279 32149 2299
rect 32105 2237 32149 2279
rect 29997 2202 30009 2222
rect 30029 2202 30041 2222
rect 29997 2164 30041 2202
rect 22047 2046 22091 2084
rect 18203 1971 18247 2013
rect 19839 1971 19883 2013
rect 19839 1951 19851 1971
rect 19871 1951 19883 1971
rect 19839 1944 19883 1951
rect 19838 1913 19883 1944
rect 19933 1971 19975 2013
rect 19933 1951 19947 1971
rect 19967 1951 19975 1971
rect 19933 1913 19975 1951
rect 20049 1971 20091 2013
rect 20049 1951 20057 1971
rect 20077 1951 20091 1971
rect 20049 1913 20091 1951
rect 20141 1971 20185 2013
rect 20141 1951 20153 1971
rect 20173 1951 20185 1971
rect 20141 1913 20185 1951
rect 20267 1971 20309 2013
rect 20267 1951 20275 1971
rect 20295 1951 20309 1971
rect 20267 1913 20309 1951
rect 20359 1971 20403 2013
rect 22047 2026 22059 2046
rect 22079 2026 22091 2046
rect 20359 1951 20371 1971
rect 20391 1951 20403 1971
rect 22047 1984 22091 2026
rect 22141 2046 22183 2084
rect 22141 2026 22155 2046
rect 22175 2026 22183 2046
rect 22141 1984 22183 2026
rect 22265 2046 22309 2084
rect 22265 2026 22277 2046
rect 22297 2026 22309 2046
rect 22265 1984 22309 2026
rect 22359 2046 22401 2084
rect 22359 2026 22373 2046
rect 22393 2026 22401 2046
rect 22359 1984 22401 2026
rect 22475 2046 22517 2084
rect 22475 2026 22483 2046
rect 22503 2026 22517 2046
rect 22475 1984 22517 2026
rect 22567 2053 22612 2084
rect 22567 2046 22611 2053
rect 22567 2026 22579 2046
rect 22599 2026 22611 2046
rect 33841 2235 33885 2277
rect 33841 2215 33853 2235
rect 33873 2215 33885 2235
rect 33841 2208 33885 2215
rect 33840 2177 33885 2208
rect 33935 2235 33977 2277
rect 33935 2215 33949 2235
rect 33969 2215 33977 2235
rect 33935 2177 33977 2215
rect 34051 2235 34093 2277
rect 34051 2215 34059 2235
rect 34079 2215 34093 2235
rect 34051 2177 34093 2215
rect 34143 2235 34187 2277
rect 34143 2215 34155 2235
rect 34175 2215 34187 2235
rect 34143 2177 34187 2215
rect 34269 2235 34311 2277
rect 34269 2215 34277 2235
rect 34297 2215 34311 2235
rect 34269 2177 34311 2215
rect 34361 2235 34405 2277
rect 34361 2215 34373 2235
rect 34393 2215 34405 2235
rect 34361 2177 34405 2215
rect 26424 2058 26468 2096
rect 22567 1984 22611 2026
rect 24203 1984 24247 2026
rect 20359 1913 20403 1951
rect 24203 1964 24215 1984
rect 24235 1964 24247 1984
rect 24203 1957 24247 1964
rect 24202 1926 24247 1957
rect 24297 1984 24339 2026
rect 24297 1964 24311 1984
rect 24331 1964 24339 1984
rect 24297 1926 24339 1964
rect 24413 1984 24455 2026
rect 24413 1964 24421 1984
rect 24441 1964 24455 1984
rect 24413 1926 24455 1964
rect 24505 1984 24549 2026
rect 24505 1964 24517 1984
rect 24537 1964 24549 1984
rect 24505 1926 24549 1964
rect 24631 1984 24673 2026
rect 24631 1964 24639 1984
rect 24659 1964 24673 1984
rect 24631 1926 24673 1964
rect 24723 1984 24767 2026
rect 26424 2038 26436 2058
rect 26456 2038 26468 2058
rect 24723 1964 24735 1984
rect 24755 1964 24767 1984
rect 26424 1996 26468 2038
rect 26518 2058 26560 2096
rect 26518 2038 26532 2058
rect 26552 2038 26560 2058
rect 26518 1996 26560 2038
rect 26642 2058 26686 2096
rect 26642 2038 26654 2058
rect 26674 2038 26686 2058
rect 26642 1996 26686 2038
rect 26736 2058 26778 2096
rect 26736 2038 26750 2058
rect 26770 2038 26778 2058
rect 26736 1996 26778 2038
rect 26852 2058 26894 2096
rect 26852 2038 26860 2058
rect 26880 2038 26894 2058
rect 26852 1996 26894 2038
rect 26944 2065 26989 2096
rect 26944 2058 26988 2065
rect 26944 2038 26956 2058
rect 26976 2038 26988 2058
rect 30788 2071 30832 2109
rect 26944 1996 26988 2038
rect 28580 1996 28624 2038
rect 24723 1926 24767 1964
rect 28580 1976 28592 1996
rect 28612 1976 28624 1996
rect 28580 1969 28624 1976
rect 28579 1938 28624 1969
rect 28674 1996 28716 2038
rect 28674 1976 28688 1996
rect 28708 1976 28716 1996
rect 28674 1938 28716 1976
rect 28790 1996 28832 2038
rect 28790 1976 28798 1996
rect 28818 1976 28832 1996
rect 28790 1938 28832 1976
rect 28882 1996 28926 2038
rect 28882 1976 28894 1996
rect 28914 1976 28926 1996
rect 28882 1938 28926 1976
rect 29008 1996 29050 2038
rect 29008 1976 29016 1996
rect 29036 1976 29050 1996
rect 29008 1938 29050 1976
rect 29100 1996 29144 2038
rect 30788 2051 30800 2071
rect 30820 2051 30832 2071
rect 29100 1976 29112 1996
rect 29132 1976 29144 1996
rect 30788 2009 30832 2051
rect 30882 2071 30924 2109
rect 30882 2051 30896 2071
rect 30916 2051 30924 2071
rect 30882 2009 30924 2051
rect 31006 2071 31050 2109
rect 31006 2051 31018 2071
rect 31038 2051 31050 2071
rect 31006 2009 31050 2051
rect 31100 2071 31142 2109
rect 31100 2051 31114 2071
rect 31134 2051 31142 2071
rect 31100 2009 31142 2051
rect 31216 2071 31258 2109
rect 31216 2051 31224 2071
rect 31244 2051 31258 2071
rect 31216 2009 31258 2051
rect 31308 2078 31353 2109
rect 31308 2071 31352 2078
rect 31308 2051 31320 2071
rect 31340 2051 31352 2071
rect 31308 2009 31352 2051
rect 32944 2009 32988 2051
rect 29100 1938 29144 1976
rect 32944 1989 32956 2009
rect 32976 1989 32988 2009
rect 32944 1982 32988 1989
rect 32943 1951 32988 1982
rect 33038 2009 33080 2051
rect 33038 1989 33052 2009
rect 33072 1989 33080 2009
rect 33038 1951 33080 1989
rect 33154 2009 33196 2051
rect 33154 1989 33162 2009
rect 33182 1989 33196 2009
rect 33154 1951 33196 1989
rect 33246 2009 33290 2051
rect 33246 1989 33258 2009
rect 33278 1989 33290 2009
rect 33246 1951 33290 1989
rect 33372 2009 33414 2051
rect 33372 1989 33380 2009
rect 33400 1989 33414 2009
rect 33372 1951 33414 1989
rect 33464 2009 33508 2051
rect 33464 1989 33476 2009
rect 33496 1989 33508 2009
rect 33464 1951 33508 1989
rect 1191 1641 1235 1679
rect 1191 1621 1203 1641
rect 1223 1621 1235 1641
rect 1191 1579 1235 1621
rect 1285 1641 1327 1679
rect 1285 1621 1299 1641
rect 1319 1621 1327 1641
rect 1285 1579 1327 1621
rect 1409 1641 1453 1679
rect 1409 1621 1421 1641
rect 1441 1621 1453 1641
rect 1409 1579 1453 1621
rect 1503 1641 1545 1679
rect 1503 1621 1517 1641
rect 1537 1621 1545 1641
rect 1503 1579 1545 1621
rect 1619 1641 1661 1679
rect 1619 1621 1627 1641
rect 1647 1621 1661 1641
rect 1619 1579 1661 1621
rect 1711 1648 1756 1679
rect 1711 1641 1755 1648
rect 1711 1621 1723 1641
rect 1743 1621 1755 1641
rect 5555 1654 5599 1692
rect 1711 1579 1755 1621
rect 3347 1579 3391 1621
rect 3347 1559 3359 1579
rect 3379 1559 3391 1579
rect 3347 1552 3391 1559
rect 3346 1521 3391 1552
rect 3441 1579 3483 1621
rect 3441 1559 3455 1579
rect 3475 1559 3483 1579
rect 3441 1521 3483 1559
rect 3557 1579 3599 1621
rect 3557 1559 3565 1579
rect 3585 1559 3599 1579
rect 3557 1521 3599 1559
rect 3649 1579 3693 1621
rect 3649 1559 3661 1579
rect 3681 1559 3693 1579
rect 3649 1521 3693 1559
rect 3775 1579 3817 1621
rect 3775 1559 3783 1579
rect 3803 1559 3817 1579
rect 3775 1521 3817 1559
rect 3867 1579 3911 1621
rect 5555 1634 5567 1654
rect 5587 1634 5599 1654
rect 3867 1559 3879 1579
rect 3899 1559 3911 1579
rect 5555 1592 5599 1634
rect 5649 1654 5691 1692
rect 5649 1634 5663 1654
rect 5683 1634 5691 1654
rect 5649 1592 5691 1634
rect 5773 1654 5817 1692
rect 5773 1634 5785 1654
rect 5805 1634 5817 1654
rect 5773 1592 5817 1634
rect 5867 1654 5909 1692
rect 5867 1634 5881 1654
rect 5901 1634 5909 1654
rect 5867 1592 5909 1634
rect 5983 1654 6025 1692
rect 5983 1634 5991 1654
rect 6011 1634 6025 1654
rect 5983 1592 6025 1634
rect 6075 1661 6120 1692
rect 6075 1654 6119 1661
rect 6075 1634 6087 1654
rect 6107 1634 6119 1654
rect 9932 1666 9976 1704
rect 6075 1592 6119 1634
rect 7711 1592 7755 1634
rect 3867 1521 3911 1559
rect 7711 1572 7723 1592
rect 7743 1572 7755 1592
rect 7711 1565 7755 1572
rect 7710 1534 7755 1565
rect 7805 1592 7847 1634
rect 7805 1572 7819 1592
rect 7839 1572 7847 1592
rect 7805 1534 7847 1572
rect 7921 1592 7963 1634
rect 7921 1572 7929 1592
rect 7949 1572 7963 1592
rect 7921 1534 7963 1572
rect 8013 1592 8057 1634
rect 8013 1572 8025 1592
rect 8045 1572 8057 1592
rect 8013 1534 8057 1572
rect 8139 1592 8181 1634
rect 8139 1572 8147 1592
rect 8167 1572 8181 1592
rect 8139 1534 8181 1572
rect 8231 1592 8275 1634
rect 9932 1646 9944 1666
rect 9964 1646 9976 1666
rect 8231 1572 8243 1592
rect 8263 1572 8275 1592
rect 9932 1604 9976 1646
rect 10026 1666 10068 1704
rect 10026 1646 10040 1666
rect 10060 1646 10068 1666
rect 10026 1604 10068 1646
rect 10150 1666 10194 1704
rect 10150 1646 10162 1666
rect 10182 1646 10194 1666
rect 10150 1604 10194 1646
rect 10244 1666 10286 1704
rect 10244 1646 10258 1666
rect 10278 1646 10286 1666
rect 10244 1604 10286 1646
rect 10360 1666 10402 1704
rect 10360 1646 10368 1666
rect 10388 1646 10402 1666
rect 10360 1604 10402 1646
rect 10452 1673 10497 1704
rect 10452 1666 10496 1673
rect 10452 1646 10464 1666
rect 10484 1646 10496 1666
rect 14296 1679 14340 1717
rect 10452 1604 10496 1646
rect 12088 1604 12132 1646
rect 8231 1534 8275 1572
rect 294 1415 338 1453
rect 294 1395 306 1415
rect 326 1395 338 1415
rect 294 1353 338 1395
rect 388 1415 430 1453
rect 388 1395 402 1415
rect 422 1395 430 1415
rect 388 1353 430 1395
rect 512 1415 556 1453
rect 512 1395 524 1415
rect 544 1395 556 1415
rect 512 1353 556 1395
rect 606 1415 648 1453
rect 606 1395 620 1415
rect 640 1395 648 1415
rect 606 1353 648 1395
rect 722 1415 764 1453
rect 722 1395 730 1415
rect 750 1395 764 1415
rect 722 1353 764 1395
rect 814 1422 859 1453
rect 814 1415 858 1422
rect 814 1395 826 1415
rect 846 1395 858 1415
rect 814 1353 858 1395
rect 12088 1584 12100 1604
rect 12120 1584 12132 1604
rect 12088 1577 12132 1584
rect 12087 1546 12132 1577
rect 12182 1604 12224 1646
rect 12182 1584 12196 1604
rect 12216 1584 12224 1604
rect 12182 1546 12224 1584
rect 12298 1604 12340 1646
rect 12298 1584 12306 1604
rect 12326 1584 12340 1604
rect 12298 1546 12340 1584
rect 12390 1604 12434 1646
rect 12390 1584 12402 1604
rect 12422 1584 12434 1604
rect 12390 1546 12434 1584
rect 12516 1604 12558 1646
rect 12516 1584 12524 1604
rect 12544 1584 12558 1604
rect 12516 1546 12558 1584
rect 12608 1604 12652 1646
rect 14296 1659 14308 1679
rect 14328 1659 14340 1679
rect 12608 1584 12620 1604
rect 12640 1584 12652 1604
rect 14296 1617 14340 1659
rect 14390 1679 14432 1717
rect 14390 1659 14404 1679
rect 14424 1659 14432 1679
rect 14390 1617 14432 1659
rect 14514 1679 14558 1717
rect 14514 1659 14526 1679
rect 14546 1659 14558 1679
rect 14514 1617 14558 1659
rect 14608 1679 14650 1717
rect 14608 1659 14622 1679
rect 14642 1659 14650 1679
rect 14608 1617 14650 1659
rect 14724 1679 14766 1717
rect 14724 1659 14732 1679
rect 14752 1659 14766 1679
rect 14724 1617 14766 1659
rect 14816 1686 14861 1717
rect 14816 1679 14860 1686
rect 14816 1659 14828 1679
rect 14848 1659 14860 1679
rect 14816 1617 14860 1659
rect 16452 1617 16496 1659
rect 12608 1546 12652 1584
rect 4658 1428 4702 1466
rect 4658 1408 4670 1428
rect 4690 1408 4702 1428
rect 2550 1351 2594 1393
rect 2550 1331 2562 1351
rect 2582 1331 2594 1351
rect 2550 1324 2594 1331
rect 2549 1293 2594 1324
rect 2644 1351 2686 1393
rect 2644 1331 2658 1351
rect 2678 1331 2686 1351
rect 2644 1293 2686 1331
rect 2760 1351 2802 1393
rect 2760 1331 2768 1351
rect 2788 1331 2802 1351
rect 2760 1293 2802 1331
rect 2852 1351 2896 1393
rect 2852 1331 2864 1351
rect 2884 1331 2896 1351
rect 2852 1293 2896 1331
rect 2978 1351 3020 1393
rect 2978 1331 2986 1351
rect 3006 1331 3020 1351
rect 2978 1293 3020 1331
rect 3070 1351 3114 1393
rect 4658 1366 4702 1408
rect 4752 1428 4794 1466
rect 4752 1408 4766 1428
rect 4786 1408 4794 1428
rect 4752 1366 4794 1408
rect 4876 1428 4920 1466
rect 4876 1408 4888 1428
rect 4908 1408 4920 1428
rect 4876 1366 4920 1408
rect 4970 1428 5012 1466
rect 4970 1408 4984 1428
rect 5004 1408 5012 1428
rect 4970 1366 5012 1408
rect 5086 1428 5128 1466
rect 5086 1408 5094 1428
rect 5114 1408 5128 1428
rect 5086 1366 5128 1408
rect 5178 1435 5223 1466
rect 5178 1428 5222 1435
rect 5178 1408 5190 1428
rect 5210 1408 5222 1428
rect 5178 1366 5222 1408
rect 16452 1597 16464 1617
rect 16484 1597 16496 1617
rect 16452 1590 16496 1597
rect 16451 1559 16496 1590
rect 16546 1617 16588 1659
rect 16546 1597 16560 1617
rect 16580 1597 16588 1617
rect 16546 1559 16588 1597
rect 16662 1617 16704 1659
rect 16662 1597 16670 1617
rect 16690 1597 16704 1617
rect 16662 1559 16704 1597
rect 16754 1617 16798 1659
rect 16754 1597 16766 1617
rect 16786 1597 16798 1617
rect 16754 1559 16798 1597
rect 16880 1617 16922 1659
rect 16880 1597 16888 1617
rect 16908 1597 16922 1617
rect 16880 1559 16922 1597
rect 16972 1617 17016 1659
rect 18562 1653 18606 1691
rect 16972 1597 16984 1617
rect 17004 1597 17016 1617
rect 16972 1559 17016 1597
rect 18562 1633 18574 1653
rect 18594 1633 18606 1653
rect 18562 1591 18606 1633
rect 18656 1653 18698 1691
rect 18656 1633 18670 1653
rect 18690 1633 18698 1653
rect 18656 1591 18698 1633
rect 18780 1653 18824 1691
rect 18780 1633 18792 1653
rect 18812 1633 18824 1653
rect 18780 1591 18824 1633
rect 18874 1653 18916 1691
rect 18874 1633 18888 1653
rect 18908 1633 18916 1653
rect 18874 1591 18916 1633
rect 18990 1653 19032 1691
rect 18990 1633 18998 1653
rect 19018 1633 19032 1653
rect 18990 1591 19032 1633
rect 19082 1660 19127 1691
rect 19082 1653 19126 1660
rect 19082 1633 19094 1653
rect 19114 1633 19126 1653
rect 22926 1666 22970 1704
rect 19082 1591 19126 1633
rect 20718 1591 20762 1633
rect 9035 1440 9079 1478
rect 9035 1420 9047 1440
rect 9067 1420 9079 1440
rect 3070 1331 3082 1351
rect 3102 1331 3114 1351
rect 3070 1293 3114 1331
rect 1092 1231 1136 1269
rect 1092 1211 1104 1231
rect 1124 1211 1136 1231
rect 1092 1169 1136 1211
rect 1186 1231 1228 1269
rect 1186 1211 1200 1231
rect 1220 1211 1228 1231
rect 1186 1169 1228 1211
rect 1310 1231 1354 1269
rect 1310 1211 1322 1231
rect 1342 1211 1354 1231
rect 1310 1169 1354 1211
rect 1404 1231 1446 1269
rect 1404 1211 1418 1231
rect 1438 1211 1446 1231
rect 1404 1169 1446 1211
rect 1520 1231 1562 1269
rect 1520 1211 1528 1231
rect 1548 1211 1562 1231
rect 1520 1169 1562 1211
rect 1612 1238 1657 1269
rect 1612 1231 1656 1238
rect 1612 1211 1624 1231
rect 1644 1211 1656 1231
rect 1612 1169 1656 1211
rect 6914 1364 6958 1406
rect 6914 1344 6926 1364
rect 6946 1344 6958 1364
rect 6914 1337 6958 1344
rect 6913 1306 6958 1337
rect 7008 1364 7050 1406
rect 7008 1344 7022 1364
rect 7042 1344 7050 1364
rect 7008 1306 7050 1344
rect 7124 1364 7166 1406
rect 7124 1344 7132 1364
rect 7152 1344 7166 1364
rect 7124 1306 7166 1344
rect 7216 1364 7260 1406
rect 7216 1344 7228 1364
rect 7248 1344 7260 1364
rect 7216 1306 7260 1344
rect 7342 1364 7384 1406
rect 7342 1344 7350 1364
rect 7370 1344 7384 1364
rect 7342 1306 7384 1344
rect 7434 1364 7478 1406
rect 9035 1378 9079 1420
rect 9129 1440 9171 1478
rect 9129 1420 9143 1440
rect 9163 1420 9171 1440
rect 9129 1378 9171 1420
rect 9253 1440 9297 1478
rect 9253 1420 9265 1440
rect 9285 1420 9297 1440
rect 9253 1378 9297 1420
rect 9347 1440 9389 1478
rect 9347 1420 9361 1440
rect 9381 1420 9389 1440
rect 9347 1378 9389 1420
rect 9463 1440 9505 1478
rect 9463 1420 9471 1440
rect 9491 1420 9505 1440
rect 9463 1378 9505 1420
rect 9555 1447 9600 1478
rect 9555 1440 9599 1447
rect 9555 1420 9567 1440
rect 9587 1420 9599 1440
rect 9555 1378 9599 1420
rect 20718 1571 20730 1591
rect 20750 1571 20762 1591
rect 20718 1564 20762 1571
rect 20717 1533 20762 1564
rect 20812 1591 20854 1633
rect 20812 1571 20826 1591
rect 20846 1571 20854 1591
rect 20812 1533 20854 1571
rect 20928 1591 20970 1633
rect 20928 1571 20936 1591
rect 20956 1571 20970 1591
rect 20928 1533 20970 1571
rect 21020 1591 21064 1633
rect 21020 1571 21032 1591
rect 21052 1571 21064 1591
rect 21020 1533 21064 1571
rect 21146 1591 21188 1633
rect 21146 1571 21154 1591
rect 21174 1571 21188 1591
rect 21146 1533 21188 1571
rect 21238 1591 21282 1633
rect 22926 1646 22938 1666
rect 22958 1646 22970 1666
rect 21238 1571 21250 1591
rect 21270 1571 21282 1591
rect 22926 1604 22970 1646
rect 23020 1666 23062 1704
rect 23020 1646 23034 1666
rect 23054 1646 23062 1666
rect 23020 1604 23062 1646
rect 23144 1666 23188 1704
rect 23144 1646 23156 1666
rect 23176 1646 23188 1666
rect 23144 1604 23188 1646
rect 23238 1666 23280 1704
rect 23238 1646 23252 1666
rect 23272 1646 23280 1666
rect 23238 1604 23280 1646
rect 23354 1666 23396 1704
rect 23354 1646 23362 1666
rect 23382 1646 23396 1666
rect 23354 1604 23396 1646
rect 23446 1673 23491 1704
rect 23446 1666 23490 1673
rect 23446 1646 23458 1666
rect 23478 1646 23490 1666
rect 27303 1678 27347 1716
rect 23446 1604 23490 1646
rect 25082 1604 25126 1646
rect 21238 1533 21282 1571
rect 13399 1453 13443 1491
rect 13399 1433 13411 1453
rect 13431 1433 13443 1453
rect 7434 1344 7446 1364
rect 7466 1344 7478 1364
rect 7434 1306 7478 1344
rect 5456 1244 5500 1282
rect 5456 1224 5468 1244
rect 5488 1224 5500 1244
rect 3348 1167 3392 1209
rect 3348 1147 3360 1167
rect 3380 1147 3392 1167
rect 3348 1140 3392 1147
rect 3347 1109 3392 1140
rect 3442 1167 3484 1209
rect 3442 1147 3456 1167
rect 3476 1147 3484 1167
rect 3442 1109 3484 1147
rect 3558 1167 3600 1209
rect 3558 1147 3566 1167
rect 3586 1147 3600 1167
rect 3558 1109 3600 1147
rect 3650 1167 3694 1209
rect 3650 1147 3662 1167
rect 3682 1147 3694 1167
rect 3650 1109 3694 1147
rect 3776 1167 3818 1209
rect 3776 1147 3784 1167
rect 3804 1147 3818 1167
rect 3776 1109 3818 1147
rect 3868 1167 3912 1209
rect 5456 1182 5500 1224
rect 5550 1244 5592 1282
rect 5550 1224 5564 1244
rect 5584 1224 5592 1244
rect 5550 1182 5592 1224
rect 5674 1244 5718 1282
rect 5674 1224 5686 1244
rect 5706 1224 5718 1244
rect 5674 1182 5718 1224
rect 5768 1244 5810 1282
rect 5768 1224 5782 1244
rect 5802 1224 5810 1244
rect 5768 1182 5810 1224
rect 5884 1244 5926 1282
rect 5884 1224 5892 1244
rect 5912 1224 5926 1244
rect 5884 1182 5926 1224
rect 5976 1251 6021 1282
rect 5976 1244 6020 1251
rect 5976 1224 5988 1244
rect 6008 1224 6020 1244
rect 5976 1182 6020 1224
rect 11291 1376 11335 1418
rect 11291 1356 11303 1376
rect 11323 1356 11335 1376
rect 11291 1349 11335 1356
rect 11290 1318 11335 1349
rect 11385 1376 11427 1418
rect 11385 1356 11399 1376
rect 11419 1356 11427 1376
rect 11385 1318 11427 1356
rect 11501 1376 11543 1418
rect 11501 1356 11509 1376
rect 11529 1356 11543 1376
rect 11501 1318 11543 1356
rect 11593 1376 11637 1418
rect 11593 1356 11605 1376
rect 11625 1356 11637 1376
rect 11593 1318 11637 1356
rect 11719 1376 11761 1418
rect 11719 1356 11727 1376
rect 11747 1356 11761 1376
rect 11719 1318 11761 1356
rect 11811 1376 11855 1418
rect 13399 1391 13443 1433
rect 13493 1453 13535 1491
rect 13493 1433 13507 1453
rect 13527 1433 13535 1453
rect 13493 1391 13535 1433
rect 13617 1453 13661 1491
rect 13617 1433 13629 1453
rect 13649 1433 13661 1453
rect 13617 1391 13661 1433
rect 13711 1453 13753 1491
rect 13711 1433 13725 1453
rect 13745 1433 13753 1453
rect 13711 1391 13753 1433
rect 13827 1453 13869 1491
rect 13827 1433 13835 1453
rect 13855 1433 13869 1453
rect 13827 1391 13869 1433
rect 13919 1460 13964 1491
rect 13919 1453 13963 1460
rect 13919 1433 13931 1453
rect 13951 1433 13963 1453
rect 13919 1391 13963 1433
rect 25082 1584 25094 1604
rect 25114 1584 25126 1604
rect 25082 1577 25126 1584
rect 25081 1546 25126 1577
rect 25176 1604 25218 1646
rect 25176 1584 25190 1604
rect 25210 1584 25218 1604
rect 25176 1546 25218 1584
rect 25292 1604 25334 1646
rect 25292 1584 25300 1604
rect 25320 1584 25334 1604
rect 25292 1546 25334 1584
rect 25384 1604 25428 1646
rect 25384 1584 25396 1604
rect 25416 1584 25428 1604
rect 25384 1546 25428 1584
rect 25510 1604 25552 1646
rect 25510 1584 25518 1604
rect 25538 1584 25552 1604
rect 25510 1546 25552 1584
rect 25602 1604 25646 1646
rect 27303 1658 27315 1678
rect 27335 1658 27347 1678
rect 25602 1584 25614 1604
rect 25634 1584 25646 1604
rect 27303 1616 27347 1658
rect 27397 1678 27439 1716
rect 27397 1658 27411 1678
rect 27431 1658 27439 1678
rect 27397 1616 27439 1658
rect 27521 1678 27565 1716
rect 27521 1658 27533 1678
rect 27553 1658 27565 1678
rect 27521 1616 27565 1658
rect 27615 1678 27657 1716
rect 27615 1658 27629 1678
rect 27649 1658 27657 1678
rect 27615 1616 27657 1658
rect 27731 1678 27773 1716
rect 27731 1658 27739 1678
rect 27759 1658 27773 1678
rect 27731 1616 27773 1658
rect 27823 1685 27868 1716
rect 27823 1678 27867 1685
rect 27823 1658 27835 1678
rect 27855 1658 27867 1678
rect 31667 1691 31711 1729
rect 27823 1616 27867 1658
rect 29459 1616 29503 1658
rect 25602 1546 25646 1584
rect 11811 1356 11823 1376
rect 11843 1356 11855 1376
rect 11811 1318 11855 1356
rect 9833 1256 9877 1294
rect 9833 1236 9845 1256
rect 9865 1236 9877 1256
rect 3868 1147 3880 1167
rect 3900 1147 3912 1167
rect 3868 1109 3912 1147
rect 7712 1180 7756 1222
rect 7712 1160 7724 1180
rect 7744 1160 7756 1180
rect 7712 1153 7756 1160
rect 7711 1122 7756 1153
rect 7806 1180 7848 1222
rect 7806 1160 7820 1180
rect 7840 1160 7848 1180
rect 7806 1122 7848 1160
rect 7922 1180 7964 1222
rect 7922 1160 7930 1180
rect 7950 1160 7964 1180
rect 7922 1122 7964 1160
rect 8014 1180 8058 1222
rect 8014 1160 8026 1180
rect 8046 1160 8058 1180
rect 8014 1122 8058 1160
rect 8140 1180 8182 1222
rect 8140 1160 8148 1180
rect 8168 1160 8182 1180
rect 8140 1122 8182 1160
rect 8232 1180 8276 1222
rect 9833 1194 9877 1236
rect 9927 1256 9969 1294
rect 9927 1236 9941 1256
rect 9961 1236 9969 1256
rect 9927 1194 9969 1236
rect 10051 1256 10095 1294
rect 10051 1236 10063 1256
rect 10083 1236 10095 1256
rect 10051 1194 10095 1236
rect 10145 1256 10187 1294
rect 10145 1236 10159 1256
rect 10179 1236 10187 1256
rect 10145 1194 10187 1236
rect 10261 1256 10303 1294
rect 10261 1236 10269 1256
rect 10289 1236 10303 1256
rect 10261 1194 10303 1236
rect 10353 1263 10398 1294
rect 10353 1256 10397 1263
rect 10353 1236 10365 1256
rect 10385 1236 10397 1256
rect 10353 1194 10397 1236
rect 15655 1389 15699 1431
rect 15655 1369 15667 1389
rect 15687 1369 15699 1389
rect 15655 1362 15699 1369
rect 15654 1331 15699 1362
rect 15749 1389 15791 1431
rect 15749 1369 15763 1389
rect 15783 1369 15791 1389
rect 15749 1331 15791 1369
rect 15865 1389 15907 1431
rect 15865 1369 15873 1389
rect 15893 1369 15907 1389
rect 15865 1331 15907 1369
rect 15957 1389 16001 1431
rect 15957 1369 15969 1389
rect 15989 1369 16001 1389
rect 15957 1331 16001 1369
rect 16083 1389 16125 1431
rect 16083 1369 16091 1389
rect 16111 1369 16125 1389
rect 16083 1331 16125 1369
rect 16175 1389 16219 1431
rect 17665 1427 17709 1465
rect 17665 1407 17677 1427
rect 17697 1407 17709 1427
rect 16175 1369 16187 1389
rect 16207 1369 16219 1389
rect 16175 1331 16219 1369
rect 17665 1365 17709 1407
rect 17759 1427 17801 1465
rect 17759 1407 17773 1427
rect 17793 1407 17801 1427
rect 17759 1365 17801 1407
rect 17883 1427 17927 1465
rect 17883 1407 17895 1427
rect 17915 1407 17927 1427
rect 17883 1365 17927 1407
rect 17977 1427 18019 1465
rect 17977 1407 17991 1427
rect 18011 1407 18019 1427
rect 17977 1365 18019 1407
rect 18093 1427 18135 1465
rect 18093 1407 18101 1427
rect 18121 1407 18135 1427
rect 18093 1365 18135 1407
rect 18185 1434 18230 1465
rect 18185 1427 18229 1434
rect 18185 1407 18197 1427
rect 18217 1407 18229 1427
rect 18185 1365 18229 1407
rect 29459 1596 29471 1616
rect 29491 1596 29503 1616
rect 29459 1589 29503 1596
rect 29458 1558 29503 1589
rect 29553 1616 29595 1658
rect 29553 1596 29567 1616
rect 29587 1596 29595 1616
rect 29553 1558 29595 1596
rect 29669 1616 29711 1658
rect 29669 1596 29677 1616
rect 29697 1596 29711 1616
rect 29669 1558 29711 1596
rect 29761 1616 29805 1658
rect 29761 1596 29773 1616
rect 29793 1596 29805 1616
rect 29761 1558 29805 1596
rect 29887 1616 29929 1658
rect 29887 1596 29895 1616
rect 29915 1596 29929 1616
rect 29887 1558 29929 1596
rect 29979 1616 30023 1658
rect 31667 1671 31679 1691
rect 31699 1671 31711 1691
rect 29979 1596 29991 1616
rect 30011 1596 30023 1616
rect 31667 1629 31711 1671
rect 31761 1691 31803 1729
rect 31761 1671 31775 1691
rect 31795 1671 31803 1691
rect 31761 1629 31803 1671
rect 31885 1691 31929 1729
rect 31885 1671 31897 1691
rect 31917 1671 31929 1691
rect 31885 1629 31929 1671
rect 31979 1691 32021 1729
rect 31979 1671 31993 1691
rect 32013 1671 32021 1691
rect 31979 1629 32021 1671
rect 32095 1691 32137 1729
rect 32095 1671 32103 1691
rect 32123 1671 32137 1691
rect 32095 1629 32137 1671
rect 32187 1698 32232 1729
rect 32187 1691 32231 1698
rect 32187 1671 32199 1691
rect 32219 1671 32231 1691
rect 32187 1629 32231 1671
rect 33823 1629 33867 1671
rect 29979 1558 30023 1596
rect 22029 1440 22073 1478
rect 22029 1420 22041 1440
rect 22061 1420 22073 1440
rect 14197 1269 14241 1307
rect 14197 1249 14209 1269
rect 14229 1249 14241 1269
rect 8232 1160 8244 1180
rect 8264 1160 8276 1180
rect 8232 1122 8276 1160
rect 12089 1192 12133 1234
rect 12089 1172 12101 1192
rect 12121 1172 12133 1192
rect 12089 1165 12133 1172
rect 12088 1134 12133 1165
rect 12183 1192 12225 1234
rect 12183 1172 12197 1192
rect 12217 1172 12225 1192
rect 12183 1134 12225 1172
rect 12299 1192 12341 1234
rect 12299 1172 12307 1192
rect 12327 1172 12341 1192
rect 12299 1134 12341 1172
rect 12391 1192 12435 1234
rect 12391 1172 12403 1192
rect 12423 1172 12435 1192
rect 12391 1134 12435 1172
rect 12517 1192 12559 1234
rect 12517 1172 12525 1192
rect 12545 1172 12559 1192
rect 12517 1134 12559 1172
rect 12609 1192 12653 1234
rect 14197 1207 14241 1249
rect 14291 1269 14333 1307
rect 14291 1249 14305 1269
rect 14325 1249 14333 1269
rect 14291 1207 14333 1249
rect 14415 1269 14459 1307
rect 14415 1249 14427 1269
rect 14447 1249 14459 1269
rect 14415 1207 14459 1249
rect 14509 1269 14551 1307
rect 14509 1249 14523 1269
rect 14543 1249 14551 1269
rect 14509 1207 14551 1249
rect 14625 1269 14667 1307
rect 14625 1249 14633 1269
rect 14653 1249 14667 1269
rect 14625 1207 14667 1249
rect 14717 1276 14762 1307
rect 14717 1269 14761 1276
rect 14717 1249 14729 1269
rect 14749 1249 14761 1269
rect 14717 1207 14761 1249
rect 19921 1363 19965 1405
rect 19921 1343 19933 1363
rect 19953 1343 19965 1363
rect 19921 1336 19965 1343
rect 19920 1305 19965 1336
rect 20015 1363 20057 1405
rect 20015 1343 20029 1363
rect 20049 1343 20057 1363
rect 20015 1305 20057 1343
rect 20131 1363 20173 1405
rect 20131 1343 20139 1363
rect 20159 1343 20173 1363
rect 20131 1305 20173 1343
rect 20223 1363 20267 1405
rect 20223 1343 20235 1363
rect 20255 1343 20267 1363
rect 20223 1305 20267 1343
rect 20349 1363 20391 1405
rect 20349 1343 20357 1363
rect 20377 1343 20391 1363
rect 20349 1305 20391 1343
rect 20441 1363 20485 1405
rect 22029 1378 22073 1420
rect 22123 1440 22165 1478
rect 22123 1420 22137 1440
rect 22157 1420 22165 1440
rect 22123 1378 22165 1420
rect 22247 1440 22291 1478
rect 22247 1420 22259 1440
rect 22279 1420 22291 1440
rect 22247 1378 22291 1420
rect 22341 1440 22383 1478
rect 22341 1420 22355 1440
rect 22375 1420 22383 1440
rect 22341 1378 22383 1420
rect 22457 1440 22499 1478
rect 22457 1420 22465 1440
rect 22485 1420 22499 1440
rect 22457 1378 22499 1420
rect 22549 1447 22594 1478
rect 22549 1440 22593 1447
rect 22549 1420 22561 1440
rect 22581 1420 22593 1440
rect 22549 1378 22593 1420
rect 33823 1609 33835 1629
rect 33855 1609 33867 1629
rect 33823 1602 33867 1609
rect 33822 1571 33867 1602
rect 33917 1629 33959 1671
rect 33917 1609 33931 1629
rect 33951 1609 33959 1629
rect 33917 1571 33959 1609
rect 34033 1629 34075 1671
rect 34033 1609 34041 1629
rect 34061 1609 34075 1629
rect 34033 1571 34075 1609
rect 34125 1629 34169 1671
rect 34125 1609 34137 1629
rect 34157 1609 34169 1629
rect 34125 1571 34169 1609
rect 34251 1629 34293 1671
rect 34251 1609 34259 1629
rect 34279 1609 34293 1629
rect 34251 1571 34293 1609
rect 34343 1629 34387 1671
rect 34343 1609 34355 1629
rect 34375 1609 34387 1629
rect 34343 1571 34387 1609
rect 26406 1452 26450 1490
rect 26406 1432 26418 1452
rect 26438 1432 26450 1452
rect 20441 1343 20453 1363
rect 20473 1343 20485 1363
rect 20441 1305 20485 1343
rect 12609 1172 12621 1192
rect 12641 1172 12653 1192
rect 12609 1134 12653 1172
rect 16453 1205 16497 1247
rect 16453 1185 16465 1205
rect 16485 1185 16497 1205
rect 16453 1178 16497 1185
rect 16452 1147 16497 1178
rect 16547 1205 16589 1247
rect 16547 1185 16561 1205
rect 16581 1185 16589 1205
rect 16547 1147 16589 1185
rect 16663 1205 16705 1247
rect 16663 1185 16671 1205
rect 16691 1185 16705 1205
rect 16663 1147 16705 1185
rect 16755 1205 16799 1247
rect 16755 1185 16767 1205
rect 16787 1185 16799 1205
rect 16755 1147 16799 1185
rect 16881 1205 16923 1247
rect 16881 1185 16889 1205
rect 16909 1185 16923 1205
rect 16881 1147 16923 1185
rect 16973 1205 17017 1247
rect 18463 1243 18507 1281
rect 18463 1223 18475 1243
rect 18495 1223 18507 1243
rect 16973 1185 16985 1205
rect 17005 1185 17017 1205
rect 16973 1147 17017 1185
rect 18463 1181 18507 1223
rect 18557 1243 18599 1281
rect 18557 1223 18571 1243
rect 18591 1223 18599 1243
rect 18557 1181 18599 1223
rect 18681 1243 18725 1281
rect 18681 1223 18693 1243
rect 18713 1223 18725 1243
rect 18681 1181 18725 1223
rect 18775 1243 18817 1281
rect 18775 1223 18789 1243
rect 18809 1223 18817 1243
rect 18775 1181 18817 1223
rect 18891 1243 18933 1281
rect 18891 1223 18899 1243
rect 18919 1223 18933 1243
rect 18891 1181 18933 1223
rect 18983 1250 19028 1281
rect 18983 1243 19027 1250
rect 18983 1223 18995 1243
rect 19015 1223 19027 1243
rect 18983 1181 19027 1223
rect 24285 1376 24329 1418
rect 24285 1356 24297 1376
rect 24317 1356 24329 1376
rect 24285 1349 24329 1356
rect 24284 1318 24329 1349
rect 24379 1376 24421 1418
rect 24379 1356 24393 1376
rect 24413 1356 24421 1376
rect 24379 1318 24421 1356
rect 24495 1376 24537 1418
rect 24495 1356 24503 1376
rect 24523 1356 24537 1376
rect 24495 1318 24537 1356
rect 24587 1376 24631 1418
rect 24587 1356 24599 1376
rect 24619 1356 24631 1376
rect 24587 1318 24631 1356
rect 24713 1376 24755 1418
rect 24713 1356 24721 1376
rect 24741 1356 24755 1376
rect 24713 1318 24755 1356
rect 24805 1376 24849 1418
rect 26406 1390 26450 1432
rect 26500 1452 26542 1490
rect 26500 1432 26514 1452
rect 26534 1432 26542 1452
rect 26500 1390 26542 1432
rect 26624 1452 26668 1490
rect 26624 1432 26636 1452
rect 26656 1432 26668 1452
rect 26624 1390 26668 1432
rect 26718 1452 26760 1490
rect 26718 1432 26732 1452
rect 26752 1432 26760 1452
rect 26718 1390 26760 1432
rect 26834 1452 26876 1490
rect 26834 1432 26842 1452
rect 26862 1432 26876 1452
rect 26834 1390 26876 1432
rect 26926 1459 26971 1490
rect 26926 1452 26970 1459
rect 26926 1432 26938 1452
rect 26958 1432 26970 1452
rect 26926 1390 26970 1432
rect 30770 1465 30814 1503
rect 30770 1445 30782 1465
rect 30802 1445 30814 1465
rect 24805 1356 24817 1376
rect 24837 1356 24849 1376
rect 24805 1318 24849 1356
rect 22827 1256 22871 1294
rect 22827 1236 22839 1256
rect 22859 1236 22871 1256
rect 295 1003 339 1041
rect 295 983 307 1003
rect 327 983 339 1003
rect 295 941 339 983
rect 389 1003 431 1041
rect 389 983 403 1003
rect 423 983 431 1003
rect 389 941 431 983
rect 513 1003 557 1041
rect 513 983 525 1003
rect 545 983 557 1003
rect 513 941 557 983
rect 607 1003 649 1041
rect 607 983 621 1003
rect 641 983 649 1003
rect 607 941 649 983
rect 723 1003 765 1041
rect 723 983 731 1003
rect 751 983 765 1003
rect 723 941 765 983
rect 815 1010 860 1041
rect 815 1003 859 1010
rect 815 983 827 1003
rect 847 983 859 1003
rect 815 941 859 983
rect 4659 1016 4703 1054
rect 4659 996 4671 1016
rect 4691 996 4703 1016
rect 4659 954 4703 996
rect 4753 1016 4795 1054
rect 4753 996 4767 1016
rect 4787 996 4795 1016
rect 4753 954 4795 996
rect 4877 1016 4921 1054
rect 4877 996 4889 1016
rect 4909 996 4921 1016
rect 4877 954 4921 996
rect 4971 1016 5013 1054
rect 4971 996 4985 1016
rect 5005 996 5013 1016
rect 4971 954 5013 996
rect 5087 1016 5129 1054
rect 5087 996 5095 1016
rect 5115 996 5129 1016
rect 5087 954 5129 996
rect 5179 1023 5224 1054
rect 5179 1016 5223 1023
rect 5179 996 5191 1016
rect 5211 996 5223 1016
rect 5179 954 5223 996
rect 9036 1028 9080 1066
rect 9036 1008 9048 1028
rect 9068 1008 9080 1028
rect 9036 966 9080 1008
rect 9130 1028 9172 1066
rect 9130 1008 9144 1028
rect 9164 1008 9172 1028
rect 9130 966 9172 1008
rect 9254 1028 9298 1066
rect 9254 1008 9266 1028
rect 9286 1008 9298 1028
rect 9254 966 9298 1008
rect 9348 1028 9390 1066
rect 9348 1008 9362 1028
rect 9382 1008 9390 1028
rect 9348 966 9390 1008
rect 9464 1028 9506 1066
rect 9464 1008 9472 1028
rect 9492 1008 9506 1028
rect 9464 966 9506 1008
rect 9556 1035 9601 1066
rect 20719 1179 20763 1221
rect 20719 1159 20731 1179
rect 20751 1159 20763 1179
rect 20719 1152 20763 1159
rect 20718 1121 20763 1152
rect 20813 1179 20855 1221
rect 20813 1159 20827 1179
rect 20847 1159 20855 1179
rect 20813 1121 20855 1159
rect 20929 1179 20971 1221
rect 20929 1159 20937 1179
rect 20957 1159 20971 1179
rect 20929 1121 20971 1159
rect 21021 1179 21065 1221
rect 21021 1159 21033 1179
rect 21053 1159 21065 1179
rect 21021 1121 21065 1159
rect 21147 1179 21189 1221
rect 21147 1159 21155 1179
rect 21175 1159 21189 1179
rect 21147 1121 21189 1159
rect 21239 1179 21283 1221
rect 22827 1194 22871 1236
rect 22921 1256 22963 1294
rect 22921 1236 22935 1256
rect 22955 1236 22963 1256
rect 22921 1194 22963 1236
rect 23045 1256 23089 1294
rect 23045 1236 23057 1256
rect 23077 1236 23089 1256
rect 23045 1194 23089 1236
rect 23139 1256 23181 1294
rect 23139 1236 23153 1256
rect 23173 1236 23181 1256
rect 23139 1194 23181 1236
rect 23255 1256 23297 1294
rect 23255 1236 23263 1256
rect 23283 1236 23297 1256
rect 23255 1194 23297 1236
rect 23347 1263 23392 1294
rect 23347 1256 23391 1263
rect 23347 1236 23359 1256
rect 23379 1236 23391 1256
rect 23347 1194 23391 1236
rect 28662 1388 28706 1430
rect 28662 1368 28674 1388
rect 28694 1368 28706 1388
rect 28662 1361 28706 1368
rect 28661 1330 28706 1361
rect 28756 1388 28798 1430
rect 28756 1368 28770 1388
rect 28790 1368 28798 1388
rect 28756 1330 28798 1368
rect 28872 1388 28914 1430
rect 28872 1368 28880 1388
rect 28900 1368 28914 1388
rect 28872 1330 28914 1368
rect 28964 1388 29008 1430
rect 28964 1368 28976 1388
rect 28996 1368 29008 1388
rect 28964 1330 29008 1368
rect 29090 1388 29132 1430
rect 29090 1368 29098 1388
rect 29118 1368 29132 1388
rect 29090 1330 29132 1368
rect 29182 1388 29226 1430
rect 30770 1403 30814 1445
rect 30864 1465 30906 1503
rect 30864 1445 30878 1465
rect 30898 1445 30906 1465
rect 30864 1403 30906 1445
rect 30988 1465 31032 1503
rect 30988 1445 31000 1465
rect 31020 1445 31032 1465
rect 30988 1403 31032 1445
rect 31082 1465 31124 1503
rect 31082 1445 31096 1465
rect 31116 1445 31124 1465
rect 31082 1403 31124 1445
rect 31198 1465 31240 1503
rect 31198 1445 31206 1465
rect 31226 1445 31240 1465
rect 31198 1403 31240 1445
rect 31290 1472 31335 1503
rect 31290 1465 31334 1472
rect 31290 1445 31302 1465
rect 31322 1445 31334 1465
rect 31290 1403 31334 1445
rect 29182 1368 29194 1388
rect 29214 1368 29226 1388
rect 29182 1330 29226 1368
rect 27204 1268 27248 1306
rect 27204 1248 27216 1268
rect 27236 1248 27248 1268
rect 21239 1159 21251 1179
rect 21271 1159 21283 1179
rect 21239 1121 21283 1159
rect 25083 1192 25127 1234
rect 25083 1172 25095 1192
rect 25115 1172 25127 1192
rect 25083 1165 25127 1172
rect 25082 1134 25127 1165
rect 25177 1192 25219 1234
rect 25177 1172 25191 1192
rect 25211 1172 25219 1192
rect 25177 1134 25219 1172
rect 25293 1192 25335 1234
rect 25293 1172 25301 1192
rect 25321 1172 25335 1192
rect 25293 1134 25335 1172
rect 25385 1192 25429 1234
rect 25385 1172 25397 1192
rect 25417 1172 25429 1192
rect 25385 1134 25429 1172
rect 25511 1192 25553 1234
rect 25511 1172 25519 1192
rect 25539 1172 25553 1192
rect 25511 1134 25553 1172
rect 25603 1192 25647 1234
rect 27204 1206 27248 1248
rect 27298 1268 27340 1306
rect 27298 1248 27312 1268
rect 27332 1248 27340 1268
rect 27298 1206 27340 1248
rect 27422 1268 27466 1306
rect 27422 1248 27434 1268
rect 27454 1248 27466 1268
rect 27422 1206 27466 1248
rect 27516 1268 27558 1306
rect 27516 1248 27530 1268
rect 27550 1248 27558 1268
rect 27516 1206 27558 1248
rect 27632 1268 27674 1306
rect 27632 1248 27640 1268
rect 27660 1248 27674 1268
rect 27632 1206 27674 1248
rect 27724 1275 27769 1306
rect 27724 1268 27768 1275
rect 27724 1248 27736 1268
rect 27756 1248 27768 1268
rect 27724 1206 27768 1248
rect 33026 1401 33070 1443
rect 33026 1381 33038 1401
rect 33058 1381 33070 1401
rect 33026 1374 33070 1381
rect 33025 1343 33070 1374
rect 33120 1401 33162 1443
rect 33120 1381 33134 1401
rect 33154 1381 33162 1401
rect 33120 1343 33162 1381
rect 33236 1401 33278 1443
rect 33236 1381 33244 1401
rect 33264 1381 33278 1401
rect 33236 1343 33278 1381
rect 33328 1401 33372 1443
rect 33328 1381 33340 1401
rect 33360 1381 33372 1401
rect 33328 1343 33372 1381
rect 33454 1401 33496 1443
rect 33454 1381 33462 1401
rect 33482 1381 33496 1401
rect 33454 1343 33496 1381
rect 33546 1401 33590 1443
rect 33546 1381 33558 1401
rect 33578 1381 33590 1401
rect 33546 1343 33590 1381
rect 31568 1281 31612 1319
rect 31568 1261 31580 1281
rect 31600 1261 31612 1281
rect 25603 1172 25615 1192
rect 25635 1172 25647 1192
rect 25603 1134 25647 1172
rect 29460 1204 29504 1246
rect 29460 1184 29472 1204
rect 29492 1184 29504 1204
rect 29460 1177 29504 1184
rect 29459 1146 29504 1177
rect 29554 1204 29596 1246
rect 29554 1184 29568 1204
rect 29588 1184 29596 1204
rect 29554 1146 29596 1184
rect 29670 1204 29712 1246
rect 29670 1184 29678 1204
rect 29698 1184 29712 1204
rect 29670 1146 29712 1184
rect 29762 1204 29806 1246
rect 29762 1184 29774 1204
rect 29794 1184 29806 1204
rect 29762 1146 29806 1184
rect 29888 1204 29930 1246
rect 29888 1184 29896 1204
rect 29916 1184 29930 1204
rect 29888 1146 29930 1184
rect 29980 1204 30024 1246
rect 31568 1219 31612 1261
rect 31662 1281 31704 1319
rect 31662 1261 31676 1281
rect 31696 1261 31704 1281
rect 31662 1219 31704 1261
rect 31786 1281 31830 1319
rect 31786 1261 31798 1281
rect 31818 1261 31830 1281
rect 31786 1219 31830 1261
rect 31880 1281 31922 1319
rect 31880 1261 31894 1281
rect 31914 1261 31922 1281
rect 31880 1219 31922 1261
rect 31996 1281 32038 1319
rect 31996 1261 32004 1281
rect 32024 1261 32038 1281
rect 31996 1219 32038 1261
rect 32088 1288 32133 1319
rect 32088 1281 32132 1288
rect 32088 1261 32100 1281
rect 32120 1261 32132 1281
rect 32088 1219 32132 1261
rect 29980 1184 29992 1204
rect 30012 1184 30024 1204
rect 29980 1146 30024 1184
rect 33824 1217 33868 1259
rect 33824 1197 33836 1217
rect 33856 1197 33868 1217
rect 33824 1190 33868 1197
rect 33823 1159 33868 1190
rect 33918 1217 33960 1259
rect 33918 1197 33932 1217
rect 33952 1197 33960 1217
rect 33918 1159 33960 1197
rect 34034 1217 34076 1259
rect 34034 1197 34042 1217
rect 34062 1197 34076 1217
rect 34034 1159 34076 1197
rect 34126 1217 34170 1259
rect 34126 1197 34138 1217
rect 34158 1197 34170 1217
rect 34126 1159 34170 1197
rect 34252 1217 34294 1259
rect 34252 1197 34260 1217
rect 34280 1197 34294 1217
rect 34252 1159 34294 1197
rect 34344 1217 34388 1259
rect 34344 1197 34356 1217
rect 34376 1197 34388 1217
rect 34344 1159 34388 1197
rect 9556 1028 9600 1035
rect 9556 1008 9568 1028
rect 9588 1008 9600 1028
rect 9556 966 9600 1008
rect 13400 1041 13444 1079
rect 13400 1021 13412 1041
rect 13432 1021 13444 1041
rect 13400 979 13444 1021
rect 13494 1041 13536 1079
rect 13494 1021 13508 1041
rect 13528 1021 13536 1041
rect 13494 979 13536 1021
rect 13618 1041 13662 1079
rect 13618 1021 13630 1041
rect 13650 1021 13662 1041
rect 13618 979 13662 1021
rect 13712 1041 13754 1079
rect 13712 1021 13726 1041
rect 13746 1021 13754 1041
rect 13712 979 13754 1021
rect 13828 1041 13870 1079
rect 13828 1021 13836 1041
rect 13856 1021 13870 1041
rect 13828 979 13870 1021
rect 13920 1048 13965 1079
rect 13920 1041 13964 1048
rect 13920 1021 13932 1041
rect 13952 1021 13964 1041
rect 13920 979 13964 1021
rect 17666 1015 17710 1053
rect 17666 995 17678 1015
rect 17698 995 17710 1015
rect 17666 953 17710 995
rect 17760 1015 17802 1053
rect 17760 995 17774 1015
rect 17794 995 17802 1015
rect 17760 953 17802 995
rect 17884 1015 17928 1053
rect 17884 995 17896 1015
rect 17916 995 17928 1015
rect 17884 953 17928 995
rect 17978 1015 18020 1053
rect 17978 995 17992 1015
rect 18012 995 18020 1015
rect 17978 953 18020 995
rect 18094 1015 18136 1053
rect 18094 995 18102 1015
rect 18122 995 18136 1015
rect 18094 953 18136 995
rect 18186 1022 18231 1053
rect 18186 1015 18230 1022
rect 18186 995 18198 1015
rect 18218 995 18230 1015
rect 18186 953 18230 995
rect 22030 1028 22074 1066
rect 22030 1008 22042 1028
rect 22062 1008 22074 1028
rect 22030 966 22074 1008
rect 22124 1028 22166 1066
rect 22124 1008 22138 1028
rect 22158 1008 22166 1028
rect 22124 966 22166 1008
rect 22248 1028 22292 1066
rect 22248 1008 22260 1028
rect 22280 1008 22292 1028
rect 22248 966 22292 1008
rect 22342 1028 22384 1066
rect 22342 1008 22356 1028
rect 22376 1008 22384 1028
rect 22342 966 22384 1008
rect 22458 1028 22500 1066
rect 22458 1008 22466 1028
rect 22486 1008 22500 1028
rect 22458 966 22500 1008
rect 22550 1035 22595 1066
rect 22550 1028 22594 1035
rect 22550 1008 22562 1028
rect 22582 1008 22594 1028
rect 22550 966 22594 1008
rect 26407 1040 26451 1078
rect 26407 1020 26419 1040
rect 26439 1020 26451 1040
rect 26407 978 26451 1020
rect 26501 1040 26543 1078
rect 26501 1020 26515 1040
rect 26535 1020 26543 1040
rect 26501 978 26543 1020
rect 26625 1040 26669 1078
rect 26625 1020 26637 1040
rect 26657 1020 26669 1040
rect 26625 978 26669 1020
rect 26719 1040 26761 1078
rect 26719 1020 26733 1040
rect 26753 1020 26761 1040
rect 26719 978 26761 1020
rect 26835 1040 26877 1078
rect 26835 1020 26843 1040
rect 26863 1020 26877 1040
rect 26835 978 26877 1020
rect 26927 1047 26972 1078
rect 26927 1040 26971 1047
rect 26927 1020 26939 1040
rect 26959 1020 26971 1040
rect 26927 978 26971 1020
rect 30771 1053 30815 1091
rect 30771 1033 30783 1053
rect 30803 1033 30815 1053
rect 30771 991 30815 1033
rect 30865 1053 30907 1091
rect 30865 1033 30879 1053
rect 30899 1033 30907 1053
rect 30865 991 30907 1033
rect 30989 1053 31033 1091
rect 30989 1033 31001 1053
rect 31021 1033 31033 1053
rect 30989 991 31033 1033
rect 31083 1053 31125 1091
rect 31083 1033 31097 1053
rect 31117 1033 31125 1053
rect 31083 991 31125 1033
rect 31199 1053 31241 1091
rect 31199 1033 31207 1053
rect 31227 1033 31241 1053
rect 31199 991 31241 1033
rect 31291 1060 31336 1091
rect 31291 1053 31335 1060
rect 31291 1033 31303 1053
rect 31323 1033 31335 1053
rect 31291 991 31335 1033
rect 1508 427 1552 465
rect 1508 407 1520 427
rect 1540 407 1552 427
rect 1508 365 1552 407
rect 1602 427 1644 465
rect 1602 407 1616 427
rect 1636 407 1644 427
rect 1602 365 1644 407
rect 1726 427 1770 465
rect 1726 407 1738 427
rect 1758 407 1770 427
rect 1726 365 1770 407
rect 1820 427 1862 465
rect 1820 407 1834 427
rect 1854 407 1862 427
rect 1820 365 1862 407
rect 1936 427 1978 465
rect 1936 407 1944 427
rect 1964 407 1978 427
rect 1936 365 1978 407
rect 2028 434 2073 465
rect 5872 440 5916 478
rect 2028 427 2072 434
rect 2028 407 2040 427
rect 2060 407 2072 427
rect 2028 365 2072 407
rect 5872 420 5884 440
rect 5904 420 5916 440
rect 3997 353 4041 391
rect 3997 333 4009 353
rect 4029 333 4041 353
rect 3997 291 4041 333
rect 4091 353 4133 391
rect 4091 333 4105 353
rect 4125 333 4133 353
rect 4091 291 4133 333
rect 4215 353 4259 391
rect 4215 333 4227 353
rect 4247 333 4259 353
rect 4215 291 4259 333
rect 4309 353 4351 391
rect 4309 333 4323 353
rect 4343 333 4351 353
rect 4309 291 4351 333
rect 4425 353 4467 391
rect 4425 333 4433 353
rect 4453 333 4467 353
rect 4425 291 4467 333
rect 4517 360 4562 391
rect 5872 378 5916 420
rect 5966 440 6008 478
rect 5966 420 5980 440
rect 6000 420 6008 440
rect 5966 378 6008 420
rect 6090 440 6134 478
rect 6090 420 6102 440
rect 6122 420 6134 440
rect 6090 378 6134 420
rect 6184 440 6226 478
rect 6184 420 6198 440
rect 6218 420 6226 440
rect 6184 378 6226 420
rect 6300 440 6342 478
rect 6300 420 6308 440
rect 6328 420 6342 440
rect 6300 378 6342 420
rect 6392 447 6437 478
rect 10249 452 10293 490
rect 6392 440 6436 447
rect 6392 420 6404 440
rect 6424 420 6436 440
rect 10249 432 10261 452
rect 10281 432 10293 452
rect 6392 378 6436 420
rect 4517 353 4561 360
rect 4517 333 4529 353
rect 4549 333 4561 353
rect 4517 291 4561 333
rect 8445 377 8489 415
rect 8445 357 8457 377
rect 8477 357 8489 377
rect 8445 315 8489 357
rect 8539 377 8581 415
rect 8539 357 8553 377
rect 8573 357 8581 377
rect 8539 315 8581 357
rect 8663 377 8707 415
rect 8663 357 8675 377
rect 8695 357 8707 377
rect 8663 315 8707 357
rect 8757 377 8799 415
rect 8757 357 8771 377
rect 8791 357 8799 377
rect 8757 315 8799 357
rect 8873 377 8915 415
rect 8873 357 8881 377
rect 8901 357 8915 377
rect 8873 315 8915 357
rect 8965 384 9010 415
rect 10249 390 10293 432
rect 10343 452 10385 490
rect 10343 432 10357 452
rect 10377 432 10385 452
rect 10343 390 10385 432
rect 10467 452 10511 490
rect 10467 432 10479 452
rect 10499 432 10511 452
rect 10467 390 10511 432
rect 10561 452 10603 490
rect 10561 432 10575 452
rect 10595 432 10603 452
rect 10561 390 10603 432
rect 10677 452 10719 490
rect 10677 432 10685 452
rect 10705 432 10719 452
rect 10677 390 10719 432
rect 10769 459 10814 490
rect 14613 465 14657 503
rect 10769 452 10813 459
rect 10769 432 10781 452
rect 10801 432 10813 452
rect 10769 390 10813 432
rect 14613 445 14625 465
rect 14645 445 14657 465
rect 8965 377 9009 384
rect 8965 357 8977 377
rect 8997 357 9009 377
rect 8965 315 9009 357
rect 12738 378 12782 416
rect 12738 358 12750 378
rect 12770 358 12782 378
rect 12738 316 12782 358
rect 12832 378 12874 416
rect 12832 358 12846 378
rect 12866 358 12874 378
rect 12832 316 12874 358
rect 12956 378 13000 416
rect 12956 358 12968 378
rect 12988 358 13000 378
rect 12956 316 13000 358
rect 13050 378 13092 416
rect 13050 358 13064 378
rect 13084 358 13092 378
rect 13050 316 13092 358
rect 13166 378 13208 416
rect 13166 358 13174 378
rect 13194 358 13208 378
rect 13166 316 13208 358
rect 13258 385 13303 416
rect 14613 403 14657 445
rect 14707 465 14749 503
rect 14707 445 14721 465
rect 14741 445 14749 465
rect 14707 403 14749 445
rect 14831 465 14875 503
rect 14831 445 14843 465
rect 14863 445 14875 465
rect 14831 403 14875 445
rect 14925 465 14967 503
rect 14925 445 14939 465
rect 14959 445 14967 465
rect 14925 403 14967 445
rect 15041 465 15083 503
rect 15041 445 15049 465
rect 15069 445 15083 465
rect 15041 403 15083 445
rect 15133 472 15178 503
rect 15133 465 15177 472
rect 15133 445 15145 465
rect 15165 445 15177 465
rect 15133 403 15177 445
rect 18879 439 18923 477
rect 18879 419 18891 439
rect 18911 419 18923 439
rect 13258 378 13302 385
rect 13258 358 13270 378
rect 13290 358 13302 378
rect 13258 316 13302 358
rect 18879 377 18923 419
rect 18973 439 19015 477
rect 18973 419 18987 439
rect 19007 419 19015 439
rect 18973 377 19015 419
rect 19097 439 19141 477
rect 19097 419 19109 439
rect 19129 419 19141 439
rect 19097 377 19141 419
rect 19191 439 19233 477
rect 19191 419 19205 439
rect 19225 419 19233 439
rect 19191 377 19233 419
rect 19307 439 19349 477
rect 19307 419 19315 439
rect 19335 419 19349 439
rect 19307 377 19349 419
rect 19399 446 19444 477
rect 23243 452 23287 490
rect 19399 439 19443 446
rect 19399 419 19411 439
rect 19431 419 19443 439
rect 19399 377 19443 419
rect 23243 432 23255 452
rect 23275 432 23287 452
rect 16935 314 16979 352
rect 16935 294 16947 314
rect 16967 294 16979 314
rect 16935 252 16979 294
rect 17029 314 17071 352
rect 17029 294 17043 314
rect 17063 294 17071 314
rect 17029 252 17071 294
rect 17153 314 17197 352
rect 17153 294 17165 314
rect 17185 294 17197 314
rect 17153 252 17197 294
rect 17247 314 17289 352
rect 17247 294 17261 314
rect 17281 294 17289 314
rect 17247 252 17289 294
rect 17363 314 17405 352
rect 17363 294 17371 314
rect 17391 294 17405 314
rect 17363 252 17405 294
rect 17455 321 17500 352
rect 17455 314 17499 321
rect 17455 294 17467 314
rect 17487 294 17499 314
rect 21368 365 21412 403
rect 21368 345 21380 365
rect 21400 345 21412 365
rect 21368 303 21412 345
rect 21462 365 21504 403
rect 21462 345 21476 365
rect 21496 345 21504 365
rect 21462 303 21504 345
rect 21586 365 21630 403
rect 21586 345 21598 365
rect 21618 345 21630 365
rect 21586 303 21630 345
rect 21680 365 21722 403
rect 21680 345 21694 365
rect 21714 345 21722 365
rect 21680 303 21722 345
rect 21796 365 21838 403
rect 21796 345 21804 365
rect 21824 345 21838 365
rect 21796 303 21838 345
rect 21888 372 21933 403
rect 23243 390 23287 432
rect 23337 452 23379 490
rect 23337 432 23351 452
rect 23371 432 23379 452
rect 23337 390 23379 432
rect 23461 452 23505 490
rect 23461 432 23473 452
rect 23493 432 23505 452
rect 23461 390 23505 432
rect 23555 452 23597 490
rect 23555 432 23569 452
rect 23589 432 23597 452
rect 23555 390 23597 432
rect 23671 452 23713 490
rect 23671 432 23679 452
rect 23699 432 23713 452
rect 23671 390 23713 432
rect 23763 459 23808 490
rect 27620 464 27664 502
rect 23763 452 23807 459
rect 23763 432 23775 452
rect 23795 432 23807 452
rect 27620 444 27632 464
rect 27652 444 27664 464
rect 23763 390 23807 432
rect 21888 365 21932 372
rect 21888 345 21900 365
rect 21920 345 21932 365
rect 21888 303 21932 345
rect 25816 389 25860 427
rect 25816 369 25828 389
rect 25848 369 25860 389
rect 25816 327 25860 369
rect 25910 389 25952 427
rect 25910 369 25924 389
rect 25944 369 25952 389
rect 25910 327 25952 369
rect 26034 389 26078 427
rect 26034 369 26046 389
rect 26066 369 26078 389
rect 26034 327 26078 369
rect 26128 389 26170 427
rect 26128 369 26142 389
rect 26162 369 26170 389
rect 26128 327 26170 369
rect 26244 389 26286 427
rect 26244 369 26252 389
rect 26272 369 26286 389
rect 26244 327 26286 369
rect 26336 396 26381 427
rect 27620 402 27664 444
rect 27714 464 27756 502
rect 27714 444 27728 464
rect 27748 444 27756 464
rect 27714 402 27756 444
rect 27838 464 27882 502
rect 27838 444 27850 464
rect 27870 444 27882 464
rect 27838 402 27882 444
rect 27932 464 27974 502
rect 27932 444 27946 464
rect 27966 444 27974 464
rect 27932 402 27974 444
rect 28048 464 28090 502
rect 28048 444 28056 464
rect 28076 444 28090 464
rect 28048 402 28090 444
rect 28140 471 28185 502
rect 31984 477 32028 515
rect 28140 464 28184 471
rect 28140 444 28152 464
rect 28172 444 28184 464
rect 28140 402 28184 444
rect 31984 457 31996 477
rect 32016 457 32028 477
rect 26336 389 26380 396
rect 26336 369 26348 389
rect 26368 369 26380 389
rect 26336 327 26380 369
rect 17455 252 17499 294
rect 30109 390 30153 428
rect 30109 370 30121 390
rect 30141 370 30153 390
rect 30109 328 30153 370
rect 30203 390 30245 428
rect 30203 370 30217 390
rect 30237 370 30245 390
rect 30203 328 30245 370
rect 30327 390 30371 428
rect 30327 370 30339 390
rect 30359 370 30371 390
rect 30327 328 30371 370
rect 30421 390 30463 428
rect 30421 370 30435 390
rect 30455 370 30463 390
rect 30421 328 30463 370
rect 30537 390 30579 428
rect 30537 370 30545 390
rect 30565 370 30579 390
rect 30537 328 30579 370
rect 30629 397 30674 428
rect 31984 415 32028 457
rect 32078 477 32120 515
rect 32078 457 32092 477
rect 32112 457 32120 477
rect 32078 415 32120 457
rect 32202 477 32246 515
rect 32202 457 32214 477
rect 32234 457 32246 477
rect 32202 415 32246 457
rect 32296 477 32338 515
rect 32296 457 32310 477
rect 32330 457 32338 477
rect 32296 415 32338 457
rect 32412 477 32454 515
rect 32412 457 32420 477
rect 32440 457 32454 477
rect 32412 415 32454 457
rect 32504 484 32549 515
rect 32504 477 32548 484
rect 32504 457 32516 477
rect 32536 457 32548 477
rect 32504 415 32548 457
rect 30629 390 30673 397
rect 30629 370 30641 390
rect 30661 370 30673 390
rect 30629 328 30673 370
<< ndiffc >>
rect 3480 8834 3500 8854
rect 3583 8830 3603 8850
rect 3691 8830 3711 8850
rect 3794 8834 3814 8854
rect 3909 8830 3929 8850
rect 4012 8834 4032 8854
rect 4199 8841 4217 8859
rect 263 8779 281 8797
rect 7844 8847 7864 8867
rect 7947 8843 7967 8863
rect 8055 8843 8075 8863
rect 8158 8847 8178 8867
rect 8273 8843 8293 8863
rect 8376 8847 8396 8867
rect 8563 8854 8581 8872
rect 4627 8792 4645 8810
rect 261 8680 279 8698
rect 4197 8742 4215 8760
rect 12221 8859 12241 8879
rect 12324 8855 12344 8875
rect 12432 8855 12452 8875
rect 12535 8859 12555 8879
rect 12650 8855 12670 8875
rect 12753 8859 12773 8879
rect 12940 8866 12958 8884
rect 9004 8804 9022 8822
rect 4625 8693 4643 8711
rect 2683 8606 2703 8626
rect 2786 8602 2806 8622
rect 2894 8602 2914 8622
rect 2997 8606 3017 8626
rect 3112 8602 3132 8622
rect 8561 8755 8579 8773
rect 16585 8872 16605 8892
rect 16688 8868 16708 8888
rect 16796 8868 16816 8888
rect 16899 8872 16919 8892
rect 17014 8868 17034 8888
rect 17117 8872 17137 8892
rect 17304 8879 17322 8897
rect 13368 8817 13386 8835
rect 9002 8705 9020 8723
rect 3215 8606 3235 8626
rect 4192 8623 4210 8641
rect 7047 8619 7067 8639
rect 7150 8615 7170 8635
rect 7258 8615 7278 8635
rect 7361 8619 7381 8639
rect 7476 8615 7496 8635
rect 12938 8767 12956 8785
rect 20851 8846 20871 8866
rect 20954 8842 20974 8862
rect 21062 8842 21082 8862
rect 21165 8846 21185 8866
rect 21280 8842 21300 8862
rect 21383 8846 21403 8866
rect 21570 8853 21588 8871
rect 13366 8718 13384 8736
rect 7579 8619 7599 8639
rect 8556 8636 8574 8654
rect 11424 8631 11444 8651
rect 11527 8627 11547 8647
rect 11635 8627 11655 8647
rect 11738 8631 11758 8651
rect 11853 8627 11873 8647
rect 17302 8780 17320 8798
rect 17634 8791 17652 8809
rect 25215 8859 25235 8879
rect 25318 8855 25338 8875
rect 25426 8855 25446 8875
rect 25529 8859 25549 8879
rect 25644 8855 25664 8875
rect 25747 8859 25767 8879
rect 25934 8866 25952 8884
rect 21998 8804 22016 8822
rect 11956 8631 11976 8651
rect 12933 8648 12951 8666
rect 15788 8644 15808 8664
rect 15891 8640 15911 8660
rect 15999 8640 16019 8660
rect 16102 8644 16122 8664
rect 16217 8640 16237 8660
rect 16320 8644 16340 8664
rect 17297 8661 17315 8679
rect 17632 8692 17650 8710
rect 21568 8754 21586 8772
rect 29592 8871 29612 8891
rect 29695 8867 29715 8887
rect 29803 8867 29823 8887
rect 29906 8871 29926 8891
rect 30021 8867 30041 8887
rect 30124 8871 30144 8891
rect 30311 8878 30329 8896
rect 26375 8816 26393 8834
rect 21996 8705 22014 8723
rect 4190 8524 4208 8542
rect 258 8455 276 8473
rect 8554 8537 8572 8555
rect 3481 8422 3501 8442
rect 256 8356 274 8374
rect 427 8372 447 8392
rect 530 8376 550 8396
rect 645 8372 665 8392
rect 748 8376 768 8396
rect 856 8376 876 8396
rect 3584 8418 3604 8438
rect 3692 8418 3712 8438
rect 3795 8422 3815 8442
rect 3910 8418 3930 8438
rect 4013 8422 4033 8442
rect 4186 8440 4204 8458
rect 4622 8468 4640 8486
rect 959 8372 979 8392
rect 12931 8549 12949 8567
rect 7845 8435 7865 8455
rect 4184 8341 4202 8359
rect 4620 8369 4638 8387
rect 4791 8385 4811 8405
rect 4894 8389 4914 8409
rect 5009 8385 5029 8405
rect 5112 8389 5132 8409
rect 5220 8389 5240 8409
rect 7948 8431 7968 8451
rect 8056 8431 8076 8451
rect 8159 8435 8179 8455
rect 8274 8431 8294 8451
rect 8377 8435 8397 8455
rect 8550 8453 8568 8471
rect 8999 8480 9017 8498
rect 5323 8385 5343 8405
rect 252 8272 270 8290
rect 20054 8618 20074 8638
rect 20157 8614 20177 8634
rect 20265 8614 20285 8634
rect 20368 8618 20388 8638
rect 20483 8614 20503 8634
rect 25932 8767 25950 8785
rect 33956 8884 33976 8904
rect 34059 8880 34079 8900
rect 34167 8880 34187 8900
rect 34270 8884 34290 8904
rect 34385 8880 34405 8900
rect 34488 8884 34508 8904
rect 34675 8891 34693 8909
rect 30739 8829 30757 8847
rect 26373 8717 26391 8735
rect 20586 8618 20606 8638
rect 21563 8635 21581 8653
rect 24418 8631 24438 8651
rect 24521 8627 24541 8647
rect 24629 8627 24649 8647
rect 24732 8631 24752 8651
rect 24847 8627 24867 8647
rect 30309 8779 30327 8797
rect 30737 8730 30755 8748
rect 24950 8631 24970 8651
rect 25927 8648 25945 8666
rect 28795 8643 28815 8663
rect 28898 8639 28918 8659
rect 29006 8639 29026 8659
rect 29109 8643 29129 8663
rect 29224 8639 29244 8659
rect 34673 8792 34691 8810
rect 29327 8643 29347 8663
rect 30304 8660 30322 8678
rect 33159 8656 33179 8676
rect 33262 8652 33282 8672
rect 33370 8652 33390 8672
rect 33473 8656 33493 8676
rect 33588 8652 33608 8672
rect 33691 8656 33711 8676
rect 34668 8673 34686 8691
rect 17295 8562 17313 8580
rect 12222 8447 12242 8467
rect 8548 8354 8566 8372
rect 8997 8381 9015 8399
rect 9168 8397 9188 8417
rect 9271 8401 9291 8421
rect 9386 8397 9406 8417
rect 9489 8401 9509 8421
rect 9597 8401 9617 8421
rect 12325 8443 12345 8463
rect 12433 8443 12453 8463
rect 12536 8447 12556 8467
rect 12651 8443 12671 8463
rect 12754 8447 12774 8467
rect 12927 8465 12945 8483
rect 13363 8493 13381 8511
rect 9700 8397 9720 8417
rect 4616 8285 4634 8303
rect 250 8173 268 8191
rect 1225 8188 1245 8208
rect 1328 8192 1348 8212
rect 1443 8188 1463 8208
rect 1546 8192 1566 8212
rect 1654 8192 1674 8212
rect 1757 8188 1777 8208
rect 2584 8196 2604 8216
rect 2687 8192 2707 8212
rect 2795 8192 2815 8212
rect 2898 8196 2918 8216
rect 3013 8192 3033 8212
rect 16586 8460 16606 8480
rect 12925 8366 12943 8384
rect 13361 8394 13379 8412
rect 13532 8410 13552 8430
rect 13635 8414 13655 8434
rect 13750 8410 13770 8430
rect 13853 8414 13873 8434
rect 13961 8414 13981 8434
rect 16689 8456 16709 8476
rect 16797 8456 16817 8476
rect 16900 8460 16920 8480
rect 17015 8456 17035 8476
rect 17118 8460 17138 8480
rect 17291 8478 17309 8496
rect 21561 8536 21579 8554
rect 14064 8410 14084 8430
rect 8993 8297 9011 8315
rect 3116 8196 3136 8216
rect 4614 8186 4632 8204
rect 5589 8201 5609 8221
rect 245 8054 263 8072
rect 5692 8205 5712 8225
rect 5807 8201 5827 8221
rect 5910 8205 5930 8225
rect 6018 8205 6038 8225
rect 6121 8201 6141 8221
rect 6948 8209 6968 8229
rect 7051 8205 7071 8225
rect 7159 8205 7179 8225
rect 7262 8209 7282 8229
rect 7377 8205 7397 8225
rect 17629 8467 17647 8485
rect 17289 8379 17307 8397
rect 25925 8549 25943 8567
rect 20852 8434 20872 8454
rect 13357 8310 13375 8328
rect 7480 8209 7500 8229
rect 4181 8116 4199 8134
rect 4609 8067 4627 8085
rect 8991 8198 9009 8216
rect 9966 8213 9986 8233
rect 10069 8217 10089 8237
rect 10184 8213 10204 8233
rect 10287 8217 10307 8237
rect 10395 8217 10415 8237
rect 10498 8213 10518 8233
rect 11325 8221 11345 8241
rect 11428 8217 11448 8237
rect 11536 8217 11556 8237
rect 11639 8221 11659 8241
rect 11754 8217 11774 8237
rect 17627 8368 17645 8386
rect 17798 8384 17818 8404
rect 17901 8388 17921 8408
rect 18016 8384 18036 8404
rect 18119 8388 18139 8408
rect 18227 8388 18247 8408
rect 20955 8430 20975 8450
rect 21063 8430 21083 8450
rect 21166 8434 21186 8454
rect 21281 8430 21301 8450
rect 21384 8434 21404 8454
rect 21557 8452 21575 8470
rect 21993 8480 22011 8498
rect 18330 8384 18350 8404
rect 30302 8561 30320 8579
rect 25216 8447 25236 8467
rect 21555 8353 21573 8371
rect 21991 8381 22009 8399
rect 22162 8397 22182 8417
rect 22265 8401 22285 8421
rect 22380 8397 22400 8417
rect 22483 8401 22503 8421
rect 22591 8401 22611 8421
rect 25319 8443 25339 8463
rect 25427 8443 25447 8463
rect 25530 8447 25550 8467
rect 25645 8443 25665 8463
rect 25748 8447 25768 8467
rect 25921 8465 25939 8483
rect 26370 8492 26388 8510
rect 22694 8397 22714 8417
rect 17623 8284 17641 8302
rect 11857 8221 11877 8241
rect 13355 8211 13373 8229
rect 14330 8226 14350 8246
rect 8545 8129 8563 8147
rect 4179 8017 4197 8035
rect 243 7955 261 7973
rect 428 7960 448 7980
rect 531 7964 551 7984
rect 646 7960 666 7980
rect 749 7964 769 7984
rect 857 7964 877 7984
rect 960 7960 980 7980
rect 8986 8079 9004 8097
rect 14433 8230 14453 8250
rect 14548 8226 14568 8246
rect 14651 8230 14671 8250
rect 14759 8230 14779 8250
rect 14862 8226 14882 8246
rect 15689 8234 15709 8254
rect 15792 8230 15812 8250
rect 15900 8230 15920 8250
rect 16003 8234 16023 8254
rect 16118 8230 16138 8250
rect 16221 8234 16241 8254
rect 34666 8574 34684 8592
rect 29593 8459 29613 8479
rect 25919 8366 25937 8384
rect 26368 8393 26386 8411
rect 26539 8409 26559 8429
rect 26642 8413 26662 8433
rect 26757 8409 26777 8429
rect 26860 8413 26880 8433
rect 26968 8413 26988 8433
rect 29696 8455 29716 8475
rect 29804 8455 29824 8475
rect 29907 8459 29927 8479
rect 30022 8455 30042 8475
rect 30125 8459 30145 8479
rect 30298 8477 30316 8495
rect 30734 8505 30752 8523
rect 27071 8409 27091 8429
rect 21987 8297 22005 8315
rect 12922 8141 12940 8159
rect 8543 8030 8561 8048
rect 4607 7968 4625 7986
rect 4792 7973 4812 7993
rect 4895 7977 4915 7997
rect 5010 7973 5030 7993
rect 5113 7977 5133 7997
rect 5221 7977 5241 7997
rect 5324 7973 5344 7993
rect 13350 8092 13368 8110
rect 17286 8154 17304 8172
rect 17621 8185 17639 8203
rect 18596 8200 18616 8220
rect 18699 8204 18719 8224
rect 18814 8200 18834 8220
rect 18917 8204 18937 8224
rect 19025 8204 19045 8224
rect 19128 8200 19148 8220
rect 19955 8208 19975 8228
rect 20058 8204 20078 8224
rect 20166 8204 20186 8224
rect 20269 8208 20289 8228
rect 20384 8204 20404 8224
rect 33957 8472 33977 8492
rect 30296 8378 30314 8396
rect 30732 8406 30750 8424
rect 30903 8422 30923 8442
rect 31006 8426 31026 8446
rect 31121 8422 31141 8442
rect 31224 8426 31244 8446
rect 31332 8426 31352 8446
rect 34060 8468 34080 8488
rect 34168 8468 34188 8488
rect 34271 8472 34291 8492
rect 34386 8468 34406 8488
rect 34489 8472 34509 8492
rect 34662 8490 34680 8508
rect 31435 8422 31455 8442
rect 26364 8309 26382 8327
rect 20487 8208 20507 8228
rect 21985 8198 22003 8216
rect 22960 8213 22980 8233
rect 12920 8042 12938 8060
rect 8984 7980 9002 7998
rect 9169 7985 9189 8005
rect 9272 7989 9292 8009
rect 9387 7985 9407 8005
rect 9490 7989 9510 8009
rect 9598 7989 9618 8009
rect 9701 7985 9721 8005
rect 17284 8055 17302 8073
rect 17616 8066 17634 8084
rect 23063 8217 23083 8237
rect 23178 8213 23198 8233
rect 23281 8217 23301 8237
rect 23389 8217 23409 8237
rect 23492 8213 23512 8233
rect 24319 8221 24339 8241
rect 24422 8217 24442 8237
rect 24530 8217 24550 8237
rect 24633 8221 24653 8241
rect 24748 8217 24768 8237
rect 34660 8391 34678 8409
rect 30728 8322 30746 8340
rect 24851 8221 24871 8241
rect 21552 8128 21570 8146
rect 13348 7993 13366 8011
rect 13533 7998 13553 8018
rect 13636 8002 13656 8022
rect 13751 7998 13771 8018
rect 13854 8002 13874 8022
rect 13962 8002 13982 8022
rect 14065 7998 14085 8018
rect 21980 8079 21998 8097
rect 26362 8210 26380 8228
rect 27337 8225 27357 8245
rect 27440 8229 27460 8249
rect 27555 8225 27575 8245
rect 27658 8229 27678 8249
rect 27766 8229 27786 8249
rect 27869 8225 27889 8245
rect 28696 8233 28716 8253
rect 28799 8229 28819 8249
rect 28907 8229 28927 8249
rect 29010 8233 29030 8253
rect 29125 8229 29145 8249
rect 29228 8233 29248 8253
rect 30726 8223 30744 8241
rect 31701 8238 31721 8258
rect 25916 8141 25934 8159
rect 21550 8029 21568 8047
rect 17614 7967 17632 7985
rect 17799 7972 17819 7992
rect 17902 7976 17922 7996
rect 18017 7972 18037 7992
rect 18120 7976 18140 7996
rect 18228 7976 18248 7996
rect 18331 7972 18351 7992
rect 26357 8091 26375 8109
rect 31804 8242 31824 8262
rect 31919 8238 31939 8258
rect 32022 8242 32042 8262
rect 32130 8242 32150 8262
rect 32233 8238 32253 8258
rect 33060 8246 33080 8266
rect 33163 8242 33183 8262
rect 33271 8242 33291 8262
rect 33374 8246 33394 8266
rect 33489 8242 33509 8262
rect 33592 8246 33612 8266
rect 30293 8153 30311 8171
rect 25914 8042 25932 8060
rect 21978 7980 21996 7998
rect 22163 7985 22183 8005
rect 22266 7989 22286 8009
rect 22381 7985 22401 8005
rect 22484 7989 22504 8009
rect 22592 7989 22612 8009
rect 22695 7985 22715 8005
rect 30721 8104 30739 8122
rect 34657 8166 34675 8184
rect 30291 8054 30309 8072
rect 26355 7992 26373 8010
rect 26540 7997 26560 8017
rect 26643 8001 26663 8021
rect 26758 7997 26778 8017
rect 26861 8001 26881 8021
rect 26969 8001 26989 8021
rect 27072 7997 27092 8017
rect 34655 8067 34673 8085
rect 30719 8005 30737 8023
rect 30904 8010 30924 8030
rect 31007 8014 31027 8034
rect 31122 8010 31142 8030
rect 31225 8014 31245 8034
rect 31333 8014 31353 8034
rect 31436 8010 31456 8030
rect 3463 7816 3483 7836
rect 3566 7812 3586 7832
rect 3674 7812 3694 7832
rect 3777 7816 3797 7836
rect 3892 7812 3912 7832
rect 3995 7816 4015 7836
rect 4182 7823 4200 7841
rect 246 7761 264 7779
rect 7827 7829 7847 7849
rect 7930 7825 7950 7845
rect 8038 7825 8058 7845
rect 8141 7829 8161 7849
rect 8256 7825 8276 7845
rect 8359 7829 8379 7849
rect 8546 7836 8564 7854
rect 4610 7774 4628 7792
rect 244 7662 262 7680
rect 4180 7724 4198 7742
rect 12204 7841 12224 7861
rect 12307 7837 12327 7857
rect 12415 7837 12435 7857
rect 12518 7841 12538 7861
rect 12633 7837 12653 7857
rect 12736 7841 12756 7861
rect 12923 7848 12941 7866
rect 8987 7786 9005 7804
rect 4608 7675 4626 7693
rect 1307 7580 1327 7600
rect 1410 7584 1430 7604
rect 1525 7580 1545 7600
rect 1628 7584 1648 7604
rect 1736 7584 1756 7604
rect 1839 7580 1859 7600
rect 2666 7588 2686 7608
rect 2769 7584 2789 7604
rect 2877 7584 2897 7604
rect 2980 7588 3000 7608
rect 3095 7584 3115 7604
rect 8544 7737 8562 7755
rect 16568 7854 16588 7874
rect 16671 7850 16691 7870
rect 16779 7850 16799 7870
rect 16882 7854 16902 7874
rect 16997 7850 17017 7870
rect 17100 7854 17120 7874
rect 17287 7861 17305 7879
rect 13351 7799 13369 7817
rect 8985 7687 9003 7705
rect 3198 7588 3218 7608
rect 4175 7605 4193 7623
rect 5671 7593 5691 7613
rect 5774 7597 5794 7617
rect 5889 7593 5909 7613
rect 5992 7597 6012 7617
rect 6100 7597 6120 7617
rect 6203 7593 6223 7613
rect 7030 7601 7050 7621
rect 7133 7597 7153 7617
rect 7241 7597 7261 7617
rect 7344 7601 7364 7621
rect 7459 7597 7479 7617
rect 7562 7601 7582 7621
rect 8539 7618 8557 7636
rect 12921 7749 12939 7767
rect 20834 7828 20854 7848
rect 20937 7824 20957 7844
rect 21045 7824 21065 7844
rect 21148 7828 21168 7848
rect 21263 7824 21283 7844
rect 21366 7828 21386 7848
rect 21553 7835 21571 7853
rect 13349 7700 13367 7718
rect 10048 7605 10068 7625
rect 4173 7506 4191 7524
rect 241 7437 259 7455
rect 10151 7609 10171 7629
rect 10266 7605 10286 7625
rect 10369 7609 10389 7629
rect 10477 7609 10497 7629
rect 10580 7605 10600 7625
rect 11407 7613 11427 7633
rect 11510 7609 11530 7629
rect 11618 7609 11638 7629
rect 11721 7613 11741 7633
rect 11836 7609 11856 7629
rect 17285 7762 17303 7780
rect 17617 7773 17635 7791
rect 25198 7841 25218 7861
rect 25301 7837 25321 7857
rect 25409 7837 25429 7857
rect 25512 7841 25532 7861
rect 25627 7837 25647 7857
rect 25730 7841 25750 7861
rect 25917 7848 25935 7866
rect 21981 7786 21999 7804
rect 11939 7613 11959 7633
rect 12916 7630 12934 7648
rect 14412 7618 14432 7638
rect 8537 7519 8555 7537
rect 3464 7404 3484 7424
rect 239 7338 257 7356
rect 410 7354 430 7374
rect 513 7358 533 7378
rect 628 7354 648 7374
rect 731 7358 751 7378
rect 839 7358 859 7378
rect 3567 7400 3587 7420
rect 3675 7400 3695 7420
rect 3778 7404 3798 7424
rect 3893 7400 3913 7420
rect 3996 7404 4016 7424
rect 4169 7422 4187 7440
rect 4605 7450 4623 7468
rect 942 7354 962 7374
rect 14515 7622 14535 7642
rect 14630 7618 14650 7638
rect 14733 7622 14753 7642
rect 14841 7622 14861 7642
rect 14944 7618 14964 7638
rect 15771 7626 15791 7646
rect 15874 7622 15894 7642
rect 15982 7622 16002 7642
rect 16085 7626 16105 7646
rect 16200 7622 16220 7642
rect 16303 7626 16323 7646
rect 17280 7643 17298 7661
rect 17615 7674 17633 7692
rect 21551 7736 21569 7754
rect 29575 7853 29595 7873
rect 29678 7849 29698 7869
rect 29786 7849 29806 7869
rect 29889 7853 29909 7873
rect 30004 7849 30024 7869
rect 30107 7853 30127 7873
rect 30294 7860 30312 7878
rect 26358 7798 26376 7816
rect 21979 7687 21997 7705
rect 12914 7531 12932 7549
rect 7828 7417 7848 7437
rect 4167 7323 4185 7341
rect 4603 7351 4621 7369
rect 4774 7367 4794 7387
rect 4877 7371 4897 7391
rect 4992 7367 5012 7387
rect 5095 7371 5115 7391
rect 5203 7371 5223 7391
rect 7931 7413 7951 7433
rect 8039 7413 8059 7433
rect 8142 7417 8162 7437
rect 8257 7413 8277 7433
rect 8360 7417 8380 7437
rect 8533 7435 8551 7453
rect 8982 7462 9000 7480
rect 5306 7367 5326 7387
rect 235 7254 253 7272
rect 18678 7592 18698 7612
rect 18781 7596 18801 7616
rect 18896 7592 18916 7612
rect 18999 7596 19019 7616
rect 19107 7596 19127 7616
rect 19210 7592 19230 7612
rect 20037 7600 20057 7620
rect 20140 7596 20160 7616
rect 20248 7596 20268 7616
rect 20351 7600 20371 7620
rect 20466 7596 20486 7616
rect 25915 7749 25933 7767
rect 33939 7866 33959 7886
rect 34042 7862 34062 7882
rect 34150 7862 34170 7882
rect 34253 7866 34273 7886
rect 34368 7862 34388 7882
rect 34471 7866 34491 7886
rect 34658 7873 34676 7891
rect 30722 7811 30740 7829
rect 26356 7699 26374 7717
rect 20569 7600 20589 7620
rect 21546 7617 21564 7635
rect 23042 7605 23062 7625
rect 17278 7544 17296 7562
rect 12205 7429 12225 7449
rect 8531 7336 8549 7354
rect 8980 7363 8998 7381
rect 9151 7379 9171 7399
rect 9254 7383 9274 7403
rect 9369 7379 9389 7399
rect 9472 7383 9492 7403
rect 9580 7383 9600 7403
rect 12308 7425 12328 7445
rect 12416 7425 12436 7445
rect 12519 7429 12539 7449
rect 12634 7425 12654 7445
rect 12737 7429 12757 7449
rect 12910 7447 12928 7465
rect 13346 7475 13364 7493
rect 9683 7379 9703 7399
rect 4599 7267 4617 7285
rect 233 7155 251 7173
rect 1208 7170 1228 7190
rect 1311 7174 1331 7194
rect 1426 7170 1446 7190
rect 1529 7174 1549 7194
rect 1637 7174 1657 7194
rect 1740 7170 1760 7190
rect 2501 7180 2521 7200
rect 2604 7176 2624 7196
rect 2712 7176 2732 7196
rect 2815 7180 2835 7200
rect 2930 7176 2950 7196
rect 16569 7442 16589 7462
rect 12908 7348 12926 7366
rect 13344 7376 13362 7394
rect 13515 7392 13535 7412
rect 13618 7396 13638 7416
rect 13733 7392 13753 7412
rect 13836 7396 13856 7416
rect 13944 7396 13964 7416
rect 16672 7438 16692 7458
rect 16780 7438 16800 7458
rect 16883 7442 16903 7462
rect 16998 7438 17018 7458
rect 17101 7442 17121 7462
rect 17274 7460 17292 7478
rect 23145 7609 23165 7629
rect 23260 7605 23280 7625
rect 23363 7609 23383 7629
rect 23471 7609 23491 7629
rect 23574 7605 23594 7625
rect 24401 7613 24421 7633
rect 24504 7609 24524 7629
rect 24612 7609 24632 7629
rect 24715 7613 24735 7633
rect 24830 7609 24850 7629
rect 24933 7613 24953 7633
rect 25910 7630 25928 7648
rect 30292 7761 30310 7779
rect 30720 7712 30738 7730
rect 27419 7617 27439 7637
rect 21544 7518 21562 7536
rect 14047 7392 14067 7412
rect 8976 7279 8994 7297
rect 3033 7180 3053 7200
rect 228 7036 246 7054
rect 4597 7168 4615 7186
rect 5572 7183 5592 7203
rect 5675 7187 5695 7207
rect 5790 7183 5810 7203
rect 5893 7187 5913 7207
rect 6001 7187 6021 7207
rect 6104 7183 6124 7203
rect 6865 7193 6885 7213
rect 6968 7189 6988 7209
rect 7076 7189 7096 7209
rect 7179 7193 7199 7213
rect 7294 7189 7314 7209
rect 17612 7449 17630 7467
rect 17272 7361 17290 7379
rect 27522 7621 27542 7641
rect 27637 7617 27657 7637
rect 27740 7621 27760 7641
rect 27848 7621 27868 7641
rect 27951 7617 27971 7637
rect 28778 7625 28798 7645
rect 28881 7621 28901 7641
rect 28989 7621 29009 7641
rect 29092 7625 29112 7645
rect 29207 7621 29227 7641
rect 34656 7774 34674 7792
rect 29310 7625 29330 7645
rect 30287 7642 30305 7660
rect 31783 7630 31803 7650
rect 25908 7531 25926 7549
rect 20835 7416 20855 7436
rect 13340 7292 13358 7310
rect 7397 7193 7417 7213
rect 4164 7098 4182 7116
rect 4592 7049 4610 7067
rect 8974 7180 8992 7198
rect 9949 7195 9969 7215
rect 10052 7199 10072 7219
rect 10167 7195 10187 7215
rect 10270 7199 10290 7219
rect 10378 7199 10398 7219
rect 10481 7195 10501 7215
rect 11242 7205 11262 7225
rect 11345 7201 11365 7221
rect 11453 7201 11473 7221
rect 11556 7205 11576 7225
rect 11671 7201 11691 7221
rect 17610 7350 17628 7368
rect 17781 7366 17801 7386
rect 17884 7370 17904 7390
rect 17999 7366 18019 7386
rect 18102 7370 18122 7390
rect 18210 7370 18230 7390
rect 20938 7412 20958 7432
rect 21046 7412 21066 7432
rect 21149 7416 21169 7436
rect 21264 7412 21284 7432
rect 21367 7416 21387 7436
rect 21540 7434 21558 7452
rect 21976 7462 21994 7480
rect 18313 7366 18333 7386
rect 31886 7634 31906 7654
rect 32001 7630 32021 7650
rect 32104 7634 32124 7654
rect 32212 7634 32232 7654
rect 32315 7630 32335 7650
rect 33142 7638 33162 7658
rect 33245 7634 33265 7654
rect 33353 7634 33373 7654
rect 33456 7638 33476 7658
rect 33571 7634 33591 7654
rect 33674 7638 33694 7658
rect 34651 7655 34669 7673
rect 30285 7543 30303 7561
rect 25199 7429 25219 7449
rect 21538 7335 21556 7353
rect 21974 7363 21992 7381
rect 22145 7379 22165 7399
rect 22248 7383 22268 7403
rect 22363 7379 22383 7399
rect 22466 7383 22486 7403
rect 22574 7383 22594 7403
rect 25302 7425 25322 7445
rect 25410 7425 25430 7445
rect 25513 7429 25533 7449
rect 25628 7425 25648 7445
rect 25731 7429 25751 7449
rect 25904 7447 25922 7465
rect 26353 7474 26371 7492
rect 22677 7379 22697 7399
rect 17606 7266 17624 7284
rect 11774 7205 11794 7225
rect 8528 7111 8546 7129
rect 4162 6999 4180 7017
rect 226 6937 244 6955
rect 411 6942 431 6962
rect 514 6946 534 6966
rect 629 6942 649 6962
rect 732 6946 752 6966
rect 840 6946 860 6966
rect 943 6942 963 6962
rect 8969 7061 8987 7079
rect 13338 7193 13356 7211
rect 14313 7208 14333 7228
rect 14416 7212 14436 7232
rect 14531 7208 14551 7228
rect 14634 7212 14654 7232
rect 14742 7212 14762 7232
rect 14845 7208 14865 7228
rect 15606 7218 15626 7238
rect 15709 7214 15729 7234
rect 15817 7214 15837 7234
rect 15920 7218 15940 7238
rect 16035 7214 16055 7234
rect 16138 7218 16158 7238
rect 34649 7556 34667 7574
rect 29576 7441 29596 7461
rect 25902 7348 25920 7366
rect 26351 7375 26369 7393
rect 26522 7391 26542 7411
rect 26625 7395 26645 7415
rect 26740 7391 26760 7411
rect 26843 7395 26863 7415
rect 26951 7395 26971 7415
rect 29679 7437 29699 7457
rect 29787 7437 29807 7457
rect 29890 7441 29910 7461
rect 30005 7437 30025 7457
rect 30108 7441 30128 7461
rect 30281 7459 30299 7477
rect 30717 7487 30735 7505
rect 27054 7391 27074 7411
rect 21970 7279 21988 7297
rect 12905 7123 12923 7141
rect 8526 7012 8544 7030
rect 4590 6950 4608 6968
rect 4775 6955 4795 6975
rect 4878 6959 4898 6979
rect 4993 6955 5013 6975
rect 5096 6959 5116 6979
rect 5204 6959 5224 6979
rect 5307 6955 5327 6975
rect 13333 7074 13351 7092
rect 17269 7136 17287 7154
rect 17604 7167 17622 7185
rect 18579 7182 18599 7202
rect 18682 7186 18702 7206
rect 18797 7182 18817 7202
rect 18900 7186 18920 7206
rect 19008 7186 19028 7206
rect 19111 7182 19131 7202
rect 19872 7192 19892 7212
rect 19975 7188 19995 7208
rect 20083 7188 20103 7208
rect 20186 7192 20206 7212
rect 20301 7188 20321 7208
rect 33940 7454 33960 7474
rect 30279 7360 30297 7378
rect 30715 7388 30733 7406
rect 30886 7404 30906 7424
rect 30989 7408 31009 7428
rect 31104 7404 31124 7424
rect 31207 7408 31227 7428
rect 31315 7408 31335 7428
rect 34043 7450 34063 7470
rect 34151 7450 34171 7470
rect 34254 7454 34274 7474
rect 34369 7450 34389 7470
rect 34472 7454 34492 7474
rect 34645 7472 34663 7490
rect 31418 7404 31438 7424
rect 26347 7291 26365 7309
rect 20404 7192 20424 7212
rect 12903 7024 12921 7042
rect 8967 6962 8985 6980
rect 9152 6967 9172 6987
rect 9255 6971 9275 6991
rect 9370 6967 9390 6987
rect 9473 6971 9493 6991
rect 9581 6971 9601 6991
rect 9684 6967 9704 6987
rect 17267 7037 17285 7055
rect 17599 7048 17617 7066
rect 21968 7180 21986 7198
rect 22943 7195 22963 7215
rect 23046 7199 23066 7219
rect 23161 7195 23181 7215
rect 23264 7199 23284 7219
rect 23372 7199 23392 7219
rect 23475 7195 23495 7215
rect 24236 7205 24256 7225
rect 24339 7201 24359 7221
rect 24447 7201 24467 7221
rect 24550 7205 24570 7225
rect 24665 7201 24685 7221
rect 34643 7373 34661 7391
rect 30711 7304 30729 7322
rect 24768 7205 24788 7225
rect 21535 7110 21553 7128
rect 13331 6975 13349 6993
rect 13516 6980 13536 7000
rect 13619 6984 13639 7004
rect 13734 6980 13754 7000
rect 13837 6984 13857 7004
rect 13945 6984 13965 7004
rect 14048 6980 14068 7000
rect 21963 7061 21981 7079
rect 26345 7192 26363 7210
rect 27320 7207 27340 7227
rect 27423 7211 27443 7231
rect 27538 7207 27558 7227
rect 27641 7211 27661 7231
rect 27749 7211 27769 7231
rect 27852 7207 27872 7227
rect 28613 7217 28633 7237
rect 28716 7213 28736 7233
rect 28824 7213 28844 7233
rect 28927 7217 28947 7237
rect 29042 7213 29062 7233
rect 29145 7217 29165 7237
rect 25899 7123 25917 7141
rect 21533 7011 21551 7029
rect 17597 6949 17615 6967
rect 17782 6954 17802 6974
rect 17885 6958 17905 6978
rect 18000 6954 18020 6974
rect 18103 6958 18123 6978
rect 18211 6958 18231 6978
rect 18314 6954 18334 6974
rect 26340 7073 26358 7091
rect 30709 7205 30727 7223
rect 31684 7220 31704 7240
rect 31787 7224 31807 7244
rect 31902 7220 31922 7240
rect 32005 7224 32025 7244
rect 32113 7224 32133 7244
rect 32216 7220 32236 7240
rect 32977 7230 32997 7250
rect 33080 7226 33100 7246
rect 33188 7226 33208 7246
rect 33291 7230 33311 7250
rect 33406 7226 33426 7246
rect 33509 7230 33529 7250
rect 30276 7135 30294 7153
rect 25897 7024 25915 7042
rect 21961 6962 21979 6980
rect 22146 6967 22166 6987
rect 22249 6971 22269 6991
rect 22364 6967 22384 6987
rect 22467 6971 22487 6991
rect 22575 6971 22595 6991
rect 22678 6967 22698 6987
rect 30704 7086 30722 7104
rect 34640 7148 34658 7166
rect 30274 7036 30292 7054
rect 26338 6974 26356 6992
rect 26523 6979 26543 6999
rect 26626 6983 26646 7003
rect 26741 6979 26761 6999
rect 26844 6983 26864 7003
rect 26952 6983 26972 7003
rect 27055 6979 27075 6999
rect 34638 7049 34656 7067
rect 30702 6987 30720 7005
rect 30887 6992 30907 7012
rect 30990 6996 31010 7016
rect 31105 6992 31125 7012
rect 31208 6996 31228 7016
rect 31316 6996 31336 7016
rect 31419 6992 31439 7012
rect 3443 6798 3463 6818
rect 3546 6794 3566 6814
rect 3654 6794 3674 6814
rect 3757 6798 3777 6818
rect 3872 6794 3892 6814
rect 3975 6798 3995 6818
rect 4162 6805 4180 6823
rect 226 6743 244 6761
rect 7807 6811 7827 6831
rect 7910 6807 7930 6827
rect 8018 6807 8038 6827
rect 8121 6811 8141 6831
rect 8236 6807 8256 6827
rect 8339 6811 8359 6831
rect 8526 6818 8544 6836
rect 4590 6756 4608 6774
rect 224 6644 242 6662
rect 4160 6706 4178 6724
rect 12184 6823 12204 6843
rect 12287 6819 12307 6839
rect 12395 6819 12415 6839
rect 12498 6823 12518 6843
rect 12613 6819 12633 6839
rect 12716 6823 12736 6843
rect 12903 6830 12921 6848
rect 8967 6768 8985 6786
rect 4588 6657 4606 6675
rect 1353 6560 1373 6580
rect 1456 6564 1476 6584
rect 1571 6560 1591 6580
rect 1674 6564 1694 6584
rect 1782 6564 1802 6584
rect 1885 6560 1905 6580
rect 2646 6570 2666 6590
rect 2749 6566 2769 6586
rect 2857 6566 2877 6586
rect 2960 6570 2980 6590
rect 3075 6566 3095 6586
rect 3178 6570 3198 6590
rect 4155 6587 4173 6605
rect 8524 6719 8542 6737
rect 16548 6836 16568 6856
rect 16651 6832 16671 6852
rect 16759 6832 16779 6852
rect 16862 6836 16882 6856
rect 16977 6832 16997 6852
rect 17080 6836 17100 6856
rect 17267 6843 17285 6861
rect 13331 6781 13349 6799
rect 8965 6669 8983 6687
rect 5717 6573 5737 6593
rect 5820 6577 5840 6597
rect 5935 6573 5955 6593
rect 6038 6577 6058 6597
rect 6146 6577 6166 6597
rect 6249 6573 6269 6593
rect 7010 6583 7030 6603
rect 7113 6579 7133 6599
rect 7221 6579 7241 6599
rect 7324 6583 7344 6603
rect 7439 6579 7459 6599
rect 7542 6583 7562 6603
rect 8519 6600 8537 6618
rect 12901 6731 12919 6749
rect 20814 6810 20834 6830
rect 20917 6806 20937 6826
rect 21025 6806 21045 6826
rect 21128 6810 21148 6830
rect 21243 6806 21263 6826
rect 21346 6810 21366 6830
rect 21533 6817 21551 6835
rect 13329 6682 13347 6700
rect 10094 6585 10114 6605
rect 4153 6488 4171 6506
rect 221 6419 239 6437
rect 10197 6589 10217 6609
rect 10312 6585 10332 6605
rect 10415 6589 10435 6609
rect 10523 6589 10543 6609
rect 10626 6585 10646 6605
rect 11387 6595 11407 6615
rect 11490 6591 11510 6611
rect 11598 6591 11618 6611
rect 11701 6595 11721 6615
rect 11816 6591 11836 6611
rect 11919 6595 11939 6615
rect 12896 6612 12914 6630
rect 17265 6744 17283 6762
rect 17597 6755 17615 6773
rect 25178 6823 25198 6843
rect 25281 6819 25301 6839
rect 25389 6819 25409 6839
rect 25492 6823 25512 6843
rect 25607 6819 25627 6839
rect 25710 6823 25730 6843
rect 25897 6830 25915 6848
rect 21961 6768 21979 6786
rect 14458 6598 14478 6618
rect 8517 6501 8535 6519
rect 3444 6386 3464 6406
rect 219 6320 237 6338
rect 390 6336 410 6356
rect 493 6340 513 6360
rect 608 6336 628 6356
rect 711 6340 731 6360
rect 819 6340 839 6360
rect 3547 6382 3567 6402
rect 3655 6382 3675 6402
rect 3758 6386 3778 6406
rect 3873 6382 3893 6402
rect 3976 6386 3996 6406
rect 4149 6404 4167 6422
rect 4585 6432 4603 6450
rect 922 6336 942 6356
rect 14561 6602 14581 6622
rect 14676 6598 14696 6618
rect 14779 6602 14799 6622
rect 14887 6602 14907 6622
rect 14990 6598 15010 6618
rect 15751 6608 15771 6628
rect 15854 6604 15874 6624
rect 15962 6604 15982 6624
rect 16065 6608 16085 6628
rect 16180 6604 16200 6624
rect 16283 6608 16303 6628
rect 17260 6625 17278 6643
rect 17595 6656 17613 6674
rect 21531 6718 21549 6736
rect 29555 6835 29575 6855
rect 29658 6831 29678 6851
rect 29766 6831 29786 6851
rect 29869 6835 29889 6855
rect 29984 6831 30004 6851
rect 30087 6835 30107 6855
rect 30274 6842 30292 6860
rect 26338 6780 26356 6798
rect 21959 6669 21977 6687
rect 12894 6513 12912 6531
rect 7808 6399 7828 6419
rect 4147 6305 4165 6323
rect 4583 6333 4601 6351
rect 4754 6349 4774 6369
rect 4857 6353 4877 6373
rect 4972 6349 4992 6369
rect 5075 6353 5095 6373
rect 5183 6353 5203 6373
rect 7911 6395 7931 6415
rect 8019 6395 8039 6415
rect 8122 6399 8142 6419
rect 8237 6395 8257 6415
rect 8340 6399 8360 6419
rect 8513 6417 8531 6435
rect 8962 6444 8980 6462
rect 5286 6349 5306 6369
rect 215 6236 233 6254
rect 18724 6572 18744 6592
rect 18827 6576 18847 6596
rect 18942 6572 18962 6592
rect 19045 6576 19065 6596
rect 19153 6576 19173 6596
rect 19256 6572 19276 6592
rect 20017 6582 20037 6602
rect 20120 6578 20140 6598
rect 20228 6578 20248 6598
rect 20331 6582 20351 6602
rect 20446 6578 20466 6598
rect 20549 6582 20569 6602
rect 21526 6599 21544 6617
rect 25895 6731 25913 6749
rect 33919 6848 33939 6868
rect 34022 6844 34042 6864
rect 34130 6844 34150 6864
rect 34233 6848 34253 6868
rect 34348 6844 34368 6864
rect 34451 6848 34471 6868
rect 34638 6855 34656 6873
rect 30702 6793 30720 6811
rect 26336 6681 26354 6699
rect 23088 6585 23108 6605
rect 17258 6526 17276 6544
rect 12185 6411 12205 6431
rect 8511 6318 8529 6336
rect 8960 6345 8978 6363
rect 9131 6361 9151 6381
rect 9234 6365 9254 6385
rect 9349 6361 9369 6381
rect 9452 6365 9472 6385
rect 9560 6365 9580 6385
rect 12288 6407 12308 6427
rect 12396 6407 12416 6427
rect 12499 6411 12519 6431
rect 12614 6407 12634 6427
rect 12717 6411 12737 6431
rect 12890 6429 12908 6447
rect 13326 6457 13344 6475
rect 9663 6361 9683 6381
rect 4579 6249 4597 6267
rect 213 6137 231 6155
rect 1188 6152 1208 6172
rect 1291 6156 1311 6176
rect 1406 6152 1426 6172
rect 1509 6156 1529 6176
rect 1617 6156 1637 6176
rect 1720 6152 1740 6172
rect 2547 6160 2567 6180
rect 2650 6156 2670 6176
rect 2758 6156 2778 6176
rect 2861 6160 2881 6180
rect 2976 6156 2996 6176
rect 16549 6424 16569 6444
rect 12888 6330 12906 6348
rect 13324 6358 13342 6376
rect 13495 6374 13515 6394
rect 13598 6378 13618 6398
rect 13713 6374 13733 6394
rect 13816 6378 13836 6398
rect 13924 6378 13944 6398
rect 16652 6420 16672 6440
rect 16760 6420 16780 6440
rect 16863 6424 16883 6444
rect 16978 6420 16998 6440
rect 17081 6424 17101 6444
rect 17254 6442 17272 6460
rect 23191 6589 23211 6609
rect 23306 6585 23326 6605
rect 23409 6589 23429 6609
rect 23517 6589 23537 6609
rect 23620 6585 23640 6605
rect 24381 6595 24401 6615
rect 24484 6591 24504 6611
rect 24592 6591 24612 6611
rect 24695 6595 24715 6615
rect 24810 6591 24830 6611
rect 24913 6595 24933 6615
rect 25890 6612 25908 6630
rect 30272 6743 30290 6761
rect 30700 6694 30718 6712
rect 27465 6597 27485 6617
rect 21524 6500 21542 6518
rect 14027 6374 14047 6394
rect 8956 6261 8974 6279
rect 3079 6160 3099 6180
rect 4577 6150 4595 6168
rect 5552 6165 5572 6185
rect 208 6018 226 6036
rect 5655 6169 5675 6189
rect 5770 6165 5790 6185
rect 5873 6169 5893 6189
rect 5981 6169 6001 6189
rect 6084 6165 6104 6185
rect 6911 6173 6931 6193
rect 7014 6169 7034 6189
rect 7122 6169 7142 6189
rect 7225 6173 7245 6193
rect 7340 6169 7360 6189
rect 17592 6431 17610 6449
rect 17252 6343 17270 6361
rect 27568 6601 27588 6621
rect 27683 6597 27703 6617
rect 27786 6601 27806 6621
rect 27894 6601 27914 6621
rect 27997 6597 28017 6617
rect 28758 6607 28778 6627
rect 28861 6603 28881 6623
rect 28969 6603 28989 6623
rect 29072 6607 29092 6627
rect 29187 6603 29207 6623
rect 29290 6607 29310 6627
rect 30267 6624 30285 6642
rect 34636 6756 34654 6774
rect 31829 6610 31849 6630
rect 25888 6513 25906 6531
rect 20815 6398 20835 6418
rect 13320 6274 13338 6292
rect 7443 6173 7463 6193
rect 4144 6080 4162 6098
rect 4572 6031 4590 6049
rect 8954 6162 8972 6180
rect 9929 6177 9949 6197
rect 10032 6181 10052 6201
rect 10147 6177 10167 6197
rect 10250 6181 10270 6201
rect 10358 6181 10378 6201
rect 10461 6177 10481 6197
rect 11288 6185 11308 6205
rect 11391 6181 11411 6201
rect 11499 6181 11519 6201
rect 11602 6185 11622 6205
rect 11717 6181 11737 6201
rect 17590 6332 17608 6350
rect 17761 6348 17781 6368
rect 17864 6352 17884 6372
rect 17979 6348 17999 6368
rect 18082 6352 18102 6372
rect 18190 6352 18210 6372
rect 20918 6394 20938 6414
rect 21026 6394 21046 6414
rect 21129 6398 21149 6418
rect 21244 6394 21264 6414
rect 21347 6398 21367 6418
rect 21520 6416 21538 6434
rect 21956 6444 21974 6462
rect 18293 6348 18313 6368
rect 31932 6614 31952 6634
rect 32047 6610 32067 6630
rect 32150 6614 32170 6634
rect 32258 6614 32278 6634
rect 32361 6610 32381 6630
rect 33122 6620 33142 6640
rect 33225 6616 33245 6636
rect 33333 6616 33353 6636
rect 33436 6620 33456 6640
rect 33551 6616 33571 6636
rect 33654 6620 33674 6640
rect 34631 6637 34649 6655
rect 30265 6525 30283 6543
rect 25179 6411 25199 6431
rect 21518 6317 21536 6335
rect 21954 6345 21972 6363
rect 22125 6361 22145 6381
rect 22228 6365 22248 6385
rect 22343 6361 22363 6381
rect 22446 6365 22466 6385
rect 22554 6365 22574 6385
rect 25282 6407 25302 6427
rect 25390 6407 25410 6427
rect 25493 6411 25513 6431
rect 25608 6407 25628 6427
rect 25711 6411 25731 6431
rect 25884 6429 25902 6447
rect 26333 6456 26351 6474
rect 22657 6361 22677 6381
rect 17586 6248 17604 6266
rect 11820 6185 11840 6205
rect 13318 6175 13336 6193
rect 14293 6190 14313 6210
rect 8508 6093 8526 6111
rect 4142 5981 4160 5999
rect 206 5919 224 5937
rect 391 5924 411 5944
rect 494 5928 514 5948
rect 609 5924 629 5944
rect 712 5928 732 5948
rect 820 5928 840 5948
rect 923 5924 943 5944
rect 8949 6043 8967 6061
rect 14396 6194 14416 6214
rect 14511 6190 14531 6210
rect 14614 6194 14634 6214
rect 14722 6194 14742 6214
rect 14825 6190 14845 6210
rect 15652 6198 15672 6218
rect 15755 6194 15775 6214
rect 15863 6194 15883 6214
rect 15966 6198 15986 6218
rect 16081 6194 16101 6214
rect 16184 6198 16204 6218
rect 34629 6538 34647 6556
rect 29556 6423 29576 6443
rect 25882 6330 25900 6348
rect 26331 6357 26349 6375
rect 26502 6373 26522 6393
rect 26605 6377 26625 6397
rect 26720 6373 26740 6393
rect 26823 6377 26843 6397
rect 26931 6377 26951 6397
rect 29659 6419 29679 6439
rect 29767 6419 29787 6439
rect 29870 6423 29890 6443
rect 29985 6419 30005 6439
rect 30088 6423 30108 6443
rect 30261 6441 30279 6459
rect 30697 6469 30715 6487
rect 27034 6373 27054 6393
rect 21950 6261 21968 6279
rect 12885 6105 12903 6123
rect 8506 5994 8524 6012
rect 4570 5932 4588 5950
rect 4755 5937 4775 5957
rect 4858 5941 4878 5961
rect 4973 5937 4993 5957
rect 5076 5941 5096 5961
rect 5184 5941 5204 5961
rect 5287 5937 5307 5957
rect 13313 6056 13331 6074
rect 17249 6118 17267 6136
rect 17584 6149 17602 6167
rect 18559 6164 18579 6184
rect 18662 6168 18682 6188
rect 18777 6164 18797 6184
rect 18880 6168 18900 6188
rect 18988 6168 19008 6188
rect 19091 6164 19111 6184
rect 19918 6172 19938 6192
rect 20021 6168 20041 6188
rect 20129 6168 20149 6188
rect 20232 6172 20252 6192
rect 20347 6168 20367 6188
rect 33920 6436 33940 6456
rect 30259 6342 30277 6360
rect 30695 6370 30713 6388
rect 30866 6386 30886 6406
rect 30969 6390 30989 6410
rect 31084 6386 31104 6406
rect 31187 6390 31207 6410
rect 31295 6390 31315 6410
rect 34023 6432 34043 6452
rect 34131 6432 34151 6452
rect 34234 6436 34254 6456
rect 34349 6432 34369 6452
rect 34452 6436 34472 6456
rect 34625 6454 34643 6472
rect 31398 6386 31418 6406
rect 26327 6273 26345 6291
rect 20450 6172 20470 6192
rect 21948 6162 21966 6180
rect 22923 6177 22943 6197
rect 12883 6006 12901 6024
rect 8947 5944 8965 5962
rect 9132 5949 9152 5969
rect 9235 5953 9255 5973
rect 9350 5949 9370 5969
rect 9453 5953 9473 5973
rect 9561 5953 9581 5973
rect 9664 5949 9684 5969
rect 17247 6019 17265 6037
rect 17579 6030 17597 6048
rect 23026 6181 23046 6201
rect 23141 6177 23161 6197
rect 23244 6181 23264 6201
rect 23352 6181 23372 6201
rect 23455 6177 23475 6197
rect 24282 6185 24302 6205
rect 24385 6181 24405 6201
rect 24493 6181 24513 6201
rect 24596 6185 24616 6205
rect 24711 6181 24731 6201
rect 34623 6355 34641 6373
rect 30691 6286 30709 6304
rect 24814 6185 24834 6205
rect 21515 6092 21533 6110
rect 13311 5957 13329 5975
rect 13496 5962 13516 5982
rect 13599 5966 13619 5986
rect 13714 5962 13734 5982
rect 13817 5966 13837 5986
rect 13925 5966 13945 5986
rect 14028 5962 14048 5982
rect 21943 6043 21961 6061
rect 26325 6174 26343 6192
rect 27300 6189 27320 6209
rect 27403 6193 27423 6213
rect 27518 6189 27538 6209
rect 27621 6193 27641 6213
rect 27729 6193 27749 6213
rect 27832 6189 27852 6209
rect 28659 6197 28679 6217
rect 28762 6193 28782 6213
rect 28870 6193 28890 6213
rect 28973 6197 28993 6217
rect 29088 6193 29108 6213
rect 29191 6197 29211 6217
rect 30689 6187 30707 6205
rect 31664 6202 31684 6222
rect 25879 6105 25897 6123
rect 21513 5993 21531 6011
rect 17577 5931 17595 5949
rect 17762 5936 17782 5956
rect 17865 5940 17885 5960
rect 17980 5936 18000 5956
rect 18083 5940 18103 5960
rect 18191 5940 18211 5960
rect 18294 5936 18314 5956
rect 26320 6055 26338 6073
rect 31767 6206 31787 6226
rect 31882 6202 31902 6222
rect 31985 6206 32005 6226
rect 32093 6206 32113 6226
rect 32196 6202 32216 6222
rect 33023 6210 33043 6230
rect 33126 6206 33146 6226
rect 33234 6206 33254 6226
rect 33337 6210 33357 6230
rect 33452 6206 33472 6226
rect 33555 6210 33575 6230
rect 30256 6117 30274 6135
rect 25877 6006 25895 6024
rect 21941 5944 21959 5962
rect 22126 5949 22146 5969
rect 22229 5953 22249 5973
rect 22344 5949 22364 5969
rect 22447 5953 22467 5973
rect 22555 5953 22575 5973
rect 22658 5949 22678 5969
rect 30684 6068 30702 6086
rect 34620 6130 34638 6148
rect 30254 6018 30272 6036
rect 26318 5956 26336 5974
rect 26503 5961 26523 5981
rect 26606 5965 26626 5985
rect 26721 5961 26741 5981
rect 26824 5965 26844 5985
rect 26932 5965 26952 5985
rect 27035 5961 27055 5981
rect 34618 6031 34636 6049
rect 30682 5969 30700 5987
rect 30867 5974 30887 5994
rect 30970 5978 30990 5998
rect 31085 5974 31105 5994
rect 31188 5978 31208 5998
rect 31296 5978 31316 5998
rect 31399 5974 31419 5994
rect 3426 5780 3446 5800
rect 3529 5776 3549 5796
rect 3637 5776 3657 5796
rect 3740 5780 3760 5800
rect 3855 5776 3875 5796
rect 3958 5780 3978 5800
rect 4145 5787 4163 5805
rect 209 5725 227 5743
rect 7790 5793 7810 5813
rect 7893 5789 7913 5809
rect 8001 5789 8021 5809
rect 8104 5793 8124 5813
rect 8219 5789 8239 5809
rect 8322 5793 8342 5813
rect 8509 5800 8527 5818
rect 4573 5738 4591 5756
rect 207 5626 225 5644
rect 4143 5688 4161 5706
rect 12167 5805 12187 5825
rect 12270 5801 12290 5821
rect 12378 5801 12398 5821
rect 12481 5805 12501 5825
rect 12596 5801 12616 5821
rect 12699 5805 12719 5825
rect 12886 5812 12904 5830
rect 8950 5750 8968 5768
rect 4571 5639 4589 5657
rect 1270 5544 1290 5564
rect 1373 5548 1393 5568
rect 1488 5544 1508 5564
rect 1591 5548 1611 5568
rect 1699 5548 1719 5568
rect 1802 5544 1822 5564
rect 2629 5552 2649 5572
rect 2732 5548 2752 5568
rect 2840 5548 2860 5568
rect 2943 5552 2963 5572
rect 3058 5548 3078 5568
rect 8507 5701 8525 5719
rect 16531 5818 16551 5838
rect 16634 5814 16654 5834
rect 16742 5814 16762 5834
rect 16845 5818 16865 5838
rect 16960 5814 16980 5834
rect 17063 5818 17083 5838
rect 17250 5825 17268 5843
rect 13314 5763 13332 5781
rect 8948 5651 8966 5669
rect 3161 5552 3181 5572
rect 4138 5569 4156 5587
rect 5634 5557 5654 5577
rect 5737 5561 5757 5581
rect 5852 5557 5872 5577
rect 5955 5561 5975 5581
rect 6063 5561 6083 5581
rect 6166 5557 6186 5577
rect 6993 5565 7013 5585
rect 7096 5561 7116 5581
rect 7204 5561 7224 5581
rect 7307 5565 7327 5585
rect 7422 5561 7442 5581
rect 7525 5565 7545 5585
rect 8502 5582 8520 5600
rect 12884 5713 12902 5731
rect 20797 5792 20817 5812
rect 20900 5788 20920 5808
rect 21008 5788 21028 5808
rect 21111 5792 21131 5812
rect 21226 5788 21246 5808
rect 21329 5792 21349 5812
rect 21516 5799 21534 5817
rect 13312 5664 13330 5682
rect 10011 5569 10031 5589
rect 4136 5470 4154 5488
rect 204 5401 222 5419
rect 10114 5573 10134 5593
rect 10229 5569 10249 5589
rect 10332 5573 10352 5593
rect 10440 5573 10460 5593
rect 10543 5569 10563 5589
rect 11370 5577 11390 5597
rect 11473 5573 11493 5593
rect 11581 5573 11601 5593
rect 11684 5577 11704 5597
rect 11799 5573 11819 5593
rect 17248 5726 17266 5744
rect 17580 5737 17598 5755
rect 25161 5805 25181 5825
rect 25264 5801 25284 5821
rect 25372 5801 25392 5821
rect 25475 5805 25495 5825
rect 25590 5801 25610 5821
rect 25693 5805 25713 5825
rect 25880 5812 25898 5830
rect 21944 5750 21962 5768
rect 11902 5577 11922 5597
rect 12879 5594 12897 5612
rect 14375 5582 14395 5602
rect 8500 5483 8518 5501
rect 3427 5368 3447 5388
rect 202 5302 220 5320
rect 373 5318 393 5338
rect 476 5322 496 5342
rect 591 5318 611 5338
rect 694 5322 714 5342
rect 802 5322 822 5342
rect 3530 5364 3550 5384
rect 3638 5364 3658 5384
rect 3741 5368 3761 5388
rect 3856 5364 3876 5384
rect 3959 5368 3979 5388
rect 4132 5386 4150 5404
rect 4568 5414 4586 5432
rect 905 5318 925 5338
rect 14478 5586 14498 5606
rect 14593 5582 14613 5602
rect 14696 5586 14716 5606
rect 14804 5586 14824 5606
rect 14907 5582 14927 5602
rect 15734 5590 15754 5610
rect 15837 5586 15857 5606
rect 15945 5586 15965 5606
rect 16048 5590 16068 5610
rect 16163 5586 16183 5606
rect 16266 5590 16286 5610
rect 17243 5607 17261 5625
rect 17578 5638 17596 5656
rect 21514 5700 21532 5718
rect 29538 5817 29558 5837
rect 29641 5813 29661 5833
rect 29749 5813 29769 5833
rect 29852 5817 29872 5837
rect 29967 5813 29987 5833
rect 30070 5817 30090 5837
rect 30257 5824 30275 5842
rect 26321 5762 26339 5780
rect 21942 5651 21960 5669
rect 12877 5495 12895 5513
rect 7791 5381 7811 5401
rect 4130 5287 4148 5305
rect 4566 5315 4584 5333
rect 4737 5331 4757 5351
rect 4840 5335 4860 5355
rect 4955 5331 4975 5351
rect 5058 5335 5078 5355
rect 5166 5335 5186 5355
rect 7894 5377 7914 5397
rect 8002 5377 8022 5397
rect 8105 5381 8125 5401
rect 8220 5377 8240 5397
rect 8323 5381 8343 5401
rect 8496 5399 8514 5417
rect 8945 5426 8963 5444
rect 5269 5331 5289 5351
rect 198 5218 216 5236
rect 18641 5556 18661 5576
rect 18744 5560 18764 5580
rect 18859 5556 18879 5576
rect 18962 5560 18982 5580
rect 19070 5560 19090 5580
rect 19173 5556 19193 5576
rect 20000 5564 20020 5584
rect 20103 5560 20123 5580
rect 20211 5560 20231 5580
rect 20314 5564 20334 5584
rect 20429 5560 20449 5580
rect 25878 5713 25896 5731
rect 33902 5830 33922 5850
rect 34005 5826 34025 5846
rect 34113 5826 34133 5846
rect 34216 5830 34236 5850
rect 34331 5826 34351 5846
rect 34434 5830 34454 5850
rect 34621 5837 34639 5855
rect 30685 5775 30703 5793
rect 26319 5663 26337 5681
rect 20532 5564 20552 5584
rect 21509 5581 21527 5599
rect 23005 5569 23025 5589
rect 17241 5508 17259 5526
rect 12168 5393 12188 5413
rect 8494 5300 8512 5318
rect 8943 5327 8961 5345
rect 9114 5343 9134 5363
rect 9217 5347 9237 5367
rect 9332 5343 9352 5363
rect 9435 5347 9455 5367
rect 9543 5347 9563 5367
rect 12271 5389 12291 5409
rect 12379 5389 12399 5409
rect 12482 5393 12502 5413
rect 12597 5389 12617 5409
rect 12700 5393 12720 5413
rect 12873 5411 12891 5429
rect 13309 5439 13327 5457
rect 9646 5343 9666 5363
rect 4562 5231 4580 5249
rect 196 5119 214 5137
rect 1171 5134 1191 5154
rect 1274 5138 1294 5158
rect 1389 5134 1409 5154
rect 1492 5138 1512 5158
rect 1600 5138 1620 5158
rect 1703 5134 1723 5154
rect 2325 5146 2345 5166
rect 2428 5142 2448 5162
rect 2536 5142 2556 5162
rect 2639 5146 2659 5166
rect 2754 5142 2774 5162
rect 16532 5406 16552 5426
rect 12871 5312 12889 5330
rect 13307 5340 13325 5358
rect 13478 5356 13498 5376
rect 13581 5360 13601 5380
rect 13696 5356 13716 5376
rect 13799 5360 13819 5380
rect 13907 5360 13927 5380
rect 16635 5402 16655 5422
rect 16743 5402 16763 5422
rect 16846 5406 16866 5426
rect 16961 5402 16981 5422
rect 17064 5406 17084 5426
rect 17237 5424 17255 5442
rect 23108 5573 23128 5593
rect 23223 5569 23243 5589
rect 23326 5573 23346 5593
rect 23434 5573 23454 5593
rect 23537 5569 23557 5589
rect 24364 5577 24384 5597
rect 24467 5573 24487 5593
rect 24575 5573 24595 5593
rect 24678 5577 24698 5597
rect 24793 5573 24813 5593
rect 24896 5577 24916 5597
rect 25873 5594 25891 5612
rect 30255 5725 30273 5743
rect 30683 5676 30701 5694
rect 27382 5581 27402 5601
rect 21507 5482 21525 5500
rect 14010 5356 14030 5376
rect 8939 5243 8957 5261
rect 2857 5146 2877 5166
rect 191 5000 209 5018
rect 4560 5132 4578 5150
rect 5535 5147 5555 5167
rect 5638 5151 5658 5171
rect 5753 5147 5773 5167
rect 5856 5151 5876 5171
rect 5964 5151 5984 5171
rect 6067 5147 6087 5167
rect 6689 5159 6709 5179
rect 6792 5155 6812 5175
rect 6900 5155 6920 5175
rect 7003 5159 7023 5179
rect 7118 5155 7138 5175
rect 17575 5413 17593 5431
rect 17235 5325 17253 5343
rect 27485 5585 27505 5605
rect 27600 5581 27620 5601
rect 27703 5585 27723 5605
rect 27811 5585 27831 5605
rect 27914 5581 27934 5601
rect 28741 5589 28761 5609
rect 28844 5585 28864 5605
rect 28952 5585 28972 5605
rect 29055 5589 29075 5609
rect 29170 5585 29190 5605
rect 34619 5738 34637 5756
rect 29273 5589 29293 5609
rect 30250 5606 30268 5624
rect 31746 5594 31766 5614
rect 25871 5495 25889 5513
rect 20798 5380 20818 5400
rect 13303 5256 13321 5274
rect 7221 5159 7241 5179
rect 4127 5062 4145 5080
rect 4555 5013 4573 5031
rect 8937 5144 8955 5162
rect 9912 5159 9932 5179
rect 10015 5163 10035 5183
rect 10130 5159 10150 5179
rect 10233 5163 10253 5183
rect 10341 5163 10361 5183
rect 10444 5159 10464 5179
rect 11066 5171 11086 5191
rect 11169 5167 11189 5187
rect 11277 5167 11297 5187
rect 11380 5171 11400 5191
rect 11495 5167 11515 5187
rect 17573 5314 17591 5332
rect 17744 5330 17764 5350
rect 17847 5334 17867 5354
rect 17962 5330 17982 5350
rect 18065 5334 18085 5354
rect 18173 5334 18193 5354
rect 20901 5376 20921 5396
rect 21009 5376 21029 5396
rect 21112 5380 21132 5400
rect 21227 5376 21247 5396
rect 21330 5380 21350 5400
rect 21503 5398 21521 5416
rect 21939 5426 21957 5444
rect 18276 5330 18296 5350
rect 31849 5598 31869 5618
rect 31964 5594 31984 5614
rect 32067 5598 32087 5618
rect 32175 5598 32195 5618
rect 32278 5594 32298 5614
rect 33105 5602 33125 5622
rect 33208 5598 33228 5618
rect 33316 5598 33336 5618
rect 33419 5602 33439 5622
rect 33534 5598 33554 5618
rect 33637 5602 33657 5622
rect 34614 5619 34632 5637
rect 30248 5507 30266 5525
rect 25162 5393 25182 5413
rect 21501 5299 21519 5317
rect 21937 5327 21955 5345
rect 22108 5343 22128 5363
rect 22211 5347 22231 5367
rect 22326 5343 22346 5363
rect 22429 5347 22449 5367
rect 22537 5347 22557 5367
rect 25265 5389 25285 5409
rect 25373 5389 25393 5409
rect 25476 5393 25496 5413
rect 25591 5389 25611 5409
rect 25694 5393 25714 5413
rect 25867 5411 25885 5429
rect 26316 5438 26334 5456
rect 22640 5343 22660 5363
rect 17569 5230 17587 5248
rect 11598 5171 11618 5191
rect 8491 5075 8509 5093
rect 4125 4963 4143 4981
rect 189 4901 207 4919
rect 374 4906 394 4926
rect 477 4910 497 4930
rect 592 4906 612 4926
rect 695 4910 715 4930
rect 803 4910 823 4930
rect 906 4906 926 4926
rect 8932 5025 8950 5043
rect 13301 5157 13319 5175
rect 14276 5172 14296 5192
rect 14379 5176 14399 5196
rect 14494 5172 14514 5192
rect 14597 5176 14617 5196
rect 14705 5176 14725 5196
rect 14808 5172 14828 5192
rect 15430 5184 15450 5204
rect 15533 5180 15553 5200
rect 15641 5180 15661 5200
rect 15744 5184 15764 5204
rect 15859 5180 15879 5200
rect 15962 5184 15982 5204
rect 12868 5087 12886 5105
rect 8489 4976 8507 4994
rect 4553 4914 4571 4932
rect 4738 4919 4758 4939
rect 4841 4923 4861 4943
rect 4956 4919 4976 4939
rect 5059 4923 5079 4943
rect 5167 4923 5187 4943
rect 5270 4919 5290 4939
rect 13296 5038 13314 5056
rect 34612 5520 34630 5538
rect 29539 5405 29559 5425
rect 25865 5312 25883 5330
rect 26314 5339 26332 5357
rect 26485 5355 26505 5375
rect 26588 5359 26608 5379
rect 26703 5355 26723 5375
rect 26806 5359 26826 5379
rect 26914 5359 26934 5379
rect 29642 5401 29662 5421
rect 29750 5401 29770 5421
rect 29853 5405 29873 5425
rect 29968 5401 29988 5421
rect 30071 5405 30091 5425
rect 30244 5423 30262 5441
rect 30680 5451 30698 5469
rect 27017 5355 27037 5375
rect 21933 5243 21951 5261
rect 17232 5100 17250 5118
rect 17567 5131 17585 5149
rect 18542 5146 18562 5166
rect 18645 5150 18665 5170
rect 18760 5146 18780 5166
rect 18863 5150 18883 5170
rect 18971 5150 18991 5170
rect 19074 5146 19094 5166
rect 19696 5158 19716 5178
rect 19799 5154 19819 5174
rect 19907 5154 19927 5174
rect 20010 5158 20030 5178
rect 20125 5154 20145 5174
rect 33903 5418 33923 5438
rect 30242 5324 30260 5342
rect 30678 5352 30696 5370
rect 30849 5368 30869 5388
rect 30952 5372 30972 5392
rect 31067 5368 31087 5388
rect 31170 5372 31190 5392
rect 31278 5372 31298 5392
rect 34006 5414 34026 5434
rect 34114 5414 34134 5434
rect 34217 5418 34237 5438
rect 34332 5414 34352 5434
rect 34435 5418 34455 5438
rect 34608 5436 34626 5454
rect 31381 5368 31401 5388
rect 26310 5255 26328 5273
rect 20228 5158 20248 5178
rect 12866 4988 12884 5006
rect 8930 4926 8948 4944
rect 9115 4931 9135 4951
rect 9218 4935 9238 4955
rect 9333 4931 9353 4951
rect 9436 4935 9456 4955
rect 9544 4935 9564 4955
rect 9647 4931 9667 4951
rect 17230 5001 17248 5019
rect 17562 5012 17580 5030
rect 21931 5144 21949 5162
rect 22906 5159 22926 5179
rect 23009 5163 23029 5183
rect 23124 5159 23144 5179
rect 23227 5163 23247 5183
rect 23335 5163 23355 5183
rect 23438 5159 23458 5179
rect 24060 5171 24080 5191
rect 24163 5167 24183 5187
rect 24271 5167 24291 5187
rect 24374 5171 24394 5191
rect 24489 5167 24509 5187
rect 34606 5337 34624 5355
rect 30674 5268 30692 5286
rect 24592 5171 24612 5191
rect 21498 5074 21516 5092
rect 13294 4939 13312 4957
rect 13479 4944 13499 4964
rect 13582 4948 13602 4968
rect 13697 4944 13717 4964
rect 13800 4948 13820 4968
rect 13908 4948 13928 4968
rect 14011 4944 14031 4964
rect 21926 5025 21944 5043
rect 26308 5156 26326 5174
rect 27283 5171 27303 5191
rect 27386 5175 27406 5195
rect 27501 5171 27521 5191
rect 27604 5175 27624 5195
rect 27712 5175 27732 5195
rect 27815 5171 27835 5191
rect 28437 5183 28457 5203
rect 28540 5179 28560 5199
rect 28648 5179 28668 5199
rect 28751 5183 28771 5203
rect 28866 5179 28886 5199
rect 28969 5183 28989 5203
rect 25862 5087 25880 5105
rect 21496 4975 21514 4993
rect 17560 4913 17578 4931
rect 17745 4918 17765 4938
rect 17848 4922 17868 4942
rect 17963 4918 17983 4938
rect 18066 4922 18086 4942
rect 18174 4922 18194 4942
rect 18277 4918 18297 4938
rect 26303 5037 26321 5055
rect 30672 5169 30690 5187
rect 31647 5184 31667 5204
rect 31750 5188 31770 5208
rect 31865 5184 31885 5204
rect 31968 5188 31988 5208
rect 32076 5188 32096 5208
rect 32179 5184 32199 5204
rect 32801 5196 32821 5216
rect 32904 5192 32924 5212
rect 33012 5192 33032 5212
rect 33115 5196 33135 5216
rect 33230 5192 33250 5212
rect 33333 5196 33353 5216
rect 30239 5099 30257 5117
rect 25860 4988 25878 5006
rect 21924 4926 21942 4944
rect 22109 4931 22129 4951
rect 22212 4935 22232 4955
rect 22327 4931 22347 4951
rect 22430 4935 22450 4955
rect 22538 4935 22558 4955
rect 22641 4931 22661 4951
rect 30667 5050 30685 5068
rect 34603 5112 34621 5130
rect 30237 5000 30255 5018
rect 26301 4938 26319 4956
rect 26486 4943 26506 4963
rect 26589 4947 26609 4967
rect 26704 4943 26724 4963
rect 26807 4947 26827 4967
rect 26915 4947 26935 4967
rect 27018 4943 27038 4963
rect 34601 5013 34619 5031
rect 30665 4951 30683 4969
rect 30850 4956 30870 4976
rect 30953 4960 30973 4980
rect 31068 4956 31088 4976
rect 31171 4960 31191 4980
rect 31279 4960 31299 4980
rect 31382 4956 31402 4976
rect 3407 4762 3427 4782
rect 3510 4758 3530 4778
rect 3618 4758 3638 4778
rect 3721 4762 3741 4782
rect 3836 4758 3856 4778
rect 3939 4762 3959 4782
rect 4126 4769 4144 4787
rect 190 4707 208 4725
rect 7771 4775 7791 4795
rect 7874 4771 7894 4791
rect 7982 4771 8002 4791
rect 8085 4775 8105 4795
rect 8200 4771 8220 4791
rect 8303 4775 8323 4795
rect 8490 4782 8508 4800
rect 4554 4720 4572 4738
rect 188 4608 206 4626
rect 4124 4670 4142 4688
rect 12148 4787 12168 4807
rect 12251 4783 12271 4803
rect 12359 4783 12379 4803
rect 12462 4787 12482 4807
rect 12577 4783 12597 4803
rect 12680 4787 12700 4807
rect 12867 4794 12885 4812
rect 8931 4732 8949 4750
rect 4552 4621 4570 4639
rect 1456 4522 1476 4542
rect 1559 4526 1579 4546
rect 1674 4522 1694 4542
rect 1777 4526 1797 4546
rect 1885 4526 1905 4546
rect 1988 4522 2008 4542
rect 2610 4534 2630 4554
rect 2713 4530 2733 4550
rect 2821 4530 2841 4550
rect 2924 4534 2944 4554
rect 3039 4530 3059 4550
rect 3142 4534 3162 4554
rect 4119 4551 4137 4569
rect 8488 4683 8506 4701
rect 16512 4800 16532 4820
rect 16615 4796 16635 4816
rect 16723 4796 16743 4816
rect 16826 4800 16846 4820
rect 16941 4796 16961 4816
rect 17044 4800 17064 4820
rect 17231 4807 17249 4825
rect 13295 4745 13313 4763
rect 8929 4633 8947 4651
rect 5820 4535 5840 4555
rect 5923 4539 5943 4559
rect 6038 4535 6058 4555
rect 6141 4539 6161 4559
rect 6249 4539 6269 4559
rect 6352 4535 6372 4555
rect 6974 4547 6994 4567
rect 7077 4543 7097 4563
rect 7185 4543 7205 4563
rect 7288 4547 7308 4567
rect 7403 4543 7423 4563
rect 7506 4547 7526 4567
rect 8483 4564 8501 4582
rect 12865 4695 12883 4713
rect 20778 4774 20798 4794
rect 20881 4770 20901 4790
rect 20989 4770 21009 4790
rect 21092 4774 21112 4794
rect 21207 4770 21227 4790
rect 21310 4774 21330 4794
rect 21497 4781 21515 4799
rect 13293 4646 13311 4664
rect 10197 4547 10217 4567
rect 4117 4452 4135 4470
rect 185 4383 203 4401
rect 10300 4551 10320 4571
rect 10415 4547 10435 4567
rect 10518 4551 10538 4571
rect 10626 4551 10646 4571
rect 10729 4547 10749 4567
rect 11351 4559 11371 4579
rect 11454 4555 11474 4575
rect 11562 4555 11582 4575
rect 11665 4559 11685 4579
rect 11780 4555 11800 4575
rect 11883 4559 11903 4579
rect 12860 4576 12878 4594
rect 17229 4708 17247 4726
rect 17561 4719 17579 4737
rect 25142 4787 25162 4807
rect 25245 4783 25265 4803
rect 25353 4783 25373 4803
rect 25456 4787 25476 4807
rect 25571 4783 25591 4803
rect 25674 4787 25694 4807
rect 25861 4794 25879 4812
rect 21925 4732 21943 4750
rect 14561 4560 14581 4580
rect 8481 4465 8499 4483
rect 3408 4350 3428 4370
rect 183 4284 201 4302
rect 354 4300 374 4320
rect 457 4304 477 4324
rect 572 4300 592 4320
rect 675 4304 695 4324
rect 783 4304 803 4324
rect 3511 4346 3531 4366
rect 3619 4346 3639 4366
rect 3722 4350 3742 4370
rect 3837 4346 3857 4366
rect 3940 4350 3960 4370
rect 4113 4368 4131 4386
rect 4549 4396 4567 4414
rect 886 4300 906 4320
rect 14664 4564 14684 4584
rect 14779 4560 14799 4580
rect 14882 4564 14902 4584
rect 14990 4564 15010 4584
rect 15093 4560 15113 4580
rect 15715 4572 15735 4592
rect 15818 4568 15838 4588
rect 15926 4568 15946 4588
rect 16029 4572 16049 4592
rect 16144 4568 16164 4588
rect 16247 4572 16267 4592
rect 17224 4589 17242 4607
rect 17559 4620 17577 4638
rect 12858 4477 12876 4495
rect 7772 4363 7792 4383
rect 4111 4269 4129 4287
rect 4547 4297 4565 4315
rect 4718 4313 4738 4333
rect 4821 4317 4841 4337
rect 4936 4313 4956 4333
rect 5039 4317 5059 4337
rect 5147 4317 5167 4337
rect 7875 4359 7895 4379
rect 7983 4359 8003 4379
rect 8086 4363 8106 4383
rect 8201 4359 8221 4379
rect 8304 4363 8324 4383
rect 8477 4381 8495 4399
rect 8926 4408 8944 4426
rect 5250 4313 5270 4333
rect 179 4200 197 4218
rect 21495 4682 21513 4700
rect 29519 4799 29539 4819
rect 29622 4795 29642 4815
rect 29730 4795 29750 4815
rect 29833 4799 29853 4819
rect 29948 4795 29968 4815
rect 30051 4799 30071 4819
rect 30238 4806 30256 4824
rect 26302 4744 26320 4762
rect 21923 4633 21941 4651
rect 18827 4534 18847 4554
rect 18930 4538 18950 4558
rect 19045 4534 19065 4554
rect 19148 4538 19168 4558
rect 19256 4538 19276 4558
rect 19359 4534 19379 4554
rect 19981 4546 20001 4566
rect 20084 4542 20104 4562
rect 20192 4542 20212 4562
rect 20295 4546 20315 4566
rect 20410 4542 20430 4562
rect 20513 4546 20533 4566
rect 21490 4563 21508 4581
rect 25859 4695 25877 4713
rect 33883 4812 33903 4832
rect 33986 4808 34006 4828
rect 34094 4808 34114 4828
rect 34197 4812 34217 4832
rect 34312 4808 34332 4828
rect 34415 4812 34435 4832
rect 34602 4819 34620 4837
rect 30666 4757 30684 4775
rect 26300 4645 26318 4663
rect 23191 4547 23211 4567
rect 17222 4490 17240 4508
rect 12149 4375 12169 4395
rect 8475 4282 8493 4300
rect 8924 4309 8942 4327
rect 9095 4325 9115 4345
rect 9198 4329 9218 4349
rect 9313 4325 9333 4345
rect 9416 4329 9436 4349
rect 9524 4329 9544 4349
rect 12252 4371 12272 4391
rect 12360 4371 12380 4391
rect 12463 4375 12483 4395
rect 12578 4371 12598 4391
rect 12681 4375 12701 4395
rect 12854 4393 12872 4411
rect 13290 4421 13308 4439
rect 9627 4325 9647 4345
rect 4543 4213 4561 4231
rect 177 4101 195 4119
rect 1152 4116 1172 4136
rect 1255 4120 1275 4140
rect 1370 4116 1390 4136
rect 1473 4120 1493 4140
rect 1581 4120 1601 4140
rect 1684 4116 1704 4136
rect 2511 4124 2531 4144
rect 2614 4120 2634 4140
rect 2722 4120 2742 4140
rect 2825 4124 2845 4144
rect 2940 4120 2960 4140
rect 16513 4388 16533 4408
rect 12852 4294 12870 4312
rect 13288 4322 13306 4340
rect 13459 4338 13479 4358
rect 13562 4342 13582 4362
rect 13677 4338 13697 4358
rect 13780 4342 13800 4362
rect 13888 4342 13908 4362
rect 16616 4384 16636 4404
rect 16724 4384 16744 4404
rect 16827 4388 16847 4408
rect 16942 4384 16962 4404
rect 17045 4388 17065 4408
rect 17218 4406 17236 4424
rect 23294 4551 23314 4571
rect 23409 4547 23429 4567
rect 23512 4551 23532 4571
rect 23620 4551 23640 4571
rect 23723 4547 23743 4567
rect 24345 4559 24365 4579
rect 24448 4555 24468 4575
rect 24556 4555 24576 4575
rect 24659 4559 24679 4579
rect 24774 4555 24794 4575
rect 24877 4559 24897 4579
rect 25854 4576 25872 4594
rect 30236 4707 30254 4725
rect 30664 4658 30682 4676
rect 27568 4559 27588 4579
rect 21488 4464 21506 4482
rect 13991 4338 14011 4358
rect 8920 4225 8938 4243
rect 3043 4124 3063 4144
rect 4541 4114 4559 4132
rect 5516 4129 5536 4149
rect 172 3982 190 4000
rect 5619 4133 5639 4153
rect 5734 4129 5754 4149
rect 5837 4133 5857 4153
rect 5945 4133 5965 4153
rect 6048 4129 6068 4149
rect 6875 4137 6895 4157
rect 6978 4133 6998 4153
rect 7086 4133 7106 4153
rect 7189 4137 7209 4157
rect 7304 4133 7324 4153
rect 17556 4395 17574 4413
rect 17216 4307 17234 4325
rect 27671 4563 27691 4583
rect 27786 4559 27806 4579
rect 27889 4563 27909 4583
rect 27997 4563 28017 4583
rect 28100 4559 28120 4579
rect 28722 4571 28742 4591
rect 28825 4567 28845 4587
rect 28933 4567 28953 4587
rect 29036 4571 29056 4591
rect 29151 4567 29171 4587
rect 29254 4571 29274 4591
rect 30231 4588 30249 4606
rect 34600 4720 34618 4738
rect 31932 4572 31952 4592
rect 25852 4477 25870 4495
rect 20779 4362 20799 4382
rect 13284 4238 13302 4256
rect 7407 4137 7427 4157
rect 4108 4044 4126 4062
rect 4536 3995 4554 4013
rect 8918 4126 8936 4144
rect 9893 4141 9913 4161
rect 9996 4145 10016 4165
rect 10111 4141 10131 4161
rect 10214 4145 10234 4165
rect 10322 4145 10342 4165
rect 10425 4141 10445 4161
rect 11252 4149 11272 4169
rect 11355 4145 11375 4165
rect 11463 4145 11483 4165
rect 11566 4149 11586 4169
rect 11681 4145 11701 4165
rect 17554 4296 17572 4314
rect 17725 4312 17745 4332
rect 17828 4316 17848 4336
rect 17943 4312 17963 4332
rect 18046 4316 18066 4336
rect 18154 4316 18174 4336
rect 20882 4358 20902 4378
rect 20990 4358 21010 4378
rect 21093 4362 21113 4382
rect 21208 4358 21228 4378
rect 21311 4362 21331 4382
rect 21484 4380 21502 4398
rect 21920 4408 21938 4426
rect 18257 4312 18277 4332
rect 32035 4576 32055 4596
rect 32150 4572 32170 4592
rect 32253 4576 32273 4596
rect 32361 4576 32381 4596
rect 32464 4572 32484 4592
rect 33086 4584 33106 4604
rect 33189 4580 33209 4600
rect 33297 4580 33317 4600
rect 33400 4584 33420 4604
rect 33515 4580 33535 4600
rect 33618 4584 33638 4604
rect 34595 4601 34613 4619
rect 30229 4489 30247 4507
rect 25143 4375 25163 4395
rect 21482 4281 21500 4299
rect 21918 4309 21936 4327
rect 22089 4325 22109 4345
rect 22192 4329 22212 4349
rect 22307 4325 22327 4345
rect 22410 4329 22430 4349
rect 22518 4329 22538 4349
rect 25246 4371 25266 4391
rect 25354 4371 25374 4391
rect 25457 4375 25477 4395
rect 25572 4371 25592 4391
rect 25675 4375 25695 4395
rect 25848 4393 25866 4411
rect 26297 4420 26315 4438
rect 22621 4325 22641 4345
rect 17550 4212 17568 4230
rect 11784 4149 11804 4169
rect 13282 4139 13300 4157
rect 14257 4154 14277 4174
rect 8472 4057 8490 4075
rect 4106 3945 4124 3963
rect 170 3883 188 3901
rect 355 3888 375 3908
rect 458 3892 478 3912
rect 573 3888 593 3908
rect 676 3892 696 3912
rect 784 3892 804 3912
rect 887 3888 907 3908
rect 8913 4007 8931 4025
rect 14360 4158 14380 4178
rect 14475 4154 14495 4174
rect 14578 4158 14598 4178
rect 14686 4158 14706 4178
rect 14789 4154 14809 4174
rect 15616 4162 15636 4182
rect 15719 4158 15739 4178
rect 15827 4158 15847 4178
rect 15930 4162 15950 4182
rect 16045 4158 16065 4178
rect 16148 4162 16168 4182
rect 34593 4502 34611 4520
rect 29520 4387 29540 4407
rect 25846 4294 25864 4312
rect 26295 4321 26313 4339
rect 26466 4337 26486 4357
rect 26569 4341 26589 4361
rect 26684 4337 26704 4357
rect 26787 4341 26807 4361
rect 26895 4341 26915 4361
rect 29623 4383 29643 4403
rect 29731 4383 29751 4403
rect 29834 4387 29854 4407
rect 29949 4383 29969 4403
rect 30052 4387 30072 4407
rect 30225 4405 30243 4423
rect 30661 4433 30679 4451
rect 26998 4337 27018 4357
rect 21914 4225 21932 4243
rect 12849 4069 12867 4087
rect 8470 3958 8488 3976
rect 4534 3896 4552 3914
rect 4719 3901 4739 3921
rect 4822 3905 4842 3925
rect 4937 3901 4957 3921
rect 5040 3905 5060 3925
rect 5148 3905 5168 3925
rect 5251 3901 5271 3921
rect 13277 4020 13295 4038
rect 17213 4082 17231 4100
rect 17548 4113 17566 4131
rect 18523 4128 18543 4148
rect 18626 4132 18646 4152
rect 18741 4128 18761 4148
rect 18844 4132 18864 4152
rect 18952 4132 18972 4152
rect 19055 4128 19075 4148
rect 19882 4136 19902 4156
rect 19985 4132 20005 4152
rect 20093 4132 20113 4152
rect 20196 4136 20216 4156
rect 20311 4132 20331 4152
rect 33884 4400 33904 4420
rect 30223 4306 30241 4324
rect 30659 4334 30677 4352
rect 30830 4350 30850 4370
rect 30933 4354 30953 4374
rect 31048 4350 31068 4370
rect 31151 4354 31171 4374
rect 31259 4354 31279 4374
rect 33987 4396 34007 4416
rect 34095 4396 34115 4416
rect 34198 4400 34218 4420
rect 34313 4396 34333 4416
rect 34416 4400 34436 4420
rect 34589 4418 34607 4436
rect 31362 4350 31382 4370
rect 26291 4237 26309 4255
rect 20414 4136 20434 4156
rect 21912 4126 21930 4144
rect 22887 4141 22907 4161
rect 12847 3970 12865 3988
rect 8911 3908 8929 3926
rect 9096 3913 9116 3933
rect 9199 3917 9219 3937
rect 9314 3913 9334 3933
rect 9417 3917 9437 3937
rect 9525 3917 9545 3937
rect 9628 3913 9648 3933
rect 17211 3983 17229 4001
rect 17543 3994 17561 4012
rect 22990 4145 23010 4165
rect 23105 4141 23125 4161
rect 23208 4145 23228 4165
rect 23316 4145 23336 4165
rect 23419 4141 23439 4161
rect 24246 4149 24266 4169
rect 24349 4145 24369 4165
rect 24457 4145 24477 4165
rect 24560 4149 24580 4169
rect 24675 4145 24695 4165
rect 34587 4319 34605 4337
rect 30655 4250 30673 4268
rect 24778 4149 24798 4169
rect 21479 4056 21497 4074
rect 13275 3921 13293 3939
rect 13460 3926 13480 3946
rect 13563 3930 13583 3950
rect 13678 3926 13698 3946
rect 13781 3930 13801 3950
rect 13889 3930 13909 3950
rect 13992 3926 14012 3946
rect 21907 4007 21925 4025
rect 26289 4138 26307 4156
rect 27264 4153 27284 4173
rect 27367 4157 27387 4177
rect 27482 4153 27502 4173
rect 27585 4157 27605 4177
rect 27693 4157 27713 4177
rect 27796 4153 27816 4173
rect 28623 4161 28643 4181
rect 28726 4157 28746 4177
rect 28834 4157 28854 4177
rect 28937 4161 28957 4181
rect 29052 4157 29072 4177
rect 29155 4161 29175 4181
rect 30653 4151 30671 4169
rect 31628 4166 31648 4186
rect 25843 4069 25861 4087
rect 21477 3957 21495 3975
rect 17541 3895 17559 3913
rect 17726 3900 17746 3920
rect 17829 3904 17849 3924
rect 17944 3900 17964 3920
rect 18047 3904 18067 3924
rect 18155 3904 18175 3924
rect 18258 3900 18278 3920
rect 26284 4019 26302 4037
rect 31731 4170 31751 4190
rect 31846 4166 31866 4186
rect 31949 4170 31969 4190
rect 32057 4170 32077 4190
rect 32160 4166 32180 4186
rect 32987 4174 33007 4194
rect 33090 4170 33110 4190
rect 33198 4170 33218 4190
rect 33301 4174 33321 4194
rect 33416 4170 33436 4190
rect 33519 4174 33539 4194
rect 30220 4081 30238 4099
rect 25841 3970 25859 3988
rect 21905 3908 21923 3926
rect 22090 3913 22110 3933
rect 22193 3917 22213 3937
rect 22308 3913 22328 3933
rect 22411 3917 22431 3937
rect 22519 3917 22539 3937
rect 22622 3913 22642 3933
rect 30648 4032 30666 4050
rect 34584 4094 34602 4112
rect 30218 3982 30236 4000
rect 26282 3920 26300 3938
rect 26467 3925 26487 3945
rect 26570 3929 26590 3949
rect 26685 3925 26705 3945
rect 26788 3929 26808 3949
rect 26896 3929 26916 3949
rect 26999 3925 27019 3945
rect 34582 3995 34600 4013
rect 30646 3933 30664 3951
rect 30831 3938 30851 3958
rect 30934 3942 30954 3962
rect 31049 3938 31069 3958
rect 31152 3942 31172 3962
rect 31260 3942 31280 3962
rect 31363 3938 31383 3958
rect 3390 3744 3410 3764
rect 3493 3740 3513 3760
rect 3601 3740 3621 3760
rect 3704 3744 3724 3764
rect 3819 3740 3839 3760
rect 3922 3744 3942 3764
rect 4109 3751 4127 3769
rect 173 3689 191 3707
rect 7754 3757 7774 3777
rect 7857 3753 7877 3773
rect 7965 3753 7985 3773
rect 8068 3757 8088 3777
rect 8183 3753 8203 3773
rect 8286 3757 8306 3777
rect 8473 3764 8491 3782
rect 4537 3702 4555 3720
rect 171 3590 189 3608
rect 4107 3652 4125 3670
rect 12131 3769 12151 3789
rect 12234 3765 12254 3785
rect 12342 3765 12362 3785
rect 12445 3769 12465 3789
rect 12560 3765 12580 3785
rect 12663 3769 12683 3789
rect 12850 3776 12868 3794
rect 8914 3714 8932 3732
rect 4535 3603 4553 3621
rect 1234 3508 1254 3528
rect 1337 3512 1357 3532
rect 1452 3508 1472 3528
rect 1555 3512 1575 3532
rect 1663 3512 1683 3532
rect 1766 3508 1786 3528
rect 2593 3516 2613 3536
rect 2696 3512 2716 3532
rect 2804 3512 2824 3532
rect 2907 3516 2927 3536
rect 3022 3512 3042 3532
rect 8471 3665 8489 3683
rect 16495 3782 16515 3802
rect 16598 3778 16618 3798
rect 16706 3778 16726 3798
rect 16809 3782 16829 3802
rect 16924 3778 16944 3798
rect 17027 3782 17047 3802
rect 17214 3789 17232 3807
rect 13278 3727 13296 3745
rect 8912 3615 8930 3633
rect 3125 3516 3145 3536
rect 4102 3533 4120 3551
rect 5598 3521 5618 3541
rect 5701 3525 5721 3545
rect 5816 3521 5836 3541
rect 5919 3525 5939 3545
rect 6027 3525 6047 3545
rect 6130 3521 6150 3541
rect 6957 3529 6977 3549
rect 7060 3525 7080 3545
rect 7168 3525 7188 3545
rect 7271 3529 7291 3549
rect 7386 3525 7406 3545
rect 7489 3529 7509 3549
rect 8466 3546 8484 3564
rect 12848 3677 12866 3695
rect 20761 3756 20781 3776
rect 20864 3752 20884 3772
rect 20972 3752 20992 3772
rect 21075 3756 21095 3776
rect 21190 3752 21210 3772
rect 21293 3756 21313 3776
rect 21480 3763 21498 3781
rect 13276 3628 13294 3646
rect 9975 3533 9995 3553
rect 4100 3434 4118 3452
rect 168 3365 186 3383
rect 10078 3537 10098 3557
rect 10193 3533 10213 3553
rect 10296 3537 10316 3557
rect 10404 3537 10424 3557
rect 10507 3533 10527 3553
rect 11334 3541 11354 3561
rect 11437 3537 11457 3557
rect 11545 3537 11565 3557
rect 11648 3541 11668 3561
rect 11763 3537 11783 3557
rect 17212 3690 17230 3708
rect 17544 3701 17562 3719
rect 25125 3769 25145 3789
rect 25228 3765 25248 3785
rect 25336 3765 25356 3785
rect 25439 3769 25459 3789
rect 25554 3765 25574 3785
rect 25657 3769 25677 3789
rect 25844 3776 25862 3794
rect 21908 3714 21926 3732
rect 11866 3541 11886 3561
rect 12843 3558 12861 3576
rect 14339 3546 14359 3566
rect 8464 3447 8482 3465
rect 3391 3332 3411 3352
rect 166 3266 184 3284
rect 337 3282 357 3302
rect 440 3286 460 3306
rect 555 3282 575 3302
rect 658 3286 678 3306
rect 766 3286 786 3306
rect 3494 3328 3514 3348
rect 3602 3328 3622 3348
rect 3705 3332 3725 3352
rect 3820 3328 3840 3348
rect 3923 3332 3943 3352
rect 4096 3350 4114 3368
rect 4532 3378 4550 3396
rect 869 3282 889 3302
rect 14442 3550 14462 3570
rect 14557 3546 14577 3566
rect 14660 3550 14680 3570
rect 14768 3550 14788 3570
rect 14871 3546 14891 3566
rect 15698 3554 15718 3574
rect 15801 3550 15821 3570
rect 15909 3550 15929 3570
rect 16012 3554 16032 3574
rect 16127 3550 16147 3570
rect 16230 3554 16250 3574
rect 17207 3571 17225 3589
rect 17542 3602 17560 3620
rect 21478 3664 21496 3682
rect 29502 3781 29522 3801
rect 29605 3777 29625 3797
rect 29713 3777 29733 3797
rect 29816 3781 29836 3801
rect 29931 3777 29951 3797
rect 30034 3781 30054 3801
rect 30221 3788 30239 3806
rect 26285 3726 26303 3744
rect 21906 3615 21924 3633
rect 12841 3459 12859 3477
rect 7755 3345 7775 3365
rect 4094 3251 4112 3269
rect 4530 3279 4548 3297
rect 4701 3295 4721 3315
rect 4804 3299 4824 3319
rect 4919 3295 4939 3315
rect 5022 3299 5042 3319
rect 5130 3299 5150 3319
rect 7858 3341 7878 3361
rect 7966 3341 7986 3361
rect 8069 3345 8089 3365
rect 8184 3341 8204 3361
rect 8287 3345 8307 3365
rect 8460 3363 8478 3381
rect 8909 3390 8927 3408
rect 5233 3295 5253 3315
rect 162 3182 180 3200
rect 18605 3520 18625 3540
rect 18708 3524 18728 3544
rect 18823 3520 18843 3540
rect 18926 3524 18946 3544
rect 19034 3524 19054 3544
rect 19137 3520 19157 3540
rect 19964 3528 19984 3548
rect 20067 3524 20087 3544
rect 20175 3524 20195 3544
rect 20278 3528 20298 3548
rect 20393 3524 20413 3544
rect 25842 3677 25860 3695
rect 33866 3794 33886 3814
rect 33969 3790 33989 3810
rect 34077 3790 34097 3810
rect 34180 3794 34200 3814
rect 34295 3790 34315 3810
rect 34398 3794 34418 3814
rect 34585 3801 34603 3819
rect 30649 3739 30667 3757
rect 26283 3627 26301 3645
rect 20496 3528 20516 3548
rect 21473 3545 21491 3563
rect 22969 3533 22989 3553
rect 17205 3472 17223 3490
rect 12132 3357 12152 3377
rect 8458 3264 8476 3282
rect 8907 3291 8925 3309
rect 9078 3307 9098 3327
rect 9181 3311 9201 3331
rect 9296 3307 9316 3327
rect 9399 3311 9419 3331
rect 9507 3311 9527 3331
rect 12235 3353 12255 3373
rect 12343 3353 12363 3373
rect 12446 3357 12466 3377
rect 12561 3353 12581 3373
rect 12664 3357 12684 3377
rect 12837 3375 12855 3393
rect 13273 3403 13291 3421
rect 9610 3307 9630 3327
rect 4526 3195 4544 3213
rect 160 3083 178 3101
rect 1135 3098 1155 3118
rect 1238 3102 1258 3122
rect 1353 3098 1373 3118
rect 1456 3102 1476 3122
rect 1564 3102 1584 3122
rect 1667 3098 1687 3118
rect 2428 3108 2448 3128
rect 2531 3104 2551 3124
rect 2639 3104 2659 3124
rect 2742 3108 2762 3128
rect 2857 3104 2877 3124
rect 16496 3370 16516 3390
rect 12835 3276 12853 3294
rect 13271 3304 13289 3322
rect 13442 3320 13462 3340
rect 13545 3324 13565 3344
rect 13660 3320 13680 3340
rect 13763 3324 13783 3344
rect 13871 3324 13891 3344
rect 16599 3366 16619 3386
rect 16707 3366 16727 3386
rect 16810 3370 16830 3390
rect 16925 3366 16945 3386
rect 17028 3370 17048 3390
rect 17201 3388 17219 3406
rect 23072 3537 23092 3557
rect 23187 3533 23207 3553
rect 23290 3537 23310 3557
rect 23398 3537 23418 3557
rect 23501 3533 23521 3553
rect 24328 3541 24348 3561
rect 24431 3537 24451 3557
rect 24539 3537 24559 3557
rect 24642 3541 24662 3561
rect 24757 3537 24777 3557
rect 24860 3541 24880 3561
rect 25837 3558 25855 3576
rect 30219 3689 30237 3707
rect 30647 3640 30665 3658
rect 27346 3545 27366 3565
rect 21471 3446 21489 3464
rect 13974 3320 13994 3340
rect 8903 3207 8921 3225
rect 2960 3108 2980 3128
rect 155 2964 173 2982
rect 4524 3096 4542 3114
rect 5499 3111 5519 3131
rect 5602 3115 5622 3135
rect 5717 3111 5737 3131
rect 5820 3115 5840 3135
rect 5928 3115 5948 3135
rect 6031 3111 6051 3131
rect 6792 3121 6812 3141
rect 6895 3117 6915 3137
rect 7003 3117 7023 3137
rect 7106 3121 7126 3141
rect 7221 3117 7241 3137
rect 17539 3377 17557 3395
rect 17199 3289 17217 3307
rect 27449 3549 27469 3569
rect 27564 3545 27584 3565
rect 27667 3549 27687 3569
rect 27775 3549 27795 3569
rect 27878 3545 27898 3565
rect 28705 3553 28725 3573
rect 28808 3549 28828 3569
rect 28916 3549 28936 3569
rect 29019 3553 29039 3573
rect 29134 3549 29154 3569
rect 34583 3702 34601 3720
rect 29237 3553 29257 3573
rect 30214 3570 30232 3588
rect 31710 3558 31730 3578
rect 25835 3459 25853 3477
rect 20762 3344 20782 3364
rect 13267 3220 13285 3238
rect 7324 3121 7344 3141
rect 4091 3026 4109 3044
rect 4519 2977 4537 2995
rect 8901 3108 8919 3126
rect 9876 3123 9896 3143
rect 9979 3127 9999 3147
rect 10094 3123 10114 3143
rect 10197 3127 10217 3147
rect 10305 3127 10325 3147
rect 10408 3123 10428 3143
rect 11169 3133 11189 3153
rect 11272 3129 11292 3149
rect 11380 3129 11400 3149
rect 11483 3133 11503 3153
rect 11598 3129 11618 3149
rect 17537 3278 17555 3296
rect 17708 3294 17728 3314
rect 17811 3298 17831 3318
rect 17926 3294 17946 3314
rect 18029 3298 18049 3318
rect 18137 3298 18157 3318
rect 20865 3340 20885 3360
rect 20973 3340 20993 3360
rect 21076 3344 21096 3364
rect 21191 3340 21211 3360
rect 21294 3344 21314 3364
rect 21467 3362 21485 3380
rect 21903 3390 21921 3408
rect 18240 3294 18260 3314
rect 31813 3562 31833 3582
rect 31928 3558 31948 3578
rect 32031 3562 32051 3582
rect 32139 3562 32159 3582
rect 32242 3558 32262 3578
rect 33069 3566 33089 3586
rect 33172 3562 33192 3582
rect 33280 3562 33300 3582
rect 33383 3566 33403 3586
rect 33498 3562 33518 3582
rect 33601 3566 33621 3586
rect 34578 3583 34596 3601
rect 30212 3471 30230 3489
rect 25126 3357 25146 3377
rect 21465 3263 21483 3281
rect 21901 3291 21919 3309
rect 22072 3307 22092 3327
rect 22175 3311 22195 3331
rect 22290 3307 22310 3327
rect 22393 3311 22413 3331
rect 22501 3311 22521 3331
rect 25229 3353 25249 3373
rect 25337 3353 25357 3373
rect 25440 3357 25460 3377
rect 25555 3353 25575 3373
rect 25658 3357 25678 3377
rect 25831 3375 25849 3393
rect 26280 3402 26298 3420
rect 22604 3307 22624 3327
rect 17533 3194 17551 3212
rect 11701 3133 11721 3153
rect 8455 3039 8473 3057
rect 4089 2927 4107 2945
rect 153 2865 171 2883
rect 338 2870 358 2890
rect 441 2874 461 2894
rect 556 2870 576 2890
rect 659 2874 679 2894
rect 767 2874 787 2894
rect 870 2870 890 2890
rect 8896 2989 8914 3007
rect 13265 3121 13283 3139
rect 14240 3136 14260 3156
rect 14343 3140 14363 3160
rect 14458 3136 14478 3156
rect 14561 3140 14581 3160
rect 14669 3140 14689 3160
rect 14772 3136 14792 3156
rect 15533 3146 15553 3166
rect 15636 3142 15656 3162
rect 15744 3142 15764 3162
rect 15847 3146 15867 3166
rect 15962 3142 15982 3162
rect 16065 3146 16085 3166
rect 34576 3484 34594 3502
rect 29503 3369 29523 3389
rect 25829 3276 25847 3294
rect 26278 3303 26296 3321
rect 26449 3319 26469 3339
rect 26552 3323 26572 3343
rect 26667 3319 26687 3339
rect 26770 3323 26790 3343
rect 26878 3323 26898 3343
rect 29606 3365 29626 3385
rect 29714 3365 29734 3385
rect 29817 3369 29837 3389
rect 29932 3365 29952 3385
rect 30035 3369 30055 3389
rect 30208 3387 30226 3405
rect 30644 3415 30662 3433
rect 26981 3319 27001 3339
rect 21897 3207 21915 3225
rect 12832 3051 12850 3069
rect 8453 2940 8471 2958
rect 4517 2878 4535 2896
rect 4702 2883 4722 2903
rect 4805 2887 4825 2907
rect 4920 2883 4940 2903
rect 5023 2887 5043 2907
rect 5131 2887 5151 2907
rect 5234 2883 5254 2903
rect 13260 3002 13278 3020
rect 17196 3064 17214 3082
rect 17531 3095 17549 3113
rect 18506 3110 18526 3130
rect 18609 3114 18629 3134
rect 18724 3110 18744 3130
rect 18827 3114 18847 3134
rect 18935 3114 18955 3134
rect 19038 3110 19058 3130
rect 19799 3120 19819 3140
rect 19902 3116 19922 3136
rect 20010 3116 20030 3136
rect 20113 3120 20133 3140
rect 20228 3116 20248 3136
rect 33867 3382 33887 3402
rect 30206 3288 30224 3306
rect 30642 3316 30660 3334
rect 30813 3332 30833 3352
rect 30916 3336 30936 3356
rect 31031 3332 31051 3352
rect 31134 3336 31154 3356
rect 31242 3336 31262 3356
rect 33970 3378 33990 3398
rect 34078 3378 34098 3398
rect 34181 3382 34201 3402
rect 34296 3378 34316 3398
rect 34399 3382 34419 3402
rect 34572 3400 34590 3418
rect 31345 3332 31365 3352
rect 26274 3219 26292 3237
rect 20331 3120 20351 3140
rect 12830 2952 12848 2970
rect 8894 2890 8912 2908
rect 9079 2895 9099 2915
rect 9182 2899 9202 2919
rect 9297 2895 9317 2915
rect 9400 2899 9420 2919
rect 9508 2899 9528 2919
rect 9611 2895 9631 2915
rect 17194 2965 17212 2983
rect 17526 2976 17544 2994
rect 21895 3108 21913 3126
rect 22870 3123 22890 3143
rect 22973 3127 22993 3147
rect 23088 3123 23108 3143
rect 23191 3127 23211 3147
rect 23299 3127 23319 3147
rect 23402 3123 23422 3143
rect 24163 3133 24183 3153
rect 24266 3129 24286 3149
rect 24374 3129 24394 3149
rect 24477 3133 24497 3153
rect 24592 3129 24612 3149
rect 34570 3301 34588 3319
rect 30638 3232 30656 3250
rect 24695 3133 24715 3153
rect 21462 3038 21480 3056
rect 13258 2903 13276 2921
rect 13443 2908 13463 2928
rect 13546 2912 13566 2932
rect 13661 2908 13681 2928
rect 13764 2912 13784 2932
rect 13872 2912 13892 2932
rect 13975 2908 13995 2928
rect 21890 2989 21908 3007
rect 26272 3120 26290 3138
rect 27247 3135 27267 3155
rect 27350 3139 27370 3159
rect 27465 3135 27485 3155
rect 27568 3139 27588 3159
rect 27676 3139 27696 3159
rect 27779 3135 27799 3155
rect 28540 3145 28560 3165
rect 28643 3141 28663 3161
rect 28751 3141 28771 3161
rect 28854 3145 28874 3165
rect 28969 3141 28989 3161
rect 29072 3145 29092 3165
rect 25826 3051 25844 3069
rect 21460 2939 21478 2957
rect 17524 2877 17542 2895
rect 17709 2882 17729 2902
rect 17812 2886 17832 2906
rect 17927 2882 17947 2902
rect 18030 2886 18050 2906
rect 18138 2886 18158 2906
rect 18241 2882 18261 2902
rect 26267 3001 26285 3019
rect 30636 3133 30654 3151
rect 31611 3148 31631 3168
rect 31714 3152 31734 3172
rect 31829 3148 31849 3168
rect 31932 3152 31952 3172
rect 32040 3152 32060 3172
rect 32143 3148 32163 3168
rect 32904 3158 32924 3178
rect 33007 3154 33027 3174
rect 33115 3154 33135 3174
rect 33218 3158 33238 3178
rect 33333 3154 33353 3174
rect 33436 3158 33456 3178
rect 30203 3063 30221 3081
rect 25824 2952 25842 2970
rect 21888 2890 21906 2908
rect 22073 2895 22093 2915
rect 22176 2899 22196 2919
rect 22291 2895 22311 2915
rect 22394 2899 22414 2919
rect 22502 2899 22522 2919
rect 22605 2895 22625 2915
rect 30631 3014 30649 3032
rect 34567 3076 34585 3094
rect 30201 2964 30219 2982
rect 26265 2902 26283 2920
rect 26450 2907 26470 2927
rect 26553 2911 26573 2931
rect 26668 2907 26688 2927
rect 26771 2911 26791 2931
rect 26879 2911 26899 2931
rect 26982 2907 27002 2927
rect 34565 2977 34583 2995
rect 30629 2915 30647 2933
rect 30814 2920 30834 2940
rect 30917 2924 30937 2944
rect 31032 2920 31052 2940
rect 31135 2924 31155 2944
rect 31243 2924 31263 2944
rect 31346 2920 31366 2940
rect 3370 2726 3390 2746
rect 3473 2722 3493 2742
rect 3581 2722 3601 2742
rect 3684 2726 3704 2746
rect 3799 2722 3819 2742
rect 3902 2726 3922 2746
rect 4089 2733 4107 2751
rect 153 2671 171 2689
rect 7734 2739 7754 2759
rect 7837 2735 7857 2755
rect 7945 2735 7965 2755
rect 8048 2739 8068 2759
rect 8163 2735 8183 2755
rect 8266 2739 8286 2759
rect 8453 2746 8471 2764
rect 4517 2684 4535 2702
rect 151 2572 169 2590
rect 4087 2634 4105 2652
rect 12111 2751 12131 2771
rect 12214 2747 12234 2767
rect 12322 2747 12342 2767
rect 12425 2751 12445 2771
rect 12540 2747 12560 2767
rect 12643 2751 12663 2771
rect 12830 2758 12848 2776
rect 8894 2696 8912 2714
rect 4515 2585 4533 2603
rect 1280 2488 1300 2508
rect 1383 2492 1403 2512
rect 1498 2488 1518 2508
rect 1601 2492 1621 2512
rect 1709 2492 1729 2512
rect 1812 2488 1832 2508
rect 2573 2498 2593 2518
rect 2676 2494 2696 2514
rect 2784 2494 2804 2514
rect 2887 2498 2907 2518
rect 3002 2494 3022 2514
rect 3105 2498 3125 2518
rect 4082 2515 4100 2533
rect 8451 2647 8469 2665
rect 16475 2764 16495 2784
rect 16578 2760 16598 2780
rect 16686 2760 16706 2780
rect 16789 2764 16809 2784
rect 16904 2760 16924 2780
rect 17007 2764 17027 2784
rect 17194 2771 17212 2789
rect 13258 2709 13276 2727
rect 8892 2597 8910 2615
rect 5644 2501 5664 2521
rect 5747 2505 5767 2525
rect 5862 2501 5882 2521
rect 5965 2505 5985 2525
rect 6073 2505 6093 2525
rect 6176 2501 6196 2521
rect 6937 2511 6957 2531
rect 7040 2507 7060 2527
rect 7148 2507 7168 2527
rect 7251 2511 7271 2531
rect 7366 2507 7386 2527
rect 7469 2511 7489 2531
rect 8446 2528 8464 2546
rect 12828 2659 12846 2677
rect 20741 2738 20761 2758
rect 20844 2734 20864 2754
rect 20952 2734 20972 2754
rect 21055 2738 21075 2758
rect 21170 2734 21190 2754
rect 21273 2738 21293 2758
rect 21460 2745 21478 2763
rect 13256 2610 13274 2628
rect 10021 2513 10041 2533
rect 4080 2416 4098 2434
rect 148 2347 166 2365
rect 10124 2517 10144 2537
rect 10239 2513 10259 2533
rect 10342 2517 10362 2537
rect 10450 2517 10470 2537
rect 10553 2513 10573 2533
rect 11314 2523 11334 2543
rect 11417 2519 11437 2539
rect 11525 2519 11545 2539
rect 11628 2523 11648 2543
rect 11743 2519 11763 2539
rect 11846 2523 11866 2543
rect 12823 2540 12841 2558
rect 17192 2672 17210 2690
rect 17524 2683 17542 2701
rect 25105 2751 25125 2771
rect 25208 2747 25228 2767
rect 25316 2747 25336 2767
rect 25419 2751 25439 2771
rect 25534 2747 25554 2767
rect 25637 2751 25657 2771
rect 25824 2758 25842 2776
rect 21888 2696 21906 2714
rect 14385 2526 14405 2546
rect 8444 2429 8462 2447
rect 3371 2314 3391 2334
rect 146 2248 164 2266
rect 317 2264 337 2284
rect 420 2268 440 2288
rect 535 2264 555 2284
rect 638 2268 658 2288
rect 746 2268 766 2288
rect 3474 2310 3494 2330
rect 3582 2310 3602 2330
rect 3685 2314 3705 2334
rect 3800 2310 3820 2330
rect 3903 2314 3923 2334
rect 4076 2332 4094 2350
rect 4512 2360 4530 2378
rect 849 2264 869 2284
rect 14488 2530 14508 2550
rect 14603 2526 14623 2546
rect 14706 2530 14726 2550
rect 14814 2530 14834 2550
rect 14917 2526 14937 2546
rect 15678 2536 15698 2556
rect 15781 2532 15801 2552
rect 15889 2532 15909 2552
rect 15992 2536 16012 2556
rect 16107 2532 16127 2552
rect 16210 2536 16230 2556
rect 17187 2553 17205 2571
rect 17522 2584 17540 2602
rect 21458 2646 21476 2664
rect 29482 2763 29502 2783
rect 29585 2759 29605 2779
rect 29693 2759 29713 2779
rect 29796 2763 29816 2783
rect 29911 2759 29931 2779
rect 30014 2763 30034 2783
rect 30201 2770 30219 2788
rect 26265 2708 26283 2726
rect 21886 2597 21904 2615
rect 12821 2441 12839 2459
rect 7735 2327 7755 2347
rect 4074 2233 4092 2251
rect 4510 2261 4528 2279
rect 4681 2277 4701 2297
rect 4784 2281 4804 2301
rect 4899 2277 4919 2297
rect 5002 2281 5022 2301
rect 5110 2281 5130 2301
rect 7838 2323 7858 2343
rect 7946 2323 7966 2343
rect 8049 2327 8069 2347
rect 8164 2323 8184 2343
rect 8267 2327 8287 2347
rect 8440 2345 8458 2363
rect 8889 2372 8907 2390
rect 5213 2277 5233 2297
rect 142 2164 160 2182
rect 18651 2500 18671 2520
rect 18754 2504 18774 2524
rect 18869 2500 18889 2520
rect 18972 2504 18992 2524
rect 19080 2504 19100 2524
rect 19183 2500 19203 2520
rect 19944 2510 19964 2530
rect 20047 2506 20067 2526
rect 20155 2506 20175 2526
rect 20258 2510 20278 2530
rect 20373 2506 20393 2526
rect 20476 2510 20496 2530
rect 21453 2527 21471 2545
rect 25822 2659 25840 2677
rect 33846 2776 33866 2796
rect 33949 2772 33969 2792
rect 34057 2772 34077 2792
rect 34160 2776 34180 2796
rect 34275 2772 34295 2792
rect 34378 2776 34398 2796
rect 34565 2783 34583 2801
rect 30629 2721 30647 2739
rect 26263 2609 26281 2627
rect 23015 2513 23035 2533
rect 17185 2454 17203 2472
rect 12112 2339 12132 2359
rect 8438 2246 8456 2264
rect 8887 2273 8905 2291
rect 9058 2289 9078 2309
rect 9161 2293 9181 2313
rect 9276 2289 9296 2309
rect 9379 2293 9399 2313
rect 9487 2293 9507 2313
rect 12215 2335 12235 2355
rect 12323 2335 12343 2355
rect 12426 2339 12446 2359
rect 12541 2335 12561 2355
rect 12644 2339 12664 2359
rect 12817 2357 12835 2375
rect 13253 2385 13271 2403
rect 9590 2289 9610 2309
rect 4506 2177 4524 2195
rect 140 2065 158 2083
rect 1115 2080 1135 2100
rect 1218 2084 1238 2104
rect 1333 2080 1353 2100
rect 1436 2084 1456 2104
rect 1544 2084 1564 2104
rect 1647 2080 1667 2100
rect 2474 2088 2494 2108
rect 2577 2084 2597 2104
rect 2685 2084 2705 2104
rect 2788 2088 2808 2108
rect 2903 2084 2923 2104
rect 16476 2352 16496 2372
rect 12815 2258 12833 2276
rect 13251 2286 13269 2304
rect 13422 2302 13442 2322
rect 13525 2306 13545 2326
rect 13640 2302 13660 2322
rect 13743 2306 13763 2326
rect 13851 2306 13871 2326
rect 16579 2348 16599 2368
rect 16687 2348 16707 2368
rect 16790 2352 16810 2372
rect 16905 2348 16925 2368
rect 17008 2352 17028 2372
rect 17181 2370 17199 2388
rect 23118 2517 23138 2537
rect 23233 2513 23253 2533
rect 23336 2517 23356 2537
rect 23444 2517 23464 2537
rect 23547 2513 23567 2533
rect 24308 2523 24328 2543
rect 24411 2519 24431 2539
rect 24519 2519 24539 2539
rect 24622 2523 24642 2543
rect 24737 2519 24757 2539
rect 24840 2523 24860 2543
rect 25817 2540 25835 2558
rect 30199 2671 30217 2689
rect 30627 2622 30645 2640
rect 27392 2525 27412 2545
rect 21451 2428 21469 2446
rect 13954 2302 13974 2322
rect 8883 2189 8901 2207
rect 3006 2088 3026 2108
rect 4504 2078 4522 2096
rect 5479 2093 5499 2113
rect 135 1946 153 1964
rect 5582 2097 5602 2117
rect 5697 2093 5717 2113
rect 5800 2097 5820 2117
rect 5908 2097 5928 2117
rect 6011 2093 6031 2113
rect 6838 2101 6858 2121
rect 6941 2097 6961 2117
rect 7049 2097 7069 2117
rect 7152 2101 7172 2121
rect 7267 2097 7287 2117
rect 17519 2359 17537 2377
rect 17179 2271 17197 2289
rect 27495 2529 27515 2549
rect 27610 2525 27630 2545
rect 27713 2529 27733 2549
rect 27821 2529 27841 2549
rect 27924 2525 27944 2545
rect 28685 2535 28705 2555
rect 28788 2531 28808 2551
rect 28896 2531 28916 2551
rect 28999 2535 29019 2555
rect 29114 2531 29134 2551
rect 29217 2535 29237 2555
rect 30194 2552 30212 2570
rect 34563 2684 34581 2702
rect 31756 2538 31776 2558
rect 25815 2441 25833 2459
rect 20742 2326 20762 2346
rect 13247 2202 13265 2220
rect 7370 2101 7390 2121
rect 4071 2008 4089 2026
rect 4499 1959 4517 1977
rect 8881 2090 8899 2108
rect 9856 2105 9876 2125
rect 9959 2109 9979 2129
rect 10074 2105 10094 2125
rect 10177 2109 10197 2129
rect 10285 2109 10305 2129
rect 10388 2105 10408 2125
rect 11215 2113 11235 2133
rect 11318 2109 11338 2129
rect 11426 2109 11446 2129
rect 11529 2113 11549 2133
rect 11644 2109 11664 2129
rect 17517 2260 17535 2278
rect 17688 2276 17708 2296
rect 17791 2280 17811 2300
rect 17906 2276 17926 2296
rect 18009 2280 18029 2300
rect 18117 2280 18137 2300
rect 20845 2322 20865 2342
rect 20953 2322 20973 2342
rect 21056 2326 21076 2346
rect 21171 2322 21191 2342
rect 21274 2326 21294 2346
rect 21447 2344 21465 2362
rect 21883 2372 21901 2390
rect 18220 2276 18240 2296
rect 31859 2542 31879 2562
rect 31974 2538 31994 2558
rect 32077 2542 32097 2562
rect 32185 2542 32205 2562
rect 32288 2538 32308 2558
rect 33049 2548 33069 2568
rect 33152 2544 33172 2564
rect 33260 2544 33280 2564
rect 33363 2548 33383 2568
rect 33478 2544 33498 2564
rect 33581 2548 33601 2568
rect 34558 2565 34576 2583
rect 30192 2453 30210 2471
rect 25106 2339 25126 2359
rect 21445 2245 21463 2263
rect 21881 2273 21899 2291
rect 22052 2289 22072 2309
rect 22155 2293 22175 2313
rect 22270 2289 22290 2309
rect 22373 2293 22393 2313
rect 22481 2293 22501 2313
rect 25209 2335 25229 2355
rect 25317 2335 25337 2355
rect 25420 2339 25440 2359
rect 25535 2335 25555 2355
rect 25638 2339 25658 2359
rect 25811 2357 25829 2375
rect 26260 2384 26278 2402
rect 22584 2289 22604 2309
rect 17513 2176 17531 2194
rect 11747 2113 11767 2133
rect 13245 2103 13263 2121
rect 14220 2118 14240 2138
rect 8435 2021 8453 2039
rect 4069 1909 4087 1927
rect 133 1847 151 1865
rect 318 1852 338 1872
rect 421 1856 441 1876
rect 536 1852 556 1872
rect 639 1856 659 1876
rect 747 1856 767 1876
rect 850 1852 870 1872
rect 8876 1971 8894 1989
rect 14323 2122 14343 2142
rect 14438 2118 14458 2138
rect 14541 2122 14561 2142
rect 14649 2122 14669 2142
rect 14752 2118 14772 2138
rect 15579 2126 15599 2146
rect 15682 2122 15702 2142
rect 15790 2122 15810 2142
rect 15893 2126 15913 2146
rect 16008 2122 16028 2142
rect 16111 2126 16131 2146
rect 34556 2466 34574 2484
rect 29483 2351 29503 2371
rect 25809 2258 25827 2276
rect 26258 2285 26276 2303
rect 26429 2301 26449 2321
rect 26532 2305 26552 2325
rect 26647 2301 26667 2321
rect 26750 2305 26770 2325
rect 26858 2305 26878 2325
rect 29586 2347 29606 2367
rect 29694 2347 29714 2367
rect 29797 2351 29817 2371
rect 29912 2347 29932 2367
rect 30015 2351 30035 2371
rect 30188 2369 30206 2387
rect 30624 2397 30642 2415
rect 26961 2301 26981 2321
rect 21877 2189 21895 2207
rect 12812 2033 12830 2051
rect 8433 1922 8451 1940
rect 4497 1860 4515 1878
rect 4682 1865 4702 1885
rect 4785 1869 4805 1889
rect 4900 1865 4920 1885
rect 5003 1869 5023 1889
rect 5111 1869 5131 1889
rect 5214 1865 5234 1885
rect 13240 1984 13258 2002
rect 17176 2046 17194 2064
rect 17511 2077 17529 2095
rect 18486 2092 18506 2112
rect 18589 2096 18609 2116
rect 18704 2092 18724 2112
rect 18807 2096 18827 2116
rect 18915 2096 18935 2116
rect 19018 2092 19038 2112
rect 19845 2100 19865 2120
rect 19948 2096 19968 2116
rect 20056 2096 20076 2116
rect 20159 2100 20179 2120
rect 20274 2096 20294 2116
rect 33847 2364 33867 2384
rect 30186 2270 30204 2288
rect 30622 2298 30640 2316
rect 30793 2314 30813 2334
rect 30896 2318 30916 2338
rect 31011 2314 31031 2334
rect 31114 2318 31134 2338
rect 31222 2318 31242 2338
rect 33950 2360 33970 2380
rect 34058 2360 34078 2380
rect 34161 2364 34181 2384
rect 34276 2360 34296 2380
rect 34379 2364 34399 2384
rect 34552 2382 34570 2400
rect 31325 2314 31345 2334
rect 26254 2201 26272 2219
rect 20377 2100 20397 2120
rect 21875 2090 21893 2108
rect 22850 2105 22870 2125
rect 12810 1934 12828 1952
rect 8874 1872 8892 1890
rect 9059 1877 9079 1897
rect 9162 1881 9182 1901
rect 9277 1877 9297 1897
rect 9380 1881 9400 1901
rect 9488 1881 9508 1901
rect 9591 1877 9611 1897
rect 17174 1947 17192 1965
rect 17506 1958 17524 1976
rect 22953 2109 22973 2129
rect 23068 2105 23088 2125
rect 23171 2109 23191 2129
rect 23279 2109 23299 2129
rect 23382 2105 23402 2125
rect 24209 2113 24229 2133
rect 24312 2109 24332 2129
rect 24420 2109 24440 2129
rect 24523 2113 24543 2133
rect 24638 2109 24658 2129
rect 34550 2283 34568 2301
rect 30618 2214 30636 2232
rect 24741 2113 24761 2133
rect 21442 2020 21460 2038
rect 13238 1885 13256 1903
rect 13423 1890 13443 1910
rect 13526 1894 13546 1914
rect 13641 1890 13661 1910
rect 13744 1894 13764 1914
rect 13852 1894 13872 1914
rect 13955 1890 13975 1910
rect 21870 1971 21888 1989
rect 26252 2102 26270 2120
rect 27227 2117 27247 2137
rect 27330 2121 27350 2141
rect 27445 2117 27465 2137
rect 27548 2121 27568 2141
rect 27656 2121 27676 2141
rect 27759 2117 27779 2137
rect 28586 2125 28606 2145
rect 28689 2121 28709 2141
rect 28797 2121 28817 2141
rect 28900 2125 28920 2145
rect 29015 2121 29035 2141
rect 29118 2125 29138 2145
rect 30616 2115 30634 2133
rect 31591 2130 31611 2150
rect 25806 2033 25824 2051
rect 21440 1921 21458 1939
rect 17504 1859 17522 1877
rect 17689 1864 17709 1884
rect 17792 1868 17812 1888
rect 17907 1864 17927 1884
rect 18010 1868 18030 1888
rect 18118 1868 18138 1888
rect 18221 1864 18241 1884
rect 26247 1983 26265 2001
rect 31694 2134 31714 2154
rect 31809 2130 31829 2150
rect 31912 2134 31932 2154
rect 32020 2134 32040 2154
rect 32123 2130 32143 2150
rect 32950 2138 32970 2158
rect 33053 2134 33073 2154
rect 33161 2134 33181 2154
rect 33264 2138 33284 2158
rect 33379 2134 33399 2154
rect 33482 2138 33502 2158
rect 30183 2045 30201 2063
rect 25804 1934 25822 1952
rect 21868 1872 21886 1890
rect 22053 1877 22073 1897
rect 22156 1881 22176 1901
rect 22271 1877 22291 1897
rect 22374 1881 22394 1901
rect 22482 1881 22502 1901
rect 22585 1877 22605 1897
rect 30611 1996 30629 2014
rect 34547 2058 34565 2076
rect 30181 1946 30199 1964
rect 26245 1884 26263 1902
rect 26430 1889 26450 1909
rect 26533 1893 26553 1913
rect 26648 1889 26668 1909
rect 26751 1893 26771 1913
rect 26859 1893 26879 1913
rect 26962 1889 26982 1909
rect 34545 1959 34563 1977
rect 30609 1897 30627 1915
rect 30794 1902 30814 1922
rect 30897 1906 30917 1926
rect 31012 1902 31032 1922
rect 31115 1906 31135 1926
rect 31223 1906 31243 1926
rect 31326 1902 31346 1922
rect 3353 1708 3373 1728
rect 3456 1704 3476 1724
rect 3564 1704 3584 1724
rect 3667 1708 3687 1728
rect 3782 1704 3802 1724
rect 3885 1708 3905 1728
rect 4072 1715 4090 1733
rect 136 1653 154 1671
rect 7717 1721 7737 1741
rect 7820 1717 7840 1737
rect 7928 1717 7948 1737
rect 8031 1721 8051 1741
rect 8146 1717 8166 1737
rect 8249 1721 8269 1741
rect 8436 1728 8454 1746
rect 4500 1666 4518 1684
rect 134 1554 152 1572
rect 4070 1616 4088 1634
rect 12094 1733 12114 1753
rect 12197 1729 12217 1749
rect 12305 1729 12325 1749
rect 12408 1733 12428 1753
rect 12523 1729 12543 1749
rect 12626 1733 12646 1753
rect 12813 1740 12831 1758
rect 8877 1678 8895 1696
rect 4498 1567 4516 1585
rect 1197 1472 1217 1492
rect 1300 1476 1320 1496
rect 1415 1472 1435 1492
rect 1518 1476 1538 1496
rect 1626 1476 1646 1496
rect 1729 1472 1749 1492
rect 2556 1480 2576 1500
rect 2659 1476 2679 1496
rect 2767 1476 2787 1496
rect 2870 1480 2890 1500
rect 2985 1476 3005 1496
rect 8434 1629 8452 1647
rect 16458 1746 16478 1766
rect 16561 1742 16581 1762
rect 16669 1742 16689 1762
rect 16772 1746 16792 1766
rect 16887 1742 16907 1762
rect 16990 1746 17010 1766
rect 17177 1753 17195 1771
rect 13241 1691 13259 1709
rect 8875 1579 8893 1597
rect 3088 1480 3108 1500
rect 4065 1497 4083 1515
rect 5561 1485 5581 1505
rect 5664 1489 5684 1509
rect 5779 1485 5799 1505
rect 5882 1489 5902 1509
rect 5990 1489 6010 1509
rect 6093 1485 6113 1505
rect 6920 1493 6940 1513
rect 7023 1489 7043 1509
rect 7131 1489 7151 1509
rect 7234 1493 7254 1513
rect 7349 1489 7369 1509
rect 7452 1493 7472 1513
rect 8429 1510 8447 1528
rect 12811 1641 12829 1659
rect 20724 1720 20744 1740
rect 20827 1716 20847 1736
rect 20935 1716 20955 1736
rect 21038 1720 21058 1740
rect 21153 1716 21173 1736
rect 21256 1720 21276 1740
rect 21443 1727 21461 1745
rect 13239 1592 13257 1610
rect 9938 1497 9958 1517
rect 4063 1398 4081 1416
rect 131 1329 149 1347
rect 10041 1501 10061 1521
rect 10156 1497 10176 1517
rect 10259 1501 10279 1521
rect 10367 1501 10387 1521
rect 10470 1497 10490 1517
rect 11297 1505 11317 1525
rect 11400 1501 11420 1521
rect 11508 1501 11528 1521
rect 11611 1505 11631 1525
rect 11726 1501 11746 1521
rect 17175 1654 17193 1672
rect 17507 1665 17525 1683
rect 25088 1733 25108 1753
rect 25191 1729 25211 1749
rect 25299 1729 25319 1749
rect 25402 1733 25422 1753
rect 25517 1729 25537 1749
rect 25620 1733 25640 1753
rect 25807 1740 25825 1758
rect 21871 1678 21889 1696
rect 11829 1505 11849 1525
rect 12806 1522 12824 1540
rect 14302 1510 14322 1530
rect 8427 1411 8445 1429
rect 3354 1296 3374 1316
rect 129 1230 147 1248
rect 300 1246 320 1266
rect 403 1250 423 1270
rect 518 1246 538 1266
rect 621 1250 641 1270
rect 729 1250 749 1270
rect 3457 1292 3477 1312
rect 3565 1292 3585 1312
rect 3668 1296 3688 1316
rect 3783 1292 3803 1312
rect 3886 1296 3906 1316
rect 4059 1314 4077 1332
rect 4495 1342 4513 1360
rect 832 1246 852 1266
rect 14405 1514 14425 1534
rect 14520 1510 14540 1530
rect 14623 1514 14643 1534
rect 14731 1514 14751 1534
rect 14834 1510 14854 1530
rect 15661 1518 15681 1538
rect 15764 1514 15784 1534
rect 15872 1514 15892 1534
rect 15975 1518 15995 1538
rect 16090 1514 16110 1534
rect 16193 1518 16213 1538
rect 17170 1535 17188 1553
rect 17505 1566 17523 1584
rect 21441 1628 21459 1646
rect 29465 1745 29485 1765
rect 29568 1741 29588 1761
rect 29676 1741 29696 1761
rect 29779 1745 29799 1765
rect 29894 1741 29914 1761
rect 29997 1745 30017 1765
rect 30184 1752 30202 1770
rect 26248 1690 26266 1708
rect 21869 1579 21887 1597
rect 12804 1423 12822 1441
rect 7718 1309 7738 1329
rect 4057 1215 4075 1233
rect 4493 1243 4511 1261
rect 4664 1259 4684 1279
rect 4767 1263 4787 1283
rect 4882 1259 4902 1279
rect 4985 1263 5005 1283
rect 5093 1263 5113 1283
rect 7821 1305 7841 1325
rect 7929 1305 7949 1325
rect 8032 1309 8052 1329
rect 8147 1305 8167 1325
rect 8250 1309 8270 1329
rect 8423 1327 8441 1345
rect 8872 1354 8890 1372
rect 5196 1259 5216 1279
rect 125 1146 143 1164
rect 18568 1484 18588 1504
rect 18671 1488 18691 1508
rect 18786 1484 18806 1504
rect 18889 1488 18909 1508
rect 18997 1488 19017 1508
rect 19100 1484 19120 1504
rect 19927 1492 19947 1512
rect 20030 1488 20050 1508
rect 20138 1488 20158 1508
rect 20241 1492 20261 1512
rect 20356 1488 20376 1508
rect 25805 1641 25823 1659
rect 33829 1758 33849 1778
rect 33932 1754 33952 1774
rect 34040 1754 34060 1774
rect 34143 1758 34163 1778
rect 34258 1754 34278 1774
rect 34361 1758 34381 1778
rect 34548 1765 34566 1783
rect 30612 1703 30630 1721
rect 26246 1591 26264 1609
rect 20459 1492 20479 1512
rect 21436 1509 21454 1527
rect 22932 1497 22952 1517
rect 17168 1436 17186 1454
rect 12095 1321 12115 1341
rect 8421 1228 8439 1246
rect 8870 1255 8888 1273
rect 9041 1271 9061 1291
rect 9144 1275 9164 1295
rect 9259 1271 9279 1291
rect 9362 1275 9382 1295
rect 9470 1275 9490 1295
rect 12198 1317 12218 1337
rect 12306 1317 12326 1337
rect 12409 1321 12429 1341
rect 12524 1317 12544 1337
rect 12627 1321 12647 1341
rect 12800 1339 12818 1357
rect 13236 1367 13254 1385
rect 9573 1271 9593 1291
rect 4489 1159 4507 1177
rect 16459 1334 16479 1354
rect 12798 1240 12816 1258
rect 13234 1268 13252 1286
rect 13405 1284 13425 1304
rect 13508 1288 13528 1308
rect 13623 1284 13643 1304
rect 13726 1288 13746 1308
rect 13834 1288 13854 1308
rect 16562 1330 16582 1350
rect 16670 1330 16690 1350
rect 16773 1334 16793 1354
rect 16888 1330 16908 1350
rect 16991 1334 17011 1354
rect 17164 1352 17182 1370
rect 23035 1501 23055 1521
rect 23150 1497 23170 1517
rect 23253 1501 23273 1521
rect 23361 1501 23381 1521
rect 23464 1497 23484 1517
rect 24291 1505 24311 1525
rect 24394 1501 24414 1521
rect 24502 1501 24522 1521
rect 24605 1505 24625 1525
rect 24720 1501 24740 1521
rect 24823 1505 24843 1525
rect 25800 1522 25818 1540
rect 30182 1653 30200 1671
rect 30610 1604 30628 1622
rect 27309 1509 27329 1529
rect 21434 1410 21452 1428
rect 13937 1284 13957 1304
rect 8866 1171 8884 1189
rect 17502 1341 17520 1359
rect 17162 1253 17180 1271
rect 27412 1513 27432 1533
rect 27527 1509 27547 1529
rect 27630 1513 27650 1533
rect 27738 1513 27758 1533
rect 27841 1509 27861 1529
rect 28668 1517 28688 1537
rect 28771 1513 28791 1533
rect 28879 1513 28899 1533
rect 28982 1517 29002 1537
rect 29097 1513 29117 1533
rect 34546 1666 34564 1684
rect 29200 1517 29220 1537
rect 30177 1534 30195 1552
rect 31673 1522 31693 1542
rect 25798 1423 25816 1441
rect 20725 1308 20745 1328
rect 13230 1184 13248 1202
rect 17500 1242 17518 1260
rect 17671 1258 17691 1278
rect 17774 1262 17794 1282
rect 17889 1258 17909 1278
rect 17992 1262 18012 1282
rect 18100 1262 18120 1282
rect 20828 1304 20848 1324
rect 20936 1304 20956 1324
rect 21039 1308 21059 1328
rect 21154 1304 21174 1324
rect 21257 1308 21277 1328
rect 21430 1326 21448 1344
rect 21866 1354 21884 1372
rect 18203 1258 18223 1278
rect 31776 1526 31796 1546
rect 31891 1522 31911 1542
rect 31994 1526 32014 1546
rect 32102 1526 32122 1546
rect 32205 1522 32225 1542
rect 33032 1530 33052 1550
rect 33135 1526 33155 1546
rect 33243 1526 33263 1546
rect 33346 1530 33366 1550
rect 33461 1526 33481 1546
rect 33564 1530 33584 1550
rect 34541 1547 34559 1565
rect 30175 1435 30193 1453
rect 25089 1321 25109 1341
rect 21428 1227 21446 1245
rect 21864 1255 21882 1273
rect 22035 1271 22055 1291
rect 22138 1275 22158 1295
rect 22253 1271 22273 1291
rect 22356 1275 22376 1295
rect 22464 1275 22484 1295
rect 25192 1317 25212 1337
rect 25300 1317 25320 1337
rect 25403 1321 25423 1341
rect 25518 1317 25538 1337
rect 25621 1321 25641 1341
rect 25794 1339 25812 1357
rect 26243 1366 26261 1384
rect 22567 1271 22587 1291
rect 17496 1158 17514 1176
rect 123 1047 141 1065
rect 1098 1062 1118 1082
rect 1201 1066 1221 1086
rect 1316 1062 1336 1082
rect 1419 1066 1439 1086
rect 1527 1066 1547 1086
rect 1630 1062 1650 1082
rect 4487 1060 4505 1078
rect 5462 1075 5482 1095
rect 118 928 136 946
rect 5565 1079 5585 1099
rect 5680 1075 5700 1095
rect 5783 1079 5803 1099
rect 5891 1079 5911 1099
rect 5994 1075 6014 1095
rect 8864 1072 8882 1090
rect 9839 1087 9859 1107
rect 4054 990 4072 1008
rect 4482 941 4500 959
rect 9942 1091 9962 1111
rect 10057 1087 10077 1107
rect 10160 1091 10180 1111
rect 10268 1091 10288 1111
rect 10371 1087 10391 1107
rect 13228 1085 13246 1103
rect 14203 1100 14223 1120
rect 8418 1003 8436 1021
rect 4052 891 4070 909
rect 116 829 134 847
rect 301 834 321 854
rect 404 838 424 858
rect 519 834 539 854
rect 622 838 642 858
rect 730 838 750 858
rect 833 834 853 854
rect 8859 953 8877 971
rect 14306 1104 14326 1124
rect 14421 1100 14441 1120
rect 14524 1104 14544 1124
rect 14632 1104 14652 1124
rect 14735 1100 14755 1120
rect 34539 1448 34557 1466
rect 29466 1333 29486 1353
rect 25792 1240 25810 1258
rect 26241 1267 26259 1285
rect 26412 1283 26432 1303
rect 26515 1287 26535 1307
rect 26630 1283 26650 1303
rect 26733 1287 26753 1307
rect 26841 1287 26861 1307
rect 29569 1329 29589 1349
rect 29677 1329 29697 1349
rect 29780 1333 29800 1353
rect 29895 1329 29915 1349
rect 29998 1333 30018 1353
rect 30171 1351 30189 1369
rect 30607 1379 30625 1397
rect 26944 1283 26964 1303
rect 21860 1171 21878 1189
rect 33830 1346 33850 1366
rect 30169 1252 30187 1270
rect 30605 1280 30623 1298
rect 30776 1296 30796 1316
rect 30879 1300 30899 1320
rect 30994 1296 31014 1316
rect 31097 1300 31117 1320
rect 31205 1300 31225 1320
rect 33933 1342 33953 1362
rect 34041 1342 34061 1362
rect 34144 1346 34164 1366
rect 34259 1342 34279 1362
rect 34362 1346 34382 1366
rect 34535 1364 34553 1382
rect 31308 1296 31328 1316
rect 26237 1183 26255 1201
rect 34533 1265 34551 1283
rect 30601 1196 30619 1214
rect 12795 1015 12813 1033
rect 8416 904 8434 922
rect 4480 842 4498 860
rect 4665 847 4685 867
rect 4768 851 4788 871
rect 4883 847 4903 867
rect 4986 851 5006 871
rect 5094 851 5114 871
rect 5197 847 5217 867
rect 13223 966 13241 984
rect 17159 1028 17177 1046
rect 17494 1059 17512 1077
rect 18469 1074 18489 1094
rect 18572 1078 18592 1098
rect 18687 1074 18707 1094
rect 18790 1078 18810 1098
rect 18898 1078 18918 1098
rect 19001 1074 19021 1094
rect 21858 1072 21876 1090
rect 22833 1087 22853 1107
rect 12793 916 12811 934
rect 8857 854 8875 872
rect 9042 859 9062 879
rect 9145 863 9165 883
rect 9260 859 9280 879
rect 9363 863 9383 883
rect 9471 863 9491 883
rect 9574 859 9594 879
rect 17157 929 17175 947
rect 17489 940 17507 958
rect 22936 1091 22956 1111
rect 23051 1087 23071 1107
rect 23154 1091 23174 1111
rect 23262 1091 23282 1111
rect 23365 1087 23385 1107
rect 26235 1084 26253 1102
rect 27210 1099 27230 1119
rect 21425 1002 21443 1020
rect 13221 867 13239 885
rect 13406 872 13426 892
rect 13509 876 13529 896
rect 13624 872 13644 892
rect 13727 876 13747 896
rect 13835 876 13855 896
rect 13938 872 13958 892
rect 21853 953 21871 971
rect 27313 1103 27333 1123
rect 27428 1099 27448 1119
rect 27531 1103 27551 1123
rect 27639 1103 27659 1123
rect 27742 1099 27762 1119
rect 30599 1097 30617 1115
rect 31574 1112 31594 1132
rect 25789 1015 25807 1033
rect 21423 903 21441 921
rect 17487 841 17505 859
rect 17672 846 17692 866
rect 17775 850 17795 870
rect 17890 846 17910 866
rect 17993 850 18013 870
rect 18101 850 18121 870
rect 18204 846 18224 866
rect 26230 965 26248 983
rect 31677 1116 31697 1136
rect 31792 1112 31812 1132
rect 31895 1116 31915 1136
rect 32003 1116 32023 1136
rect 32106 1112 32126 1132
rect 30166 1027 30184 1045
rect 25787 916 25805 934
rect 21851 854 21869 872
rect 22036 859 22056 879
rect 22139 863 22159 883
rect 22254 859 22274 879
rect 22357 863 22377 883
rect 22465 863 22485 883
rect 22568 859 22588 879
rect 30594 978 30612 996
rect 34530 1040 34548 1058
rect 30164 928 30182 946
rect 26228 866 26246 884
rect 26413 871 26433 891
rect 26516 875 26536 895
rect 26631 871 26651 891
rect 26734 875 26754 895
rect 26842 875 26862 895
rect 26945 871 26965 891
rect 34528 941 34546 959
rect 30592 879 30610 897
rect 30777 884 30797 904
rect 30880 888 30900 908
rect 30995 884 31015 904
rect 31098 888 31118 908
rect 31206 888 31226 908
rect 31309 884 31329 904
rect 1514 258 1534 278
rect 1617 262 1637 282
rect 1732 258 1752 278
rect 1835 262 1855 282
rect 1943 262 1963 282
rect 2046 258 2066 278
rect 5878 271 5898 291
rect 5981 275 6001 295
rect 6096 271 6116 291
rect 6199 275 6219 295
rect 6307 275 6327 295
rect 6410 271 6430 291
rect 10255 283 10275 303
rect 10358 287 10378 307
rect 10473 283 10493 303
rect 10576 287 10596 307
rect 10684 287 10704 307
rect 10787 283 10807 303
rect 14619 296 14639 316
rect 14722 300 14742 320
rect 14837 296 14857 316
rect 14940 300 14960 320
rect 15048 300 15068 320
rect 15151 296 15171 316
rect 18885 270 18905 290
rect 18988 274 19008 294
rect 19103 270 19123 290
rect 19206 274 19226 294
rect 19314 274 19334 294
rect 19417 270 19437 290
rect 4003 184 4023 204
rect 4106 188 4126 208
rect 4221 184 4241 204
rect 4324 188 4344 208
rect 4432 188 4452 208
rect 4535 184 4555 204
rect 8451 208 8471 228
rect 8554 212 8574 232
rect 8669 208 8689 228
rect 8772 212 8792 232
rect 8880 212 8900 232
rect 8983 208 9003 228
rect 12744 209 12764 229
rect 12847 213 12867 233
rect 12962 209 12982 229
rect 13065 213 13085 233
rect 13173 213 13193 233
rect 13276 209 13296 229
rect 23249 283 23269 303
rect 23352 287 23372 307
rect 23467 283 23487 303
rect 23570 287 23590 307
rect 23678 287 23698 307
rect 23781 283 23801 303
rect 27626 295 27646 315
rect 27729 299 27749 319
rect 27844 295 27864 315
rect 27947 299 27967 319
rect 28055 299 28075 319
rect 28158 295 28178 315
rect 31990 308 32010 328
rect 32093 312 32113 332
rect 32208 308 32228 328
rect 32311 312 32331 332
rect 32419 312 32439 332
rect 32522 308 32542 328
rect 21374 196 21394 216
rect 21477 200 21497 220
rect 21592 196 21612 216
rect 21695 200 21715 220
rect 21803 200 21823 220
rect 21906 196 21926 216
rect 25822 220 25842 240
rect 25925 224 25945 244
rect 26040 220 26060 240
rect 26143 224 26163 244
rect 26251 224 26271 244
rect 26354 220 26374 240
rect 30115 221 30135 241
rect 30218 225 30238 245
rect 30333 221 30353 241
rect 30436 225 30456 245
rect 30544 225 30564 245
rect 30647 221 30667 241
rect 16941 145 16961 165
rect 17044 149 17064 169
rect 17159 145 17179 165
rect 17262 149 17282 169
rect 17370 149 17390 169
rect 17473 145 17493 165
<< pdiffc >>
rect 3486 8685 3506 8705
rect 3582 8685 3602 8705
rect 3692 8685 3712 8705
rect 3788 8685 3808 8705
rect 3910 8685 3930 8705
rect 4006 8685 4026 8705
rect 7850 8698 7870 8718
rect 7946 8698 7966 8718
rect 8056 8698 8076 8718
rect 8152 8698 8172 8718
rect 8274 8698 8294 8718
rect 8370 8698 8390 8718
rect 12227 8710 12247 8730
rect 12323 8710 12343 8730
rect 12433 8710 12453 8730
rect 12529 8710 12549 8730
rect 12651 8710 12671 8730
rect 12747 8710 12767 8730
rect 16591 8723 16611 8743
rect 16687 8723 16707 8743
rect 16797 8723 16817 8743
rect 16893 8723 16913 8743
rect 17015 8723 17035 8743
rect 17111 8723 17131 8743
rect 20857 8697 20877 8717
rect 20953 8697 20973 8717
rect 21063 8697 21083 8717
rect 21159 8697 21179 8717
rect 21281 8697 21301 8717
rect 21377 8697 21397 8717
rect 25221 8710 25241 8730
rect 433 8521 453 8541
rect 529 8521 549 8541
rect 651 8521 671 8541
rect 747 8521 767 8541
rect 857 8521 877 8541
rect 953 8521 973 8541
rect 4797 8534 4817 8554
rect 2689 8457 2709 8477
rect 2785 8457 2805 8477
rect 2895 8457 2915 8477
rect 2991 8457 3011 8477
rect 3113 8457 3133 8477
rect 4893 8534 4913 8554
rect 5015 8534 5035 8554
rect 5111 8534 5131 8554
rect 5221 8534 5241 8554
rect 5317 8534 5337 8554
rect 9174 8546 9194 8566
rect 3209 8457 3229 8477
rect 1231 8337 1251 8357
rect 1327 8337 1347 8357
rect 1449 8337 1469 8357
rect 1545 8337 1565 8357
rect 1655 8337 1675 8357
rect 1751 8337 1771 8357
rect 7053 8470 7073 8490
rect 7149 8470 7169 8490
rect 7259 8470 7279 8490
rect 7355 8470 7375 8490
rect 7477 8470 7497 8490
rect 9270 8546 9290 8566
rect 9392 8546 9412 8566
rect 9488 8546 9508 8566
rect 9598 8546 9618 8566
rect 9694 8546 9714 8566
rect 13538 8559 13558 8579
rect 7573 8470 7593 8490
rect 5595 8350 5615 8370
rect 3487 8273 3507 8293
rect 3583 8273 3603 8293
rect 3693 8273 3713 8293
rect 3789 8273 3809 8293
rect 3911 8273 3931 8293
rect 5691 8350 5711 8370
rect 5813 8350 5833 8370
rect 5909 8350 5929 8370
rect 6019 8350 6039 8370
rect 6115 8350 6135 8370
rect 11430 8482 11450 8502
rect 11526 8482 11546 8502
rect 11636 8482 11656 8502
rect 11732 8482 11752 8502
rect 11854 8482 11874 8502
rect 13634 8559 13654 8579
rect 13756 8559 13776 8579
rect 13852 8559 13872 8579
rect 13962 8559 13982 8579
rect 14058 8559 14078 8579
rect 25317 8710 25337 8730
rect 25427 8710 25447 8730
rect 25523 8710 25543 8730
rect 25645 8710 25665 8730
rect 25741 8710 25761 8730
rect 29598 8722 29618 8742
rect 29694 8722 29714 8742
rect 29804 8722 29824 8742
rect 29900 8722 29920 8742
rect 30022 8722 30042 8742
rect 30118 8722 30138 8742
rect 33962 8735 33982 8755
rect 34058 8735 34078 8755
rect 34168 8735 34188 8755
rect 34264 8735 34284 8755
rect 34386 8735 34406 8755
rect 34482 8735 34502 8755
rect 11950 8482 11970 8502
rect 9972 8362 9992 8382
rect 4007 8273 4027 8293
rect 7851 8286 7871 8306
rect 7947 8286 7967 8306
rect 8057 8286 8077 8306
rect 8153 8286 8173 8306
rect 8275 8286 8295 8306
rect 10068 8362 10088 8382
rect 10190 8362 10210 8382
rect 10286 8362 10306 8382
rect 10396 8362 10416 8382
rect 10492 8362 10512 8382
rect 15794 8495 15814 8515
rect 15890 8495 15910 8515
rect 16000 8495 16020 8515
rect 16096 8495 16116 8515
rect 16218 8495 16238 8515
rect 17804 8533 17824 8553
rect 16314 8495 16334 8515
rect 17900 8533 17920 8553
rect 18022 8533 18042 8553
rect 18118 8533 18138 8553
rect 18228 8533 18248 8553
rect 18324 8533 18344 8553
rect 22168 8546 22188 8566
rect 14336 8375 14356 8395
rect 8371 8286 8391 8306
rect 434 8109 454 8129
rect 530 8109 550 8129
rect 652 8109 672 8129
rect 748 8109 768 8129
rect 858 8109 878 8129
rect 954 8109 974 8129
rect 12228 8298 12248 8318
rect 12324 8298 12344 8318
rect 12434 8298 12454 8318
rect 12530 8298 12550 8318
rect 12652 8298 12672 8318
rect 14432 8375 14452 8395
rect 14554 8375 14574 8395
rect 14650 8375 14670 8395
rect 14760 8375 14780 8395
rect 14856 8375 14876 8395
rect 20060 8469 20080 8489
rect 20156 8469 20176 8489
rect 20266 8469 20286 8489
rect 20362 8469 20382 8489
rect 20484 8469 20504 8489
rect 22264 8546 22284 8566
rect 22386 8546 22406 8566
rect 22482 8546 22502 8566
rect 22592 8546 22612 8566
rect 22688 8546 22708 8566
rect 26545 8558 26565 8578
rect 20580 8469 20600 8489
rect 12748 8298 12768 8318
rect 2590 8047 2610 8067
rect 2686 8047 2706 8067
rect 2796 8047 2816 8067
rect 2892 8047 2912 8067
rect 3014 8047 3034 8067
rect 4798 8122 4818 8142
rect 3110 8047 3130 8067
rect 4894 8122 4914 8142
rect 5016 8122 5036 8142
rect 5112 8122 5132 8142
rect 5222 8122 5242 8142
rect 5318 8122 5338 8142
rect 16592 8311 16612 8331
rect 16688 8311 16708 8331
rect 16798 8311 16818 8331
rect 16894 8311 16914 8331
rect 17016 8311 17036 8331
rect 18602 8349 18622 8369
rect 17112 8311 17132 8331
rect 18698 8349 18718 8369
rect 18820 8349 18840 8369
rect 18916 8349 18936 8369
rect 19026 8349 19046 8369
rect 19122 8349 19142 8369
rect 24424 8482 24444 8502
rect 24520 8482 24540 8502
rect 24630 8482 24650 8502
rect 24726 8482 24746 8502
rect 24848 8482 24868 8502
rect 26641 8558 26661 8578
rect 26763 8558 26783 8578
rect 26859 8558 26879 8578
rect 26969 8558 26989 8578
rect 27065 8558 27085 8578
rect 30909 8571 30929 8591
rect 24944 8482 24964 8502
rect 22966 8362 22986 8382
rect 6954 8060 6974 8080
rect 7050 8060 7070 8080
rect 7160 8060 7180 8080
rect 7256 8060 7276 8080
rect 7378 8060 7398 8080
rect 9175 8134 9195 8154
rect 7474 8060 7494 8080
rect 9271 8134 9291 8154
rect 9393 8134 9413 8154
rect 9489 8134 9509 8154
rect 9599 8134 9619 8154
rect 9695 8134 9715 8154
rect 20858 8285 20878 8305
rect 20954 8285 20974 8305
rect 21064 8285 21084 8305
rect 21160 8285 21180 8305
rect 21282 8285 21302 8305
rect 23062 8362 23082 8382
rect 23184 8362 23204 8382
rect 23280 8362 23300 8382
rect 23390 8362 23410 8382
rect 23486 8362 23506 8382
rect 28801 8494 28821 8514
rect 28897 8494 28917 8514
rect 29007 8494 29027 8514
rect 29103 8494 29123 8514
rect 29225 8494 29245 8514
rect 31005 8571 31025 8591
rect 31127 8571 31147 8591
rect 31223 8571 31243 8591
rect 31333 8571 31353 8591
rect 31429 8571 31449 8591
rect 29321 8494 29341 8514
rect 27343 8374 27363 8394
rect 21378 8285 21398 8305
rect 11331 8072 11351 8092
rect 11427 8072 11447 8092
rect 11537 8072 11557 8092
rect 11633 8072 11653 8092
rect 11755 8072 11775 8092
rect 13539 8147 13559 8167
rect 11851 8072 11871 8092
rect 13635 8147 13655 8167
rect 13757 8147 13777 8167
rect 13853 8147 13873 8167
rect 13963 8147 13983 8167
rect 14059 8147 14079 8167
rect 25222 8298 25242 8318
rect 25318 8298 25338 8318
rect 25428 8298 25448 8318
rect 25524 8298 25544 8318
rect 25646 8298 25666 8318
rect 27439 8374 27459 8394
rect 27561 8374 27581 8394
rect 27657 8374 27677 8394
rect 27767 8374 27787 8394
rect 27863 8374 27883 8394
rect 33165 8507 33185 8527
rect 33261 8507 33281 8527
rect 33371 8507 33391 8527
rect 33467 8507 33487 8527
rect 33589 8507 33609 8527
rect 33685 8507 33705 8527
rect 31707 8387 31727 8407
rect 25742 8298 25762 8318
rect 15695 8085 15715 8105
rect 15791 8085 15811 8105
rect 15901 8085 15921 8105
rect 15997 8085 16017 8105
rect 16119 8085 16139 8105
rect 16215 8085 16235 8105
rect 17805 8121 17825 8141
rect 17901 8121 17921 8141
rect 18023 8121 18043 8141
rect 18119 8121 18139 8141
rect 18229 8121 18249 8141
rect 18325 8121 18345 8141
rect 29599 8310 29619 8330
rect 29695 8310 29715 8330
rect 29805 8310 29825 8330
rect 29901 8310 29921 8330
rect 30023 8310 30043 8330
rect 31803 8387 31823 8407
rect 31925 8387 31945 8407
rect 32021 8387 32041 8407
rect 32131 8387 32151 8407
rect 32227 8387 32247 8407
rect 30119 8310 30139 8330
rect 19961 8059 19981 8079
rect 20057 8059 20077 8079
rect 20167 8059 20187 8079
rect 20263 8059 20283 8079
rect 20385 8059 20405 8079
rect 22169 8134 22189 8154
rect 20481 8059 20501 8079
rect 22265 8134 22285 8154
rect 22387 8134 22407 8154
rect 22483 8134 22503 8154
rect 22593 8134 22613 8154
rect 22689 8134 22709 8154
rect 33963 8323 33983 8343
rect 34059 8323 34079 8343
rect 34169 8323 34189 8343
rect 34265 8323 34285 8343
rect 34387 8323 34407 8343
rect 34483 8323 34503 8343
rect 24325 8072 24345 8092
rect 24421 8072 24441 8092
rect 24531 8072 24551 8092
rect 24627 8072 24647 8092
rect 24749 8072 24769 8092
rect 26546 8146 26566 8166
rect 24845 8072 24865 8092
rect 26642 8146 26662 8166
rect 26764 8146 26784 8166
rect 26860 8146 26880 8166
rect 26970 8146 26990 8166
rect 27066 8146 27086 8166
rect 28702 8084 28722 8104
rect 28798 8084 28818 8104
rect 28908 8084 28928 8104
rect 29004 8084 29024 8104
rect 29126 8084 29146 8104
rect 30910 8159 30930 8179
rect 29222 8084 29242 8104
rect 31006 8159 31026 8179
rect 31128 8159 31148 8179
rect 31224 8159 31244 8179
rect 31334 8159 31354 8179
rect 31430 8159 31450 8179
rect 33066 8097 33086 8117
rect 33162 8097 33182 8117
rect 33272 8097 33292 8117
rect 33368 8097 33388 8117
rect 33490 8097 33510 8117
rect 33586 8097 33606 8117
rect 1313 7729 1333 7749
rect 1409 7729 1429 7749
rect 1531 7729 1551 7749
rect 1627 7729 1647 7749
rect 1737 7729 1757 7749
rect 1833 7729 1853 7749
rect 3469 7667 3489 7687
rect 3565 7667 3585 7687
rect 3675 7667 3695 7687
rect 3771 7667 3791 7687
rect 3893 7667 3913 7687
rect 5677 7742 5697 7762
rect 3989 7667 4009 7687
rect 5773 7742 5793 7762
rect 5895 7742 5915 7762
rect 5991 7742 6011 7762
rect 6101 7742 6121 7762
rect 6197 7742 6217 7762
rect 7833 7680 7853 7700
rect 7929 7680 7949 7700
rect 8039 7680 8059 7700
rect 8135 7680 8155 7700
rect 8257 7680 8277 7700
rect 10054 7754 10074 7774
rect 8353 7680 8373 7700
rect 10150 7754 10170 7774
rect 10272 7754 10292 7774
rect 10368 7754 10388 7774
rect 10478 7754 10498 7774
rect 10574 7754 10594 7774
rect 416 7503 436 7523
rect 512 7503 532 7523
rect 634 7503 654 7523
rect 730 7503 750 7523
rect 840 7503 860 7523
rect 936 7503 956 7523
rect 12210 7692 12230 7712
rect 12306 7692 12326 7712
rect 12416 7692 12436 7712
rect 12512 7692 12532 7712
rect 12634 7692 12654 7712
rect 14418 7767 14438 7787
rect 12730 7692 12750 7712
rect 14514 7767 14534 7787
rect 14636 7767 14656 7787
rect 14732 7767 14752 7787
rect 14842 7767 14862 7787
rect 14938 7767 14958 7787
rect 4780 7516 4800 7536
rect 2672 7439 2692 7459
rect 2768 7439 2788 7459
rect 2878 7439 2898 7459
rect 2974 7439 2994 7459
rect 3096 7439 3116 7459
rect 4876 7516 4896 7536
rect 4998 7516 5018 7536
rect 5094 7516 5114 7536
rect 5204 7516 5224 7536
rect 5300 7516 5320 7536
rect 16574 7705 16594 7725
rect 16670 7705 16690 7725
rect 16780 7705 16800 7725
rect 16876 7705 16896 7725
rect 16998 7705 17018 7725
rect 17094 7705 17114 7725
rect 18684 7741 18704 7761
rect 18780 7741 18800 7761
rect 18902 7741 18922 7761
rect 18998 7741 19018 7761
rect 19108 7741 19128 7761
rect 19204 7741 19224 7761
rect 9157 7528 9177 7548
rect 3192 7439 3212 7459
rect 1214 7319 1234 7339
rect 1310 7319 1330 7339
rect 1432 7319 1452 7339
rect 1528 7319 1548 7339
rect 1638 7319 1658 7339
rect 1734 7319 1754 7339
rect 7036 7452 7056 7472
rect 7132 7452 7152 7472
rect 7242 7452 7262 7472
rect 7338 7452 7358 7472
rect 7460 7452 7480 7472
rect 9253 7528 9273 7548
rect 9375 7528 9395 7548
rect 9471 7528 9491 7548
rect 9581 7528 9601 7548
rect 9677 7528 9697 7548
rect 20840 7679 20860 7699
rect 20936 7679 20956 7699
rect 21046 7679 21066 7699
rect 21142 7679 21162 7699
rect 21264 7679 21284 7699
rect 23048 7754 23068 7774
rect 21360 7679 21380 7699
rect 23144 7754 23164 7774
rect 23266 7754 23286 7774
rect 23362 7754 23382 7774
rect 23472 7754 23492 7774
rect 23568 7754 23588 7774
rect 13521 7541 13541 7561
rect 7556 7452 7576 7472
rect 5578 7332 5598 7352
rect 3470 7255 3490 7275
rect 3566 7255 3586 7275
rect 3676 7255 3696 7275
rect 3772 7255 3792 7275
rect 3894 7255 3914 7275
rect 5674 7332 5694 7352
rect 5796 7332 5816 7352
rect 5892 7332 5912 7352
rect 6002 7332 6022 7352
rect 6098 7332 6118 7352
rect 11413 7464 11433 7484
rect 11509 7464 11529 7484
rect 11619 7464 11639 7484
rect 11715 7464 11735 7484
rect 11837 7464 11857 7484
rect 13617 7541 13637 7561
rect 13739 7541 13759 7561
rect 13835 7541 13855 7561
rect 13945 7541 13965 7561
rect 14041 7541 14061 7561
rect 25204 7692 25224 7712
rect 25300 7692 25320 7712
rect 25410 7692 25430 7712
rect 25506 7692 25526 7712
rect 25628 7692 25648 7712
rect 27425 7766 27445 7786
rect 25724 7692 25744 7712
rect 27521 7766 27541 7786
rect 27643 7766 27663 7786
rect 27739 7766 27759 7786
rect 27849 7766 27869 7786
rect 27945 7766 27965 7786
rect 11933 7464 11953 7484
rect 9955 7344 9975 7364
rect 3990 7255 4010 7275
rect 7834 7268 7854 7288
rect 7930 7268 7950 7288
rect 8040 7268 8060 7288
rect 8136 7268 8156 7288
rect 8258 7268 8278 7288
rect 10051 7344 10071 7364
rect 10173 7344 10193 7364
rect 10269 7344 10289 7364
rect 10379 7344 10399 7364
rect 10475 7344 10495 7364
rect 15777 7477 15797 7497
rect 15873 7477 15893 7497
rect 15983 7477 16003 7497
rect 16079 7477 16099 7497
rect 16201 7477 16221 7497
rect 17787 7515 17807 7535
rect 16297 7477 16317 7497
rect 17883 7515 17903 7535
rect 18005 7515 18025 7535
rect 18101 7515 18121 7535
rect 18211 7515 18231 7535
rect 18307 7515 18327 7535
rect 29581 7704 29601 7724
rect 29677 7704 29697 7724
rect 29787 7704 29807 7724
rect 29883 7704 29903 7724
rect 30005 7704 30025 7724
rect 31789 7779 31809 7799
rect 30101 7704 30121 7724
rect 31885 7779 31905 7799
rect 32007 7779 32027 7799
rect 32103 7779 32123 7799
rect 32213 7779 32233 7799
rect 32309 7779 32329 7799
rect 22151 7528 22171 7548
rect 14319 7357 14339 7377
rect 8354 7268 8374 7288
rect 417 7091 437 7111
rect 513 7091 533 7111
rect 635 7091 655 7111
rect 731 7091 751 7111
rect 841 7091 861 7111
rect 937 7091 957 7111
rect 12211 7280 12231 7300
rect 12307 7280 12327 7300
rect 12417 7280 12437 7300
rect 12513 7280 12533 7300
rect 12635 7280 12655 7300
rect 14415 7357 14435 7377
rect 14537 7357 14557 7377
rect 14633 7357 14653 7377
rect 14743 7357 14763 7377
rect 14839 7357 14859 7377
rect 20043 7451 20063 7471
rect 20139 7451 20159 7471
rect 20249 7451 20269 7471
rect 20345 7451 20365 7471
rect 20467 7451 20487 7471
rect 22247 7528 22267 7548
rect 22369 7528 22389 7548
rect 22465 7528 22485 7548
rect 22575 7528 22595 7548
rect 22671 7528 22691 7548
rect 33945 7717 33965 7737
rect 34041 7717 34061 7737
rect 34151 7717 34171 7737
rect 34247 7717 34267 7737
rect 34369 7717 34389 7737
rect 34465 7717 34485 7737
rect 26528 7540 26548 7560
rect 20563 7451 20583 7471
rect 12731 7280 12751 7300
rect 2507 7031 2527 7051
rect 2603 7031 2623 7051
rect 2713 7031 2733 7051
rect 2809 7031 2829 7051
rect 2931 7031 2951 7051
rect 4781 7104 4801 7124
rect 3027 7031 3047 7051
rect 4877 7104 4897 7124
rect 4999 7104 5019 7124
rect 5095 7104 5115 7124
rect 5205 7104 5225 7124
rect 5301 7104 5321 7124
rect 16575 7293 16595 7313
rect 16671 7293 16691 7313
rect 16781 7293 16801 7313
rect 16877 7293 16897 7313
rect 16999 7293 17019 7313
rect 18585 7331 18605 7351
rect 17095 7293 17115 7313
rect 18681 7331 18701 7351
rect 18803 7331 18823 7351
rect 18899 7331 18919 7351
rect 19009 7331 19029 7351
rect 19105 7331 19125 7351
rect 24407 7464 24427 7484
rect 24503 7464 24523 7484
rect 24613 7464 24633 7484
rect 24709 7464 24729 7484
rect 24831 7464 24851 7484
rect 26624 7540 26644 7560
rect 26746 7540 26766 7560
rect 26842 7540 26862 7560
rect 26952 7540 26972 7560
rect 27048 7540 27068 7560
rect 30892 7553 30912 7573
rect 24927 7464 24947 7484
rect 22949 7344 22969 7364
rect 6871 7044 6891 7064
rect 6967 7044 6987 7064
rect 7077 7044 7097 7064
rect 7173 7044 7193 7064
rect 7295 7044 7315 7064
rect 9158 7116 9178 7136
rect 7391 7044 7411 7064
rect 9254 7116 9274 7136
rect 9376 7116 9396 7136
rect 9472 7116 9492 7136
rect 9582 7116 9602 7136
rect 9678 7116 9698 7136
rect 20841 7267 20861 7287
rect 20937 7267 20957 7287
rect 21047 7267 21067 7287
rect 21143 7267 21163 7287
rect 21265 7267 21285 7287
rect 23045 7344 23065 7364
rect 23167 7344 23187 7364
rect 23263 7344 23283 7364
rect 23373 7344 23393 7364
rect 23469 7344 23489 7364
rect 28784 7476 28804 7496
rect 28880 7476 28900 7496
rect 28990 7476 29010 7496
rect 29086 7476 29106 7496
rect 29208 7476 29228 7496
rect 30988 7553 31008 7573
rect 31110 7553 31130 7573
rect 31206 7553 31226 7573
rect 31316 7553 31336 7573
rect 31412 7553 31432 7573
rect 29304 7476 29324 7496
rect 27326 7356 27346 7376
rect 21361 7267 21381 7287
rect 11248 7056 11268 7076
rect 11344 7056 11364 7076
rect 11454 7056 11474 7076
rect 11550 7056 11570 7076
rect 11672 7056 11692 7076
rect 13522 7129 13542 7149
rect 11768 7056 11788 7076
rect 13618 7129 13638 7149
rect 13740 7129 13760 7149
rect 13836 7129 13856 7149
rect 13946 7129 13966 7149
rect 14042 7129 14062 7149
rect 25205 7280 25225 7300
rect 25301 7280 25321 7300
rect 25411 7280 25431 7300
rect 25507 7280 25527 7300
rect 25629 7280 25649 7300
rect 27422 7356 27442 7376
rect 27544 7356 27564 7376
rect 27640 7356 27660 7376
rect 27750 7356 27770 7376
rect 27846 7356 27866 7376
rect 33148 7489 33168 7509
rect 33244 7489 33264 7509
rect 33354 7489 33374 7509
rect 33450 7489 33470 7509
rect 33572 7489 33592 7509
rect 33668 7489 33688 7509
rect 31690 7369 31710 7389
rect 25725 7280 25745 7300
rect 15612 7069 15632 7089
rect 15708 7069 15728 7089
rect 15818 7069 15838 7089
rect 15914 7069 15934 7089
rect 16036 7069 16056 7089
rect 16132 7069 16152 7089
rect 17788 7103 17808 7123
rect 17884 7103 17904 7123
rect 18006 7103 18026 7123
rect 18102 7103 18122 7123
rect 18212 7103 18232 7123
rect 18308 7103 18328 7123
rect 29582 7292 29602 7312
rect 29678 7292 29698 7312
rect 29788 7292 29808 7312
rect 29884 7292 29904 7312
rect 30006 7292 30026 7312
rect 31786 7369 31806 7389
rect 31908 7369 31928 7389
rect 32004 7369 32024 7389
rect 32114 7369 32134 7389
rect 32210 7369 32230 7389
rect 30102 7292 30122 7312
rect 19878 7043 19898 7063
rect 19974 7043 19994 7063
rect 20084 7043 20104 7063
rect 20180 7043 20200 7063
rect 20302 7043 20322 7063
rect 22152 7116 22172 7136
rect 20398 7043 20418 7063
rect 22248 7116 22268 7136
rect 22370 7116 22390 7136
rect 22466 7116 22486 7136
rect 22576 7116 22596 7136
rect 22672 7116 22692 7136
rect 33946 7305 33966 7325
rect 34042 7305 34062 7325
rect 34152 7305 34172 7325
rect 34248 7305 34268 7325
rect 34370 7305 34390 7325
rect 34466 7305 34486 7325
rect 24242 7056 24262 7076
rect 24338 7056 24358 7076
rect 24448 7056 24468 7076
rect 24544 7056 24564 7076
rect 24666 7056 24686 7076
rect 26529 7128 26549 7148
rect 24762 7056 24782 7076
rect 26625 7128 26645 7148
rect 26747 7128 26767 7148
rect 26843 7128 26863 7148
rect 26953 7128 26973 7148
rect 27049 7128 27069 7148
rect 28619 7068 28639 7088
rect 28715 7068 28735 7088
rect 28825 7068 28845 7088
rect 28921 7068 28941 7088
rect 29043 7068 29063 7088
rect 30893 7141 30913 7161
rect 29139 7068 29159 7088
rect 30989 7141 31009 7161
rect 31111 7141 31131 7161
rect 31207 7141 31227 7161
rect 31317 7141 31337 7161
rect 31413 7141 31433 7161
rect 32983 7081 33003 7101
rect 33079 7081 33099 7101
rect 33189 7081 33209 7101
rect 33285 7081 33305 7101
rect 33407 7081 33427 7101
rect 33503 7081 33523 7101
rect 1359 6709 1379 6729
rect 1455 6709 1475 6729
rect 1577 6709 1597 6729
rect 1673 6709 1693 6729
rect 1783 6709 1803 6729
rect 1879 6709 1899 6729
rect 3449 6649 3469 6669
rect 3545 6649 3565 6669
rect 3655 6649 3675 6669
rect 3751 6649 3771 6669
rect 3873 6649 3893 6669
rect 5723 6722 5743 6742
rect 3969 6649 3989 6669
rect 5819 6722 5839 6742
rect 5941 6722 5961 6742
rect 6037 6722 6057 6742
rect 6147 6722 6167 6742
rect 6243 6722 6263 6742
rect 7813 6662 7833 6682
rect 7909 6662 7929 6682
rect 8019 6662 8039 6682
rect 8115 6662 8135 6682
rect 8237 6662 8257 6682
rect 10100 6734 10120 6754
rect 8333 6662 8353 6682
rect 10196 6734 10216 6754
rect 10318 6734 10338 6754
rect 10414 6734 10434 6754
rect 10524 6734 10544 6754
rect 10620 6734 10640 6754
rect 396 6485 416 6505
rect 492 6485 512 6505
rect 614 6485 634 6505
rect 710 6485 730 6505
rect 820 6485 840 6505
rect 916 6485 936 6505
rect 12190 6674 12210 6694
rect 12286 6674 12306 6694
rect 12396 6674 12416 6694
rect 12492 6674 12512 6694
rect 12614 6674 12634 6694
rect 14464 6747 14484 6767
rect 12710 6674 12730 6694
rect 14560 6747 14580 6767
rect 14682 6747 14702 6767
rect 14778 6747 14798 6767
rect 14888 6747 14908 6767
rect 14984 6747 15004 6767
rect 4760 6498 4780 6518
rect 2652 6421 2672 6441
rect 2748 6421 2768 6441
rect 2858 6421 2878 6441
rect 2954 6421 2974 6441
rect 3076 6421 3096 6441
rect 4856 6498 4876 6518
rect 4978 6498 4998 6518
rect 5074 6498 5094 6518
rect 5184 6498 5204 6518
rect 5280 6498 5300 6518
rect 16554 6687 16574 6707
rect 16650 6687 16670 6707
rect 16760 6687 16780 6707
rect 16856 6687 16876 6707
rect 16978 6687 16998 6707
rect 17074 6687 17094 6707
rect 18730 6721 18750 6741
rect 18826 6721 18846 6741
rect 18948 6721 18968 6741
rect 19044 6721 19064 6741
rect 19154 6721 19174 6741
rect 19250 6721 19270 6741
rect 9137 6510 9157 6530
rect 3172 6421 3192 6441
rect 1194 6301 1214 6321
rect 1290 6301 1310 6321
rect 1412 6301 1432 6321
rect 1508 6301 1528 6321
rect 1618 6301 1638 6321
rect 1714 6301 1734 6321
rect 7016 6434 7036 6454
rect 7112 6434 7132 6454
rect 7222 6434 7242 6454
rect 7318 6434 7338 6454
rect 7440 6434 7460 6454
rect 9233 6510 9253 6530
rect 9355 6510 9375 6530
rect 9451 6510 9471 6530
rect 9561 6510 9581 6530
rect 9657 6510 9677 6530
rect 20820 6661 20840 6681
rect 20916 6661 20936 6681
rect 21026 6661 21046 6681
rect 21122 6661 21142 6681
rect 21244 6661 21264 6681
rect 23094 6734 23114 6754
rect 21340 6661 21360 6681
rect 23190 6734 23210 6754
rect 23312 6734 23332 6754
rect 23408 6734 23428 6754
rect 23518 6734 23538 6754
rect 23614 6734 23634 6754
rect 13501 6523 13521 6543
rect 7536 6434 7556 6454
rect 5558 6314 5578 6334
rect 3450 6237 3470 6257
rect 3546 6237 3566 6257
rect 3656 6237 3676 6257
rect 3752 6237 3772 6257
rect 3874 6237 3894 6257
rect 5654 6314 5674 6334
rect 5776 6314 5796 6334
rect 5872 6314 5892 6334
rect 5982 6314 6002 6334
rect 6078 6314 6098 6334
rect 11393 6446 11413 6466
rect 11489 6446 11509 6466
rect 11599 6446 11619 6466
rect 11695 6446 11715 6466
rect 11817 6446 11837 6466
rect 13597 6523 13617 6543
rect 13719 6523 13739 6543
rect 13815 6523 13835 6543
rect 13925 6523 13945 6543
rect 14021 6523 14041 6543
rect 25184 6674 25204 6694
rect 25280 6674 25300 6694
rect 25390 6674 25410 6694
rect 25486 6674 25506 6694
rect 25608 6674 25628 6694
rect 27471 6746 27491 6766
rect 25704 6674 25724 6694
rect 27567 6746 27587 6766
rect 27689 6746 27709 6766
rect 27785 6746 27805 6766
rect 27895 6746 27915 6766
rect 27991 6746 28011 6766
rect 11913 6446 11933 6466
rect 9935 6326 9955 6346
rect 3970 6237 3990 6257
rect 7814 6250 7834 6270
rect 7910 6250 7930 6270
rect 8020 6250 8040 6270
rect 8116 6250 8136 6270
rect 8238 6250 8258 6270
rect 10031 6326 10051 6346
rect 10153 6326 10173 6346
rect 10249 6326 10269 6346
rect 10359 6326 10379 6346
rect 10455 6326 10475 6346
rect 15757 6459 15777 6479
rect 15853 6459 15873 6479
rect 15963 6459 15983 6479
rect 16059 6459 16079 6479
rect 16181 6459 16201 6479
rect 17767 6497 17787 6517
rect 16277 6459 16297 6479
rect 17863 6497 17883 6517
rect 17985 6497 18005 6517
rect 18081 6497 18101 6517
rect 18191 6497 18211 6517
rect 18287 6497 18307 6517
rect 29561 6686 29581 6706
rect 29657 6686 29677 6706
rect 29767 6686 29787 6706
rect 29863 6686 29883 6706
rect 29985 6686 30005 6706
rect 31835 6759 31855 6779
rect 30081 6686 30101 6706
rect 31931 6759 31951 6779
rect 32053 6759 32073 6779
rect 32149 6759 32169 6779
rect 32259 6759 32279 6779
rect 32355 6759 32375 6779
rect 22131 6510 22151 6530
rect 14299 6339 14319 6359
rect 8334 6250 8354 6270
rect 397 6073 417 6093
rect 493 6073 513 6093
rect 615 6073 635 6093
rect 711 6073 731 6093
rect 821 6073 841 6093
rect 917 6073 937 6093
rect 12191 6262 12211 6282
rect 12287 6262 12307 6282
rect 12397 6262 12417 6282
rect 12493 6262 12513 6282
rect 12615 6262 12635 6282
rect 14395 6339 14415 6359
rect 14517 6339 14537 6359
rect 14613 6339 14633 6359
rect 14723 6339 14743 6359
rect 14819 6339 14839 6359
rect 20023 6433 20043 6453
rect 20119 6433 20139 6453
rect 20229 6433 20249 6453
rect 20325 6433 20345 6453
rect 20447 6433 20467 6453
rect 22227 6510 22247 6530
rect 22349 6510 22369 6530
rect 22445 6510 22465 6530
rect 22555 6510 22575 6530
rect 22651 6510 22671 6530
rect 33925 6699 33945 6719
rect 34021 6699 34041 6719
rect 34131 6699 34151 6719
rect 34227 6699 34247 6719
rect 34349 6699 34369 6719
rect 34445 6699 34465 6719
rect 26508 6522 26528 6542
rect 20543 6433 20563 6453
rect 12711 6262 12731 6282
rect 2553 6011 2573 6031
rect 2649 6011 2669 6031
rect 2759 6011 2779 6031
rect 2855 6011 2875 6031
rect 2977 6011 2997 6031
rect 4761 6086 4781 6106
rect 3073 6011 3093 6031
rect 4857 6086 4877 6106
rect 4979 6086 4999 6106
rect 5075 6086 5095 6106
rect 5185 6086 5205 6106
rect 5281 6086 5301 6106
rect 16555 6275 16575 6295
rect 16651 6275 16671 6295
rect 16761 6275 16781 6295
rect 16857 6275 16877 6295
rect 16979 6275 16999 6295
rect 18565 6313 18585 6333
rect 17075 6275 17095 6295
rect 18661 6313 18681 6333
rect 18783 6313 18803 6333
rect 18879 6313 18899 6333
rect 18989 6313 19009 6333
rect 19085 6313 19105 6333
rect 24387 6446 24407 6466
rect 24483 6446 24503 6466
rect 24593 6446 24613 6466
rect 24689 6446 24709 6466
rect 24811 6446 24831 6466
rect 26604 6522 26624 6542
rect 26726 6522 26746 6542
rect 26822 6522 26842 6542
rect 26932 6522 26952 6542
rect 27028 6522 27048 6542
rect 30872 6535 30892 6555
rect 24907 6446 24927 6466
rect 22929 6326 22949 6346
rect 6917 6024 6937 6044
rect 7013 6024 7033 6044
rect 7123 6024 7143 6044
rect 7219 6024 7239 6044
rect 7341 6024 7361 6044
rect 9138 6098 9158 6118
rect 7437 6024 7457 6044
rect 9234 6098 9254 6118
rect 9356 6098 9376 6118
rect 9452 6098 9472 6118
rect 9562 6098 9582 6118
rect 9658 6098 9678 6118
rect 20821 6249 20841 6269
rect 20917 6249 20937 6269
rect 21027 6249 21047 6269
rect 21123 6249 21143 6269
rect 21245 6249 21265 6269
rect 23025 6326 23045 6346
rect 23147 6326 23167 6346
rect 23243 6326 23263 6346
rect 23353 6326 23373 6346
rect 23449 6326 23469 6346
rect 28764 6458 28784 6478
rect 28860 6458 28880 6478
rect 28970 6458 28990 6478
rect 29066 6458 29086 6478
rect 29188 6458 29208 6478
rect 30968 6535 30988 6555
rect 31090 6535 31110 6555
rect 31186 6535 31206 6555
rect 31296 6535 31316 6555
rect 31392 6535 31412 6555
rect 29284 6458 29304 6478
rect 27306 6338 27326 6358
rect 21341 6249 21361 6269
rect 11294 6036 11314 6056
rect 11390 6036 11410 6056
rect 11500 6036 11520 6056
rect 11596 6036 11616 6056
rect 11718 6036 11738 6056
rect 13502 6111 13522 6131
rect 11814 6036 11834 6056
rect 13598 6111 13618 6131
rect 13720 6111 13740 6131
rect 13816 6111 13836 6131
rect 13926 6111 13946 6131
rect 14022 6111 14042 6131
rect 25185 6262 25205 6282
rect 25281 6262 25301 6282
rect 25391 6262 25411 6282
rect 25487 6262 25507 6282
rect 25609 6262 25629 6282
rect 27402 6338 27422 6358
rect 27524 6338 27544 6358
rect 27620 6338 27640 6358
rect 27730 6338 27750 6358
rect 27826 6338 27846 6358
rect 33128 6471 33148 6491
rect 33224 6471 33244 6491
rect 33334 6471 33354 6491
rect 33430 6471 33450 6491
rect 33552 6471 33572 6491
rect 33648 6471 33668 6491
rect 31670 6351 31690 6371
rect 25705 6262 25725 6282
rect 15658 6049 15678 6069
rect 15754 6049 15774 6069
rect 15864 6049 15884 6069
rect 15960 6049 15980 6069
rect 16082 6049 16102 6069
rect 16178 6049 16198 6069
rect 17768 6085 17788 6105
rect 17864 6085 17884 6105
rect 17986 6085 18006 6105
rect 18082 6085 18102 6105
rect 18192 6085 18212 6105
rect 18288 6085 18308 6105
rect 29562 6274 29582 6294
rect 29658 6274 29678 6294
rect 29768 6274 29788 6294
rect 29864 6274 29884 6294
rect 29986 6274 30006 6294
rect 31766 6351 31786 6371
rect 31888 6351 31908 6371
rect 31984 6351 32004 6371
rect 32094 6351 32114 6371
rect 32190 6351 32210 6371
rect 30082 6274 30102 6294
rect 19924 6023 19944 6043
rect 20020 6023 20040 6043
rect 20130 6023 20150 6043
rect 20226 6023 20246 6043
rect 20348 6023 20368 6043
rect 22132 6098 22152 6118
rect 20444 6023 20464 6043
rect 22228 6098 22248 6118
rect 22350 6098 22370 6118
rect 22446 6098 22466 6118
rect 22556 6098 22576 6118
rect 22652 6098 22672 6118
rect 33926 6287 33946 6307
rect 34022 6287 34042 6307
rect 34132 6287 34152 6307
rect 34228 6287 34248 6307
rect 34350 6287 34370 6307
rect 34446 6287 34466 6307
rect 24288 6036 24308 6056
rect 24384 6036 24404 6056
rect 24494 6036 24514 6056
rect 24590 6036 24610 6056
rect 24712 6036 24732 6056
rect 26509 6110 26529 6130
rect 24808 6036 24828 6056
rect 26605 6110 26625 6130
rect 26727 6110 26747 6130
rect 26823 6110 26843 6130
rect 26933 6110 26953 6130
rect 27029 6110 27049 6130
rect 28665 6048 28685 6068
rect 28761 6048 28781 6068
rect 28871 6048 28891 6068
rect 28967 6048 28987 6068
rect 29089 6048 29109 6068
rect 30873 6123 30893 6143
rect 29185 6048 29205 6068
rect 30969 6123 30989 6143
rect 31091 6123 31111 6143
rect 31187 6123 31207 6143
rect 31297 6123 31317 6143
rect 31393 6123 31413 6143
rect 33029 6061 33049 6081
rect 33125 6061 33145 6081
rect 33235 6061 33255 6081
rect 33331 6061 33351 6081
rect 33453 6061 33473 6081
rect 33549 6061 33569 6081
rect 1276 5693 1296 5713
rect 1372 5693 1392 5713
rect 1494 5693 1514 5713
rect 1590 5693 1610 5713
rect 1700 5693 1720 5713
rect 1796 5693 1816 5713
rect 3432 5631 3452 5651
rect 3528 5631 3548 5651
rect 3638 5631 3658 5651
rect 3734 5631 3754 5651
rect 3856 5631 3876 5651
rect 5640 5706 5660 5726
rect 3952 5631 3972 5651
rect 5736 5706 5756 5726
rect 5858 5706 5878 5726
rect 5954 5706 5974 5726
rect 6064 5706 6084 5726
rect 6160 5706 6180 5726
rect 7796 5644 7816 5664
rect 7892 5644 7912 5664
rect 8002 5644 8022 5664
rect 8098 5644 8118 5664
rect 8220 5644 8240 5664
rect 10017 5718 10037 5738
rect 8316 5644 8336 5664
rect 10113 5718 10133 5738
rect 10235 5718 10255 5738
rect 10331 5718 10351 5738
rect 10441 5718 10461 5738
rect 10537 5718 10557 5738
rect 379 5467 399 5487
rect 475 5467 495 5487
rect 597 5467 617 5487
rect 693 5467 713 5487
rect 803 5467 823 5487
rect 899 5467 919 5487
rect 12173 5656 12193 5676
rect 12269 5656 12289 5676
rect 12379 5656 12399 5676
rect 12475 5656 12495 5676
rect 12597 5656 12617 5676
rect 14381 5731 14401 5751
rect 12693 5656 12713 5676
rect 14477 5731 14497 5751
rect 14599 5731 14619 5751
rect 14695 5731 14715 5751
rect 14805 5731 14825 5751
rect 14901 5731 14921 5751
rect 4743 5480 4763 5500
rect 2635 5403 2655 5423
rect 2731 5403 2751 5423
rect 2841 5403 2861 5423
rect 2937 5403 2957 5423
rect 3059 5403 3079 5423
rect 4839 5480 4859 5500
rect 4961 5480 4981 5500
rect 5057 5480 5077 5500
rect 5167 5480 5187 5500
rect 5263 5480 5283 5500
rect 16537 5669 16557 5689
rect 16633 5669 16653 5689
rect 16743 5669 16763 5689
rect 16839 5669 16859 5689
rect 16961 5669 16981 5689
rect 17057 5669 17077 5689
rect 18647 5705 18667 5725
rect 18743 5705 18763 5725
rect 18865 5705 18885 5725
rect 18961 5705 18981 5725
rect 19071 5705 19091 5725
rect 19167 5705 19187 5725
rect 9120 5492 9140 5512
rect 3155 5403 3175 5423
rect 1177 5283 1197 5303
rect 1273 5283 1293 5303
rect 1395 5283 1415 5303
rect 1491 5283 1511 5303
rect 1601 5283 1621 5303
rect 1697 5283 1717 5303
rect 6999 5416 7019 5436
rect 7095 5416 7115 5436
rect 7205 5416 7225 5436
rect 7301 5416 7321 5436
rect 7423 5416 7443 5436
rect 9216 5492 9236 5512
rect 9338 5492 9358 5512
rect 9434 5492 9454 5512
rect 9544 5492 9564 5512
rect 9640 5492 9660 5512
rect 20803 5643 20823 5663
rect 20899 5643 20919 5663
rect 21009 5643 21029 5663
rect 21105 5643 21125 5663
rect 21227 5643 21247 5663
rect 23011 5718 23031 5738
rect 21323 5643 21343 5663
rect 23107 5718 23127 5738
rect 23229 5718 23249 5738
rect 23325 5718 23345 5738
rect 23435 5718 23455 5738
rect 23531 5718 23551 5738
rect 13484 5505 13504 5525
rect 7519 5416 7539 5436
rect 5541 5296 5561 5316
rect 3433 5219 3453 5239
rect 3529 5219 3549 5239
rect 3639 5219 3659 5239
rect 3735 5219 3755 5239
rect 3857 5219 3877 5239
rect 5637 5296 5657 5316
rect 5759 5296 5779 5316
rect 5855 5296 5875 5316
rect 5965 5296 5985 5316
rect 6061 5296 6081 5316
rect 11376 5428 11396 5448
rect 11472 5428 11492 5448
rect 11582 5428 11602 5448
rect 11678 5428 11698 5448
rect 11800 5428 11820 5448
rect 13580 5505 13600 5525
rect 13702 5505 13722 5525
rect 13798 5505 13818 5525
rect 13908 5505 13928 5525
rect 14004 5505 14024 5525
rect 25167 5656 25187 5676
rect 25263 5656 25283 5676
rect 25373 5656 25393 5676
rect 25469 5656 25489 5676
rect 25591 5656 25611 5676
rect 27388 5730 27408 5750
rect 25687 5656 25707 5676
rect 27484 5730 27504 5750
rect 27606 5730 27626 5750
rect 27702 5730 27722 5750
rect 27812 5730 27832 5750
rect 27908 5730 27928 5750
rect 11896 5428 11916 5448
rect 9918 5308 9938 5328
rect 3953 5219 3973 5239
rect 7797 5232 7817 5252
rect 7893 5232 7913 5252
rect 8003 5232 8023 5252
rect 8099 5232 8119 5252
rect 8221 5232 8241 5252
rect 10014 5308 10034 5328
rect 10136 5308 10156 5328
rect 10232 5308 10252 5328
rect 10342 5308 10362 5328
rect 10438 5308 10458 5328
rect 15740 5441 15760 5461
rect 15836 5441 15856 5461
rect 15946 5441 15966 5461
rect 16042 5441 16062 5461
rect 16164 5441 16184 5461
rect 17750 5479 17770 5499
rect 16260 5441 16280 5461
rect 17846 5479 17866 5499
rect 17968 5479 17988 5499
rect 18064 5479 18084 5499
rect 18174 5479 18194 5499
rect 18270 5479 18290 5499
rect 29544 5668 29564 5688
rect 29640 5668 29660 5688
rect 29750 5668 29770 5688
rect 29846 5668 29866 5688
rect 29968 5668 29988 5688
rect 31752 5743 31772 5763
rect 30064 5668 30084 5688
rect 31848 5743 31868 5763
rect 31970 5743 31990 5763
rect 32066 5743 32086 5763
rect 32176 5743 32196 5763
rect 32272 5743 32292 5763
rect 22114 5492 22134 5512
rect 14282 5321 14302 5341
rect 8317 5232 8337 5252
rect 380 5055 400 5075
rect 476 5055 496 5075
rect 598 5055 618 5075
rect 694 5055 714 5075
rect 804 5055 824 5075
rect 900 5055 920 5075
rect 12174 5244 12194 5264
rect 12270 5244 12290 5264
rect 12380 5244 12400 5264
rect 12476 5244 12496 5264
rect 12598 5244 12618 5264
rect 14378 5321 14398 5341
rect 14500 5321 14520 5341
rect 14596 5321 14616 5341
rect 14706 5321 14726 5341
rect 14802 5321 14822 5341
rect 20006 5415 20026 5435
rect 20102 5415 20122 5435
rect 20212 5415 20232 5435
rect 20308 5415 20328 5435
rect 20430 5415 20450 5435
rect 22210 5492 22230 5512
rect 22332 5492 22352 5512
rect 22428 5492 22448 5512
rect 22538 5492 22558 5512
rect 22634 5492 22654 5512
rect 33908 5681 33928 5701
rect 34004 5681 34024 5701
rect 34114 5681 34134 5701
rect 34210 5681 34230 5701
rect 34332 5681 34352 5701
rect 34428 5681 34448 5701
rect 26491 5504 26511 5524
rect 20526 5415 20546 5435
rect 12694 5244 12714 5264
rect 2331 4997 2351 5017
rect 2427 4997 2447 5017
rect 2537 4997 2557 5017
rect 2633 4997 2653 5017
rect 2755 4997 2775 5017
rect 4744 5068 4764 5088
rect 2851 4997 2871 5017
rect 4840 5068 4860 5088
rect 4962 5068 4982 5088
rect 5058 5068 5078 5088
rect 5168 5068 5188 5088
rect 5264 5068 5284 5088
rect 16538 5257 16558 5277
rect 16634 5257 16654 5277
rect 16744 5257 16764 5277
rect 16840 5257 16860 5277
rect 16962 5257 16982 5277
rect 18548 5295 18568 5315
rect 17058 5257 17078 5277
rect 18644 5295 18664 5315
rect 18766 5295 18786 5315
rect 18862 5295 18882 5315
rect 18972 5295 18992 5315
rect 19068 5295 19088 5315
rect 24370 5428 24390 5448
rect 24466 5428 24486 5448
rect 24576 5428 24596 5448
rect 24672 5428 24692 5448
rect 24794 5428 24814 5448
rect 26587 5504 26607 5524
rect 26709 5504 26729 5524
rect 26805 5504 26825 5524
rect 26915 5504 26935 5524
rect 27011 5504 27031 5524
rect 30855 5517 30875 5537
rect 24890 5428 24910 5448
rect 22912 5308 22932 5328
rect 6695 5010 6715 5030
rect 6791 5010 6811 5030
rect 6901 5010 6921 5030
rect 6997 5010 7017 5030
rect 7119 5010 7139 5030
rect 9121 5080 9141 5100
rect 7215 5010 7235 5030
rect 9217 5080 9237 5100
rect 9339 5080 9359 5100
rect 9435 5080 9455 5100
rect 9545 5080 9565 5100
rect 9641 5080 9661 5100
rect 11072 5022 11092 5042
rect 11168 5022 11188 5042
rect 11278 5022 11298 5042
rect 11374 5022 11394 5042
rect 11496 5022 11516 5042
rect 13485 5093 13505 5113
rect 11592 5022 11612 5042
rect 13581 5093 13601 5113
rect 13703 5093 13723 5113
rect 13799 5093 13819 5113
rect 13909 5093 13929 5113
rect 14005 5093 14025 5113
rect 20804 5231 20824 5251
rect 20900 5231 20920 5251
rect 21010 5231 21030 5251
rect 21106 5231 21126 5251
rect 21228 5231 21248 5251
rect 23008 5308 23028 5328
rect 23130 5308 23150 5328
rect 23226 5308 23246 5328
rect 23336 5308 23356 5328
rect 23432 5308 23452 5328
rect 28747 5440 28767 5460
rect 28843 5440 28863 5460
rect 28953 5440 28973 5460
rect 29049 5440 29069 5460
rect 29171 5440 29191 5460
rect 30951 5517 30971 5537
rect 31073 5517 31093 5537
rect 31169 5517 31189 5537
rect 31279 5517 31299 5537
rect 31375 5517 31395 5537
rect 29267 5440 29287 5460
rect 27289 5320 27309 5340
rect 21324 5231 21344 5251
rect 25168 5244 25188 5264
rect 25264 5244 25284 5264
rect 25374 5244 25394 5264
rect 25470 5244 25490 5264
rect 25592 5244 25612 5264
rect 27385 5320 27405 5340
rect 27507 5320 27527 5340
rect 27603 5320 27623 5340
rect 27713 5320 27733 5340
rect 27809 5320 27829 5340
rect 33111 5453 33131 5473
rect 33207 5453 33227 5473
rect 33317 5453 33337 5473
rect 33413 5453 33433 5473
rect 33535 5453 33555 5473
rect 33631 5453 33651 5473
rect 31653 5333 31673 5353
rect 25688 5244 25708 5264
rect 15436 5035 15456 5055
rect 15532 5035 15552 5055
rect 15642 5035 15662 5055
rect 15738 5035 15758 5055
rect 15860 5035 15880 5055
rect 15956 5035 15976 5055
rect 17751 5067 17771 5087
rect 17847 5067 17867 5087
rect 17969 5067 17989 5087
rect 18065 5067 18085 5087
rect 18175 5067 18195 5087
rect 18271 5067 18291 5087
rect 29545 5256 29565 5276
rect 29641 5256 29661 5276
rect 29751 5256 29771 5276
rect 29847 5256 29867 5276
rect 29969 5256 29989 5276
rect 31749 5333 31769 5353
rect 31871 5333 31891 5353
rect 31967 5333 31987 5353
rect 32077 5333 32097 5353
rect 32173 5333 32193 5353
rect 30065 5256 30085 5276
rect 19702 5009 19722 5029
rect 19798 5009 19818 5029
rect 19908 5009 19928 5029
rect 20004 5009 20024 5029
rect 20126 5009 20146 5029
rect 22115 5080 22135 5100
rect 20222 5009 20242 5029
rect 22211 5080 22231 5100
rect 22333 5080 22353 5100
rect 22429 5080 22449 5100
rect 22539 5080 22559 5100
rect 22635 5080 22655 5100
rect 33909 5269 33929 5289
rect 34005 5269 34025 5289
rect 34115 5269 34135 5289
rect 34211 5269 34231 5289
rect 34333 5269 34353 5289
rect 34429 5269 34449 5289
rect 24066 5022 24086 5042
rect 24162 5022 24182 5042
rect 24272 5022 24292 5042
rect 24368 5022 24388 5042
rect 24490 5022 24510 5042
rect 26492 5092 26512 5112
rect 24586 5022 24606 5042
rect 26588 5092 26608 5112
rect 26710 5092 26730 5112
rect 26806 5092 26826 5112
rect 26916 5092 26936 5112
rect 27012 5092 27032 5112
rect 28443 5034 28463 5054
rect 28539 5034 28559 5054
rect 28649 5034 28669 5054
rect 28745 5034 28765 5054
rect 28867 5034 28887 5054
rect 30856 5105 30876 5125
rect 28963 5034 28983 5054
rect 30952 5105 30972 5125
rect 31074 5105 31094 5125
rect 31170 5105 31190 5125
rect 31280 5105 31300 5125
rect 31376 5105 31396 5125
rect 32807 5047 32827 5067
rect 32903 5047 32923 5067
rect 33013 5047 33033 5067
rect 33109 5047 33129 5067
rect 33231 5047 33251 5067
rect 33327 5047 33347 5067
rect 1462 4671 1482 4691
rect 1558 4671 1578 4691
rect 1680 4671 1700 4691
rect 1776 4671 1796 4691
rect 1886 4671 1906 4691
rect 1982 4671 2002 4691
rect 3413 4613 3433 4633
rect 3509 4613 3529 4633
rect 3619 4613 3639 4633
rect 3715 4613 3735 4633
rect 3837 4613 3857 4633
rect 5826 4684 5846 4704
rect 3933 4613 3953 4633
rect 5922 4684 5942 4704
rect 6044 4684 6064 4704
rect 6140 4684 6160 4704
rect 6250 4684 6270 4704
rect 6346 4684 6366 4704
rect 7777 4626 7797 4646
rect 7873 4626 7893 4646
rect 7983 4626 8003 4646
rect 8079 4626 8099 4646
rect 8201 4626 8221 4646
rect 10203 4696 10223 4716
rect 8297 4626 8317 4646
rect 10299 4696 10319 4716
rect 10421 4696 10441 4716
rect 10517 4696 10537 4716
rect 10627 4696 10647 4716
rect 10723 4696 10743 4716
rect 360 4449 380 4469
rect 456 4449 476 4469
rect 578 4449 598 4469
rect 674 4449 694 4469
rect 784 4449 804 4469
rect 880 4449 900 4469
rect 12154 4638 12174 4658
rect 12250 4638 12270 4658
rect 12360 4638 12380 4658
rect 12456 4638 12476 4658
rect 12578 4638 12598 4658
rect 14567 4709 14587 4729
rect 12674 4638 12694 4658
rect 14663 4709 14683 4729
rect 14785 4709 14805 4729
rect 14881 4709 14901 4729
rect 14991 4709 15011 4729
rect 15087 4709 15107 4729
rect 4724 4462 4744 4482
rect 2616 4385 2636 4405
rect 2712 4385 2732 4405
rect 2822 4385 2842 4405
rect 2918 4385 2938 4405
rect 3040 4385 3060 4405
rect 4820 4462 4840 4482
rect 4942 4462 4962 4482
rect 5038 4462 5058 4482
rect 5148 4462 5168 4482
rect 5244 4462 5264 4482
rect 16518 4651 16538 4671
rect 16614 4651 16634 4671
rect 16724 4651 16744 4671
rect 16820 4651 16840 4671
rect 16942 4651 16962 4671
rect 17038 4651 17058 4671
rect 18833 4683 18853 4703
rect 18929 4683 18949 4703
rect 19051 4683 19071 4703
rect 19147 4683 19167 4703
rect 19257 4683 19277 4703
rect 19353 4683 19373 4703
rect 9101 4474 9121 4494
rect 3136 4385 3156 4405
rect 1158 4265 1178 4285
rect 1254 4265 1274 4285
rect 1376 4265 1396 4285
rect 1472 4265 1492 4285
rect 1582 4265 1602 4285
rect 1678 4265 1698 4285
rect 6980 4398 7000 4418
rect 7076 4398 7096 4418
rect 7186 4398 7206 4418
rect 7282 4398 7302 4418
rect 7404 4398 7424 4418
rect 9197 4474 9217 4494
rect 9319 4474 9339 4494
rect 9415 4474 9435 4494
rect 9525 4474 9545 4494
rect 9621 4474 9641 4494
rect 13465 4487 13485 4507
rect 7500 4398 7520 4418
rect 5522 4278 5542 4298
rect 3414 4201 3434 4221
rect 3510 4201 3530 4221
rect 3620 4201 3640 4221
rect 3716 4201 3736 4221
rect 3838 4201 3858 4221
rect 5618 4278 5638 4298
rect 5740 4278 5760 4298
rect 5836 4278 5856 4298
rect 5946 4278 5966 4298
rect 6042 4278 6062 4298
rect 11357 4410 11377 4430
rect 11453 4410 11473 4430
rect 11563 4410 11583 4430
rect 11659 4410 11679 4430
rect 11781 4410 11801 4430
rect 13561 4487 13581 4507
rect 13683 4487 13703 4507
rect 13779 4487 13799 4507
rect 13889 4487 13909 4507
rect 13985 4487 14005 4507
rect 20784 4625 20804 4645
rect 20880 4625 20900 4645
rect 20990 4625 21010 4645
rect 21086 4625 21106 4645
rect 21208 4625 21228 4645
rect 23197 4696 23217 4716
rect 21304 4625 21324 4645
rect 23293 4696 23313 4716
rect 23415 4696 23435 4716
rect 23511 4696 23531 4716
rect 23621 4696 23641 4716
rect 23717 4696 23737 4716
rect 25148 4638 25168 4658
rect 25244 4638 25264 4658
rect 25354 4638 25374 4658
rect 25450 4638 25470 4658
rect 25572 4638 25592 4658
rect 27574 4708 27594 4728
rect 25668 4638 25688 4658
rect 27670 4708 27690 4728
rect 27792 4708 27812 4728
rect 27888 4708 27908 4728
rect 27998 4708 28018 4728
rect 28094 4708 28114 4728
rect 11877 4410 11897 4430
rect 9899 4290 9919 4310
rect 3934 4201 3954 4221
rect 7778 4214 7798 4234
rect 7874 4214 7894 4234
rect 7984 4214 8004 4234
rect 8080 4214 8100 4234
rect 8202 4214 8222 4234
rect 9995 4290 10015 4310
rect 10117 4290 10137 4310
rect 10213 4290 10233 4310
rect 10323 4290 10343 4310
rect 10419 4290 10439 4310
rect 15721 4423 15741 4443
rect 15817 4423 15837 4443
rect 15927 4423 15947 4443
rect 16023 4423 16043 4443
rect 16145 4423 16165 4443
rect 17731 4461 17751 4481
rect 16241 4423 16261 4443
rect 17827 4461 17847 4481
rect 17949 4461 17969 4481
rect 18045 4461 18065 4481
rect 18155 4461 18175 4481
rect 18251 4461 18271 4481
rect 29525 4650 29545 4670
rect 29621 4650 29641 4670
rect 29731 4650 29751 4670
rect 29827 4650 29847 4670
rect 29949 4650 29969 4670
rect 31938 4721 31958 4741
rect 30045 4650 30065 4670
rect 32034 4721 32054 4741
rect 32156 4721 32176 4741
rect 32252 4721 32272 4741
rect 32362 4721 32382 4741
rect 32458 4721 32478 4741
rect 22095 4474 22115 4494
rect 14263 4303 14283 4323
rect 8298 4214 8318 4234
rect 361 4037 381 4057
rect 457 4037 477 4057
rect 579 4037 599 4057
rect 675 4037 695 4057
rect 785 4037 805 4057
rect 881 4037 901 4057
rect 12155 4226 12175 4246
rect 12251 4226 12271 4246
rect 12361 4226 12381 4246
rect 12457 4226 12477 4246
rect 12579 4226 12599 4246
rect 14359 4303 14379 4323
rect 14481 4303 14501 4323
rect 14577 4303 14597 4323
rect 14687 4303 14707 4323
rect 14783 4303 14803 4323
rect 19987 4397 20007 4417
rect 20083 4397 20103 4417
rect 20193 4397 20213 4417
rect 20289 4397 20309 4417
rect 20411 4397 20431 4417
rect 22191 4474 22211 4494
rect 22313 4474 22333 4494
rect 22409 4474 22429 4494
rect 22519 4474 22539 4494
rect 22615 4474 22635 4494
rect 33889 4663 33909 4683
rect 33985 4663 34005 4683
rect 34095 4663 34115 4683
rect 34191 4663 34211 4683
rect 34313 4663 34333 4683
rect 34409 4663 34429 4683
rect 26472 4486 26492 4506
rect 20507 4397 20527 4417
rect 12675 4226 12695 4246
rect 2517 3975 2537 3995
rect 2613 3975 2633 3995
rect 2723 3975 2743 3995
rect 2819 3975 2839 3995
rect 2941 3975 2961 3995
rect 4725 4050 4745 4070
rect 3037 3975 3057 3995
rect 4821 4050 4841 4070
rect 4943 4050 4963 4070
rect 5039 4050 5059 4070
rect 5149 4050 5169 4070
rect 5245 4050 5265 4070
rect 16519 4239 16539 4259
rect 16615 4239 16635 4259
rect 16725 4239 16745 4259
rect 16821 4239 16841 4259
rect 16943 4239 16963 4259
rect 18529 4277 18549 4297
rect 17039 4239 17059 4259
rect 18625 4277 18645 4297
rect 18747 4277 18767 4297
rect 18843 4277 18863 4297
rect 18953 4277 18973 4297
rect 19049 4277 19069 4297
rect 24351 4410 24371 4430
rect 24447 4410 24467 4430
rect 24557 4410 24577 4430
rect 24653 4410 24673 4430
rect 24775 4410 24795 4430
rect 26568 4486 26588 4506
rect 26690 4486 26710 4506
rect 26786 4486 26806 4506
rect 26896 4486 26916 4506
rect 26992 4486 27012 4506
rect 30836 4499 30856 4519
rect 24871 4410 24891 4430
rect 22893 4290 22913 4310
rect 6881 3988 6901 4008
rect 6977 3988 6997 4008
rect 7087 3988 7107 4008
rect 7183 3988 7203 4008
rect 7305 3988 7325 4008
rect 9102 4062 9122 4082
rect 7401 3988 7421 4008
rect 9198 4062 9218 4082
rect 9320 4062 9340 4082
rect 9416 4062 9436 4082
rect 9526 4062 9546 4082
rect 9622 4062 9642 4082
rect 20785 4213 20805 4233
rect 20881 4213 20901 4233
rect 20991 4213 21011 4233
rect 21087 4213 21107 4233
rect 21209 4213 21229 4233
rect 22989 4290 23009 4310
rect 23111 4290 23131 4310
rect 23207 4290 23227 4310
rect 23317 4290 23337 4310
rect 23413 4290 23433 4310
rect 28728 4422 28748 4442
rect 28824 4422 28844 4442
rect 28934 4422 28954 4442
rect 29030 4422 29050 4442
rect 29152 4422 29172 4442
rect 30932 4499 30952 4519
rect 31054 4499 31074 4519
rect 31150 4499 31170 4519
rect 31260 4499 31280 4519
rect 31356 4499 31376 4519
rect 29248 4422 29268 4442
rect 27270 4302 27290 4322
rect 21305 4213 21325 4233
rect 11258 4000 11278 4020
rect 11354 4000 11374 4020
rect 11464 4000 11484 4020
rect 11560 4000 11580 4020
rect 11682 4000 11702 4020
rect 13466 4075 13486 4095
rect 11778 4000 11798 4020
rect 13562 4075 13582 4095
rect 13684 4075 13704 4095
rect 13780 4075 13800 4095
rect 13890 4075 13910 4095
rect 13986 4075 14006 4095
rect 25149 4226 25169 4246
rect 25245 4226 25265 4246
rect 25355 4226 25375 4246
rect 25451 4226 25471 4246
rect 25573 4226 25593 4246
rect 27366 4302 27386 4322
rect 27488 4302 27508 4322
rect 27584 4302 27604 4322
rect 27694 4302 27714 4322
rect 27790 4302 27810 4322
rect 33092 4435 33112 4455
rect 33188 4435 33208 4455
rect 33298 4435 33318 4455
rect 33394 4435 33414 4455
rect 33516 4435 33536 4455
rect 33612 4435 33632 4455
rect 31634 4315 31654 4335
rect 25669 4226 25689 4246
rect 15622 4013 15642 4033
rect 15718 4013 15738 4033
rect 15828 4013 15848 4033
rect 15924 4013 15944 4033
rect 16046 4013 16066 4033
rect 16142 4013 16162 4033
rect 17732 4049 17752 4069
rect 17828 4049 17848 4069
rect 17950 4049 17970 4069
rect 18046 4049 18066 4069
rect 18156 4049 18176 4069
rect 18252 4049 18272 4069
rect 29526 4238 29546 4258
rect 29622 4238 29642 4258
rect 29732 4238 29752 4258
rect 29828 4238 29848 4258
rect 29950 4238 29970 4258
rect 31730 4315 31750 4335
rect 31852 4315 31872 4335
rect 31948 4315 31968 4335
rect 32058 4315 32078 4335
rect 32154 4315 32174 4335
rect 30046 4238 30066 4258
rect 19888 3987 19908 4007
rect 19984 3987 20004 4007
rect 20094 3987 20114 4007
rect 20190 3987 20210 4007
rect 20312 3987 20332 4007
rect 22096 4062 22116 4082
rect 20408 3987 20428 4007
rect 22192 4062 22212 4082
rect 22314 4062 22334 4082
rect 22410 4062 22430 4082
rect 22520 4062 22540 4082
rect 22616 4062 22636 4082
rect 33890 4251 33910 4271
rect 33986 4251 34006 4271
rect 34096 4251 34116 4271
rect 34192 4251 34212 4271
rect 34314 4251 34334 4271
rect 34410 4251 34430 4271
rect 24252 4000 24272 4020
rect 24348 4000 24368 4020
rect 24458 4000 24478 4020
rect 24554 4000 24574 4020
rect 24676 4000 24696 4020
rect 26473 4074 26493 4094
rect 24772 4000 24792 4020
rect 26569 4074 26589 4094
rect 26691 4074 26711 4094
rect 26787 4074 26807 4094
rect 26897 4074 26917 4094
rect 26993 4074 27013 4094
rect 28629 4012 28649 4032
rect 28725 4012 28745 4032
rect 28835 4012 28855 4032
rect 28931 4012 28951 4032
rect 29053 4012 29073 4032
rect 30837 4087 30857 4107
rect 29149 4012 29169 4032
rect 30933 4087 30953 4107
rect 31055 4087 31075 4107
rect 31151 4087 31171 4107
rect 31261 4087 31281 4107
rect 31357 4087 31377 4107
rect 32993 4025 33013 4045
rect 33089 4025 33109 4045
rect 33199 4025 33219 4045
rect 33295 4025 33315 4045
rect 33417 4025 33437 4045
rect 33513 4025 33533 4045
rect 1240 3657 1260 3677
rect 1336 3657 1356 3677
rect 1458 3657 1478 3677
rect 1554 3657 1574 3677
rect 1664 3657 1684 3677
rect 1760 3657 1780 3677
rect 3396 3595 3416 3615
rect 3492 3595 3512 3615
rect 3602 3595 3622 3615
rect 3698 3595 3718 3615
rect 3820 3595 3840 3615
rect 5604 3670 5624 3690
rect 3916 3595 3936 3615
rect 5700 3670 5720 3690
rect 5822 3670 5842 3690
rect 5918 3670 5938 3690
rect 6028 3670 6048 3690
rect 6124 3670 6144 3690
rect 7760 3608 7780 3628
rect 7856 3608 7876 3628
rect 7966 3608 7986 3628
rect 8062 3608 8082 3628
rect 8184 3608 8204 3628
rect 9981 3682 10001 3702
rect 8280 3608 8300 3628
rect 10077 3682 10097 3702
rect 10199 3682 10219 3702
rect 10295 3682 10315 3702
rect 10405 3682 10425 3702
rect 10501 3682 10521 3702
rect 343 3431 363 3451
rect 439 3431 459 3451
rect 561 3431 581 3451
rect 657 3431 677 3451
rect 767 3431 787 3451
rect 863 3431 883 3451
rect 12137 3620 12157 3640
rect 12233 3620 12253 3640
rect 12343 3620 12363 3640
rect 12439 3620 12459 3640
rect 12561 3620 12581 3640
rect 14345 3695 14365 3715
rect 12657 3620 12677 3640
rect 14441 3695 14461 3715
rect 14563 3695 14583 3715
rect 14659 3695 14679 3715
rect 14769 3695 14789 3715
rect 14865 3695 14885 3715
rect 4707 3444 4727 3464
rect 2599 3367 2619 3387
rect 2695 3367 2715 3387
rect 2805 3367 2825 3387
rect 2901 3367 2921 3387
rect 3023 3367 3043 3387
rect 4803 3444 4823 3464
rect 4925 3444 4945 3464
rect 5021 3444 5041 3464
rect 5131 3444 5151 3464
rect 5227 3444 5247 3464
rect 16501 3633 16521 3653
rect 16597 3633 16617 3653
rect 16707 3633 16727 3653
rect 16803 3633 16823 3653
rect 16925 3633 16945 3653
rect 17021 3633 17041 3653
rect 18611 3669 18631 3689
rect 18707 3669 18727 3689
rect 18829 3669 18849 3689
rect 18925 3669 18945 3689
rect 19035 3669 19055 3689
rect 19131 3669 19151 3689
rect 9084 3456 9104 3476
rect 3119 3367 3139 3387
rect 1141 3247 1161 3267
rect 1237 3247 1257 3267
rect 1359 3247 1379 3267
rect 1455 3247 1475 3267
rect 1565 3247 1585 3267
rect 1661 3247 1681 3267
rect 6963 3380 6983 3400
rect 7059 3380 7079 3400
rect 7169 3380 7189 3400
rect 7265 3380 7285 3400
rect 7387 3380 7407 3400
rect 9180 3456 9200 3476
rect 9302 3456 9322 3476
rect 9398 3456 9418 3476
rect 9508 3456 9528 3476
rect 9604 3456 9624 3476
rect 20767 3607 20787 3627
rect 20863 3607 20883 3627
rect 20973 3607 20993 3627
rect 21069 3607 21089 3627
rect 21191 3607 21211 3627
rect 22975 3682 22995 3702
rect 21287 3607 21307 3627
rect 23071 3682 23091 3702
rect 23193 3682 23213 3702
rect 23289 3682 23309 3702
rect 23399 3682 23419 3702
rect 23495 3682 23515 3702
rect 13448 3469 13468 3489
rect 7483 3380 7503 3400
rect 5505 3260 5525 3280
rect 3397 3183 3417 3203
rect 3493 3183 3513 3203
rect 3603 3183 3623 3203
rect 3699 3183 3719 3203
rect 3821 3183 3841 3203
rect 5601 3260 5621 3280
rect 5723 3260 5743 3280
rect 5819 3260 5839 3280
rect 5929 3260 5949 3280
rect 6025 3260 6045 3280
rect 11340 3392 11360 3412
rect 11436 3392 11456 3412
rect 11546 3392 11566 3412
rect 11642 3392 11662 3412
rect 11764 3392 11784 3412
rect 13544 3469 13564 3489
rect 13666 3469 13686 3489
rect 13762 3469 13782 3489
rect 13872 3469 13892 3489
rect 13968 3469 13988 3489
rect 25131 3620 25151 3640
rect 25227 3620 25247 3640
rect 25337 3620 25357 3640
rect 25433 3620 25453 3640
rect 25555 3620 25575 3640
rect 27352 3694 27372 3714
rect 25651 3620 25671 3640
rect 27448 3694 27468 3714
rect 27570 3694 27590 3714
rect 27666 3694 27686 3714
rect 27776 3694 27796 3714
rect 27872 3694 27892 3714
rect 11860 3392 11880 3412
rect 9882 3272 9902 3292
rect 3917 3183 3937 3203
rect 7761 3196 7781 3216
rect 7857 3196 7877 3216
rect 7967 3196 7987 3216
rect 8063 3196 8083 3216
rect 8185 3196 8205 3216
rect 9978 3272 9998 3292
rect 10100 3272 10120 3292
rect 10196 3272 10216 3292
rect 10306 3272 10326 3292
rect 10402 3272 10422 3292
rect 15704 3405 15724 3425
rect 15800 3405 15820 3425
rect 15910 3405 15930 3425
rect 16006 3405 16026 3425
rect 16128 3405 16148 3425
rect 17714 3443 17734 3463
rect 16224 3405 16244 3425
rect 17810 3443 17830 3463
rect 17932 3443 17952 3463
rect 18028 3443 18048 3463
rect 18138 3443 18158 3463
rect 18234 3443 18254 3463
rect 29508 3632 29528 3652
rect 29604 3632 29624 3652
rect 29714 3632 29734 3652
rect 29810 3632 29830 3652
rect 29932 3632 29952 3652
rect 31716 3707 31736 3727
rect 30028 3632 30048 3652
rect 31812 3707 31832 3727
rect 31934 3707 31954 3727
rect 32030 3707 32050 3727
rect 32140 3707 32160 3727
rect 32236 3707 32256 3727
rect 22078 3456 22098 3476
rect 14246 3285 14266 3305
rect 8281 3196 8301 3216
rect 344 3019 364 3039
rect 440 3019 460 3039
rect 562 3019 582 3039
rect 658 3019 678 3039
rect 768 3019 788 3039
rect 864 3019 884 3039
rect 12138 3208 12158 3228
rect 12234 3208 12254 3228
rect 12344 3208 12364 3228
rect 12440 3208 12460 3228
rect 12562 3208 12582 3228
rect 14342 3285 14362 3305
rect 14464 3285 14484 3305
rect 14560 3285 14580 3305
rect 14670 3285 14690 3305
rect 14766 3285 14786 3305
rect 19970 3379 19990 3399
rect 20066 3379 20086 3399
rect 20176 3379 20196 3399
rect 20272 3379 20292 3399
rect 20394 3379 20414 3399
rect 22174 3456 22194 3476
rect 22296 3456 22316 3476
rect 22392 3456 22412 3476
rect 22502 3456 22522 3476
rect 22598 3456 22618 3476
rect 33872 3645 33892 3665
rect 33968 3645 33988 3665
rect 34078 3645 34098 3665
rect 34174 3645 34194 3665
rect 34296 3645 34316 3665
rect 34392 3645 34412 3665
rect 26455 3468 26475 3488
rect 20490 3379 20510 3399
rect 12658 3208 12678 3228
rect 2434 2959 2454 2979
rect 2530 2959 2550 2979
rect 2640 2959 2660 2979
rect 2736 2959 2756 2979
rect 2858 2959 2878 2979
rect 4708 3032 4728 3052
rect 2954 2959 2974 2979
rect 4804 3032 4824 3052
rect 4926 3032 4946 3052
rect 5022 3032 5042 3052
rect 5132 3032 5152 3052
rect 5228 3032 5248 3052
rect 16502 3221 16522 3241
rect 16598 3221 16618 3241
rect 16708 3221 16728 3241
rect 16804 3221 16824 3241
rect 16926 3221 16946 3241
rect 18512 3259 18532 3279
rect 17022 3221 17042 3241
rect 18608 3259 18628 3279
rect 18730 3259 18750 3279
rect 18826 3259 18846 3279
rect 18936 3259 18956 3279
rect 19032 3259 19052 3279
rect 24334 3392 24354 3412
rect 24430 3392 24450 3412
rect 24540 3392 24560 3412
rect 24636 3392 24656 3412
rect 24758 3392 24778 3412
rect 26551 3468 26571 3488
rect 26673 3468 26693 3488
rect 26769 3468 26789 3488
rect 26879 3468 26899 3488
rect 26975 3468 26995 3488
rect 30819 3481 30839 3501
rect 24854 3392 24874 3412
rect 22876 3272 22896 3292
rect 6798 2972 6818 2992
rect 6894 2972 6914 2992
rect 7004 2972 7024 2992
rect 7100 2972 7120 2992
rect 7222 2972 7242 2992
rect 9085 3044 9105 3064
rect 7318 2972 7338 2992
rect 9181 3044 9201 3064
rect 9303 3044 9323 3064
rect 9399 3044 9419 3064
rect 9509 3044 9529 3064
rect 9605 3044 9625 3064
rect 20768 3195 20788 3215
rect 20864 3195 20884 3215
rect 20974 3195 20994 3215
rect 21070 3195 21090 3215
rect 21192 3195 21212 3215
rect 22972 3272 22992 3292
rect 23094 3272 23114 3292
rect 23190 3272 23210 3292
rect 23300 3272 23320 3292
rect 23396 3272 23416 3292
rect 28711 3404 28731 3424
rect 28807 3404 28827 3424
rect 28917 3404 28937 3424
rect 29013 3404 29033 3424
rect 29135 3404 29155 3424
rect 30915 3481 30935 3501
rect 31037 3481 31057 3501
rect 31133 3481 31153 3501
rect 31243 3481 31263 3501
rect 31339 3481 31359 3501
rect 29231 3404 29251 3424
rect 27253 3284 27273 3304
rect 21288 3195 21308 3215
rect 11175 2984 11195 3004
rect 11271 2984 11291 3004
rect 11381 2984 11401 3004
rect 11477 2984 11497 3004
rect 11599 2984 11619 3004
rect 13449 3057 13469 3077
rect 11695 2984 11715 3004
rect 13545 3057 13565 3077
rect 13667 3057 13687 3077
rect 13763 3057 13783 3077
rect 13873 3057 13893 3077
rect 13969 3057 13989 3077
rect 25132 3208 25152 3228
rect 25228 3208 25248 3228
rect 25338 3208 25358 3228
rect 25434 3208 25454 3228
rect 25556 3208 25576 3228
rect 27349 3284 27369 3304
rect 27471 3284 27491 3304
rect 27567 3284 27587 3304
rect 27677 3284 27697 3304
rect 27773 3284 27793 3304
rect 33075 3417 33095 3437
rect 33171 3417 33191 3437
rect 33281 3417 33301 3437
rect 33377 3417 33397 3437
rect 33499 3417 33519 3437
rect 33595 3417 33615 3437
rect 31617 3297 31637 3317
rect 25652 3208 25672 3228
rect 15539 2997 15559 3017
rect 15635 2997 15655 3017
rect 15745 2997 15765 3017
rect 15841 2997 15861 3017
rect 15963 2997 15983 3017
rect 16059 2997 16079 3017
rect 17715 3031 17735 3051
rect 17811 3031 17831 3051
rect 17933 3031 17953 3051
rect 18029 3031 18049 3051
rect 18139 3031 18159 3051
rect 18235 3031 18255 3051
rect 29509 3220 29529 3240
rect 29605 3220 29625 3240
rect 29715 3220 29735 3240
rect 29811 3220 29831 3240
rect 29933 3220 29953 3240
rect 31713 3297 31733 3317
rect 31835 3297 31855 3317
rect 31931 3297 31951 3317
rect 32041 3297 32061 3317
rect 32137 3297 32157 3317
rect 30029 3220 30049 3240
rect 19805 2971 19825 2991
rect 19901 2971 19921 2991
rect 20011 2971 20031 2991
rect 20107 2971 20127 2991
rect 20229 2971 20249 2991
rect 22079 3044 22099 3064
rect 20325 2971 20345 2991
rect 22175 3044 22195 3064
rect 22297 3044 22317 3064
rect 22393 3044 22413 3064
rect 22503 3044 22523 3064
rect 22599 3044 22619 3064
rect 33873 3233 33893 3253
rect 33969 3233 33989 3253
rect 34079 3233 34099 3253
rect 34175 3233 34195 3253
rect 34297 3233 34317 3253
rect 34393 3233 34413 3253
rect 24169 2984 24189 3004
rect 24265 2984 24285 3004
rect 24375 2984 24395 3004
rect 24471 2984 24491 3004
rect 24593 2984 24613 3004
rect 26456 3056 26476 3076
rect 24689 2984 24709 3004
rect 26552 3056 26572 3076
rect 26674 3056 26694 3076
rect 26770 3056 26790 3076
rect 26880 3056 26900 3076
rect 26976 3056 26996 3076
rect 28546 2996 28566 3016
rect 28642 2996 28662 3016
rect 28752 2996 28772 3016
rect 28848 2996 28868 3016
rect 28970 2996 28990 3016
rect 30820 3069 30840 3089
rect 29066 2996 29086 3016
rect 30916 3069 30936 3089
rect 31038 3069 31058 3089
rect 31134 3069 31154 3089
rect 31244 3069 31264 3089
rect 31340 3069 31360 3089
rect 32910 3009 32930 3029
rect 33006 3009 33026 3029
rect 33116 3009 33136 3029
rect 33212 3009 33232 3029
rect 33334 3009 33354 3029
rect 33430 3009 33450 3029
rect 1286 2637 1306 2657
rect 1382 2637 1402 2657
rect 1504 2637 1524 2657
rect 1600 2637 1620 2657
rect 1710 2637 1730 2657
rect 1806 2637 1826 2657
rect 3376 2577 3396 2597
rect 3472 2577 3492 2597
rect 3582 2577 3602 2597
rect 3678 2577 3698 2597
rect 3800 2577 3820 2597
rect 5650 2650 5670 2670
rect 3896 2577 3916 2597
rect 5746 2650 5766 2670
rect 5868 2650 5888 2670
rect 5964 2650 5984 2670
rect 6074 2650 6094 2670
rect 6170 2650 6190 2670
rect 7740 2590 7760 2610
rect 7836 2590 7856 2610
rect 7946 2590 7966 2610
rect 8042 2590 8062 2610
rect 8164 2590 8184 2610
rect 10027 2662 10047 2682
rect 8260 2590 8280 2610
rect 10123 2662 10143 2682
rect 10245 2662 10265 2682
rect 10341 2662 10361 2682
rect 10451 2662 10471 2682
rect 10547 2662 10567 2682
rect 323 2413 343 2433
rect 419 2413 439 2433
rect 541 2413 561 2433
rect 637 2413 657 2433
rect 747 2413 767 2433
rect 843 2413 863 2433
rect 12117 2602 12137 2622
rect 12213 2602 12233 2622
rect 12323 2602 12343 2622
rect 12419 2602 12439 2622
rect 12541 2602 12561 2622
rect 14391 2675 14411 2695
rect 12637 2602 12657 2622
rect 14487 2675 14507 2695
rect 14609 2675 14629 2695
rect 14705 2675 14725 2695
rect 14815 2675 14835 2695
rect 14911 2675 14931 2695
rect 4687 2426 4707 2446
rect 2579 2349 2599 2369
rect 2675 2349 2695 2369
rect 2785 2349 2805 2369
rect 2881 2349 2901 2369
rect 3003 2349 3023 2369
rect 4783 2426 4803 2446
rect 4905 2426 4925 2446
rect 5001 2426 5021 2446
rect 5111 2426 5131 2446
rect 5207 2426 5227 2446
rect 16481 2615 16501 2635
rect 16577 2615 16597 2635
rect 16687 2615 16707 2635
rect 16783 2615 16803 2635
rect 16905 2615 16925 2635
rect 17001 2615 17021 2635
rect 18657 2649 18677 2669
rect 18753 2649 18773 2669
rect 18875 2649 18895 2669
rect 18971 2649 18991 2669
rect 19081 2649 19101 2669
rect 19177 2649 19197 2669
rect 9064 2438 9084 2458
rect 3099 2349 3119 2369
rect 1121 2229 1141 2249
rect 1217 2229 1237 2249
rect 1339 2229 1359 2249
rect 1435 2229 1455 2249
rect 1545 2229 1565 2249
rect 1641 2229 1661 2249
rect 6943 2362 6963 2382
rect 7039 2362 7059 2382
rect 7149 2362 7169 2382
rect 7245 2362 7265 2382
rect 7367 2362 7387 2382
rect 9160 2438 9180 2458
rect 9282 2438 9302 2458
rect 9378 2438 9398 2458
rect 9488 2438 9508 2458
rect 9584 2438 9604 2458
rect 20747 2589 20767 2609
rect 20843 2589 20863 2609
rect 20953 2589 20973 2609
rect 21049 2589 21069 2609
rect 21171 2589 21191 2609
rect 23021 2662 23041 2682
rect 21267 2589 21287 2609
rect 23117 2662 23137 2682
rect 23239 2662 23259 2682
rect 23335 2662 23355 2682
rect 23445 2662 23465 2682
rect 23541 2662 23561 2682
rect 13428 2451 13448 2471
rect 7463 2362 7483 2382
rect 5485 2242 5505 2262
rect 3377 2165 3397 2185
rect 3473 2165 3493 2185
rect 3583 2165 3603 2185
rect 3679 2165 3699 2185
rect 3801 2165 3821 2185
rect 5581 2242 5601 2262
rect 5703 2242 5723 2262
rect 5799 2242 5819 2262
rect 5909 2242 5929 2262
rect 6005 2242 6025 2262
rect 11320 2374 11340 2394
rect 11416 2374 11436 2394
rect 11526 2374 11546 2394
rect 11622 2374 11642 2394
rect 11744 2374 11764 2394
rect 13524 2451 13544 2471
rect 13646 2451 13666 2471
rect 13742 2451 13762 2471
rect 13852 2451 13872 2471
rect 13948 2451 13968 2471
rect 25111 2602 25131 2622
rect 25207 2602 25227 2622
rect 25317 2602 25337 2622
rect 25413 2602 25433 2622
rect 25535 2602 25555 2622
rect 27398 2674 27418 2694
rect 25631 2602 25651 2622
rect 27494 2674 27514 2694
rect 27616 2674 27636 2694
rect 27712 2674 27732 2694
rect 27822 2674 27842 2694
rect 27918 2674 27938 2694
rect 11840 2374 11860 2394
rect 9862 2254 9882 2274
rect 3897 2165 3917 2185
rect 7741 2178 7761 2198
rect 7837 2178 7857 2198
rect 7947 2178 7967 2198
rect 8043 2178 8063 2198
rect 8165 2178 8185 2198
rect 9958 2254 9978 2274
rect 10080 2254 10100 2274
rect 10176 2254 10196 2274
rect 10286 2254 10306 2274
rect 10382 2254 10402 2274
rect 15684 2387 15704 2407
rect 15780 2387 15800 2407
rect 15890 2387 15910 2407
rect 15986 2387 16006 2407
rect 16108 2387 16128 2407
rect 17694 2425 17714 2445
rect 16204 2387 16224 2407
rect 17790 2425 17810 2445
rect 17912 2425 17932 2445
rect 18008 2425 18028 2445
rect 18118 2425 18138 2445
rect 18214 2425 18234 2445
rect 29488 2614 29508 2634
rect 29584 2614 29604 2634
rect 29694 2614 29714 2634
rect 29790 2614 29810 2634
rect 29912 2614 29932 2634
rect 31762 2687 31782 2707
rect 30008 2614 30028 2634
rect 31858 2687 31878 2707
rect 31980 2687 32000 2707
rect 32076 2687 32096 2707
rect 32186 2687 32206 2707
rect 32282 2687 32302 2707
rect 22058 2438 22078 2458
rect 14226 2267 14246 2287
rect 8261 2178 8281 2198
rect 324 2001 344 2021
rect 420 2001 440 2021
rect 542 2001 562 2021
rect 638 2001 658 2021
rect 748 2001 768 2021
rect 844 2001 864 2021
rect 12118 2190 12138 2210
rect 12214 2190 12234 2210
rect 12324 2190 12344 2210
rect 12420 2190 12440 2210
rect 12542 2190 12562 2210
rect 14322 2267 14342 2287
rect 14444 2267 14464 2287
rect 14540 2267 14560 2287
rect 14650 2267 14670 2287
rect 14746 2267 14766 2287
rect 19950 2361 19970 2381
rect 20046 2361 20066 2381
rect 20156 2361 20176 2381
rect 20252 2361 20272 2381
rect 20374 2361 20394 2381
rect 22154 2438 22174 2458
rect 22276 2438 22296 2458
rect 22372 2438 22392 2458
rect 22482 2438 22502 2458
rect 22578 2438 22598 2458
rect 33852 2627 33872 2647
rect 33948 2627 33968 2647
rect 34058 2627 34078 2647
rect 34154 2627 34174 2647
rect 34276 2627 34296 2647
rect 34372 2627 34392 2647
rect 26435 2450 26455 2470
rect 20470 2361 20490 2381
rect 12638 2190 12658 2210
rect 2480 1939 2500 1959
rect 2576 1939 2596 1959
rect 2686 1939 2706 1959
rect 2782 1939 2802 1959
rect 2904 1939 2924 1959
rect 4688 2014 4708 2034
rect 3000 1939 3020 1959
rect 4784 2014 4804 2034
rect 4906 2014 4926 2034
rect 5002 2014 5022 2034
rect 5112 2014 5132 2034
rect 5208 2014 5228 2034
rect 16482 2203 16502 2223
rect 16578 2203 16598 2223
rect 16688 2203 16708 2223
rect 16784 2203 16804 2223
rect 16906 2203 16926 2223
rect 18492 2241 18512 2261
rect 17002 2203 17022 2223
rect 18588 2241 18608 2261
rect 18710 2241 18730 2261
rect 18806 2241 18826 2261
rect 18916 2241 18936 2261
rect 19012 2241 19032 2261
rect 24314 2374 24334 2394
rect 24410 2374 24430 2394
rect 24520 2374 24540 2394
rect 24616 2374 24636 2394
rect 24738 2374 24758 2394
rect 26531 2450 26551 2470
rect 26653 2450 26673 2470
rect 26749 2450 26769 2470
rect 26859 2450 26879 2470
rect 26955 2450 26975 2470
rect 30799 2463 30819 2483
rect 24834 2374 24854 2394
rect 22856 2254 22876 2274
rect 6844 1952 6864 1972
rect 6940 1952 6960 1972
rect 7050 1952 7070 1972
rect 7146 1952 7166 1972
rect 7268 1952 7288 1972
rect 9065 2026 9085 2046
rect 7364 1952 7384 1972
rect 9161 2026 9181 2046
rect 9283 2026 9303 2046
rect 9379 2026 9399 2046
rect 9489 2026 9509 2046
rect 9585 2026 9605 2046
rect 20748 2177 20768 2197
rect 20844 2177 20864 2197
rect 20954 2177 20974 2197
rect 21050 2177 21070 2197
rect 21172 2177 21192 2197
rect 22952 2254 22972 2274
rect 23074 2254 23094 2274
rect 23170 2254 23190 2274
rect 23280 2254 23300 2274
rect 23376 2254 23396 2274
rect 28691 2386 28711 2406
rect 28787 2386 28807 2406
rect 28897 2386 28917 2406
rect 28993 2386 29013 2406
rect 29115 2386 29135 2406
rect 30895 2463 30915 2483
rect 31017 2463 31037 2483
rect 31113 2463 31133 2483
rect 31223 2463 31243 2483
rect 31319 2463 31339 2483
rect 29211 2386 29231 2406
rect 27233 2266 27253 2286
rect 21268 2177 21288 2197
rect 11221 1964 11241 1984
rect 11317 1964 11337 1984
rect 11427 1964 11447 1984
rect 11523 1964 11543 1984
rect 11645 1964 11665 1984
rect 13429 2039 13449 2059
rect 11741 1964 11761 1984
rect 13525 2039 13545 2059
rect 13647 2039 13667 2059
rect 13743 2039 13763 2059
rect 13853 2039 13873 2059
rect 13949 2039 13969 2059
rect 25112 2190 25132 2210
rect 25208 2190 25228 2210
rect 25318 2190 25338 2210
rect 25414 2190 25434 2210
rect 25536 2190 25556 2210
rect 27329 2266 27349 2286
rect 27451 2266 27471 2286
rect 27547 2266 27567 2286
rect 27657 2266 27677 2286
rect 27753 2266 27773 2286
rect 33055 2399 33075 2419
rect 33151 2399 33171 2419
rect 33261 2399 33281 2419
rect 33357 2399 33377 2419
rect 33479 2399 33499 2419
rect 33575 2399 33595 2419
rect 31597 2279 31617 2299
rect 25632 2190 25652 2210
rect 15585 1977 15605 1997
rect 15681 1977 15701 1997
rect 15791 1977 15811 1997
rect 15887 1977 15907 1997
rect 16009 1977 16029 1997
rect 16105 1977 16125 1997
rect 17695 2013 17715 2033
rect 17791 2013 17811 2033
rect 17913 2013 17933 2033
rect 18009 2013 18029 2033
rect 18119 2013 18139 2033
rect 18215 2013 18235 2033
rect 29489 2202 29509 2222
rect 29585 2202 29605 2222
rect 29695 2202 29715 2222
rect 29791 2202 29811 2222
rect 29913 2202 29933 2222
rect 31693 2279 31713 2299
rect 31815 2279 31835 2299
rect 31911 2279 31931 2299
rect 32021 2279 32041 2299
rect 32117 2279 32137 2299
rect 30009 2202 30029 2222
rect 19851 1951 19871 1971
rect 19947 1951 19967 1971
rect 20057 1951 20077 1971
rect 20153 1951 20173 1971
rect 20275 1951 20295 1971
rect 22059 2026 22079 2046
rect 20371 1951 20391 1971
rect 22155 2026 22175 2046
rect 22277 2026 22297 2046
rect 22373 2026 22393 2046
rect 22483 2026 22503 2046
rect 22579 2026 22599 2046
rect 33853 2215 33873 2235
rect 33949 2215 33969 2235
rect 34059 2215 34079 2235
rect 34155 2215 34175 2235
rect 34277 2215 34297 2235
rect 34373 2215 34393 2235
rect 24215 1964 24235 1984
rect 24311 1964 24331 1984
rect 24421 1964 24441 1984
rect 24517 1964 24537 1984
rect 24639 1964 24659 1984
rect 26436 2038 26456 2058
rect 24735 1964 24755 1984
rect 26532 2038 26552 2058
rect 26654 2038 26674 2058
rect 26750 2038 26770 2058
rect 26860 2038 26880 2058
rect 26956 2038 26976 2058
rect 28592 1976 28612 1996
rect 28688 1976 28708 1996
rect 28798 1976 28818 1996
rect 28894 1976 28914 1996
rect 29016 1976 29036 1996
rect 30800 2051 30820 2071
rect 29112 1976 29132 1996
rect 30896 2051 30916 2071
rect 31018 2051 31038 2071
rect 31114 2051 31134 2071
rect 31224 2051 31244 2071
rect 31320 2051 31340 2071
rect 32956 1989 32976 2009
rect 33052 1989 33072 2009
rect 33162 1989 33182 2009
rect 33258 1989 33278 2009
rect 33380 1989 33400 2009
rect 33476 1989 33496 2009
rect 1203 1621 1223 1641
rect 1299 1621 1319 1641
rect 1421 1621 1441 1641
rect 1517 1621 1537 1641
rect 1627 1621 1647 1641
rect 1723 1621 1743 1641
rect 3359 1559 3379 1579
rect 3455 1559 3475 1579
rect 3565 1559 3585 1579
rect 3661 1559 3681 1579
rect 3783 1559 3803 1579
rect 5567 1634 5587 1654
rect 3879 1559 3899 1579
rect 5663 1634 5683 1654
rect 5785 1634 5805 1654
rect 5881 1634 5901 1654
rect 5991 1634 6011 1654
rect 6087 1634 6107 1654
rect 7723 1572 7743 1592
rect 7819 1572 7839 1592
rect 7929 1572 7949 1592
rect 8025 1572 8045 1592
rect 8147 1572 8167 1592
rect 9944 1646 9964 1666
rect 8243 1572 8263 1592
rect 10040 1646 10060 1666
rect 10162 1646 10182 1666
rect 10258 1646 10278 1666
rect 10368 1646 10388 1666
rect 10464 1646 10484 1666
rect 306 1395 326 1415
rect 402 1395 422 1415
rect 524 1395 544 1415
rect 620 1395 640 1415
rect 730 1395 750 1415
rect 826 1395 846 1415
rect 12100 1584 12120 1604
rect 12196 1584 12216 1604
rect 12306 1584 12326 1604
rect 12402 1584 12422 1604
rect 12524 1584 12544 1604
rect 14308 1659 14328 1679
rect 12620 1584 12640 1604
rect 14404 1659 14424 1679
rect 14526 1659 14546 1679
rect 14622 1659 14642 1679
rect 14732 1659 14752 1679
rect 14828 1659 14848 1679
rect 4670 1408 4690 1428
rect 2562 1331 2582 1351
rect 2658 1331 2678 1351
rect 2768 1331 2788 1351
rect 2864 1331 2884 1351
rect 2986 1331 3006 1351
rect 4766 1408 4786 1428
rect 4888 1408 4908 1428
rect 4984 1408 5004 1428
rect 5094 1408 5114 1428
rect 5190 1408 5210 1428
rect 16464 1597 16484 1617
rect 16560 1597 16580 1617
rect 16670 1597 16690 1617
rect 16766 1597 16786 1617
rect 16888 1597 16908 1617
rect 16984 1597 17004 1617
rect 18574 1633 18594 1653
rect 18670 1633 18690 1653
rect 18792 1633 18812 1653
rect 18888 1633 18908 1653
rect 18998 1633 19018 1653
rect 19094 1633 19114 1653
rect 9047 1420 9067 1440
rect 3082 1331 3102 1351
rect 1104 1211 1124 1231
rect 1200 1211 1220 1231
rect 1322 1211 1342 1231
rect 1418 1211 1438 1231
rect 1528 1211 1548 1231
rect 1624 1211 1644 1231
rect 6926 1344 6946 1364
rect 7022 1344 7042 1364
rect 7132 1344 7152 1364
rect 7228 1344 7248 1364
rect 7350 1344 7370 1364
rect 9143 1420 9163 1440
rect 9265 1420 9285 1440
rect 9361 1420 9381 1440
rect 9471 1420 9491 1440
rect 9567 1420 9587 1440
rect 20730 1571 20750 1591
rect 20826 1571 20846 1591
rect 20936 1571 20956 1591
rect 21032 1571 21052 1591
rect 21154 1571 21174 1591
rect 22938 1646 22958 1666
rect 21250 1571 21270 1591
rect 23034 1646 23054 1666
rect 23156 1646 23176 1666
rect 23252 1646 23272 1666
rect 23362 1646 23382 1666
rect 23458 1646 23478 1666
rect 13411 1433 13431 1453
rect 7446 1344 7466 1364
rect 5468 1224 5488 1244
rect 3360 1147 3380 1167
rect 3456 1147 3476 1167
rect 3566 1147 3586 1167
rect 3662 1147 3682 1167
rect 3784 1147 3804 1167
rect 5564 1224 5584 1244
rect 5686 1224 5706 1244
rect 5782 1224 5802 1244
rect 5892 1224 5912 1244
rect 5988 1224 6008 1244
rect 11303 1356 11323 1376
rect 11399 1356 11419 1376
rect 11509 1356 11529 1376
rect 11605 1356 11625 1376
rect 11727 1356 11747 1376
rect 13507 1433 13527 1453
rect 13629 1433 13649 1453
rect 13725 1433 13745 1453
rect 13835 1433 13855 1453
rect 13931 1433 13951 1453
rect 25094 1584 25114 1604
rect 25190 1584 25210 1604
rect 25300 1584 25320 1604
rect 25396 1584 25416 1604
rect 25518 1584 25538 1604
rect 27315 1658 27335 1678
rect 25614 1584 25634 1604
rect 27411 1658 27431 1678
rect 27533 1658 27553 1678
rect 27629 1658 27649 1678
rect 27739 1658 27759 1678
rect 27835 1658 27855 1678
rect 11823 1356 11843 1376
rect 9845 1236 9865 1256
rect 3880 1147 3900 1167
rect 7724 1160 7744 1180
rect 7820 1160 7840 1180
rect 7930 1160 7950 1180
rect 8026 1160 8046 1180
rect 8148 1160 8168 1180
rect 9941 1236 9961 1256
rect 10063 1236 10083 1256
rect 10159 1236 10179 1256
rect 10269 1236 10289 1256
rect 10365 1236 10385 1256
rect 15667 1369 15687 1389
rect 15763 1369 15783 1389
rect 15873 1369 15893 1389
rect 15969 1369 15989 1389
rect 16091 1369 16111 1389
rect 17677 1407 17697 1427
rect 16187 1369 16207 1389
rect 17773 1407 17793 1427
rect 17895 1407 17915 1427
rect 17991 1407 18011 1427
rect 18101 1407 18121 1427
rect 18197 1407 18217 1427
rect 29471 1596 29491 1616
rect 29567 1596 29587 1616
rect 29677 1596 29697 1616
rect 29773 1596 29793 1616
rect 29895 1596 29915 1616
rect 31679 1671 31699 1691
rect 29991 1596 30011 1616
rect 31775 1671 31795 1691
rect 31897 1671 31917 1691
rect 31993 1671 32013 1691
rect 32103 1671 32123 1691
rect 32199 1671 32219 1691
rect 22041 1420 22061 1440
rect 14209 1249 14229 1269
rect 8244 1160 8264 1180
rect 12101 1172 12121 1192
rect 12197 1172 12217 1192
rect 12307 1172 12327 1192
rect 12403 1172 12423 1192
rect 12525 1172 12545 1192
rect 14305 1249 14325 1269
rect 14427 1249 14447 1269
rect 14523 1249 14543 1269
rect 14633 1249 14653 1269
rect 14729 1249 14749 1269
rect 19933 1343 19953 1363
rect 20029 1343 20049 1363
rect 20139 1343 20159 1363
rect 20235 1343 20255 1363
rect 20357 1343 20377 1363
rect 22137 1420 22157 1440
rect 22259 1420 22279 1440
rect 22355 1420 22375 1440
rect 22465 1420 22485 1440
rect 22561 1420 22581 1440
rect 33835 1609 33855 1629
rect 33931 1609 33951 1629
rect 34041 1609 34061 1629
rect 34137 1609 34157 1629
rect 34259 1609 34279 1629
rect 34355 1609 34375 1629
rect 26418 1432 26438 1452
rect 20453 1343 20473 1363
rect 12621 1172 12641 1192
rect 16465 1185 16485 1205
rect 16561 1185 16581 1205
rect 16671 1185 16691 1205
rect 16767 1185 16787 1205
rect 16889 1185 16909 1205
rect 18475 1223 18495 1243
rect 16985 1185 17005 1205
rect 18571 1223 18591 1243
rect 18693 1223 18713 1243
rect 18789 1223 18809 1243
rect 18899 1223 18919 1243
rect 18995 1223 19015 1243
rect 24297 1356 24317 1376
rect 24393 1356 24413 1376
rect 24503 1356 24523 1376
rect 24599 1356 24619 1376
rect 24721 1356 24741 1376
rect 26514 1432 26534 1452
rect 26636 1432 26656 1452
rect 26732 1432 26752 1452
rect 26842 1432 26862 1452
rect 26938 1432 26958 1452
rect 30782 1445 30802 1465
rect 24817 1356 24837 1376
rect 22839 1236 22859 1256
rect 307 983 327 1003
rect 403 983 423 1003
rect 525 983 545 1003
rect 621 983 641 1003
rect 731 983 751 1003
rect 827 983 847 1003
rect 4671 996 4691 1016
rect 4767 996 4787 1016
rect 4889 996 4909 1016
rect 4985 996 5005 1016
rect 5095 996 5115 1016
rect 5191 996 5211 1016
rect 9048 1008 9068 1028
rect 9144 1008 9164 1028
rect 9266 1008 9286 1028
rect 9362 1008 9382 1028
rect 9472 1008 9492 1028
rect 20731 1159 20751 1179
rect 20827 1159 20847 1179
rect 20937 1159 20957 1179
rect 21033 1159 21053 1179
rect 21155 1159 21175 1179
rect 22935 1236 22955 1256
rect 23057 1236 23077 1256
rect 23153 1236 23173 1256
rect 23263 1236 23283 1256
rect 23359 1236 23379 1256
rect 28674 1368 28694 1388
rect 28770 1368 28790 1388
rect 28880 1368 28900 1388
rect 28976 1368 28996 1388
rect 29098 1368 29118 1388
rect 30878 1445 30898 1465
rect 31000 1445 31020 1465
rect 31096 1445 31116 1465
rect 31206 1445 31226 1465
rect 31302 1445 31322 1465
rect 29194 1368 29214 1388
rect 27216 1248 27236 1268
rect 21251 1159 21271 1179
rect 25095 1172 25115 1192
rect 25191 1172 25211 1192
rect 25301 1172 25321 1192
rect 25397 1172 25417 1192
rect 25519 1172 25539 1192
rect 27312 1248 27332 1268
rect 27434 1248 27454 1268
rect 27530 1248 27550 1268
rect 27640 1248 27660 1268
rect 27736 1248 27756 1268
rect 33038 1381 33058 1401
rect 33134 1381 33154 1401
rect 33244 1381 33264 1401
rect 33340 1381 33360 1401
rect 33462 1381 33482 1401
rect 33558 1381 33578 1401
rect 31580 1261 31600 1281
rect 25615 1172 25635 1192
rect 29472 1184 29492 1204
rect 29568 1184 29588 1204
rect 29678 1184 29698 1204
rect 29774 1184 29794 1204
rect 29896 1184 29916 1204
rect 31676 1261 31696 1281
rect 31798 1261 31818 1281
rect 31894 1261 31914 1281
rect 32004 1261 32024 1281
rect 32100 1261 32120 1281
rect 29992 1184 30012 1204
rect 33836 1197 33856 1217
rect 33932 1197 33952 1217
rect 34042 1197 34062 1217
rect 34138 1197 34158 1217
rect 34260 1197 34280 1217
rect 34356 1197 34376 1217
rect 9568 1008 9588 1028
rect 13412 1021 13432 1041
rect 13508 1021 13528 1041
rect 13630 1021 13650 1041
rect 13726 1021 13746 1041
rect 13836 1021 13856 1041
rect 13932 1021 13952 1041
rect 17678 995 17698 1015
rect 17774 995 17794 1015
rect 17896 995 17916 1015
rect 17992 995 18012 1015
rect 18102 995 18122 1015
rect 18198 995 18218 1015
rect 22042 1008 22062 1028
rect 22138 1008 22158 1028
rect 22260 1008 22280 1028
rect 22356 1008 22376 1028
rect 22466 1008 22486 1028
rect 22562 1008 22582 1028
rect 26419 1020 26439 1040
rect 26515 1020 26535 1040
rect 26637 1020 26657 1040
rect 26733 1020 26753 1040
rect 26843 1020 26863 1040
rect 26939 1020 26959 1040
rect 30783 1033 30803 1053
rect 30879 1033 30899 1053
rect 31001 1033 31021 1053
rect 31097 1033 31117 1053
rect 31207 1033 31227 1053
rect 31303 1033 31323 1053
rect 1520 407 1540 427
rect 1616 407 1636 427
rect 1738 407 1758 427
rect 1834 407 1854 427
rect 1944 407 1964 427
rect 2040 407 2060 427
rect 5884 420 5904 440
rect 4009 333 4029 353
rect 4105 333 4125 353
rect 4227 333 4247 353
rect 4323 333 4343 353
rect 4433 333 4453 353
rect 5980 420 6000 440
rect 6102 420 6122 440
rect 6198 420 6218 440
rect 6308 420 6328 440
rect 6404 420 6424 440
rect 10261 432 10281 452
rect 4529 333 4549 353
rect 8457 357 8477 377
rect 8553 357 8573 377
rect 8675 357 8695 377
rect 8771 357 8791 377
rect 8881 357 8901 377
rect 10357 432 10377 452
rect 10479 432 10499 452
rect 10575 432 10595 452
rect 10685 432 10705 452
rect 10781 432 10801 452
rect 14625 445 14645 465
rect 8977 357 8997 377
rect 12750 358 12770 378
rect 12846 358 12866 378
rect 12968 358 12988 378
rect 13064 358 13084 378
rect 13174 358 13194 378
rect 14721 445 14741 465
rect 14843 445 14863 465
rect 14939 445 14959 465
rect 15049 445 15069 465
rect 15145 445 15165 465
rect 18891 419 18911 439
rect 13270 358 13290 378
rect 18987 419 19007 439
rect 19109 419 19129 439
rect 19205 419 19225 439
rect 19315 419 19335 439
rect 19411 419 19431 439
rect 23255 432 23275 452
rect 16947 294 16967 314
rect 17043 294 17063 314
rect 17165 294 17185 314
rect 17261 294 17281 314
rect 17371 294 17391 314
rect 17467 294 17487 314
rect 21380 345 21400 365
rect 21476 345 21496 365
rect 21598 345 21618 365
rect 21694 345 21714 365
rect 21804 345 21824 365
rect 23351 432 23371 452
rect 23473 432 23493 452
rect 23569 432 23589 452
rect 23679 432 23699 452
rect 23775 432 23795 452
rect 27632 444 27652 464
rect 21900 345 21920 365
rect 25828 369 25848 389
rect 25924 369 25944 389
rect 26046 369 26066 389
rect 26142 369 26162 389
rect 26252 369 26272 389
rect 27728 444 27748 464
rect 27850 444 27870 464
rect 27946 444 27966 464
rect 28056 444 28076 464
rect 28152 444 28172 464
rect 31996 457 32016 477
rect 26348 369 26368 389
rect 30121 370 30141 390
rect 30217 370 30237 390
rect 30339 370 30359 390
rect 30435 370 30455 390
rect 30545 370 30565 390
rect 32092 457 32112 477
rect 32214 457 32234 477
rect 32310 457 32330 477
rect 32420 457 32440 477
rect 32516 457 32536 477
rect 30641 370 30661 390
<< poly >>
rect 3518 8866 3568 8882
rect 3726 8866 3776 8882
rect 3944 8866 3994 8882
rect 7882 8879 7932 8895
rect 8090 8879 8140 8895
rect 8308 8879 8358 8895
rect 12259 8891 12309 8907
rect 12467 8891 12517 8907
rect 12685 8891 12735 8907
rect 16623 8904 16673 8920
rect 16831 8904 16881 8920
rect 17049 8904 17099 8920
rect 3518 8794 3568 8824
rect 3518 8774 3525 8794
rect 3545 8774 3568 8794
rect 3518 8747 3568 8774
rect 3726 8792 3776 8824
rect 3726 8772 3743 8792
rect 3763 8772 3776 8792
rect 3726 8747 3776 8772
rect 3944 8795 3994 8824
rect 3944 8775 3961 8795
rect 3981 8775 3994 8795
rect 3944 8747 3994 8775
rect 7882 8807 7932 8837
rect 7882 8787 7889 8807
rect 7909 8787 7932 8807
rect 2721 8638 2771 8654
rect 2929 8638 2979 8654
rect 3147 8638 3197 8654
rect 7882 8760 7932 8787
rect 8090 8805 8140 8837
rect 8090 8785 8107 8805
rect 8127 8785 8140 8805
rect 8090 8760 8140 8785
rect 8308 8808 8358 8837
rect 8308 8788 8325 8808
rect 8345 8788 8358 8808
rect 8308 8760 8358 8788
rect 12259 8819 12309 8849
rect 12259 8799 12266 8819
rect 12286 8799 12309 8819
rect 3518 8634 3568 8647
rect 3726 8634 3776 8647
rect 3944 8634 3994 8647
rect 7085 8651 7135 8667
rect 7293 8651 7343 8667
rect 7511 8651 7561 8667
rect 12259 8772 12309 8799
rect 12467 8817 12517 8849
rect 12467 8797 12484 8817
rect 12504 8797 12517 8817
rect 12467 8772 12517 8797
rect 12685 8820 12735 8849
rect 12685 8800 12702 8820
rect 12722 8800 12735 8820
rect 12685 8772 12735 8800
rect 16623 8832 16673 8862
rect 16623 8812 16630 8832
rect 16650 8812 16673 8832
rect 7882 8647 7932 8660
rect 8090 8647 8140 8660
rect 8308 8647 8358 8660
rect 11462 8663 11512 8679
rect 11670 8663 11720 8679
rect 11888 8663 11938 8679
rect 16623 8785 16673 8812
rect 16831 8830 16881 8862
rect 16831 8810 16848 8830
rect 16868 8810 16881 8830
rect 16831 8785 16881 8810
rect 17049 8833 17099 8862
rect 20889 8878 20939 8894
rect 21097 8878 21147 8894
rect 21315 8878 21365 8894
rect 25253 8891 25303 8907
rect 25461 8891 25511 8907
rect 25679 8891 25729 8907
rect 29630 8903 29680 8919
rect 29838 8903 29888 8919
rect 30056 8903 30106 8919
rect 33994 8916 34044 8932
rect 34202 8916 34252 8932
rect 34420 8916 34470 8932
rect 17049 8813 17066 8833
rect 17086 8813 17099 8833
rect 17049 8785 17099 8813
rect 12259 8659 12309 8672
rect 12467 8659 12517 8672
rect 12685 8659 12735 8672
rect 15826 8676 15876 8692
rect 16034 8676 16084 8692
rect 16252 8676 16302 8692
rect 20889 8806 20939 8836
rect 20889 8786 20896 8806
rect 20916 8786 20939 8806
rect 20889 8759 20939 8786
rect 21097 8804 21147 8836
rect 21097 8784 21114 8804
rect 21134 8784 21147 8804
rect 21097 8759 21147 8784
rect 21315 8807 21365 8836
rect 21315 8787 21332 8807
rect 21352 8787 21365 8807
rect 21315 8759 21365 8787
rect 25253 8819 25303 8849
rect 25253 8799 25260 8819
rect 25280 8799 25303 8819
rect 16623 8672 16673 8685
rect 16831 8672 16881 8685
rect 17049 8672 17099 8685
rect 20092 8650 20142 8666
rect 20300 8650 20350 8666
rect 20518 8650 20568 8666
rect 25253 8772 25303 8799
rect 25461 8817 25511 8849
rect 25461 8797 25478 8817
rect 25498 8797 25511 8817
rect 25461 8772 25511 8797
rect 25679 8820 25729 8849
rect 25679 8800 25696 8820
rect 25716 8800 25729 8820
rect 25679 8772 25729 8800
rect 29630 8831 29680 8861
rect 29630 8811 29637 8831
rect 29657 8811 29680 8831
rect 465 8579 515 8592
rect 683 8579 733 8592
rect 891 8579 941 8592
rect 2721 8566 2771 8596
rect 2721 8546 2728 8566
rect 2748 8546 2771 8566
rect 2721 8519 2771 8546
rect 2929 8564 2979 8596
rect 2929 8544 2946 8564
rect 2966 8544 2979 8564
rect 2929 8519 2979 8544
rect 3147 8567 3197 8596
rect 3147 8547 3164 8567
rect 3184 8547 3197 8567
rect 4829 8592 4879 8605
rect 5047 8592 5097 8605
rect 5255 8592 5305 8605
rect 3147 8519 3197 8547
rect 465 8451 515 8479
rect 465 8431 478 8451
rect 498 8431 515 8451
rect 465 8402 515 8431
rect 683 8454 733 8479
rect 683 8434 696 8454
rect 716 8434 733 8454
rect 683 8402 733 8434
rect 891 8452 941 8479
rect 891 8432 914 8452
rect 934 8432 941 8452
rect 891 8402 941 8432
rect 7085 8579 7135 8609
rect 7085 8559 7092 8579
rect 7112 8559 7135 8579
rect 7085 8532 7135 8559
rect 7293 8577 7343 8609
rect 7293 8557 7310 8577
rect 7330 8557 7343 8577
rect 7293 8532 7343 8557
rect 7511 8580 7561 8609
rect 7511 8560 7528 8580
rect 7548 8560 7561 8580
rect 9206 8604 9256 8617
rect 9424 8604 9474 8617
rect 9632 8604 9682 8617
rect 7511 8532 7561 8560
rect 3519 8454 3569 8470
rect 3727 8454 3777 8470
rect 3945 8454 3995 8470
rect 1263 8395 1313 8408
rect 1481 8395 1531 8408
rect 1689 8395 1739 8408
rect 2721 8406 2771 8419
rect 2929 8406 2979 8419
rect 3147 8406 3197 8419
rect 4829 8464 4879 8492
rect 465 8344 515 8360
rect 683 8344 733 8360
rect 891 8344 941 8360
rect 3519 8382 3569 8412
rect 3519 8362 3526 8382
rect 3546 8362 3569 8382
rect 3519 8335 3569 8362
rect 3727 8380 3777 8412
rect 3727 8360 3744 8380
rect 3764 8360 3777 8380
rect 3727 8335 3777 8360
rect 3945 8383 3995 8412
rect 3945 8363 3962 8383
rect 3982 8363 3995 8383
rect 4829 8444 4842 8464
rect 4862 8444 4879 8464
rect 4829 8415 4879 8444
rect 5047 8467 5097 8492
rect 5047 8447 5060 8467
rect 5080 8447 5097 8467
rect 5047 8415 5097 8447
rect 5255 8465 5305 8492
rect 5255 8445 5278 8465
rect 5298 8445 5305 8465
rect 5255 8415 5305 8445
rect 11462 8591 11512 8621
rect 11462 8571 11469 8591
rect 11489 8571 11512 8591
rect 11462 8544 11512 8571
rect 11670 8589 11720 8621
rect 11670 8569 11687 8589
rect 11707 8569 11720 8589
rect 11670 8544 11720 8569
rect 11888 8592 11938 8621
rect 11888 8572 11905 8592
rect 11925 8572 11938 8592
rect 13570 8617 13620 8630
rect 13788 8617 13838 8630
rect 13996 8617 14046 8630
rect 11888 8544 11938 8572
rect 7883 8467 7933 8483
rect 8091 8467 8141 8483
rect 8309 8467 8359 8483
rect 3945 8335 3995 8363
rect 5627 8408 5677 8421
rect 5845 8408 5895 8421
rect 6053 8408 6103 8421
rect 7085 8419 7135 8432
rect 7293 8419 7343 8432
rect 7511 8419 7561 8432
rect 9206 8476 9256 8504
rect 4829 8357 4879 8373
rect 5047 8357 5097 8373
rect 5255 8357 5305 8373
rect 1263 8267 1313 8295
rect 1263 8247 1276 8267
rect 1296 8247 1313 8267
rect 1263 8218 1313 8247
rect 1481 8270 1531 8295
rect 1481 8250 1494 8270
rect 1514 8250 1531 8270
rect 1481 8218 1531 8250
rect 1689 8268 1739 8295
rect 1689 8248 1712 8268
rect 1732 8248 1739 8268
rect 1689 8218 1739 8248
rect 2622 8228 2672 8244
rect 2830 8228 2880 8244
rect 3048 8228 3098 8244
rect 7883 8395 7933 8425
rect 7883 8375 7890 8395
rect 7910 8375 7933 8395
rect 7883 8348 7933 8375
rect 8091 8393 8141 8425
rect 8091 8373 8108 8393
rect 8128 8373 8141 8393
rect 8091 8348 8141 8373
rect 8309 8396 8359 8425
rect 8309 8376 8326 8396
rect 8346 8376 8359 8396
rect 9206 8456 9219 8476
rect 9239 8456 9256 8476
rect 9206 8427 9256 8456
rect 9424 8479 9474 8504
rect 9424 8459 9437 8479
rect 9457 8459 9474 8479
rect 9424 8427 9474 8459
rect 9632 8477 9682 8504
rect 9632 8457 9655 8477
rect 9675 8457 9682 8477
rect 9632 8427 9682 8457
rect 15826 8604 15876 8634
rect 15826 8584 15833 8604
rect 15853 8584 15876 8604
rect 15826 8557 15876 8584
rect 16034 8602 16084 8634
rect 16034 8582 16051 8602
rect 16071 8582 16084 8602
rect 16034 8557 16084 8582
rect 16252 8605 16302 8634
rect 16252 8585 16269 8605
rect 16289 8585 16302 8605
rect 20889 8646 20939 8659
rect 21097 8646 21147 8659
rect 21315 8646 21365 8659
rect 24456 8663 24506 8679
rect 24664 8663 24714 8679
rect 24882 8663 24932 8679
rect 29630 8784 29680 8811
rect 29838 8829 29888 8861
rect 29838 8809 29855 8829
rect 29875 8809 29888 8829
rect 29838 8784 29888 8809
rect 30056 8832 30106 8861
rect 30056 8812 30073 8832
rect 30093 8812 30106 8832
rect 30056 8784 30106 8812
rect 33994 8844 34044 8874
rect 33994 8824 34001 8844
rect 34021 8824 34044 8844
rect 25253 8659 25303 8672
rect 25461 8659 25511 8672
rect 25679 8659 25729 8672
rect 28833 8675 28883 8691
rect 29041 8675 29091 8691
rect 29259 8675 29309 8691
rect 33994 8797 34044 8824
rect 34202 8842 34252 8874
rect 34202 8822 34219 8842
rect 34239 8822 34252 8842
rect 34202 8797 34252 8822
rect 34420 8845 34470 8874
rect 34420 8825 34437 8845
rect 34457 8825 34470 8845
rect 34420 8797 34470 8825
rect 29630 8671 29680 8684
rect 29838 8671 29888 8684
rect 30056 8671 30106 8684
rect 33197 8688 33247 8704
rect 33405 8688 33455 8704
rect 33623 8688 33673 8704
rect 33994 8684 34044 8697
rect 34202 8684 34252 8697
rect 34420 8684 34470 8697
rect 16252 8557 16302 8585
rect 17836 8591 17886 8604
rect 18054 8591 18104 8604
rect 18262 8591 18312 8604
rect 12260 8479 12310 8495
rect 12468 8479 12518 8495
rect 12686 8479 12736 8495
rect 8309 8348 8359 8376
rect 10004 8420 10054 8433
rect 10222 8420 10272 8433
rect 10430 8420 10480 8433
rect 11462 8431 11512 8444
rect 11670 8431 11720 8444
rect 11888 8431 11938 8444
rect 13570 8489 13620 8517
rect 9206 8369 9256 8385
rect 9424 8369 9474 8385
rect 9632 8369 9682 8385
rect 5627 8280 5677 8308
rect 466 8167 516 8180
rect 684 8167 734 8180
rect 892 8167 942 8180
rect 3519 8222 3569 8235
rect 3727 8222 3777 8235
rect 3945 8222 3995 8235
rect 5627 8260 5640 8280
rect 5660 8260 5677 8280
rect 5627 8231 5677 8260
rect 5845 8283 5895 8308
rect 5845 8263 5858 8283
rect 5878 8263 5895 8283
rect 5845 8231 5895 8263
rect 6053 8281 6103 8308
rect 6053 8261 6076 8281
rect 6096 8261 6103 8281
rect 6053 8231 6103 8261
rect 6986 8241 7036 8257
rect 7194 8241 7244 8257
rect 7412 8241 7462 8257
rect 12260 8407 12310 8437
rect 12260 8387 12267 8407
rect 12287 8387 12310 8407
rect 12260 8360 12310 8387
rect 12468 8405 12518 8437
rect 12468 8385 12485 8405
rect 12505 8385 12518 8405
rect 12468 8360 12518 8385
rect 12686 8408 12736 8437
rect 12686 8388 12703 8408
rect 12723 8388 12736 8408
rect 13570 8469 13583 8489
rect 13603 8469 13620 8489
rect 13570 8440 13620 8469
rect 13788 8492 13838 8517
rect 13788 8472 13801 8492
rect 13821 8472 13838 8492
rect 13788 8440 13838 8472
rect 13996 8490 14046 8517
rect 13996 8470 14019 8490
rect 14039 8470 14046 8490
rect 13996 8440 14046 8470
rect 16624 8492 16674 8508
rect 16832 8492 16882 8508
rect 17050 8492 17100 8508
rect 12686 8360 12736 8388
rect 14368 8433 14418 8446
rect 14586 8433 14636 8446
rect 14794 8433 14844 8446
rect 15826 8444 15876 8457
rect 16034 8444 16084 8457
rect 16252 8444 16302 8457
rect 20092 8578 20142 8608
rect 20092 8558 20099 8578
rect 20119 8558 20142 8578
rect 20092 8531 20142 8558
rect 20300 8576 20350 8608
rect 20300 8556 20317 8576
rect 20337 8556 20350 8576
rect 20300 8531 20350 8556
rect 20518 8579 20568 8608
rect 20518 8559 20535 8579
rect 20555 8559 20568 8579
rect 22200 8604 22250 8617
rect 22418 8604 22468 8617
rect 22626 8604 22676 8617
rect 20518 8531 20568 8559
rect 13570 8382 13620 8398
rect 13788 8382 13838 8398
rect 13996 8382 14046 8398
rect 10004 8292 10054 8320
rect 1263 8160 1313 8176
rect 1481 8160 1531 8176
rect 1689 8160 1739 8176
rect 2622 8156 2672 8186
rect 2622 8136 2629 8156
rect 2649 8136 2672 8156
rect 2622 8109 2672 8136
rect 2830 8154 2880 8186
rect 2830 8134 2847 8154
rect 2867 8134 2880 8154
rect 2830 8109 2880 8134
rect 3048 8157 3098 8186
rect 4830 8180 4880 8193
rect 5048 8180 5098 8193
rect 5256 8180 5306 8193
rect 7883 8235 7933 8248
rect 8091 8235 8141 8248
rect 8309 8235 8359 8248
rect 10004 8272 10017 8292
rect 10037 8272 10054 8292
rect 10004 8243 10054 8272
rect 10222 8295 10272 8320
rect 10222 8275 10235 8295
rect 10255 8275 10272 8295
rect 10222 8243 10272 8275
rect 10430 8293 10480 8320
rect 10430 8273 10453 8293
rect 10473 8273 10480 8293
rect 10430 8243 10480 8273
rect 11363 8253 11413 8269
rect 11571 8253 11621 8269
rect 11789 8253 11839 8269
rect 16624 8420 16674 8450
rect 16624 8400 16631 8420
rect 16651 8400 16674 8420
rect 16624 8373 16674 8400
rect 16832 8418 16882 8450
rect 16832 8398 16849 8418
rect 16869 8398 16882 8418
rect 16832 8373 16882 8398
rect 17050 8421 17100 8450
rect 17050 8401 17067 8421
rect 17087 8401 17100 8421
rect 17836 8463 17886 8491
rect 17050 8373 17100 8401
rect 17836 8443 17849 8463
rect 17869 8443 17886 8463
rect 17836 8414 17886 8443
rect 18054 8466 18104 8491
rect 18054 8446 18067 8466
rect 18087 8446 18104 8466
rect 18054 8414 18104 8446
rect 18262 8464 18312 8491
rect 18262 8444 18285 8464
rect 18305 8444 18312 8464
rect 18262 8414 18312 8444
rect 24456 8591 24506 8621
rect 24456 8571 24463 8591
rect 24483 8571 24506 8591
rect 24456 8544 24506 8571
rect 24664 8589 24714 8621
rect 24664 8569 24681 8589
rect 24701 8569 24714 8589
rect 24664 8544 24714 8569
rect 24882 8592 24932 8621
rect 24882 8572 24899 8592
rect 24919 8572 24932 8592
rect 26577 8616 26627 8629
rect 26795 8616 26845 8629
rect 27003 8616 27053 8629
rect 24882 8544 24932 8572
rect 20890 8466 20940 8482
rect 21098 8466 21148 8482
rect 21316 8466 21366 8482
rect 14368 8305 14418 8333
rect 3048 8137 3065 8157
rect 3085 8137 3098 8157
rect 3048 8109 3098 8137
rect 466 8039 516 8067
rect 466 8019 479 8039
rect 499 8019 516 8039
rect 466 7990 516 8019
rect 684 8042 734 8067
rect 684 8022 697 8042
rect 717 8022 734 8042
rect 684 7990 734 8022
rect 892 8040 942 8067
rect 892 8020 915 8040
rect 935 8020 942 8040
rect 892 7990 942 8020
rect 5627 8173 5677 8189
rect 5845 8173 5895 8189
rect 6053 8173 6103 8189
rect 6986 8169 7036 8199
rect 6986 8149 6993 8169
rect 7013 8149 7036 8169
rect 6986 8122 7036 8149
rect 7194 8167 7244 8199
rect 7194 8147 7211 8167
rect 7231 8147 7244 8167
rect 7194 8122 7244 8147
rect 7412 8170 7462 8199
rect 9207 8192 9257 8205
rect 9425 8192 9475 8205
rect 9633 8192 9683 8205
rect 12260 8247 12310 8260
rect 12468 8247 12518 8260
rect 12686 8247 12736 8260
rect 14368 8285 14381 8305
rect 14401 8285 14418 8305
rect 14368 8256 14418 8285
rect 14586 8308 14636 8333
rect 14586 8288 14599 8308
rect 14619 8288 14636 8308
rect 14586 8256 14636 8288
rect 14794 8306 14844 8333
rect 14794 8286 14817 8306
rect 14837 8286 14844 8306
rect 14794 8256 14844 8286
rect 15727 8266 15777 8282
rect 15935 8266 15985 8282
rect 16153 8266 16203 8282
rect 18634 8407 18684 8420
rect 18852 8407 18902 8420
rect 19060 8407 19110 8420
rect 20092 8418 20142 8431
rect 20300 8418 20350 8431
rect 20518 8418 20568 8431
rect 22200 8476 22250 8504
rect 17836 8356 17886 8372
rect 18054 8356 18104 8372
rect 18262 8356 18312 8372
rect 20890 8394 20940 8424
rect 20890 8374 20897 8394
rect 20917 8374 20940 8394
rect 20890 8347 20940 8374
rect 21098 8392 21148 8424
rect 21098 8372 21115 8392
rect 21135 8372 21148 8392
rect 21098 8347 21148 8372
rect 21316 8395 21366 8424
rect 21316 8375 21333 8395
rect 21353 8375 21366 8395
rect 22200 8456 22213 8476
rect 22233 8456 22250 8476
rect 22200 8427 22250 8456
rect 22418 8479 22468 8504
rect 22418 8459 22431 8479
rect 22451 8459 22468 8479
rect 22418 8427 22468 8459
rect 22626 8477 22676 8504
rect 22626 8457 22649 8477
rect 22669 8457 22676 8477
rect 22626 8427 22676 8457
rect 28833 8603 28883 8633
rect 28833 8583 28840 8603
rect 28860 8583 28883 8603
rect 28833 8556 28883 8583
rect 29041 8601 29091 8633
rect 29041 8581 29058 8601
rect 29078 8581 29091 8601
rect 29041 8556 29091 8581
rect 29259 8604 29309 8633
rect 29259 8584 29276 8604
rect 29296 8584 29309 8604
rect 30941 8629 30991 8642
rect 31159 8629 31209 8642
rect 31367 8629 31417 8642
rect 29259 8556 29309 8584
rect 25254 8479 25304 8495
rect 25462 8479 25512 8495
rect 25680 8479 25730 8495
rect 21316 8347 21366 8375
rect 22998 8420 23048 8433
rect 23216 8420 23266 8433
rect 23424 8420 23474 8433
rect 24456 8431 24506 8444
rect 24664 8431 24714 8444
rect 24882 8431 24932 8444
rect 26577 8488 26627 8516
rect 22200 8369 22250 8385
rect 22418 8369 22468 8385
rect 22626 8369 22676 8385
rect 7412 8150 7429 8170
rect 7449 8150 7462 8170
rect 7412 8122 7462 8150
rect 4830 8052 4880 8080
rect 2622 7996 2672 8009
rect 2830 7996 2880 8009
rect 3048 7996 3098 8009
rect 4830 8032 4843 8052
rect 4863 8032 4880 8052
rect 4830 8003 4880 8032
rect 5048 8055 5098 8080
rect 5048 8035 5061 8055
rect 5081 8035 5098 8055
rect 5048 8003 5098 8035
rect 5256 8053 5306 8080
rect 5256 8033 5279 8053
rect 5299 8033 5306 8053
rect 5256 8003 5306 8033
rect 10004 8185 10054 8201
rect 10222 8185 10272 8201
rect 10430 8185 10480 8201
rect 11363 8181 11413 8211
rect 11363 8161 11370 8181
rect 11390 8161 11413 8181
rect 11363 8134 11413 8161
rect 11571 8179 11621 8211
rect 11571 8159 11588 8179
rect 11608 8159 11621 8179
rect 11571 8134 11621 8159
rect 11789 8182 11839 8211
rect 13571 8205 13621 8218
rect 13789 8205 13839 8218
rect 13997 8205 14047 8218
rect 16624 8260 16674 8273
rect 16832 8260 16882 8273
rect 17050 8260 17100 8273
rect 18634 8279 18684 8307
rect 18634 8259 18647 8279
rect 18667 8259 18684 8279
rect 18634 8230 18684 8259
rect 18852 8282 18902 8307
rect 18852 8262 18865 8282
rect 18885 8262 18902 8282
rect 18852 8230 18902 8262
rect 19060 8280 19110 8307
rect 19060 8260 19083 8280
rect 19103 8260 19110 8280
rect 19060 8230 19110 8260
rect 19993 8240 20043 8256
rect 20201 8240 20251 8256
rect 20419 8240 20469 8256
rect 25254 8407 25304 8437
rect 25254 8387 25261 8407
rect 25281 8387 25304 8407
rect 25254 8360 25304 8387
rect 25462 8405 25512 8437
rect 25462 8385 25479 8405
rect 25499 8385 25512 8405
rect 25462 8360 25512 8385
rect 25680 8408 25730 8437
rect 25680 8388 25697 8408
rect 25717 8388 25730 8408
rect 26577 8468 26590 8488
rect 26610 8468 26627 8488
rect 26577 8439 26627 8468
rect 26795 8491 26845 8516
rect 26795 8471 26808 8491
rect 26828 8471 26845 8491
rect 26795 8439 26845 8471
rect 27003 8489 27053 8516
rect 27003 8469 27026 8489
rect 27046 8469 27053 8489
rect 27003 8439 27053 8469
rect 33197 8616 33247 8646
rect 33197 8596 33204 8616
rect 33224 8596 33247 8616
rect 33197 8569 33247 8596
rect 33405 8614 33455 8646
rect 33405 8594 33422 8614
rect 33442 8594 33455 8614
rect 33405 8569 33455 8594
rect 33623 8617 33673 8646
rect 33623 8597 33640 8617
rect 33660 8597 33673 8617
rect 33623 8569 33673 8597
rect 29631 8491 29681 8507
rect 29839 8491 29889 8507
rect 30057 8491 30107 8507
rect 25680 8360 25730 8388
rect 27375 8432 27425 8445
rect 27593 8432 27643 8445
rect 27801 8432 27851 8445
rect 28833 8443 28883 8456
rect 29041 8443 29091 8456
rect 29259 8443 29309 8456
rect 30941 8501 30991 8529
rect 26577 8381 26627 8397
rect 26795 8381 26845 8397
rect 27003 8381 27053 8397
rect 22998 8292 23048 8320
rect 11789 8162 11806 8182
rect 11826 8162 11839 8182
rect 11789 8134 11839 8162
rect 9207 8064 9257 8092
rect 6986 8009 7036 8022
rect 7194 8009 7244 8022
rect 7412 8009 7462 8022
rect 9207 8044 9220 8064
rect 9240 8044 9257 8064
rect 9207 8015 9257 8044
rect 9425 8067 9475 8092
rect 9425 8047 9438 8067
rect 9458 8047 9475 8067
rect 9425 8015 9475 8047
rect 9633 8065 9683 8092
rect 9633 8045 9656 8065
rect 9676 8045 9683 8065
rect 9633 8015 9683 8045
rect 14368 8198 14418 8214
rect 14586 8198 14636 8214
rect 14794 8198 14844 8214
rect 15727 8194 15777 8224
rect 15727 8174 15734 8194
rect 15754 8174 15777 8194
rect 15727 8147 15777 8174
rect 15935 8192 15985 8224
rect 15935 8172 15952 8192
rect 15972 8172 15985 8192
rect 15935 8147 15985 8172
rect 16153 8195 16203 8224
rect 16153 8175 16170 8195
rect 16190 8175 16203 8195
rect 16153 8147 16203 8175
rect 17837 8179 17887 8192
rect 18055 8179 18105 8192
rect 18263 8179 18313 8192
rect 20890 8234 20940 8247
rect 21098 8234 21148 8247
rect 21316 8234 21366 8247
rect 22998 8272 23011 8292
rect 23031 8272 23048 8292
rect 22998 8243 23048 8272
rect 23216 8295 23266 8320
rect 23216 8275 23229 8295
rect 23249 8275 23266 8295
rect 23216 8243 23266 8275
rect 23424 8293 23474 8320
rect 23424 8273 23447 8293
rect 23467 8273 23474 8293
rect 23424 8243 23474 8273
rect 24357 8253 24407 8269
rect 24565 8253 24615 8269
rect 24783 8253 24833 8269
rect 29631 8419 29681 8449
rect 29631 8399 29638 8419
rect 29658 8399 29681 8419
rect 29631 8372 29681 8399
rect 29839 8417 29889 8449
rect 29839 8397 29856 8417
rect 29876 8397 29889 8417
rect 29839 8372 29889 8397
rect 30057 8420 30107 8449
rect 30057 8400 30074 8420
rect 30094 8400 30107 8420
rect 30941 8481 30954 8501
rect 30974 8481 30991 8501
rect 30941 8452 30991 8481
rect 31159 8504 31209 8529
rect 31159 8484 31172 8504
rect 31192 8484 31209 8504
rect 31159 8452 31209 8484
rect 31367 8502 31417 8529
rect 31367 8482 31390 8502
rect 31410 8482 31417 8502
rect 31367 8452 31417 8482
rect 33995 8504 34045 8520
rect 34203 8504 34253 8520
rect 34421 8504 34471 8520
rect 30057 8372 30107 8400
rect 31739 8445 31789 8458
rect 31957 8445 32007 8458
rect 32165 8445 32215 8458
rect 33197 8456 33247 8469
rect 33405 8456 33455 8469
rect 33623 8456 33673 8469
rect 30941 8394 30991 8410
rect 31159 8394 31209 8410
rect 31367 8394 31417 8410
rect 27375 8304 27425 8332
rect 13571 8077 13621 8105
rect 11363 8021 11413 8034
rect 11571 8021 11621 8034
rect 11789 8021 11839 8034
rect 13571 8057 13584 8077
rect 13604 8057 13621 8077
rect 13571 8028 13621 8057
rect 13789 8080 13839 8105
rect 13789 8060 13802 8080
rect 13822 8060 13839 8080
rect 13789 8028 13839 8060
rect 13997 8078 14047 8105
rect 13997 8058 14020 8078
rect 14040 8058 14047 8078
rect 13997 8028 14047 8058
rect 18634 8172 18684 8188
rect 18852 8172 18902 8188
rect 19060 8172 19110 8188
rect 19993 8168 20043 8198
rect 19993 8148 20000 8168
rect 20020 8148 20043 8168
rect 19993 8121 20043 8148
rect 20201 8166 20251 8198
rect 20201 8146 20218 8166
rect 20238 8146 20251 8166
rect 20201 8121 20251 8146
rect 20419 8169 20469 8198
rect 22201 8192 22251 8205
rect 22419 8192 22469 8205
rect 22627 8192 22677 8205
rect 25254 8247 25304 8260
rect 25462 8247 25512 8260
rect 25680 8247 25730 8260
rect 27375 8284 27388 8304
rect 27408 8284 27425 8304
rect 27375 8255 27425 8284
rect 27593 8307 27643 8332
rect 27593 8287 27606 8307
rect 27626 8287 27643 8307
rect 27593 8255 27643 8287
rect 27801 8305 27851 8332
rect 27801 8285 27824 8305
rect 27844 8285 27851 8305
rect 27801 8255 27851 8285
rect 28734 8265 28784 8281
rect 28942 8265 28992 8281
rect 29160 8265 29210 8281
rect 33995 8432 34045 8462
rect 33995 8412 34002 8432
rect 34022 8412 34045 8432
rect 33995 8385 34045 8412
rect 34203 8430 34253 8462
rect 34203 8410 34220 8430
rect 34240 8410 34253 8430
rect 34203 8385 34253 8410
rect 34421 8433 34471 8462
rect 34421 8413 34438 8433
rect 34458 8413 34471 8433
rect 34421 8385 34471 8413
rect 31739 8317 31789 8345
rect 20419 8149 20436 8169
rect 20456 8149 20469 8169
rect 20419 8121 20469 8149
rect 15727 8034 15777 8047
rect 15935 8034 15985 8047
rect 16153 8034 16203 8047
rect 17837 8051 17887 8079
rect 17837 8031 17850 8051
rect 17870 8031 17887 8051
rect 466 7932 516 7948
rect 684 7932 734 7948
rect 892 7932 942 7948
rect 4830 7945 4880 7961
rect 5048 7945 5098 7961
rect 5256 7945 5306 7961
rect 9207 7957 9257 7973
rect 9425 7957 9475 7973
rect 9633 7957 9683 7973
rect 13571 7970 13621 7986
rect 13789 7970 13839 7986
rect 13997 7970 14047 7986
rect 17837 8002 17887 8031
rect 18055 8054 18105 8079
rect 18055 8034 18068 8054
rect 18088 8034 18105 8054
rect 18055 8002 18105 8034
rect 18263 8052 18313 8079
rect 18263 8032 18286 8052
rect 18306 8032 18313 8052
rect 18263 8002 18313 8032
rect 22998 8185 23048 8201
rect 23216 8185 23266 8201
rect 23424 8185 23474 8201
rect 24357 8181 24407 8211
rect 24357 8161 24364 8181
rect 24384 8161 24407 8181
rect 24357 8134 24407 8161
rect 24565 8179 24615 8211
rect 24565 8159 24582 8179
rect 24602 8159 24615 8179
rect 24565 8134 24615 8159
rect 24783 8182 24833 8211
rect 26578 8204 26628 8217
rect 26796 8204 26846 8217
rect 27004 8204 27054 8217
rect 29631 8259 29681 8272
rect 29839 8259 29889 8272
rect 30057 8259 30107 8272
rect 31739 8297 31752 8317
rect 31772 8297 31789 8317
rect 31739 8268 31789 8297
rect 31957 8320 32007 8345
rect 31957 8300 31970 8320
rect 31990 8300 32007 8320
rect 31957 8268 32007 8300
rect 32165 8318 32215 8345
rect 32165 8298 32188 8318
rect 32208 8298 32215 8318
rect 32165 8268 32215 8298
rect 33098 8278 33148 8294
rect 33306 8278 33356 8294
rect 33524 8278 33574 8294
rect 24783 8162 24800 8182
rect 24820 8162 24833 8182
rect 24783 8134 24833 8162
rect 22201 8064 22251 8092
rect 19993 8008 20043 8021
rect 20201 8008 20251 8021
rect 20419 8008 20469 8021
rect 22201 8044 22214 8064
rect 22234 8044 22251 8064
rect 22201 8015 22251 8044
rect 22419 8067 22469 8092
rect 22419 8047 22432 8067
rect 22452 8047 22469 8067
rect 22419 8015 22469 8047
rect 22627 8065 22677 8092
rect 22627 8045 22650 8065
rect 22670 8045 22677 8065
rect 22627 8015 22677 8045
rect 27375 8197 27425 8213
rect 27593 8197 27643 8213
rect 27801 8197 27851 8213
rect 28734 8193 28784 8223
rect 28734 8173 28741 8193
rect 28761 8173 28784 8193
rect 28734 8146 28784 8173
rect 28942 8191 28992 8223
rect 28942 8171 28959 8191
rect 28979 8171 28992 8191
rect 28942 8146 28992 8171
rect 29160 8194 29210 8223
rect 30942 8217 30992 8230
rect 31160 8217 31210 8230
rect 31368 8217 31418 8230
rect 33995 8272 34045 8285
rect 34203 8272 34253 8285
rect 34421 8272 34471 8285
rect 29160 8174 29177 8194
rect 29197 8174 29210 8194
rect 29160 8146 29210 8174
rect 26578 8076 26628 8104
rect 24357 8021 24407 8034
rect 24565 8021 24615 8034
rect 24783 8021 24833 8034
rect 26578 8056 26591 8076
rect 26611 8056 26628 8076
rect 26578 8027 26628 8056
rect 26796 8079 26846 8104
rect 26796 8059 26809 8079
rect 26829 8059 26846 8079
rect 26796 8027 26846 8059
rect 27004 8077 27054 8104
rect 27004 8057 27027 8077
rect 27047 8057 27054 8077
rect 27004 8027 27054 8057
rect 31739 8210 31789 8226
rect 31957 8210 32007 8226
rect 32165 8210 32215 8226
rect 33098 8206 33148 8236
rect 33098 8186 33105 8206
rect 33125 8186 33148 8206
rect 33098 8159 33148 8186
rect 33306 8204 33356 8236
rect 33306 8184 33323 8204
rect 33343 8184 33356 8204
rect 33306 8159 33356 8184
rect 33524 8207 33574 8236
rect 33524 8187 33541 8207
rect 33561 8187 33574 8207
rect 33524 8159 33574 8187
rect 30942 8089 30992 8117
rect 28734 8033 28784 8046
rect 28942 8033 28992 8046
rect 29160 8033 29210 8046
rect 30942 8069 30955 8089
rect 30975 8069 30992 8089
rect 30942 8040 30992 8069
rect 31160 8092 31210 8117
rect 31160 8072 31173 8092
rect 31193 8072 31210 8092
rect 31160 8040 31210 8072
rect 31368 8090 31418 8117
rect 31368 8070 31391 8090
rect 31411 8070 31418 8090
rect 31368 8040 31418 8070
rect 33098 8046 33148 8059
rect 33306 8046 33356 8059
rect 33524 8046 33574 8059
rect 17837 7944 17887 7960
rect 18055 7944 18105 7960
rect 18263 7944 18313 7960
rect 22201 7957 22251 7973
rect 22419 7957 22469 7973
rect 22627 7957 22677 7973
rect 26578 7969 26628 7985
rect 26796 7969 26846 7985
rect 27004 7969 27054 7985
rect 30942 7982 30992 7998
rect 31160 7982 31210 7998
rect 31368 7982 31418 7998
rect 3501 7848 3551 7864
rect 3709 7848 3759 7864
rect 3927 7848 3977 7864
rect 7865 7861 7915 7877
rect 8073 7861 8123 7877
rect 8291 7861 8341 7877
rect 12242 7873 12292 7889
rect 12450 7873 12500 7889
rect 12668 7873 12718 7889
rect 16606 7886 16656 7902
rect 16814 7886 16864 7902
rect 17032 7886 17082 7902
rect 1345 7787 1395 7800
rect 1563 7787 1613 7800
rect 1771 7787 1821 7800
rect 3501 7776 3551 7806
rect 3501 7756 3508 7776
rect 3528 7756 3551 7776
rect 3501 7729 3551 7756
rect 3709 7774 3759 7806
rect 3709 7754 3726 7774
rect 3746 7754 3759 7774
rect 3709 7729 3759 7754
rect 3927 7777 3977 7806
rect 3927 7757 3944 7777
rect 3964 7757 3977 7777
rect 5709 7800 5759 7813
rect 5927 7800 5977 7813
rect 6135 7800 6185 7813
rect 3927 7729 3977 7757
rect 1345 7659 1395 7687
rect 1345 7639 1358 7659
rect 1378 7639 1395 7659
rect 1345 7610 1395 7639
rect 1563 7662 1613 7687
rect 1563 7642 1576 7662
rect 1596 7642 1613 7662
rect 1563 7610 1613 7642
rect 1771 7660 1821 7687
rect 1771 7640 1794 7660
rect 1814 7640 1821 7660
rect 1771 7610 1821 7640
rect 2704 7620 2754 7636
rect 2912 7620 2962 7636
rect 3130 7620 3180 7636
rect 7865 7789 7915 7819
rect 7865 7769 7872 7789
rect 7892 7769 7915 7789
rect 7865 7742 7915 7769
rect 8073 7787 8123 7819
rect 8073 7767 8090 7787
rect 8110 7767 8123 7787
rect 8073 7742 8123 7767
rect 8291 7790 8341 7819
rect 8291 7770 8308 7790
rect 8328 7770 8341 7790
rect 10086 7812 10136 7825
rect 10304 7812 10354 7825
rect 10512 7812 10562 7825
rect 8291 7742 8341 7770
rect 5709 7672 5759 7700
rect 5709 7652 5722 7672
rect 5742 7652 5759 7672
rect 448 7561 498 7574
rect 666 7561 716 7574
rect 874 7561 924 7574
rect 3501 7616 3551 7629
rect 3709 7616 3759 7629
rect 3927 7616 3977 7629
rect 5709 7623 5759 7652
rect 5927 7675 5977 7700
rect 5927 7655 5940 7675
rect 5960 7655 5977 7675
rect 5927 7623 5977 7655
rect 6135 7673 6185 7700
rect 6135 7653 6158 7673
rect 6178 7653 6185 7673
rect 6135 7623 6185 7653
rect 7068 7633 7118 7649
rect 7276 7633 7326 7649
rect 7494 7633 7544 7649
rect 12242 7801 12292 7831
rect 12242 7781 12249 7801
rect 12269 7781 12292 7801
rect 12242 7754 12292 7781
rect 12450 7799 12500 7831
rect 12450 7779 12467 7799
rect 12487 7779 12500 7799
rect 12450 7754 12500 7779
rect 12668 7802 12718 7831
rect 12668 7782 12685 7802
rect 12705 7782 12718 7802
rect 14450 7825 14500 7838
rect 14668 7825 14718 7838
rect 14876 7825 14926 7838
rect 12668 7754 12718 7782
rect 10086 7684 10136 7712
rect 10086 7664 10099 7684
rect 10119 7664 10136 7684
rect 1345 7552 1395 7568
rect 1563 7552 1613 7568
rect 1771 7552 1821 7568
rect 2704 7548 2754 7578
rect 2704 7528 2711 7548
rect 2731 7528 2754 7548
rect 2704 7501 2754 7528
rect 2912 7546 2962 7578
rect 2912 7526 2929 7546
rect 2949 7526 2962 7546
rect 2912 7501 2962 7526
rect 3130 7549 3180 7578
rect 3130 7529 3147 7549
rect 3167 7529 3180 7549
rect 4812 7574 4862 7587
rect 5030 7574 5080 7587
rect 5238 7574 5288 7587
rect 7865 7629 7915 7642
rect 8073 7629 8123 7642
rect 8291 7629 8341 7642
rect 10086 7635 10136 7664
rect 10304 7687 10354 7712
rect 10304 7667 10317 7687
rect 10337 7667 10354 7687
rect 10304 7635 10354 7667
rect 10512 7685 10562 7712
rect 10512 7665 10535 7685
rect 10555 7665 10562 7685
rect 10512 7635 10562 7665
rect 11445 7645 11495 7661
rect 11653 7645 11703 7661
rect 11871 7645 11921 7661
rect 16606 7814 16656 7844
rect 16606 7794 16613 7814
rect 16633 7794 16656 7814
rect 16606 7767 16656 7794
rect 16814 7812 16864 7844
rect 16814 7792 16831 7812
rect 16851 7792 16864 7812
rect 16814 7767 16864 7792
rect 17032 7815 17082 7844
rect 20872 7860 20922 7876
rect 21080 7860 21130 7876
rect 21298 7860 21348 7876
rect 25236 7873 25286 7889
rect 25444 7873 25494 7889
rect 25662 7873 25712 7889
rect 29613 7885 29663 7901
rect 29821 7885 29871 7901
rect 30039 7885 30089 7901
rect 33977 7898 34027 7914
rect 34185 7898 34235 7914
rect 34403 7898 34453 7914
rect 17032 7795 17049 7815
rect 17069 7795 17082 7815
rect 17032 7767 17082 7795
rect 18716 7799 18766 7812
rect 18934 7799 18984 7812
rect 19142 7799 19192 7812
rect 14450 7697 14500 7725
rect 14450 7677 14463 7697
rect 14483 7677 14500 7697
rect 3130 7501 3180 7529
rect 448 7433 498 7461
rect 448 7413 461 7433
rect 481 7413 498 7433
rect 448 7384 498 7413
rect 666 7436 716 7461
rect 666 7416 679 7436
rect 699 7416 716 7436
rect 666 7384 716 7416
rect 874 7434 924 7461
rect 874 7414 897 7434
rect 917 7414 924 7434
rect 874 7384 924 7414
rect 5709 7565 5759 7581
rect 5927 7565 5977 7581
rect 6135 7565 6185 7581
rect 7068 7561 7118 7591
rect 7068 7541 7075 7561
rect 7095 7541 7118 7561
rect 7068 7514 7118 7541
rect 7276 7559 7326 7591
rect 7276 7539 7293 7559
rect 7313 7539 7326 7559
rect 7276 7514 7326 7539
rect 7494 7562 7544 7591
rect 7494 7542 7511 7562
rect 7531 7542 7544 7562
rect 9189 7586 9239 7599
rect 9407 7586 9457 7599
rect 9615 7586 9665 7599
rect 12242 7641 12292 7654
rect 12450 7641 12500 7654
rect 12668 7641 12718 7654
rect 14450 7648 14500 7677
rect 14668 7700 14718 7725
rect 14668 7680 14681 7700
rect 14701 7680 14718 7700
rect 14668 7648 14718 7680
rect 14876 7698 14926 7725
rect 14876 7678 14899 7698
rect 14919 7678 14926 7698
rect 14876 7648 14926 7678
rect 15809 7658 15859 7674
rect 16017 7658 16067 7674
rect 16235 7658 16285 7674
rect 20872 7788 20922 7818
rect 20872 7768 20879 7788
rect 20899 7768 20922 7788
rect 20872 7741 20922 7768
rect 21080 7786 21130 7818
rect 21080 7766 21097 7786
rect 21117 7766 21130 7786
rect 21080 7741 21130 7766
rect 21298 7789 21348 7818
rect 21298 7769 21315 7789
rect 21335 7769 21348 7789
rect 23080 7812 23130 7825
rect 23298 7812 23348 7825
rect 23506 7812 23556 7825
rect 21298 7741 21348 7769
rect 7494 7514 7544 7542
rect 3502 7436 3552 7452
rect 3710 7436 3760 7452
rect 3928 7436 3978 7452
rect 1246 7377 1296 7390
rect 1464 7377 1514 7390
rect 1672 7377 1722 7390
rect 2704 7388 2754 7401
rect 2912 7388 2962 7401
rect 3130 7388 3180 7401
rect 4812 7446 4862 7474
rect 448 7326 498 7342
rect 666 7326 716 7342
rect 874 7326 924 7342
rect 3502 7364 3552 7394
rect 3502 7344 3509 7364
rect 3529 7344 3552 7364
rect 3502 7317 3552 7344
rect 3710 7362 3760 7394
rect 3710 7342 3727 7362
rect 3747 7342 3760 7362
rect 3710 7317 3760 7342
rect 3928 7365 3978 7394
rect 3928 7345 3945 7365
rect 3965 7345 3978 7365
rect 4812 7426 4825 7446
rect 4845 7426 4862 7446
rect 4812 7397 4862 7426
rect 5030 7449 5080 7474
rect 5030 7429 5043 7449
rect 5063 7429 5080 7449
rect 5030 7397 5080 7429
rect 5238 7447 5288 7474
rect 5238 7427 5261 7447
rect 5281 7427 5288 7447
rect 5238 7397 5288 7427
rect 10086 7577 10136 7593
rect 10304 7577 10354 7593
rect 10512 7577 10562 7593
rect 11445 7573 11495 7603
rect 11445 7553 11452 7573
rect 11472 7553 11495 7573
rect 11445 7526 11495 7553
rect 11653 7571 11703 7603
rect 11653 7551 11670 7571
rect 11690 7551 11703 7571
rect 11653 7526 11703 7551
rect 11871 7574 11921 7603
rect 11871 7554 11888 7574
rect 11908 7554 11921 7574
rect 13553 7599 13603 7612
rect 13771 7599 13821 7612
rect 13979 7599 14029 7612
rect 16606 7654 16656 7667
rect 16814 7654 16864 7667
rect 17032 7654 17082 7667
rect 18716 7671 18766 7699
rect 18716 7651 18729 7671
rect 18749 7651 18766 7671
rect 18716 7622 18766 7651
rect 18934 7674 18984 7699
rect 18934 7654 18947 7674
rect 18967 7654 18984 7674
rect 18934 7622 18984 7654
rect 19142 7672 19192 7699
rect 19142 7652 19165 7672
rect 19185 7652 19192 7672
rect 19142 7622 19192 7652
rect 20075 7632 20125 7648
rect 20283 7632 20333 7648
rect 20501 7632 20551 7648
rect 25236 7801 25286 7831
rect 25236 7781 25243 7801
rect 25263 7781 25286 7801
rect 25236 7754 25286 7781
rect 25444 7799 25494 7831
rect 25444 7779 25461 7799
rect 25481 7779 25494 7799
rect 25444 7754 25494 7779
rect 25662 7802 25712 7831
rect 25662 7782 25679 7802
rect 25699 7782 25712 7802
rect 27457 7824 27507 7837
rect 27675 7824 27725 7837
rect 27883 7824 27933 7837
rect 25662 7754 25712 7782
rect 23080 7684 23130 7712
rect 23080 7664 23093 7684
rect 23113 7664 23130 7684
rect 11871 7526 11921 7554
rect 7866 7449 7916 7465
rect 8074 7449 8124 7465
rect 8292 7449 8342 7465
rect 3928 7317 3978 7345
rect 5610 7390 5660 7403
rect 5828 7390 5878 7403
rect 6036 7390 6086 7403
rect 7068 7401 7118 7414
rect 7276 7401 7326 7414
rect 7494 7401 7544 7414
rect 9189 7458 9239 7486
rect 4812 7339 4862 7355
rect 5030 7339 5080 7355
rect 5238 7339 5288 7355
rect 1246 7249 1296 7277
rect 1246 7229 1259 7249
rect 1279 7229 1296 7249
rect 1246 7200 1296 7229
rect 1464 7252 1514 7277
rect 1464 7232 1477 7252
rect 1497 7232 1514 7252
rect 1464 7200 1514 7232
rect 1672 7250 1722 7277
rect 1672 7230 1695 7250
rect 1715 7230 1722 7250
rect 1672 7200 1722 7230
rect 2539 7212 2589 7228
rect 2747 7212 2797 7228
rect 2965 7212 3015 7228
rect 7866 7377 7916 7407
rect 7866 7357 7873 7377
rect 7893 7357 7916 7377
rect 7866 7330 7916 7357
rect 8074 7375 8124 7407
rect 8074 7355 8091 7375
rect 8111 7355 8124 7375
rect 8074 7330 8124 7355
rect 8292 7378 8342 7407
rect 8292 7358 8309 7378
rect 8329 7358 8342 7378
rect 9189 7438 9202 7458
rect 9222 7438 9239 7458
rect 9189 7409 9239 7438
rect 9407 7461 9457 7486
rect 9407 7441 9420 7461
rect 9440 7441 9457 7461
rect 9407 7409 9457 7441
rect 9615 7459 9665 7486
rect 9615 7439 9638 7459
rect 9658 7439 9665 7459
rect 9615 7409 9665 7439
rect 14450 7590 14500 7606
rect 14668 7590 14718 7606
rect 14876 7590 14926 7606
rect 15809 7586 15859 7616
rect 15809 7566 15816 7586
rect 15836 7566 15859 7586
rect 15809 7539 15859 7566
rect 16017 7584 16067 7616
rect 16017 7564 16034 7584
rect 16054 7564 16067 7584
rect 16017 7539 16067 7564
rect 16235 7587 16285 7616
rect 16235 7567 16252 7587
rect 16272 7567 16285 7587
rect 16235 7539 16285 7567
rect 17819 7573 17869 7586
rect 18037 7573 18087 7586
rect 18245 7573 18295 7586
rect 20872 7628 20922 7641
rect 21080 7628 21130 7641
rect 21298 7628 21348 7641
rect 23080 7635 23130 7664
rect 23298 7687 23348 7712
rect 23298 7667 23311 7687
rect 23331 7667 23348 7687
rect 23298 7635 23348 7667
rect 23506 7685 23556 7712
rect 23506 7665 23529 7685
rect 23549 7665 23556 7685
rect 23506 7635 23556 7665
rect 24439 7645 24489 7661
rect 24647 7645 24697 7661
rect 24865 7645 24915 7661
rect 29613 7813 29663 7843
rect 29613 7793 29620 7813
rect 29640 7793 29663 7813
rect 29613 7766 29663 7793
rect 29821 7811 29871 7843
rect 29821 7791 29838 7811
rect 29858 7791 29871 7811
rect 29821 7766 29871 7791
rect 30039 7814 30089 7843
rect 30039 7794 30056 7814
rect 30076 7794 30089 7814
rect 31821 7837 31871 7850
rect 32039 7837 32089 7850
rect 32247 7837 32297 7850
rect 30039 7766 30089 7794
rect 27457 7696 27507 7724
rect 27457 7676 27470 7696
rect 27490 7676 27507 7696
rect 12243 7461 12293 7477
rect 12451 7461 12501 7477
rect 12669 7461 12719 7477
rect 8292 7330 8342 7358
rect 9987 7402 10037 7415
rect 10205 7402 10255 7415
rect 10413 7402 10463 7415
rect 11445 7413 11495 7426
rect 11653 7413 11703 7426
rect 11871 7413 11921 7426
rect 13553 7471 13603 7499
rect 9189 7351 9239 7367
rect 9407 7351 9457 7367
rect 9615 7351 9665 7367
rect 5610 7262 5660 7290
rect 449 7149 499 7162
rect 667 7149 717 7162
rect 875 7149 925 7162
rect 3502 7204 3552 7217
rect 3710 7204 3760 7217
rect 3928 7204 3978 7217
rect 5610 7242 5623 7262
rect 5643 7242 5660 7262
rect 5610 7213 5660 7242
rect 5828 7265 5878 7290
rect 5828 7245 5841 7265
rect 5861 7245 5878 7265
rect 5828 7213 5878 7245
rect 6036 7263 6086 7290
rect 6036 7243 6059 7263
rect 6079 7243 6086 7263
rect 6036 7213 6086 7243
rect 6903 7225 6953 7241
rect 7111 7225 7161 7241
rect 7329 7225 7379 7241
rect 12243 7389 12293 7419
rect 12243 7369 12250 7389
rect 12270 7369 12293 7389
rect 12243 7342 12293 7369
rect 12451 7387 12501 7419
rect 12451 7367 12468 7387
rect 12488 7367 12501 7387
rect 12451 7342 12501 7367
rect 12669 7390 12719 7419
rect 12669 7370 12686 7390
rect 12706 7370 12719 7390
rect 13553 7451 13566 7471
rect 13586 7451 13603 7471
rect 13553 7422 13603 7451
rect 13771 7474 13821 7499
rect 13771 7454 13784 7474
rect 13804 7454 13821 7474
rect 13771 7422 13821 7454
rect 13979 7472 14029 7499
rect 13979 7452 14002 7472
rect 14022 7452 14029 7472
rect 13979 7422 14029 7452
rect 16607 7474 16657 7490
rect 16815 7474 16865 7490
rect 17033 7474 17083 7490
rect 12669 7342 12719 7370
rect 14351 7415 14401 7428
rect 14569 7415 14619 7428
rect 14777 7415 14827 7428
rect 15809 7426 15859 7439
rect 16017 7426 16067 7439
rect 16235 7426 16285 7439
rect 18716 7564 18766 7580
rect 18934 7564 18984 7580
rect 19142 7564 19192 7580
rect 20075 7560 20125 7590
rect 20075 7540 20082 7560
rect 20102 7540 20125 7560
rect 20075 7513 20125 7540
rect 20283 7558 20333 7590
rect 20283 7538 20300 7558
rect 20320 7538 20333 7558
rect 20283 7513 20333 7538
rect 20501 7561 20551 7590
rect 20501 7541 20518 7561
rect 20538 7541 20551 7561
rect 22183 7586 22233 7599
rect 22401 7586 22451 7599
rect 22609 7586 22659 7599
rect 25236 7641 25286 7654
rect 25444 7641 25494 7654
rect 25662 7641 25712 7654
rect 27457 7647 27507 7676
rect 27675 7699 27725 7724
rect 27675 7679 27688 7699
rect 27708 7679 27725 7699
rect 27675 7647 27725 7679
rect 27883 7697 27933 7724
rect 27883 7677 27906 7697
rect 27926 7677 27933 7697
rect 27883 7647 27933 7677
rect 28816 7657 28866 7673
rect 29024 7657 29074 7673
rect 29242 7657 29292 7673
rect 33977 7826 34027 7856
rect 33977 7806 33984 7826
rect 34004 7806 34027 7826
rect 33977 7779 34027 7806
rect 34185 7824 34235 7856
rect 34185 7804 34202 7824
rect 34222 7804 34235 7824
rect 34185 7779 34235 7804
rect 34403 7827 34453 7856
rect 34403 7807 34420 7827
rect 34440 7807 34453 7827
rect 34403 7779 34453 7807
rect 31821 7709 31871 7737
rect 31821 7689 31834 7709
rect 31854 7689 31871 7709
rect 20501 7513 20551 7541
rect 13553 7364 13603 7380
rect 13771 7364 13821 7380
rect 13979 7364 14029 7380
rect 9987 7274 10037 7302
rect 1246 7142 1296 7158
rect 1464 7142 1514 7158
rect 1672 7142 1722 7158
rect 2539 7140 2589 7170
rect 2539 7120 2546 7140
rect 2566 7120 2589 7140
rect 2539 7093 2589 7120
rect 2747 7138 2797 7170
rect 2747 7118 2764 7138
rect 2784 7118 2797 7138
rect 2747 7093 2797 7118
rect 2965 7141 3015 7170
rect 4813 7162 4863 7175
rect 5031 7162 5081 7175
rect 5239 7162 5289 7175
rect 7866 7217 7916 7230
rect 8074 7217 8124 7230
rect 8292 7217 8342 7230
rect 9987 7254 10000 7274
rect 10020 7254 10037 7274
rect 9987 7225 10037 7254
rect 10205 7277 10255 7302
rect 10205 7257 10218 7277
rect 10238 7257 10255 7277
rect 10205 7225 10255 7257
rect 10413 7275 10463 7302
rect 10413 7255 10436 7275
rect 10456 7255 10463 7275
rect 10413 7225 10463 7255
rect 11280 7237 11330 7253
rect 11488 7237 11538 7253
rect 11706 7237 11756 7253
rect 16607 7402 16657 7432
rect 16607 7382 16614 7402
rect 16634 7382 16657 7402
rect 16607 7355 16657 7382
rect 16815 7400 16865 7432
rect 16815 7380 16832 7400
rect 16852 7380 16865 7400
rect 16815 7355 16865 7380
rect 17033 7403 17083 7432
rect 17033 7383 17050 7403
rect 17070 7383 17083 7403
rect 17819 7445 17869 7473
rect 17033 7355 17083 7383
rect 17819 7425 17832 7445
rect 17852 7425 17869 7445
rect 17819 7396 17869 7425
rect 18037 7448 18087 7473
rect 18037 7428 18050 7448
rect 18070 7428 18087 7448
rect 18037 7396 18087 7428
rect 18245 7446 18295 7473
rect 18245 7426 18268 7446
rect 18288 7426 18295 7446
rect 18245 7396 18295 7426
rect 23080 7577 23130 7593
rect 23298 7577 23348 7593
rect 23506 7577 23556 7593
rect 24439 7573 24489 7603
rect 24439 7553 24446 7573
rect 24466 7553 24489 7573
rect 24439 7526 24489 7553
rect 24647 7571 24697 7603
rect 24647 7551 24664 7571
rect 24684 7551 24697 7571
rect 24647 7526 24697 7551
rect 24865 7574 24915 7603
rect 24865 7554 24882 7574
rect 24902 7554 24915 7574
rect 26560 7598 26610 7611
rect 26778 7598 26828 7611
rect 26986 7598 27036 7611
rect 29613 7653 29663 7666
rect 29821 7653 29871 7666
rect 30039 7653 30089 7666
rect 31821 7660 31871 7689
rect 32039 7712 32089 7737
rect 32039 7692 32052 7712
rect 32072 7692 32089 7712
rect 32039 7660 32089 7692
rect 32247 7710 32297 7737
rect 32247 7690 32270 7710
rect 32290 7690 32297 7710
rect 32247 7660 32297 7690
rect 33180 7670 33230 7686
rect 33388 7670 33438 7686
rect 33606 7670 33656 7686
rect 24865 7526 24915 7554
rect 20873 7448 20923 7464
rect 21081 7448 21131 7464
rect 21299 7448 21349 7464
rect 14351 7287 14401 7315
rect 2965 7121 2982 7141
rect 3002 7121 3015 7141
rect 2965 7093 3015 7121
rect 449 7021 499 7049
rect 449 7001 462 7021
rect 482 7001 499 7021
rect 449 6972 499 7001
rect 667 7024 717 7049
rect 667 7004 680 7024
rect 700 7004 717 7024
rect 667 6972 717 7004
rect 875 7022 925 7049
rect 875 7002 898 7022
rect 918 7002 925 7022
rect 875 6972 925 7002
rect 5610 7155 5660 7171
rect 5828 7155 5878 7171
rect 6036 7155 6086 7171
rect 6903 7153 6953 7183
rect 6903 7133 6910 7153
rect 6930 7133 6953 7153
rect 6903 7106 6953 7133
rect 7111 7151 7161 7183
rect 7111 7131 7128 7151
rect 7148 7131 7161 7151
rect 7111 7106 7161 7131
rect 7329 7154 7379 7183
rect 9190 7174 9240 7187
rect 9408 7174 9458 7187
rect 9616 7174 9666 7187
rect 12243 7229 12293 7242
rect 12451 7229 12501 7242
rect 12669 7229 12719 7242
rect 14351 7267 14364 7287
rect 14384 7267 14401 7287
rect 14351 7238 14401 7267
rect 14569 7290 14619 7315
rect 14569 7270 14582 7290
rect 14602 7270 14619 7290
rect 14569 7238 14619 7270
rect 14777 7288 14827 7315
rect 14777 7268 14800 7288
rect 14820 7268 14827 7288
rect 14777 7238 14827 7268
rect 15644 7250 15694 7266
rect 15852 7250 15902 7266
rect 16070 7250 16120 7266
rect 18617 7389 18667 7402
rect 18835 7389 18885 7402
rect 19043 7389 19093 7402
rect 20075 7400 20125 7413
rect 20283 7400 20333 7413
rect 20501 7400 20551 7413
rect 22183 7458 22233 7486
rect 17819 7338 17869 7354
rect 18037 7338 18087 7354
rect 18245 7338 18295 7354
rect 20873 7376 20923 7406
rect 20873 7356 20880 7376
rect 20900 7356 20923 7376
rect 20873 7329 20923 7356
rect 21081 7374 21131 7406
rect 21081 7354 21098 7374
rect 21118 7354 21131 7374
rect 21081 7329 21131 7354
rect 21299 7377 21349 7406
rect 21299 7357 21316 7377
rect 21336 7357 21349 7377
rect 22183 7438 22196 7458
rect 22216 7438 22233 7458
rect 22183 7409 22233 7438
rect 22401 7461 22451 7486
rect 22401 7441 22414 7461
rect 22434 7441 22451 7461
rect 22401 7409 22451 7441
rect 22609 7459 22659 7486
rect 22609 7439 22632 7459
rect 22652 7439 22659 7459
rect 22609 7409 22659 7439
rect 27457 7589 27507 7605
rect 27675 7589 27725 7605
rect 27883 7589 27933 7605
rect 28816 7585 28866 7615
rect 28816 7565 28823 7585
rect 28843 7565 28866 7585
rect 28816 7538 28866 7565
rect 29024 7583 29074 7615
rect 29024 7563 29041 7583
rect 29061 7563 29074 7583
rect 29024 7538 29074 7563
rect 29242 7586 29292 7615
rect 29242 7566 29259 7586
rect 29279 7566 29292 7586
rect 30924 7611 30974 7624
rect 31142 7611 31192 7624
rect 31350 7611 31400 7624
rect 33977 7666 34027 7679
rect 34185 7666 34235 7679
rect 34403 7666 34453 7679
rect 29242 7538 29292 7566
rect 25237 7461 25287 7477
rect 25445 7461 25495 7477
rect 25663 7461 25713 7477
rect 21299 7329 21349 7357
rect 22981 7402 23031 7415
rect 23199 7402 23249 7415
rect 23407 7402 23457 7415
rect 24439 7413 24489 7426
rect 24647 7413 24697 7426
rect 24865 7413 24915 7426
rect 26560 7470 26610 7498
rect 22183 7351 22233 7367
rect 22401 7351 22451 7367
rect 22609 7351 22659 7367
rect 7329 7134 7346 7154
rect 7366 7134 7379 7154
rect 7329 7106 7379 7134
rect 4813 7034 4863 7062
rect 2539 6980 2589 6993
rect 2747 6980 2797 6993
rect 2965 6980 3015 6993
rect 4813 7014 4826 7034
rect 4846 7014 4863 7034
rect 4813 6985 4863 7014
rect 5031 7037 5081 7062
rect 5031 7017 5044 7037
rect 5064 7017 5081 7037
rect 5031 6985 5081 7017
rect 5239 7035 5289 7062
rect 5239 7015 5262 7035
rect 5282 7015 5289 7035
rect 5239 6985 5289 7015
rect 9987 7167 10037 7183
rect 10205 7167 10255 7183
rect 10413 7167 10463 7183
rect 11280 7165 11330 7195
rect 11280 7145 11287 7165
rect 11307 7145 11330 7165
rect 11280 7118 11330 7145
rect 11488 7163 11538 7195
rect 11488 7143 11505 7163
rect 11525 7143 11538 7163
rect 11488 7118 11538 7143
rect 11706 7166 11756 7195
rect 13554 7187 13604 7200
rect 13772 7187 13822 7200
rect 13980 7187 14030 7200
rect 16607 7242 16657 7255
rect 16815 7242 16865 7255
rect 17033 7242 17083 7255
rect 18617 7261 18667 7289
rect 18617 7241 18630 7261
rect 18650 7241 18667 7261
rect 18617 7212 18667 7241
rect 18835 7264 18885 7289
rect 18835 7244 18848 7264
rect 18868 7244 18885 7264
rect 18835 7212 18885 7244
rect 19043 7262 19093 7289
rect 19043 7242 19066 7262
rect 19086 7242 19093 7262
rect 19043 7212 19093 7242
rect 19910 7224 19960 7240
rect 20118 7224 20168 7240
rect 20336 7224 20386 7240
rect 25237 7389 25287 7419
rect 25237 7369 25244 7389
rect 25264 7369 25287 7389
rect 25237 7342 25287 7369
rect 25445 7387 25495 7419
rect 25445 7367 25462 7387
rect 25482 7367 25495 7387
rect 25445 7342 25495 7367
rect 25663 7390 25713 7419
rect 25663 7370 25680 7390
rect 25700 7370 25713 7390
rect 26560 7450 26573 7470
rect 26593 7450 26610 7470
rect 26560 7421 26610 7450
rect 26778 7473 26828 7498
rect 26778 7453 26791 7473
rect 26811 7453 26828 7473
rect 26778 7421 26828 7453
rect 26986 7471 27036 7498
rect 26986 7451 27009 7471
rect 27029 7451 27036 7471
rect 26986 7421 27036 7451
rect 31821 7602 31871 7618
rect 32039 7602 32089 7618
rect 32247 7602 32297 7618
rect 33180 7598 33230 7628
rect 33180 7578 33187 7598
rect 33207 7578 33230 7598
rect 33180 7551 33230 7578
rect 33388 7596 33438 7628
rect 33388 7576 33405 7596
rect 33425 7576 33438 7596
rect 33388 7551 33438 7576
rect 33606 7599 33656 7628
rect 33606 7579 33623 7599
rect 33643 7579 33656 7599
rect 33606 7551 33656 7579
rect 29614 7473 29664 7489
rect 29822 7473 29872 7489
rect 30040 7473 30090 7489
rect 25663 7342 25713 7370
rect 27358 7414 27408 7427
rect 27576 7414 27626 7427
rect 27784 7414 27834 7427
rect 28816 7425 28866 7438
rect 29024 7425 29074 7438
rect 29242 7425 29292 7438
rect 30924 7483 30974 7511
rect 26560 7363 26610 7379
rect 26778 7363 26828 7379
rect 26986 7363 27036 7379
rect 22981 7274 23031 7302
rect 11706 7146 11723 7166
rect 11743 7146 11756 7166
rect 11706 7118 11756 7146
rect 9190 7046 9240 7074
rect 6903 6993 6953 7006
rect 7111 6993 7161 7006
rect 7329 6993 7379 7006
rect 9190 7026 9203 7046
rect 9223 7026 9240 7046
rect 9190 6997 9240 7026
rect 9408 7049 9458 7074
rect 9408 7029 9421 7049
rect 9441 7029 9458 7049
rect 9408 6997 9458 7029
rect 9616 7047 9666 7074
rect 9616 7027 9639 7047
rect 9659 7027 9666 7047
rect 9616 6997 9666 7027
rect 14351 7180 14401 7196
rect 14569 7180 14619 7196
rect 14777 7180 14827 7196
rect 15644 7178 15694 7208
rect 15644 7158 15651 7178
rect 15671 7158 15694 7178
rect 15644 7131 15694 7158
rect 15852 7176 15902 7208
rect 15852 7156 15869 7176
rect 15889 7156 15902 7176
rect 15852 7131 15902 7156
rect 16070 7179 16120 7208
rect 16070 7159 16087 7179
rect 16107 7159 16120 7179
rect 16070 7131 16120 7159
rect 17820 7161 17870 7174
rect 18038 7161 18088 7174
rect 18246 7161 18296 7174
rect 20873 7216 20923 7229
rect 21081 7216 21131 7229
rect 21299 7216 21349 7229
rect 22981 7254 22994 7274
rect 23014 7254 23031 7274
rect 22981 7225 23031 7254
rect 23199 7277 23249 7302
rect 23199 7257 23212 7277
rect 23232 7257 23249 7277
rect 23199 7225 23249 7257
rect 23407 7275 23457 7302
rect 23407 7255 23430 7275
rect 23450 7255 23457 7275
rect 23407 7225 23457 7255
rect 24274 7237 24324 7253
rect 24482 7237 24532 7253
rect 24700 7237 24750 7253
rect 29614 7401 29664 7431
rect 29614 7381 29621 7401
rect 29641 7381 29664 7401
rect 29614 7354 29664 7381
rect 29822 7399 29872 7431
rect 29822 7379 29839 7399
rect 29859 7379 29872 7399
rect 29822 7354 29872 7379
rect 30040 7402 30090 7431
rect 30040 7382 30057 7402
rect 30077 7382 30090 7402
rect 30924 7463 30937 7483
rect 30957 7463 30974 7483
rect 30924 7434 30974 7463
rect 31142 7486 31192 7511
rect 31142 7466 31155 7486
rect 31175 7466 31192 7486
rect 31142 7434 31192 7466
rect 31350 7484 31400 7511
rect 31350 7464 31373 7484
rect 31393 7464 31400 7484
rect 31350 7434 31400 7464
rect 33978 7486 34028 7502
rect 34186 7486 34236 7502
rect 34404 7486 34454 7502
rect 30040 7354 30090 7382
rect 31722 7427 31772 7440
rect 31940 7427 31990 7440
rect 32148 7427 32198 7440
rect 33180 7438 33230 7451
rect 33388 7438 33438 7451
rect 33606 7438 33656 7451
rect 30924 7376 30974 7392
rect 31142 7376 31192 7392
rect 31350 7376 31400 7392
rect 27358 7286 27408 7314
rect 13554 7059 13604 7087
rect 11280 7005 11330 7018
rect 11488 7005 11538 7018
rect 11706 7005 11756 7018
rect 13554 7039 13567 7059
rect 13587 7039 13604 7059
rect 13554 7010 13604 7039
rect 13772 7062 13822 7087
rect 13772 7042 13785 7062
rect 13805 7042 13822 7062
rect 13772 7010 13822 7042
rect 13980 7060 14030 7087
rect 13980 7040 14003 7060
rect 14023 7040 14030 7060
rect 13980 7010 14030 7040
rect 18617 7154 18667 7170
rect 18835 7154 18885 7170
rect 19043 7154 19093 7170
rect 19910 7152 19960 7182
rect 19910 7132 19917 7152
rect 19937 7132 19960 7152
rect 19910 7105 19960 7132
rect 20118 7150 20168 7182
rect 20118 7130 20135 7150
rect 20155 7130 20168 7150
rect 20118 7105 20168 7130
rect 20336 7153 20386 7182
rect 22184 7174 22234 7187
rect 22402 7174 22452 7187
rect 22610 7174 22660 7187
rect 25237 7229 25287 7242
rect 25445 7229 25495 7242
rect 25663 7229 25713 7242
rect 27358 7266 27371 7286
rect 27391 7266 27408 7286
rect 27358 7237 27408 7266
rect 27576 7289 27626 7314
rect 27576 7269 27589 7289
rect 27609 7269 27626 7289
rect 27576 7237 27626 7269
rect 27784 7287 27834 7314
rect 27784 7267 27807 7287
rect 27827 7267 27834 7287
rect 27784 7237 27834 7267
rect 28651 7249 28701 7265
rect 28859 7249 28909 7265
rect 29077 7249 29127 7265
rect 33978 7414 34028 7444
rect 33978 7394 33985 7414
rect 34005 7394 34028 7414
rect 33978 7367 34028 7394
rect 34186 7412 34236 7444
rect 34186 7392 34203 7412
rect 34223 7392 34236 7412
rect 34186 7367 34236 7392
rect 34404 7415 34454 7444
rect 34404 7395 34421 7415
rect 34441 7395 34454 7415
rect 34404 7367 34454 7395
rect 31722 7299 31772 7327
rect 20336 7133 20353 7153
rect 20373 7133 20386 7153
rect 20336 7105 20386 7133
rect 15644 7018 15694 7031
rect 15852 7018 15902 7031
rect 16070 7018 16120 7031
rect 17820 7033 17870 7061
rect 17820 7013 17833 7033
rect 17853 7013 17870 7033
rect 449 6914 499 6930
rect 667 6914 717 6930
rect 875 6914 925 6930
rect 4813 6927 4863 6943
rect 5031 6927 5081 6943
rect 5239 6927 5289 6943
rect 9190 6939 9240 6955
rect 9408 6939 9458 6955
rect 9616 6939 9666 6955
rect 13554 6952 13604 6968
rect 13772 6952 13822 6968
rect 13980 6952 14030 6968
rect 17820 6984 17870 7013
rect 18038 7036 18088 7061
rect 18038 7016 18051 7036
rect 18071 7016 18088 7036
rect 18038 6984 18088 7016
rect 18246 7034 18296 7061
rect 18246 7014 18269 7034
rect 18289 7014 18296 7034
rect 18246 6984 18296 7014
rect 22981 7167 23031 7183
rect 23199 7167 23249 7183
rect 23407 7167 23457 7183
rect 24274 7165 24324 7195
rect 24274 7145 24281 7165
rect 24301 7145 24324 7165
rect 24274 7118 24324 7145
rect 24482 7163 24532 7195
rect 24482 7143 24499 7163
rect 24519 7143 24532 7163
rect 24482 7118 24532 7143
rect 24700 7166 24750 7195
rect 26561 7186 26611 7199
rect 26779 7186 26829 7199
rect 26987 7186 27037 7199
rect 29614 7241 29664 7254
rect 29822 7241 29872 7254
rect 30040 7241 30090 7254
rect 31722 7279 31735 7299
rect 31755 7279 31772 7299
rect 31722 7250 31772 7279
rect 31940 7302 31990 7327
rect 31940 7282 31953 7302
rect 31973 7282 31990 7302
rect 31940 7250 31990 7282
rect 32148 7300 32198 7327
rect 32148 7280 32171 7300
rect 32191 7280 32198 7300
rect 32148 7250 32198 7280
rect 33015 7262 33065 7278
rect 33223 7262 33273 7278
rect 33441 7262 33491 7278
rect 24700 7146 24717 7166
rect 24737 7146 24750 7166
rect 24700 7118 24750 7146
rect 22184 7046 22234 7074
rect 19910 6992 19960 7005
rect 20118 6992 20168 7005
rect 20336 6992 20386 7005
rect 22184 7026 22197 7046
rect 22217 7026 22234 7046
rect 22184 6997 22234 7026
rect 22402 7049 22452 7074
rect 22402 7029 22415 7049
rect 22435 7029 22452 7049
rect 22402 6997 22452 7029
rect 22610 7047 22660 7074
rect 22610 7027 22633 7047
rect 22653 7027 22660 7047
rect 22610 6997 22660 7027
rect 27358 7179 27408 7195
rect 27576 7179 27626 7195
rect 27784 7179 27834 7195
rect 28651 7177 28701 7207
rect 28651 7157 28658 7177
rect 28678 7157 28701 7177
rect 28651 7130 28701 7157
rect 28859 7175 28909 7207
rect 28859 7155 28876 7175
rect 28896 7155 28909 7175
rect 28859 7130 28909 7155
rect 29077 7178 29127 7207
rect 30925 7199 30975 7212
rect 31143 7199 31193 7212
rect 31351 7199 31401 7212
rect 33978 7254 34028 7267
rect 34186 7254 34236 7267
rect 34404 7254 34454 7267
rect 29077 7158 29094 7178
rect 29114 7158 29127 7178
rect 29077 7130 29127 7158
rect 26561 7058 26611 7086
rect 24274 7005 24324 7018
rect 24482 7005 24532 7018
rect 24700 7005 24750 7018
rect 26561 7038 26574 7058
rect 26594 7038 26611 7058
rect 26561 7009 26611 7038
rect 26779 7061 26829 7086
rect 26779 7041 26792 7061
rect 26812 7041 26829 7061
rect 26779 7009 26829 7041
rect 26987 7059 27037 7086
rect 26987 7039 27010 7059
rect 27030 7039 27037 7059
rect 26987 7009 27037 7039
rect 31722 7192 31772 7208
rect 31940 7192 31990 7208
rect 32148 7192 32198 7208
rect 33015 7190 33065 7220
rect 33015 7170 33022 7190
rect 33042 7170 33065 7190
rect 33015 7143 33065 7170
rect 33223 7188 33273 7220
rect 33223 7168 33240 7188
rect 33260 7168 33273 7188
rect 33223 7143 33273 7168
rect 33441 7191 33491 7220
rect 33441 7171 33458 7191
rect 33478 7171 33491 7191
rect 33441 7143 33491 7171
rect 30925 7071 30975 7099
rect 28651 7017 28701 7030
rect 28859 7017 28909 7030
rect 29077 7017 29127 7030
rect 30925 7051 30938 7071
rect 30958 7051 30975 7071
rect 30925 7022 30975 7051
rect 31143 7074 31193 7099
rect 31143 7054 31156 7074
rect 31176 7054 31193 7074
rect 31143 7022 31193 7054
rect 31351 7072 31401 7099
rect 31351 7052 31374 7072
rect 31394 7052 31401 7072
rect 31351 7022 31401 7052
rect 33015 7030 33065 7043
rect 33223 7030 33273 7043
rect 33441 7030 33491 7043
rect 17820 6926 17870 6942
rect 18038 6926 18088 6942
rect 18246 6926 18296 6942
rect 22184 6939 22234 6955
rect 22402 6939 22452 6955
rect 22610 6939 22660 6955
rect 26561 6951 26611 6967
rect 26779 6951 26829 6967
rect 26987 6951 27037 6967
rect 30925 6964 30975 6980
rect 31143 6964 31193 6980
rect 31351 6964 31401 6980
rect 3481 6830 3531 6846
rect 3689 6830 3739 6846
rect 3907 6830 3957 6846
rect 7845 6843 7895 6859
rect 8053 6843 8103 6859
rect 8271 6843 8321 6859
rect 12222 6855 12272 6871
rect 12430 6855 12480 6871
rect 12648 6855 12698 6871
rect 16586 6868 16636 6884
rect 16794 6868 16844 6884
rect 17012 6868 17062 6884
rect 1391 6767 1441 6780
rect 1609 6767 1659 6780
rect 1817 6767 1867 6780
rect 3481 6758 3531 6788
rect 3481 6738 3488 6758
rect 3508 6738 3531 6758
rect 3481 6711 3531 6738
rect 3689 6756 3739 6788
rect 3689 6736 3706 6756
rect 3726 6736 3739 6756
rect 3689 6711 3739 6736
rect 3907 6759 3957 6788
rect 3907 6739 3924 6759
rect 3944 6739 3957 6759
rect 5755 6780 5805 6793
rect 5973 6780 6023 6793
rect 6181 6780 6231 6793
rect 3907 6711 3957 6739
rect 1391 6639 1441 6667
rect 1391 6619 1404 6639
rect 1424 6619 1441 6639
rect 1391 6590 1441 6619
rect 1609 6642 1659 6667
rect 1609 6622 1622 6642
rect 1642 6622 1659 6642
rect 1609 6590 1659 6622
rect 1817 6640 1867 6667
rect 1817 6620 1840 6640
rect 1860 6620 1867 6640
rect 1817 6590 1867 6620
rect 2684 6602 2734 6618
rect 2892 6602 2942 6618
rect 3110 6602 3160 6618
rect 7845 6771 7895 6801
rect 7845 6751 7852 6771
rect 7872 6751 7895 6771
rect 7845 6724 7895 6751
rect 8053 6769 8103 6801
rect 8053 6749 8070 6769
rect 8090 6749 8103 6769
rect 8053 6724 8103 6749
rect 8271 6772 8321 6801
rect 8271 6752 8288 6772
rect 8308 6752 8321 6772
rect 10132 6792 10182 6805
rect 10350 6792 10400 6805
rect 10558 6792 10608 6805
rect 8271 6724 8321 6752
rect 5755 6652 5805 6680
rect 5755 6632 5768 6652
rect 5788 6632 5805 6652
rect 428 6543 478 6556
rect 646 6543 696 6556
rect 854 6543 904 6556
rect 3481 6598 3531 6611
rect 3689 6598 3739 6611
rect 3907 6598 3957 6611
rect 5755 6603 5805 6632
rect 5973 6655 6023 6680
rect 5973 6635 5986 6655
rect 6006 6635 6023 6655
rect 5973 6603 6023 6635
rect 6181 6653 6231 6680
rect 6181 6633 6204 6653
rect 6224 6633 6231 6653
rect 6181 6603 6231 6633
rect 7048 6615 7098 6631
rect 7256 6615 7306 6631
rect 7474 6615 7524 6631
rect 12222 6783 12272 6813
rect 12222 6763 12229 6783
rect 12249 6763 12272 6783
rect 12222 6736 12272 6763
rect 12430 6781 12480 6813
rect 12430 6761 12447 6781
rect 12467 6761 12480 6781
rect 12430 6736 12480 6761
rect 12648 6784 12698 6813
rect 12648 6764 12665 6784
rect 12685 6764 12698 6784
rect 14496 6805 14546 6818
rect 14714 6805 14764 6818
rect 14922 6805 14972 6818
rect 12648 6736 12698 6764
rect 10132 6664 10182 6692
rect 10132 6644 10145 6664
rect 10165 6644 10182 6664
rect 1391 6532 1441 6548
rect 1609 6532 1659 6548
rect 1817 6532 1867 6548
rect 2684 6530 2734 6560
rect 2684 6510 2691 6530
rect 2711 6510 2734 6530
rect 2684 6483 2734 6510
rect 2892 6528 2942 6560
rect 2892 6508 2909 6528
rect 2929 6508 2942 6528
rect 2892 6483 2942 6508
rect 3110 6531 3160 6560
rect 3110 6511 3127 6531
rect 3147 6511 3160 6531
rect 4792 6556 4842 6569
rect 5010 6556 5060 6569
rect 5218 6556 5268 6569
rect 7845 6611 7895 6624
rect 8053 6611 8103 6624
rect 8271 6611 8321 6624
rect 10132 6615 10182 6644
rect 10350 6667 10400 6692
rect 10350 6647 10363 6667
rect 10383 6647 10400 6667
rect 10350 6615 10400 6647
rect 10558 6665 10608 6692
rect 10558 6645 10581 6665
rect 10601 6645 10608 6665
rect 10558 6615 10608 6645
rect 11425 6627 11475 6643
rect 11633 6627 11683 6643
rect 11851 6627 11901 6643
rect 16586 6796 16636 6826
rect 16586 6776 16593 6796
rect 16613 6776 16636 6796
rect 16586 6749 16636 6776
rect 16794 6794 16844 6826
rect 16794 6774 16811 6794
rect 16831 6774 16844 6794
rect 16794 6749 16844 6774
rect 17012 6797 17062 6826
rect 20852 6842 20902 6858
rect 21060 6842 21110 6858
rect 21278 6842 21328 6858
rect 25216 6855 25266 6871
rect 25424 6855 25474 6871
rect 25642 6855 25692 6871
rect 29593 6867 29643 6883
rect 29801 6867 29851 6883
rect 30019 6867 30069 6883
rect 33957 6880 34007 6896
rect 34165 6880 34215 6896
rect 34383 6880 34433 6896
rect 17012 6777 17029 6797
rect 17049 6777 17062 6797
rect 17012 6749 17062 6777
rect 18762 6779 18812 6792
rect 18980 6779 19030 6792
rect 19188 6779 19238 6792
rect 14496 6677 14546 6705
rect 14496 6657 14509 6677
rect 14529 6657 14546 6677
rect 3110 6483 3160 6511
rect 428 6415 478 6443
rect 428 6395 441 6415
rect 461 6395 478 6415
rect 428 6366 478 6395
rect 646 6418 696 6443
rect 646 6398 659 6418
rect 679 6398 696 6418
rect 646 6366 696 6398
rect 854 6416 904 6443
rect 854 6396 877 6416
rect 897 6396 904 6416
rect 854 6366 904 6396
rect 5755 6545 5805 6561
rect 5973 6545 6023 6561
rect 6181 6545 6231 6561
rect 7048 6543 7098 6573
rect 7048 6523 7055 6543
rect 7075 6523 7098 6543
rect 7048 6496 7098 6523
rect 7256 6541 7306 6573
rect 7256 6521 7273 6541
rect 7293 6521 7306 6541
rect 7256 6496 7306 6521
rect 7474 6544 7524 6573
rect 7474 6524 7491 6544
rect 7511 6524 7524 6544
rect 9169 6568 9219 6581
rect 9387 6568 9437 6581
rect 9595 6568 9645 6581
rect 12222 6623 12272 6636
rect 12430 6623 12480 6636
rect 12648 6623 12698 6636
rect 14496 6628 14546 6657
rect 14714 6680 14764 6705
rect 14714 6660 14727 6680
rect 14747 6660 14764 6680
rect 14714 6628 14764 6660
rect 14922 6678 14972 6705
rect 14922 6658 14945 6678
rect 14965 6658 14972 6678
rect 14922 6628 14972 6658
rect 15789 6640 15839 6656
rect 15997 6640 16047 6656
rect 16215 6640 16265 6656
rect 20852 6770 20902 6800
rect 20852 6750 20859 6770
rect 20879 6750 20902 6770
rect 20852 6723 20902 6750
rect 21060 6768 21110 6800
rect 21060 6748 21077 6768
rect 21097 6748 21110 6768
rect 21060 6723 21110 6748
rect 21278 6771 21328 6800
rect 21278 6751 21295 6771
rect 21315 6751 21328 6771
rect 23126 6792 23176 6805
rect 23344 6792 23394 6805
rect 23552 6792 23602 6805
rect 21278 6723 21328 6751
rect 7474 6496 7524 6524
rect 3482 6418 3532 6434
rect 3690 6418 3740 6434
rect 3908 6418 3958 6434
rect 1226 6359 1276 6372
rect 1444 6359 1494 6372
rect 1652 6359 1702 6372
rect 2684 6370 2734 6383
rect 2892 6370 2942 6383
rect 3110 6370 3160 6383
rect 4792 6428 4842 6456
rect 428 6308 478 6324
rect 646 6308 696 6324
rect 854 6308 904 6324
rect 3482 6346 3532 6376
rect 3482 6326 3489 6346
rect 3509 6326 3532 6346
rect 3482 6299 3532 6326
rect 3690 6344 3740 6376
rect 3690 6324 3707 6344
rect 3727 6324 3740 6344
rect 3690 6299 3740 6324
rect 3908 6347 3958 6376
rect 3908 6327 3925 6347
rect 3945 6327 3958 6347
rect 4792 6408 4805 6428
rect 4825 6408 4842 6428
rect 4792 6379 4842 6408
rect 5010 6431 5060 6456
rect 5010 6411 5023 6431
rect 5043 6411 5060 6431
rect 5010 6379 5060 6411
rect 5218 6429 5268 6456
rect 5218 6409 5241 6429
rect 5261 6409 5268 6429
rect 5218 6379 5268 6409
rect 10132 6557 10182 6573
rect 10350 6557 10400 6573
rect 10558 6557 10608 6573
rect 11425 6555 11475 6585
rect 11425 6535 11432 6555
rect 11452 6535 11475 6555
rect 11425 6508 11475 6535
rect 11633 6553 11683 6585
rect 11633 6533 11650 6553
rect 11670 6533 11683 6553
rect 11633 6508 11683 6533
rect 11851 6556 11901 6585
rect 11851 6536 11868 6556
rect 11888 6536 11901 6556
rect 13533 6581 13583 6594
rect 13751 6581 13801 6594
rect 13959 6581 14009 6594
rect 16586 6636 16636 6649
rect 16794 6636 16844 6649
rect 17012 6636 17062 6649
rect 18762 6651 18812 6679
rect 18762 6631 18775 6651
rect 18795 6631 18812 6651
rect 18762 6602 18812 6631
rect 18980 6654 19030 6679
rect 18980 6634 18993 6654
rect 19013 6634 19030 6654
rect 18980 6602 19030 6634
rect 19188 6652 19238 6679
rect 19188 6632 19211 6652
rect 19231 6632 19238 6652
rect 19188 6602 19238 6632
rect 20055 6614 20105 6630
rect 20263 6614 20313 6630
rect 20481 6614 20531 6630
rect 25216 6783 25266 6813
rect 25216 6763 25223 6783
rect 25243 6763 25266 6783
rect 25216 6736 25266 6763
rect 25424 6781 25474 6813
rect 25424 6761 25441 6781
rect 25461 6761 25474 6781
rect 25424 6736 25474 6761
rect 25642 6784 25692 6813
rect 25642 6764 25659 6784
rect 25679 6764 25692 6784
rect 27503 6804 27553 6817
rect 27721 6804 27771 6817
rect 27929 6804 27979 6817
rect 25642 6736 25692 6764
rect 23126 6664 23176 6692
rect 23126 6644 23139 6664
rect 23159 6644 23176 6664
rect 11851 6508 11901 6536
rect 7846 6431 7896 6447
rect 8054 6431 8104 6447
rect 8272 6431 8322 6447
rect 3908 6299 3958 6327
rect 5590 6372 5640 6385
rect 5808 6372 5858 6385
rect 6016 6372 6066 6385
rect 7048 6383 7098 6396
rect 7256 6383 7306 6396
rect 7474 6383 7524 6396
rect 9169 6440 9219 6468
rect 4792 6321 4842 6337
rect 5010 6321 5060 6337
rect 5218 6321 5268 6337
rect 1226 6231 1276 6259
rect 1226 6211 1239 6231
rect 1259 6211 1276 6231
rect 1226 6182 1276 6211
rect 1444 6234 1494 6259
rect 1444 6214 1457 6234
rect 1477 6214 1494 6234
rect 1444 6182 1494 6214
rect 1652 6232 1702 6259
rect 1652 6212 1675 6232
rect 1695 6212 1702 6232
rect 1652 6182 1702 6212
rect 2585 6192 2635 6208
rect 2793 6192 2843 6208
rect 3011 6192 3061 6208
rect 7846 6359 7896 6389
rect 7846 6339 7853 6359
rect 7873 6339 7896 6359
rect 7846 6312 7896 6339
rect 8054 6357 8104 6389
rect 8054 6337 8071 6357
rect 8091 6337 8104 6357
rect 8054 6312 8104 6337
rect 8272 6360 8322 6389
rect 8272 6340 8289 6360
rect 8309 6340 8322 6360
rect 9169 6420 9182 6440
rect 9202 6420 9219 6440
rect 9169 6391 9219 6420
rect 9387 6443 9437 6468
rect 9387 6423 9400 6443
rect 9420 6423 9437 6443
rect 9387 6391 9437 6423
rect 9595 6441 9645 6468
rect 9595 6421 9618 6441
rect 9638 6421 9645 6441
rect 9595 6391 9645 6421
rect 14496 6570 14546 6586
rect 14714 6570 14764 6586
rect 14922 6570 14972 6586
rect 15789 6568 15839 6598
rect 15789 6548 15796 6568
rect 15816 6548 15839 6568
rect 15789 6521 15839 6548
rect 15997 6566 16047 6598
rect 15997 6546 16014 6566
rect 16034 6546 16047 6566
rect 15997 6521 16047 6546
rect 16215 6569 16265 6598
rect 16215 6549 16232 6569
rect 16252 6549 16265 6569
rect 16215 6521 16265 6549
rect 17799 6555 17849 6568
rect 18017 6555 18067 6568
rect 18225 6555 18275 6568
rect 20852 6610 20902 6623
rect 21060 6610 21110 6623
rect 21278 6610 21328 6623
rect 23126 6615 23176 6644
rect 23344 6667 23394 6692
rect 23344 6647 23357 6667
rect 23377 6647 23394 6667
rect 23344 6615 23394 6647
rect 23552 6665 23602 6692
rect 23552 6645 23575 6665
rect 23595 6645 23602 6665
rect 23552 6615 23602 6645
rect 24419 6627 24469 6643
rect 24627 6627 24677 6643
rect 24845 6627 24895 6643
rect 29593 6795 29643 6825
rect 29593 6775 29600 6795
rect 29620 6775 29643 6795
rect 29593 6748 29643 6775
rect 29801 6793 29851 6825
rect 29801 6773 29818 6793
rect 29838 6773 29851 6793
rect 29801 6748 29851 6773
rect 30019 6796 30069 6825
rect 30019 6776 30036 6796
rect 30056 6776 30069 6796
rect 31867 6817 31917 6830
rect 32085 6817 32135 6830
rect 32293 6817 32343 6830
rect 30019 6748 30069 6776
rect 27503 6676 27553 6704
rect 27503 6656 27516 6676
rect 27536 6656 27553 6676
rect 12223 6443 12273 6459
rect 12431 6443 12481 6459
rect 12649 6443 12699 6459
rect 8272 6312 8322 6340
rect 9967 6384 10017 6397
rect 10185 6384 10235 6397
rect 10393 6384 10443 6397
rect 11425 6395 11475 6408
rect 11633 6395 11683 6408
rect 11851 6395 11901 6408
rect 13533 6453 13583 6481
rect 9169 6333 9219 6349
rect 9387 6333 9437 6349
rect 9595 6333 9645 6349
rect 5590 6244 5640 6272
rect 429 6131 479 6144
rect 647 6131 697 6144
rect 855 6131 905 6144
rect 3482 6186 3532 6199
rect 3690 6186 3740 6199
rect 3908 6186 3958 6199
rect 5590 6224 5603 6244
rect 5623 6224 5640 6244
rect 5590 6195 5640 6224
rect 5808 6247 5858 6272
rect 5808 6227 5821 6247
rect 5841 6227 5858 6247
rect 5808 6195 5858 6227
rect 6016 6245 6066 6272
rect 6016 6225 6039 6245
rect 6059 6225 6066 6245
rect 6016 6195 6066 6225
rect 6949 6205 6999 6221
rect 7157 6205 7207 6221
rect 7375 6205 7425 6221
rect 12223 6371 12273 6401
rect 12223 6351 12230 6371
rect 12250 6351 12273 6371
rect 12223 6324 12273 6351
rect 12431 6369 12481 6401
rect 12431 6349 12448 6369
rect 12468 6349 12481 6369
rect 12431 6324 12481 6349
rect 12649 6372 12699 6401
rect 12649 6352 12666 6372
rect 12686 6352 12699 6372
rect 13533 6433 13546 6453
rect 13566 6433 13583 6453
rect 13533 6404 13583 6433
rect 13751 6456 13801 6481
rect 13751 6436 13764 6456
rect 13784 6436 13801 6456
rect 13751 6404 13801 6436
rect 13959 6454 14009 6481
rect 13959 6434 13982 6454
rect 14002 6434 14009 6454
rect 13959 6404 14009 6434
rect 16587 6456 16637 6472
rect 16795 6456 16845 6472
rect 17013 6456 17063 6472
rect 12649 6324 12699 6352
rect 14331 6397 14381 6410
rect 14549 6397 14599 6410
rect 14757 6397 14807 6410
rect 15789 6408 15839 6421
rect 15997 6408 16047 6421
rect 16215 6408 16265 6421
rect 18762 6544 18812 6560
rect 18980 6544 19030 6560
rect 19188 6544 19238 6560
rect 20055 6542 20105 6572
rect 20055 6522 20062 6542
rect 20082 6522 20105 6542
rect 20055 6495 20105 6522
rect 20263 6540 20313 6572
rect 20263 6520 20280 6540
rect 20300 6520 20313 6540
rect 20263 6495 20313 6520
rect 20481 6543 20531 6572
rect 20481 6523 20498 6543
rect 20518 6523 20531 6543
rect 22163 6568 22213 6581
rect 22381 6568 22431 6581
rect 22589 6568 22639 6581
rect 25216 6623 25266 6636
rect 25424 6623 25474 6636
rect 25642 6623 25692 6636
rect 27503 6627 27553 6656
rect 27721 6679 27771 6704
rect 27721 6659 27734 6679
rect 27754 6659 27771 6679
rect 27721 6627 27771 6659
rect 27929 6677 27979 6704
rect 27929 6657 27952 6677
rect 27972 6657 27979 6677
rect 27929 6627 27979 6657
rect 28796 6639 28846 6655
rect 29004 6639 29054 6655
rect 29222 6639 29272 6655
rect 33957 6808 34007 6838
rect 33957 6788 33964 6808
rect 33984 6788 34007 6808
rect 33957 6761 34007 6788
rect 34165 6806 34215 6838
rect 34165 6786 34182 6806
rect 34202 6786 34215 6806
rect 34165 6761 34215 6786
rect 34383 6809 34433 6838
rect 34383 6789 34400 6809
rect 34420 6789 34433 6809
rect 34383 6761 34433 6789
rect 31867 6689 31917 6717
rect 31867 6669 31880 6689
rect 31900 6669 31917 6689
rect 20481 6495 20531 6523
rect 13533 6346 13583 6362
rect 13751 6346 13801 6362
rect 13959 6346 14009 6362
rect 9967 6256 10017 6284
rect 1226 6124 1276 6140
rect 1444 6124 1494 6140
rect 1652 6124 1702 6140
rect 2585 6120 2635 6150
rect 2585 6100 2592 6120
rect 2612 6100 2635 6120
rect 2585 6073 2635 6100
rect 2793 6118 2843 6150
rect 2793 6098 2810 6118
rect 2830 6098 2843 6118
rect 2793 6073 2843 6098
rect 3011 6121 3061 6150
rect 4793 6144 4843 6157
rect 5011 6144 5061 6157
rect 5219 6144 5269 6157
rect 7846 6199 7896 6212
rect 8054 6199 8104 6212
rect 8272 6199 8322 6212
rect 9967 6236 9980 6256
rect 10000 6236 10017 6256
rect 9967 6207 10017 6236
rect 10185 6259 10235 6284
rect 10185 6239 10198 6259
rect 10218 6239 10235 6259
rect 10185 6207 10235 6239
rect 10393 6257 10443 6284
rect 10393 6237 10416 6257
rect 10436 6237 10443 6257
rect 10393 6207 10443 6237
rect 11326 6217 11376 6233
rect 11534 6217 11584 6233
rect 11752 6217 11802 6233
rect 16587 6384 16637 6414
rect 16587 6364 16594 6384
rect 16614 6364 16637 6384
rect 16587 6337 16637 6364
rect 16795 6382 16845 6414
rect 16795 6362 16812 6382
rect 16832 6362 16845 6382
rect 16795 6337 16845 6362
rect 17013 6385 17063 6414
rect 17013 6365 17030 6385
rect 17050 6365 17063 6385
rect 17799 6427 17849 6455
rect 17013 6337 17063 6365
rect 17799 6407 17812 6427
rect 17832 6407 17849 6427
rect 17799 6378 17849 6407
rect 18017 6430 18067 6455
rect 18017 6410 18030 6430
rect 18050 6410 18067 6430
rect 18017 6378 18067 6410
rect 18225 6428 18275 6455
rect 18225 6408 18248 6428
rect 18268 6408 18275 6428
rect 18225 6378 18275 6408
rect 23126 6557 23176 6573
rect 23344 6557 23394 6573
rect 23552 6557 23602 6573
rect 24419 6555 24469 6585
rect 24419 6535 24426 6555
rect 24446 6535 24469 6555
rect 24419 6508 24469 6535
rect 24627 6553 24677 6585
rect 24627 6533 24644 6553
rect 24664 6533 24677 6553
rect 24627 6508 24677 6533
rect 24845 6556 24895 6585
rect 24845 6536 24862 6556
rect 24882 6536 24895 6556
rect 26540 6580 26590 6593
rect 26758 6580 26808 6593
rect 26966 6580 27016 6593
rect 29593 6635 29643 6648
rect 29801 6635 29851 6648
rect 30019 6635 30069 6648
rect 31867 6640 31917 6669
rect 32085 6692 32135 6717
rect 32085 6672 32098 6692
rect 32118 6672 32135 6692
rect 32085 6640 32135 6672
rect 32293 6690 32343 6717
rect 32293 6670 32316 6690
rect 32336 6670 32343 6690
rect 32293 6640 32343 6670
rect 33160 6652 33210 6668
rect 33368 6652 33418 6668
rect 33586 6652 33636 6668
rect 24845 6508 24895 6536
rect 20853 6430 20903 6446
rect 21061 6430 21111 6446
rect 21279 6430 21329 6446
rect 14331 6269 14381 6297
rect 3011 6101 3028 6121
rect 3048 6101 3061 6121
rect 3011 6073 3061 6101
rect 429 6003 479 6031
rect 429 5983 442 6003
rect 462 5983 479 6003
rect 429 5954 479 5983
rect 647 6006 697 6031
rect 647 5986 660 6006
rect 680 5986 697 6006
rect 647 5954 697 5986
rect 855 6004 905 6031
rect 855 5984 878 6004
rect 898 5984 905 6004
rect 855 5954 905 5984
rect 5590 6137 5640 6153
rect 5808 6137 5858 6153
rect 6016 6137 6066 6153
rect 6949 6133 6999 6163
rect 6949 6113 6956 6133
rect 6976 6113 6999 6133
rect 6949 6086 6999 6113
rect 7157 6131 7207 6163
rect 7157 6111 7174 6131
rect 7194 6111 7207 6131
rect 7157 6086 7207 6111
rect 7375 6134 7425 6163
rect 9170 6156 9220 6169
rect 9388 6156 9438 6169
rect 9596 6156 9646 6169
rect 12223 6211 12273 6224
rect 12431 6211 12481 6224
rect 12649 6211 12699 6224
rect 14331 6249 14344 6269
rect 14364 6249 14381 6269
rect 14331 6220 14381 6249
rect 14549 6272 14599 6297
rect 14549 6252 14562 6272
rect 14582 6252 14599 6272
rect 14549 6220 14599 6252
rect 14757 6270 14807 6297
rect 14757 6250 14780 6270
rect 14800 6250 14807 6270
rect 14757 6220 14807 6250
rect 15690 6230 15740 6246
rect 15898 6230 15948 6246
rect 16116 6230 16166 6246
rect 18597 6371 18647 6384
rect 18815 6371 18865 6384
rect 19023 6371 19073 6384
rect 20055 6382 20105 6395
rect 20263 6382 20313 6395
rect 20481 6382 20531 6395
rect 22163 6440 22213 6468
rect 17799 6320 17849 6336
rect 18017 6320 18067 6336
rect 18225 6320 18275 6336
rect 20853 6358 20903 6388
rect 20853 6338 20860 6358
rect 20880 6338 20903 6358
rect 20853 6311 20903 6338
rect 21061 6356 21111 6388
rect 21061 6336 21078 6356
rect 21098 6336 21111 6356
rect 21061 6311 21111 6336
rect 21279 6359 21329 6388
rect 21279 6339 21296 6359
rect 21316 6339 21329 6359
rect 22163 6420 22176 6440
rect 22196 6420 22213 6440
rect 22163 6391 22213 6420
rect 22381 6443 22431 6468
rect 22381 6423 22394 6443
rect 22414 6423 22431 6443
rect 22381 6391 22431 6423
rect 22589 6441 22639 6468
rect 22589 6421 22612 6441
rect 22632 6421 22639 6441
rect 22589 6391 22639 6421
rect 27503 6569 27553 6585
rect 27721 6569 27771 6585
rect 27929 6569 27979 6585
rect 28796 6567 28846 6597
rect 28796 6547 28803 6567
rect 28823 6547 28846 6567
rect 28796 6520 28846 6547
rect 29004 6565 29054 6597
rect 29004 6545 29021 6565
rect 29041 6545 29054 6565
rect 29004 6520 29054 6545
rect 29222 6568 29272 6597
rect 29222 6548 29239 6568
rect 29259 6548 29272 6568
rect 30904 6593 30954 6606
rect 31122 6593 31172 6606
rect 31330 6593 31380 6606
rect 33957 6648 34007 6661
rect 34165 6648 34215 6661
rect 34383 6648 34433 6661
rect 29222 6520 29272 6548
rect 25217 6443 25267 6459
rect 25425 6443 25475 6459
rect 25643 6443 25693 6459
rect 21279 6311 21329 6339
rect 22961 6384 23011 6397
rect 23179 6384 23229 6397
rect 23387 6384 23437 6397
rect 24419 6395 24469 6408
rect 24627 6395 24677 6408
rect 24845 6395 24895 6408
rect 26540 6452 26590 6480
rect 22163 6333 22213 6349
rect 22381 6333 22431 6349
rect 22589 6333 22639 6349
rect 7375 6114 7392 6134
rect 7412 6114 7425 6134
rect 7375 6086 7425 6114
rect 4793 6016 4843 6044
rect 2585 5960 2635 5973
rect 2793 5960 2843 5973
rect 3011 5960 3061 5973
rect 4793 5996 4806 6016
rect 4826 5996 4843 6016
rect 4793 5967 4843 5996
rect 5011 6019 5061 6044
rect 5011 5999 5024 6019
rect 5044 5999 5061 6019
rect 5011 5967 5061 5999
rect 5219 6017 5269 6044
rect 5219 5997 5242 6017
rect 5262 5997 5269 6017
rect 5219 5967 5269 5997
rect 9967 6149 10017 6165
rect 10185 6149 10235 6165
rect 10393 6149 10443 6165
rect 11326 6145 11376 6175
rect 11326 6125 11333 6145
rect 11353 6125 11376 6145
rect 11326 6098 11376 6125
rect 11534 6143 11584 6175
rect 11534 6123 11551 6143
rect 11571 6123 11584 6143
rect 11534 6098 11584 6123
rect 11752 6146 11802 6175
rect 13534 6169 13584 6182
rect 13752 6169 13802 6182
rect 13960 6169 14010 6182
rect 16587 6224 16637 6237
rect 16795 6224 16845 6237
rect 17013 6224 17063 6237
rect 18597 6243 18647 6271
rect 18597 6223 18610 6243
rect 18630 6223 18647 6243
rect 18597 6194 18647 6223
rect 18815 6246 18865 6271
rect 18815 6226 18828 6246
rect 18848 6226 18865 6246
rect 18815 6194 18865 6226
rect 19023 6244 19073 6271
rect 19023 6224 19046 6244
rect 19066 6224 19073 6244
rect 19023 6194 19073 6224
rect 19956 6204 20006 6220
rect 20164 6204 20214 6220
rect 20382 6204 20432 6220
rect 25217 6371 25267 6401
rect 25217 6351 25224 6371
rect 25244 6351 25267 6371
rect 25217 6324 25267 6351
rect 25425 6369 25475 6401
rect 25425 6349 25442 6369
rect 25462 6349 25475 6369
rect 25425 6324 25475 6349
rect 25643 6372 25693 6401
rect 25643 6352 25660 6372
rect 25680 6352 25693 6372
rect 26540 6432 26553 6452
rect 26573 6432 26590 6452
rect 26540 6403 26590 6432
rect 26758 6455 26808 6480
rect 26758 6435 26771 6455
rect 26791 6435 26808 6455
rect 26758 6403 26808 6435
rect 26966 6453 27016 6480
rect 26966 6433 26989 6453
rect 27009 6433 27016 6453
rect 26966 6403 27016 6433
rect 31867 6582 31917 6598
rect 32085 6582 32135 6598
rect 32293 6582 32343 6598
rect 33160 6580 33210 6610
rect 33160 6560 33167 6580
rect 33187 6560 33210 6580
rect 33160 6533 33210 6560
rect 33368 6578 33418 6610
rect 33368 6558 33385 6578
rect 33405 6558 33418 6578
rect 33368 6533 33418 6558
rect 33586 6581 33636 6610
rect 33586 6561 33603 6581
rect 33623 6561 33636 6581
rect 33586 6533 33636 6561
rect 29594 6455 29644 6471
rect 29802 6455 29852 6471
rect 30020 6455 30070 6471
rect 25643 6324 25693 6352
rect 27338 6396 27388 6409
rect 27556 6396 27606 6409
rect 27764 6396 27814 6409
rect 28796 6407 28846 6420
rect 29004 6407 29054 6420
rect 29222 6407 29272 6420
rect 30904 6465 30954 6493
rect 26540 6345 26590 6361
rect 26758 6345 26808 6361
rect 26966 6345 27016 6361
rect 22961 6256 23011 6284
rect 11752 6126 11769 6146
rect 11789 6126 11802 6146
rect 11752 6098 11802 6126
rect 9170 6028 9220 6056
rect 6949 5973 6999 5986
rect 7157 5973 7207 5986
rect 7375 5973 7425 5986
rect 9170 6008 9183 6028
rect 9203 6008 9220 6028
rect 9170 5979 9220 6008
rect 9388 6031 9438 6056
rect 9388 6011 9401 6031
rect 9421 6011 9438 6031
rect 9388 5979 9438 6011
rect 9596 6029 9646 6056
rect 9596 6009 9619 6029
rect 9639 6009 9646 6029
rect 9596 5979 9646 6009
rect 14331 6162 14381 6178
rect 14549 6162 14599 6178
rect 14757 6162 14807 6178
rect 15690 6158 15740 6188
rect 15690 6138 15697 6158
rect 15717 6138 15740 6158
rect 15690 6111 15740 6138
rect 15898 6156 15948 6188
rect 15898 6136 15915 6156
rect 15935 6136 15948 6156
rect 15898 6111 15948 6136
rect 16116 6159 16166 6188
rect 16116 6139 16133 6159
rect 16153 6139 16166 6159
rect 16116 6111 16166 6139
rect 17800 6143 17850 6156
rect 18018 6143 18068 6156
rect 18226 6143 18276 6156
rect 20853 6198 20903 6211
rect 21061 6198 21111 6211
rect 21279 6198 21329 6211
rect 22961 6236 22974 6256
rect 22994 6236 23011 6256
rect 22961 6207 23011 6236
rect 23179 6259 23229 6284
rect 23179 6239 23192 6259
rect 23212 6239 23229 6259
rect 23179 6207 23229 6239
rect 23387 6257 23437 6284
rect 23387 6237 23410 6257
rect 23430 6237 23437 6257
rect 23387 6207 23437 6237
rect 24320 6217 24370 6233
rect 24528 6217 24578 6233
rect 24746 6217 24796 6233
rect 29594 6383 29644 6413
rect 29594 6363 29601 6383
rect 29621 6363 29644 6383
rect 29594 6336 29644 6363
rect 29802 6381 29852 6413
rect 29802 6361 29819 6381
rect 29839 6361 29852 6381
rect 29802 6336 29852 6361
rect 30020 6384 30070 6413
rect 30020 6364 30037 6384
rect 30057 6364 30070 6384
rect 30904 6445 30917 6465
rect 30937 6445 30954 6465
rect 30904 6416 30954 6445
rect 31122 6468 31172 6493
rect 31122 6448 31135 6468
rect 31155 6448 31172 6468
rect 31122 6416 31172 6448
rect 31330 6466 31380 6493
rect 31330 6446 31353 6466
rect 31373 6446 31380 6466
rect 31330 6416 31380 6446
rect 33958 6468 34008 6484
rect 34166 6468 34216 6484
rect 34384 6468 34434 6484
rect 30020 6336 30070 6364
rect 31702 6409 31752 6422
rect 31920 6409 31970 6422
rect 32128 6409 32178 6422
rect 33160 6420 33210 6433
rect 33368 6420 33418 6433
rect 33586 6420 33636 6433
rect 30904 6358 30954 6374
rect 31122 6358 31172 6374
rect 31330 6358 31380 6374
rect 27338 6268 27388 6296
rect 13534 6041 13584 6069
rect 11326 5985 11376 5998
rect 11534 5985 11584 5998
rect 11752 5985 11802 5998
rect 13534 6021 13547 6041
rect 13567 6021 13584 6041
rect 13534 5992 13584 6021
rect 13752 6044 13802 6069
rect 13752 6024 13765 6044
rect 13785 6024 13802 6044
rect 13752 5992 13802 6024
rect 13960 6042 14010 6069
rect 13960 6022 13983 6042
rect 14003 6022 14010 6042
rect 13960 5992 14010 6022
rect 18597 6136 18647 6152
rect 18815 6136 18865 6152
rect 19023 6136 19073 6152
rect 19956 6132 20006 6162
rect 19956 6112 19963 6132
rect 19983 6112 20006 6132
rect 19956 6085 20006 6112
rect 20164 6130 20214 6162
rect 20164 6110 20181 6130
rect 20201 6110 20214 6130
rect 20164 6085 20214 6110
rect 20382 6133 20432 6162
rect 22164 6156 22214 6169
rect 22382 6156 22432 6169
rect 22590 6156 22640 6169
rect 25217 6211 25267 6224
rect 25425 6211 25475 6224
rect 25643 6211 25693 6224
rect 27338 6248 27351 6268
rect 27371 6248 27388 6268
rect 27338 6219 27388 6248
rect 27556 6271 27606 6296
rect 27556 6251 27569 6271
rect 27589 6251 27606 6271
rect 27556 6219 27606 6251
rect 27764 6269 27814 6296
rect 27764 6249 27787 6269
rect 27807 6249 27814 6269
rect 27764 6219 27814 6249
rect 28697 6229 28747 6245
rect 28905 6229 28955 6245
rect 29123 6229 29173 6245
rect 33958 6396 34008 6426
rect 33958 6376 33965 6396
rect 33985 6376 34008 6396
rect 33958 6349 34008 6376
rect 34166 6394 34216 6426
rect 34166 6374 34183 6394
rect 34203 6374 34216 6394
rect 34166 6349 34216 6374
rect 34384 6397 34434 6426
rect 34384 6377 34401 6397
rect 34421 6377 34434 6397
rect 34384 6349 34434 6377
rect 31702 6281 31752 6309
rect 20382 6113 20399 6133
rect 20419 6113 20432 6133
rect 20382 6085 20432 6113
rect 15690 5998 15740 6011
rect 15898 5998 15948 6011
rect 16116 5998 16166 6011
rect 17800 6015 17850 6043
rect 17800 5995 17813 6015
rect 17833 5995 17850 6015
rect 429 5896 479 5912
rect 647 5896 697 5912
rect 855 5896 905 5912
rect 4793 5909 4843 5925
rect 5011 5909 5061 5925
rect 5219 5909 5269 5925
rect 9170 5921 9220 5937
rect 9388 5921 9438 5937
rect 9596 5921 9646 5937
rect 13534 5934 13584 5950
rect 13752 5934 13802 5950
rect 13960 5934 14010 5950
rect 17800 5966 17850 5995
rect 18018 6018 18068 6043
rect 18018 5998 18031 6018
rect 18051 5998 18068 6018
rect 18018 5966 18068 5998
rect 18226 6016 18276 6043
rect 18226 5996 18249 6016
rect 18269 5996 18276 6016
rect 18226 5966 18276 5996
rect 22961 6149 23011 6165
rect 23179 6149 23229 6165
rect 23387 6149 23437 6165
rect 24320 6145 24370 6175
rect 24320 6125 24327 6145
rect 24347 6125 24370 6145
rect 24320 6098 24370 6125
rect 24528 6143 24578 6175
rect 24528 6123 24545 6143
rect 24565 6123 24578 6143
rect 24528 6098 24578 6123
rect 24746 6146 24796 6175
rect 26541 6168 26591 6181
rect 26759 6168 26809 6181
rect 26967 6168 27017 6181
rect 29594 6223 29644 6236
rect 29802 6223 29852 6236
rect 30020 6223 30070 6236
rect 31702 6261 31715 6281
rect 31735 6261 31752 6281
rect 31702 6232 31752 6261
rect 31920 6284 31970 6309
rect 31920 6264 31933 6284
rect 31953 6264 31970 6284
rect 31920 6232 31970 6264
rect 32128 6282 32178 6309
rect 32128 6262 32151 6282
rect 32171 6262 32178 6282
rect 32128 6232 32178 6262
rect 33061 6242 33111 6258
rect 33269 6242 33319 6258
rect 33487 6242 33537 6258
rect 24746 6126 24763 6146
rect 24783 6126 24796 6146
rect 24746 6098 24796 6126
rect 22164 6028 22214 6056
rect 19956 5972 20006 5985
rect 20164 5972 20214 5985
rect 20382 5972 20432 5985
rect 22164 6008 22177 6028
rect 22197 6008 22214 6028
rect 22164 5979 22214 6008
rect 22382 6031 22432 6056
rect 22382 6011 22395 6031
rect 22415 6011 22432 6031
rect 22382 5979 22432 6011
rect 22590 6029 22640 6056
rect 22590 6009 22613 6029
rect 22633 6009 22640 6029
rect 22590 5979 22640 6009
rect 27338 6161 27388 6177
rect 27556 6161 27606 6177
rect 27764 6161 27814 6177
rect 28697 6157 28747 6187
rect 28697 6137 28704 6157
rect 28724 6137 28747 6157
rect 28697 6110 28747 6137
rect 28905 6155 28955 6187
rect 28905 6135 28922 6155
rect 28942 6135 28955 6155
rect 28905 6110 28955 6135
rect 29123 6158 29173 6187
rect 30905 6181 30955 6194
rect 31123 6181 31173 6194
rect 31331 6181 31381 6194
rect 33958 6236 34008 6249
rect 34166 6236 34216 6249
rect 34384 6236 34434 6249
rect 29123 6138 29140 6158
rect 29160 6138 29173 6158
rect 29123 6110 29173 6138
rect 26541 6040 26591 6068
rect 24320 5985 24370 5998
rect 24528 5985 24578 5998
rect 24746 5985 24796 5998
rect 26541 6020 26554 6040
rect 26574 6020 26591 6040
rect 26541 5991 26591 6020
rect 26759 6043 26809 6068
rect 26759 6023 26772 6043
rect 26792 6023 26809 6043
rect 26759 5991 26809 6023
rect 26967 6041 27017 6068
rect 26967 6021 26990 6041
rect 27010 6021 27017 6041
rect 26967 5991 27017 6021
rect 31702 6174 31752 6190
rect 31920 6174 31970 6190
rect 32128 6174 32178 6190
rect 33061 6170 33111 6200
rect 33061 6150 33068 6170
rect 33088 6150 33111 6170
rect 33061 6123 33111 6150
rect 33269 6168 33319 6200
rect 33269 6148 33286 6168
rect 33306 6148 33319 6168
rect 33269 6123 33319 6148
rect 33487 6171 33537 6200
rect 33487 6151 33504 6171
rect 33524 6151 33537 6171
rect 33487 6123 33537 6151
rect 30905 6053 30955 6081
rect 28697 5997 28747 6010
rect 28905 5997 28955 6010
rect 29123 5997 29173 6010
rect 30905 6033 30918 6053
rect 30938 6033 30955 6053
rect 30905 6004 30955 6033
rect 31123 6056 31173 6081
rect 31123 6036 31136 6056
rect 31156 6036 31173 6056
rect 31123 6004 31173 6036
rect 31331 6054 31381 6081
rect 31331 6034 31354 6054
rect 31374 6034 31381 6054
rect 31331 6004 31381 6034
rect 33061 6010 33111 6023
rect 33269 6010 33319 6023
rect 33487 6010 33537 6023
rect 17800 5908 17850 5924
rect 18018 5908 18068 5924
rect 18226 5908 18276 5924
rect 22164 5921 22214 5937
rect 22382 5921 22432 5937
rect 22590 5921 22640 5937
rect 26541 5933 26591 5949
rect 26759 5933 26809 5949
rect 26967 5933 27017 5949
rect 30905 5946 30955 5962
rect 31123 5946 31173 5962
rect 31331 5946 31381 5962
rect 3464 5812 3514 5828
rect 3672 5812 3722 5828
rect 3890 5812 3940 5828
rect 7828 5825 7878 5841
rect 8036 5825 8086 5841
rect 8254 5825 8304 5841
rect 12205 5837 12255 5853
rect 12413 5837 12463 5853
rect 12631 5837 12681 5853
rect 16569 5850 16619 5866
rect 16777 5850 16827 5866
rect 16995 5850 17045 5866
rect 1308 5751 1358 5764
rect 1526 5751 1576 5764
rect 1734 5751 1784 5764
rect 3464 5740 3514 5770
rect 3464 5720 3471 5740
rect 3491 5720 3514 5740
rect 3464 5693 3514 5720
rect 3672 5738 3722 5770
rect 3672 5718 3689 5738
rect 3709 5718 3722 5738
rect 3672 5693 3722 5718
rect 3890 5741 3940 5770
rect 3890 5721 3907 5741
rect 3927 5721 3940 5741
rect 5672 5764 5722 5777
rect 5890 5764 5940 5777
rect 6098 5764 6148 5777
rect 3890 5693 3940 5721
rect 1308 5623 1358 5651
rect 1308 5603 1321 5623
rect 1341 5603 1358 5623
rect 1308 5574 1358 5603
rect 1526 5626 1576 5651
rect 1526 5606 1539 5626
rect 1559 5606 1576 5626
rect 1526 5574 1576 5606
rect 1734 5624 1784 5651
rect 1734 5604 1757 5624
rect 1777 5604 1784 5624
rect 1734 5574 1784 5604
rect 2667 5584 2717 5600
rect 2875 5584 2925 5600
rect 3093 5584 3143 5600
rect 7828 5753 7878 5783
rect 7828 5733 7835 5753
rect 7855 5733 7878 5753
rect 7828 5706 7878 5733
rect 8036 5751 8086 5783
rect 8036 5731 8053 5751
rect 8073 5731 8086 5751
rect 8036 5706 8086 5731
rect 8254 5754 8304 5783
rect 8254 5734 8271 5754
rect 8291 5734 8304 5754
rect 10049 5776 10099 5789
rect 10267 5776 10317 5789
rect 10475 5776 10525 5789
rect 8254 5706 8304 5734
rect 5672 5636 5722 5664
rect 5672 5616 5685 5636
rect 5705 5616 5722 5636
rect 411 5525 461 5538
rect 629 5525 679 5538
rect 837 5525 887 5538
rect 3464 5580 3514 5593
rect 3672 5580 3722 5593
rect 3890 5580 3940 5593
rect 5672 5587 5722 5616
rect 5890 5639 5940 5664
rect 5890 5619 5903 5639
rect 5923 5619 5940 5639
rect 5890 5587 5940 5619
rect 6098 5637 6148 5664
rect 6098 5617 6121 5637
rect 6141 5617 6148 5637
rect 6098 5587 6148 5617
rect 7031 5597 7081 5613
rect 7239 5597 7289 5613
rect 7457 5597 7507 5613
rect 12205 5765 12255 5795
rect 12205 5745 12212 5765
rect 12232 5745 12255 5765
rect 12205 5718 12255 5745
rect 12413 5763 12463 5795
rect 12413 5743 12430 5763
rect 12450 5743 12463 5763
rect 12413 5718 12463 5743
rect 12631 5766 12681 5795
rect 12631 5746 12648 5766
rect 12668 5746 12681 5766
rect 14413 5789 14463 5802
rect 14631 5789 14681 5802
rect 14839 5789 14889 5802
rect 12631 5718 12681 5746
rect 10049 5648 10099 5676
rect 10049 5628 10062 5648
rect 10082 5628 10099 5648
rect 1308 5516 1358 5532
rect 1526 5516 1576 5532
rect 1734 5516 1784 5532
rect 2667 5512 2717 5542
rect 2667 5492 2674 5512
rect 2694 5492 2717 5512
rect 2667 5465 2717 5492
rect 2875 5510 2925 5542
rect 2875 5490 2892 5510
rect 2912 5490 2925 5510
rect 2875 5465 2925 5490
rect 3093 5513 3143 5542
rect 3093 5493 3110 5513
rect 3130 5493 3143 5513
rect 4775 5538 4825 5551
rect 4993 5538 5043 5551
rect 5201 5538 5251 5551
rect 7828 5593 7878 5606
rect 8036 5593 8086 5606
rect 8254 5593 8304 5606
rect 10049 5599 10099 5628
rect 10267 5651 10317 5676
rect 10267 5631 10280 5651
rect 10300 5631 10317 5651
rect 10267 5599 10317 5631
rect 10475 5649 10525 5676
rect 10475 5629 10498 5649
rect 10518 5629 10525 5649
rect 10475 5599 10525 5629
rect 11408 5609 11458 5625
rect 11616 5609 11666 5625
rect 11834 5609 11884 5625
rect 16569 5778 16619 5808
rect 16569 5758 16576 5778
rect 16596 5758 16619 5778
rect 16569 5731 16619 5758
rect 16777 5776 16827 5808
rect 16777 5756 16794 5776
rect 16814 5756 16827 5776
rect 16777 5731 16827 5756
rect 16995 5779 17045 5808
rect 20835 5824 20885 5840
rect 21043 5824 21093 5840
rect 21261 5824 21311 5840
rect 25199 5837 25249 5853
rect 25407 5837 25457 5853
rect 25625 5837 25675 5853
rect 29576 5849 29626 5865
rect 29784 5849 29834 5865
rect 30002 5849 30052 5865
rect 33940 5862 33990 5878
rect 34148 5862 34198 5878
rect 34366 5862 34416 5878
rect 16995 5759 17012 5779
rect 17032 5759 17045 5779
rect 16995 5731 17045 5759
rect 18679 5763 18729 5776
rect 18897 5763 18947 5776
rect 19105 5763 19155 5776
rect 14413 5661 14463 5689
rect 14413 5641 14426 5661
rect 14446 5641 14463 5661
rect 3093 5465 3143 5493
rect 411 5397 461 5425
rect 411 5377 424 5397
rect 444 5377 461 5397
rect 411 5348 461 5377
rect 629 5400 679 5425
rect 629 5380 642 5400
rect 662 5380 679 5400
rect 629 5348 679 5380
rect 837 5398 887 5425
rect 837 5378 860 5398
rect 880 5378 887 5398
rect 837 5348 887 5378
rect 5672 5529 5722 5545
rect 5890 5529 5940 5545
rect 6098 5529 6148 5545
rect 7031 5525 7081 5555
rect 7031 5505 7038 5525
rect 7058 5505 7081 5525
rect 7031 5478 7081 5505
rect 7239 5523 7289 5555
rect 7239 5503 7256 5523
rect 7276 5503 7289 5523
rect 7239 5478 7289 5503
rect 7457 5526 7507 5555
rect 7457 5506 7474 5526
rect 7494 5506 7507 5526
rect 9152 5550 9202 5563
rect 9370 5550 9420 5563
rect 9578 5550 9628 5563
rect 12205 5605 12255 5618
rect 12413 5605 12463 5618
rect 12631 5605 12681 5618
rect 14413 5612 14463 5641
rect 14631 5664 14681 5689
rect 14631 5644 14644 5664
rect 14664 5644 14681 5664
rect 14631 5612 14681 5644
rect 14839 5662 14889 5689
rect 14839 5642 14862 5662
rect 14882 5642 14889 5662
rect 14839 5612 14889 5642
rect 15772 5622 15822 5638
rect 15980 5622 16030 5638
rect 16198 5622 16248 5638
rect 20835 5752 20885 5782
rect 20835 5732 20842 5752
rect 20862 5732 20885 5752
rect 20835 5705 20885 5732
rect 21043 5750 21093 5782
rect 21043 5730 21060 5750
rect 21080 5730 21093 5750
rect 21043 5705 21093 5730
rect 21261 5753 21311 5782
rect 21261 5733 21278 5753
rect 21298 5733 21311 5753
rect 23043 5776 23093 5789
rect 23261 5776 23311 5789
rect 23469 5776 23519 5789
rect 21261 5705 21311 5733
rect 7457 5478 7507 5506
rect 3465 5400 3515 5416
rect 3673 5400 3723 5416
rect 3891 5400 3941 5416
rect 1209 5341 1259 5354
rect 1427 5341 1477 5354
rect 1635 5341 1685 5354
rect 2667 5352 2717 5365
rect 2875 5352 2925 5365
rect 3093 5352 3143 5365
rect 4775 5410 4825 5438
rect 411 5290 461 5306
rect 629 5290 679 5306
rect 837 5290 887 5306
rect 3465 5328 3515 5358
rect 3465 5308 3472 5328
rect 3492 5308 3515 5328
rect 3465 5281 3515 5308
rect 3673 5326 3723 5358
rect 3673 5306 3690 5326
rect 3710 5306 3723 5326
rect 3673 5281 3723 5306
rect 3891 5329 3941 5358
rect 3891 5309 3908 5329
rect 3928 5309 3941 5329
rect 4775 5390 4788 5410
rect 4808 5390 4825 5410
rect 4775 5361 4825 5390
rect 4993 5413 5043 5438
rect 4993 5393 5006 5413
rect 5026 5393 5043 5413
rect 4993 5361 5043 5393
rect 5201 5411 5251 5438
rect 5201 5391 5224 5411
rect 5244 5391 5251 5411
rect 5201 5361 5251 5391
rect 10049 5541 10099 5557
rect 10267 5541 10317 5557
rect 10475 5541 10525 5557
rect 11408 5537 11458 5567
rect 11408 5517 11415 5537
rect 11435 5517 11458 5537
rect 11408 5490 11458 5517
rect 11616 5535 11666 5567
rect 11616 5515 11633 5535
rect 11653 5515 11666 5535
rect 11616 5490 11666 5515
rect 11834 5538 11884 5567
rect 11834 5518 11851 5538
rect 11871 5518 11884 5538
rect 13516 5563 13566 5576
rect 13734 5563 13784 5576
rect 13942 5563 13992 5576
rect 16569 5618 16619 5631
rect 16777 5618 16827 5631
rect 16995 5618 17045 5631
rect 18679 5635 18729 5663
rect 18679 5615 18692 5635
rect 18712 5615 18729 5635
rect 18679 5586 18729 5615
rect 18897 5638 18947 5663
rect 18897 5618 18910 5638
rect 18930 5618 18947 5638
rect 18897 5586 18947 5618
rect 19105 5636 19155 5663
rect 19105 5616 19128 5636
rect 19148 5616 19155 5636
rect 19105 5586 19155 5616
rect 20038 5596 20088 5612
rect 20246 5596 20296 5612
rect 20464 5596 20514 5612
rect 25199 5765 25249 5795
rect 25199 5745 25206 5765
rect 25226 5745 25249 5765
rect 25199 5718 25249 5745
rect 25407 5763 25457 5795
rect 25407 5743 25424 5763
rect 25444 5743 25457 5763
rect 25407 5718 25457 5743
rect 25625 5766 25675 5795
rect 25625 5746 25642 5766
rect 25662 5746 25675 5766
rect 27420 5788 27470 5801
rect 27638 5788 27688 5801
rect 27846 5788 27896 5801
rect 25625 5718 25675 5746
rect 23043 5648 23093 5676
rect 23043 5628 23056 5648
rect 23076 5628 23093 5648
rect 11834 5490 11884 5518
rect 7829 5413 7879 5429
rect 8037 5413 8087 5429
rect 8255 5413 8305 5429
rect 3891 5281 3941 5309
rect 5573 5354 5623 5367
rect 5791 5354 5841 5367
rect 5999 5354 6049 5367
rect 7031 5365 7081 5378
rect 7239 5365 7289 5378
rect 7457 5365 7507 5378
rect 9152 5422 9202 5450
rect 4775 5303 4825 5319
rect 4993 5303 5043 5319
rect 5201 5303 5251 5319
rect 1209 5213 1259 5241
rect 1209 5193 1222 5213
rect 1242 5193 1259 5213
rect 1209 5164 1259 5193
rect 1427 5216 1477 5241
rect 1427 5196 1440 5216
rect 1460 5196 1477 5216
rect 1427 5164 1477 5196
rect 1635 5214 1685 5241
rect 1635 5194 1658 5214
rect 1678 5194 1685 5214
rect 1635 5164 1685 5194
rect 2363 5178 2413 5194
rect 2571 5178 2621 5194
rect 2789 5178 2839 5194
rect 7829 5341 7879 5371
rect 7829 5321 7836 5341
rect 7856 5321 7879 5341
rect 7829 5294 7879 5321
rect 8037 5339 8087 5371
rect 8037 5319 8054 5339
rect 8074 5319 8087 5339
rect 8037 5294 8087 5319
rect 8255 5342 8305 5371
rect 8255 5322 8272 5342
rect 8292 5322 8305 5342
rect 9152 5402 9165 5422
rect 9185 5402 9202 5422
rect 9152 5373 9202 5402
rect 9370 5425 9420 5450
rect 9370 5405 9383 5425
rect 9403 5405 9420 5425
rect 9370 5373 9420 5405
rect 9578 5423 9628 5450
rect 9578 5403 9601 5423
rect 9621 5403 9628 5423
rect 9578 5373 9628 5403
rect 14413 5554 14463 5570
rect 14631 5554 14681 5570
rect 14839 5554 14889 5570
rect 15772 5550 15822 5580
rect 15772 5530 15779 5550
rect 15799 5530 15822 5550
rect 15772 5503 15822 5530
rect 15980 5548 16030 5580
rect 15980 5528 15997 5548
rect 16017 5528 16030 5548
rect 15980 5503 16030 5528
rect 16198 5551 16248 5580
rect 16198 5531 16215 5551
rect 16235 5531 16248 5551
rect 16198 5503 16248 5531
rect 17782 5537 17832 5550
rect 18000 5537 18050 5550
rect 18208 5537 18258 5550
rect 20835 5592 20885 5605
rect 21043 5592 21093 5605
rect 21261 5592 21311 5605
rect 23043 5599 23093 5628
rect 23261 5651 23311 5676
rect 23261 5631 23274 5651
rect 23294 5631 23311 5651
rect 23261 5599 23311 5631
rect 23469 5649 23519 5676
rect 23469 5629 23492 5649
rect 23512 5629 23519 5649
rect 23469 5599 23519 5629
rect 24402 5609 24452 5625
rect 24610 5609 24660 5625
rect 24828 5609 24878 5625
rect 29576 5777 29626 5807
rect 29576 5757 29583 5777
rect 29603 5757 29626 5777
rect 29576 5730 29626 5757
rect 29784 5775 29834 5807
rect 29784 5755 29801 5775
rect 29821 5755 29834 5775
rect 29784 5730 29834 5755
rect 30002 5778 30052 5807
rect 30002 5758 30019 5778
rect 30039 5758 30052 5778
rect 31784 5801 31834 5814
rect 32002 5801 32052 5814
rect 32210 5801 32260 5814
rect 30002 5730 30052 5758
rect 27420 5660 27470 5688
rect 27420 5640 27433 5660
rect 27453 5640 27470 5660
rect 12206 5425 12256 5441
rect 12414 5425 12464 5441
rect 12632 5425 12682 5441
rect 8255 5294 8305 5322
rect 9950 5366 10000 5379
rect 10168 5366 10218 5379
rect 10376 5366 10426 5379
rect 11408 5377 11458 5390
rect 11616 5377 11666 5390
rect 11834 5377 11884 5390
rect 13516 5435 13566 5463
rect 9152 5315 9202 5331
rect 9370 5315 9420 5331
rect 9578 5315 9628 5331
rect 5573 5226 5623 5254
rect 412 5113 462 5126
rect 630 5113 680 5126
rect 838 5113 888 5126
rect 3465 5168 3515 5181
rect 3673 5168 3723 5181
rect 3891 5168 3941 5181
rect 5573 5206 5586 5226
rect 5606 5206 5623 5226
rect 5573 5177 5623 5206
rect 5791 5229 5841 5254
rect 5791 5209 5804 5229
rect 5824 5209 5841 5229
rect 5791 5177 5841 5209
rect 5999 5227 6049 5254
rect 5999 5207 6022 5227
rect 6042 5207 6049 5227
rect 5999 5177 6049 5207
rect 6727 5191 6777 5207
rect 6935 5191 6985 5207
rect 7153 5191 7203 5207
rect 12206 5353 12256 5383
rect 12206 5333 12213 5353
rect 12233 5333 12256 5353
rect 12206 5306 12256 5333
rect 12414 5351 12464 5383
rect 12414 5331 12431 5351
rect 12451 5331 12464 5351
rect 12414 5306 12464 5331
rect 12632 5354 12682 5383
rect 12632 5334 12649 5354
rect 12669 5334 12682 5354
rect 13516 5415 13529 5435
rect 13549 5415 13566 5435
rect 13516 5386 13566 5415
rect 13734 5438 13784 5463
rect 13734 5418 13747 5438
rect 13767 5418 13784 5438
rect 13734 5386 13784 5418
rect 13942 5436 13992 5463
rect 13942 5416 13965 5436
rect 13985 5416 13992 5436
rect 13942 5386 13992 5416
rect 16570 5438 16620 5454
rect 16778 5438 16828 5454
rect 16996 5438 17046 5454
rect 12632 5306 12682 5334
rect 14314 5379 14364 5392
rect 14532 5379 14582 5392
rect 14740 5379 14790 5392
rect 15772 5390 15822 5403
rect 15980 5390 16030 5403
rect 16198 5390 16248 5403
rect 18679 5528 18729 5544
rect 18897 5528 18947 5544
rect 19105 5528 19155 5544
rect 20038 5524 20088 5554
rect 20038 5504 20045 5524
rect 20065 5504 20088 5524
rect 20038 5477 20088 5504
rect 20246 5522 20296 5554
rect 20246 5502 20263 5522
rect 20283 5502 20296 5522
rect 20246 5477 20296 5502
rect 20464 5525 20514 5554
rect 20464 5505 20481 5525
rect 20501 5505 20514 5525
rect 22146 5550 22196 5563
rect 22364 5550 22414 5563
rect 22572 5550 22622 5563
rect 25199 5605 25249 5618
rect 25407 5605 25457 5618
rect 25625 5605 25675 5618
rect 27420 5611 27470 5640
rect 27638 5663 27688 5688
rect 27638 5643 27651 5663
rect 27671 5643 27688 5663
rect 27638 5611 27688 5643
rect 27846 5661 27896 5688
rect 27846 5641 27869 5661
rect 27889 5641 27896 5661
rect 27846 5611 27896 5641
rect 28779 5621 28829 5637
rect 28987 5621 29037 5637
rect 29205 5621 29255 5637
rect 33940 5790 33990 5820
rect 33940 5770 33947 5790
rect 33967 5770 33990 5790
rect 33940 5743 33990 5770
rect 34148 5788 34198 5820
rect 34148 5768 34165 5788
rect 34185 5768 34198 5788
rect 34148 5743 34198 5768
rect 34366 5791 34416 5820
rect 34366 5771 34383 5791
rect 34403 5771 34416 5791
rect 34366 5743 34416 5771
rect 31784 5673 31834 5701
rect 31784 5653 31797 5673
rect 31817 5653 31834 5673
rect 20464 5477 20514 5505
rect 13516 5328 13566 5344
rect 13734 5328 13784 5344
rect 13942 5328 13992 5344
rect 9950 5238 10000 5266
rect 1209 5106 1259 5122
rect 1427 5106 1477 5122
rect 1635 5106 1685 5122
rect 2363 5106 2413 5136
rect 2363 5086 2370 5106
rect 2390 5086 2413 5106
rect 2363 5059 2413 5086
rect 2571 5104 2621 5136
rect 2571 5084 2588 5104
rect 2608 5084 2621 5104
rect 2571 5059 2621 5084
rect 2789 5107 2839 5136
rect 4776 5126 4826 5139
rect 4994 5126 5044 5139
rect 5202 5126 5252 5139
rect 7829 5181 7879 5194
rect 8037 5181 8087 5194
rect 8255 5181 8305 5194
rect 9950 5218 9963 5238
rect 9983 5218 10000 5238
rect 9950 5189 10000 5218
rect 10168 5241 10218 5266
rect 10168 5221 10181 5241
rect 10201 5221 10218 5241
rect 10168 5189 10218 5221
rect 10376 5239 10426 5266
rect 10376 5219 10399 5239
rect 10419 5219 10426 5239
rect 10376 5189 10426 5219
rect 11104 5203 11154 5219
rect 11312 5203 11362 5219
rect 11530 5203 11580 5219
rect 16570 5366 16620 5396
rect 16570 5346 16577 5366
rect 16597 5346 16620 5366
rect 16570 5319 16620 5346
rect 16778 5364 16828 5396
rect 16778 5344 16795 5364
rect 16815 5344 16828 5364
rect 16778 5319 16828 5344
rect 16996 5367 17046 5396
rect 16996 5347 17013 5367
rect 17033 5347 17046 5367
rect 17782 5409 17832 5437
rect 16996 5319 17046 5347
rect 17782 5389 17795 5409
rect 17815 5389 17832 5409
rect 17782 5360 17832 5389
rect 18000 5412 18050 5437
rect 18000 5392 18013 5412
rect 18033 5392 18050 5412
rect 18000 5360 18050 5392
rect 18208 5410 18258 5437
rect 18208 5390 18231 5410
rect 18251 5390 18258 5410
rect 18208 5360 18258 5390
rect 23043 5541 23093 5557
rect 23261 5541 23311 5557
rect 23469 5541 23519 5557
rect 24402 5537 24452 5567
rect 24402 5517 24409 5537
rect 24429 5517 24452 5537
rect 24402 5490 24452 5517
rect 24610 5535 24660 5567
rect 24610 5515 24627 5535
rect 24647 5515 24660 5535
rect 24610 5490 24660 5515
rect 24828 5538 24878 5567
rect 24828 5518 24845 5538
rect 24865 5518 24878 5538
rect 26523 5562 26573 5575
rect 26741 5562 26791 5575
rect 26949 5562 26999 5575
rect 29576 5617 29626 5630
rect 29784 5617 29834 5630
rect 30002 5617 30052 5630
rect 31784 5624 31834 5653
rect 32002 5676 32052 5701
rect 32002 5656 32015 5676
rect 32035 5656 32052 5676
rect 32002 5624 32052 5656
rect 32210 5674 32260 5701
rect 32210 5654 32233 5674
rect 32253 5654 32260 5674
rect 32210 5624 32260 5654
rect 33143 5634 33193 5650
rect 33351 5634 33401 5650
rect 33569 5634 33619 5650
rect 24828 5490 24878 5518
rect 20836 5412 20886 5428
rect 21044 5412 21094 5428
rect 21262 5412 21312 5428
rect 14314 5251 14364 5279
rect 2789 5087 2806 5107
rect 2826 5087 2839 5107
rect 2789 5059 2839 5087
rect 412 4985 462 5013
rect 412 4965 425 4985
rect 445 4965 462 4985
rect 412 4936 462 4965
rect 630 4988 680 5013
rect 630 4968 643 4988
rect 663 4968 680 4988
rect 630 4936 680 4968
rect 838 4986 888 5013
rect 838 4966 861 4986
rect 881 4966 888 4986
rect 838 4936 888 4966
rect 5573 5119 5623 5135
rect 5791 5119 5841 5135
rect 5999 5119 6049 5135
rect 6727 5119 6777 5149
rect 6727 5099 6734 5119
rect 6754 5099 6777 5119
rect 6727 5072 6777 5099
rect 6935 5117 6985 5149
rect 6935 5097 6952 5117
rect 6972 5097 6985 5117
rect 6935 5072 6985 5097
rect 7153 5120 7203 5149
rect 9153 5138 9203 5151
rect 9371 5138 9421 5151
rect 9579 5138 9629 5151
rect 12206 5193 12256 5206
rect 12414 5193 12464 5206
rect 12632 5193 12682 5206
rect 14314 5231 14327 5251
rect 14347 5231 14364 5251
rect 14314 5202 14364 5231
rect 14532 5254 14582 5279
rect 14532 5234 14545 5254
rect 14565 5234 14582 5254
rect 14532 5202 14582 5234
rect 14740 5252 14790 5279
rect 14740 5232 14763 5252
rect 14783 5232 14790 5252
rect 14740 5202 14790 5232
rect 15468 5216 15518 5232
rect 15676 5216 15726 5232
rect 15894 5216 15944 5232
rect 18580 5353 18630 5366
rect 18798 5353 18848 5366
rect 19006 5353 19056 5366
rect 20038 5364 20088 5377
rect 20246 5364 20296 5377
rect 20464 5364 20514 5377
rect 22146 5422 22196 5450
rect 17782 5302 17832 5318
rect 18000 5302 18050 5318
rect 18208 5302 18258 5318
rect 20836 5340 20886 5370
rect 20836 5320 20843 5340
rect 20863 5320 20886 5340
rect 20836 5293 20886 5320
rect 21044 5338 21094 5370
rect 21044 5318 21061 5338
rect 21081 5318 21094 5338
rect 21044 5293 21094 5318
rect 21262 5341 21312 5370
rect 21262 5321 21279 5341
rect 21299 5321 21312 5341
rect 22146 5402 22159 5422
rect 22179 5402 22196 5422
rect 22146 5373 22196 5402
rect 22364 5425 22414 5450
rect 22364 5405 22377 5425
rect 22397 5405 22414 5425
rect 22364 5373 22414 5405
rect 22572 5423 22622 5450
rect 22572 5403 22595 5423
rect 22615 5403 22622 5423
rect 22572 5373 22622 5403
rect 27420 5553 27470 5569
rect 27638 5553 27688 5569
rect 27846 5553 27896 5569
rect 28779 5549 28829 5579
rect 28779 5529 28786 5549
rect 28806 5529 28829 5549
rect 28779 5502 28829 5529
rect 28987 5547 29037 5579
rect 28987 5527 29004 5547
rect 29024 5527 29037 5547
rect 28987 5502 29037 5527
rect 29205 5550 29255 5579
rect 29205 5530 29222 5550
rect 29242 5530 29255 5550
rect 30887 5575 30937 5588
rect 31105 5575 31155 5588
rect 31313 5575 31363 5588
rect 33940 5630 33990 5643
rect 34148 5630 34198 5643
rect 34366 5630 34416 5643
rect 29205 5502 29255 5530
rect 25200 5425 25250 5441
rect 25408 5425 25458 5441
rect 25626 5425 25676 5441
rect 21262 5293 21312 5321
rect 22944 5366 22994 5379
rect 23162 5366 23212 5379
rect 23370 5366 23420 5379
rect 24402 5377 24452 5390
rect 24610 5377 24660 5390
rect 24828 5377 24878 5390
rect 26523 5434 26573 5462
rect 22146 5315 22196 5331
rect 22364 5315 22414 5331
rect 22572 5315 22622 5331
rect 7153 5100 7170 5120
rect 7190 5100 7203 5120
rect 7153 5072 7203 5100
rect 4776 4998 4826 5026
rect 2363 4946 2413 4959
rect 2571 4946 2621 4959
rect 2789 4946 2839 4959
rect 4776 4978 4789 4998
rect 4809 4978 4826 4998
rect 4776 4949 4826 4978
rect 4994 5001 5044 5026
rect 4994 4981 5007 5001
rect 5027 4981 5044 5001
rect 4994 4949 5044 4981
rect 5202 4999 5252 5026
rect 5202 4979 5225 4999
rect 5245 4979 5252 4999
rect 5202 4949 5252 4979
rect 9950 5131 10000 5147
rect 10168 5131 10218 5147
rect 10376 5131 10426 5147
rect 11104 5131 11154 5161
rect 11104 5111 11111 5131
rect 11131 5111 11154 5131
rect 11104 5084 11154 5111
rect 11312 5129 11362 5161
rect 11312 5109 11329 5129
rect 11349 5109 11362 5129
rect 11312 5084 11362 5109
rect 11530 5132 11580 5161
rect 13517 5151 13567 5164
rect 13735 5151 13785 5164
rect 13943 5151 13993 5164
rect 16570 5206 16620 5219
rect 16778 5206 16828 5219
rect 16996 5206 17046 5219
rect 18580 5225 18630 5253
rect 11530 5112 11547 5132
rect 11567 5112 11580 5132
rect 11530 5084 11580 5112
rect 9153 5010 9203 5038
rect 6727 4959 6777 4972
rect 6935 4959 6985 4972
rect 7153 4959 7203 4972
rect 9153 4990 9166 5010
rect 9186 4990 9203 5010
rect 9153 4961 9203 4990
rect 9371 5013 9421 5038
rect 9371 4993 9384 5013
rect 9404 4993 9421 5013
rect 9371 4961 9421 4993
rect 9579 5011 9629 5038
rect 9579 4991 9602 5011
rect 9622 4991 9629 5011
rect 9579 4961 9629 4991
rect 14314 5144 14364 5160
rect 14532 5144 14582 5160
rect 14740 5144 14790 5160
rect 15468 5144 15518 5174
rect 15468 5124 15475 5144
rect 15495 5124 15518 5144
rect 15468 5097 15518 5124
rect 15676 5142 15726 5174
rect 15676 5122 15693 5142
rect 15713 5122 15726 5142
rect 15676 5097 15726 5122
rect 15894 5145 15944 5174
rect 15894 5125 15911 5145
rect 15931 5125 15944 5145
rect 18580 5205 18593 5225
rect 18613 5205 18630 5225
rect 18580 5176 18630 5205
rect 18798 5228 18848 5253
rect 18798 5208 18811 5228
rect 18831 5208 18848 5228
rect 18798 5176 18848 5208
rect 19006 5226 19056 5253
rect 19006 5206 19029 5226
rect 19049 5206 19056 5226
rect 19006 5176 19056 5206
rect 19734 5190 19784 5206
rect 19942 5190 19992 5206
rect 20160 5190 20210 5206
rect 25200 5353 25250 5383
rect 25200 5333 25207 5353
rect 25227 5333 25250 5353
rect 25200 5306 25250 5333
rect 25408 5351 25458 5383
rect 25408 5331 25425 5351
rect 25445 5331 25458 5351
rect 25408 5306 25458 5331
rect 25626 5354 25676 5383
rect 25626 5334 25643 5354
rect 25663 5334 25676 5354
rect 26523 5414 26536 5434
rect 26556 5414 26573 5434
rect 26523 5385 26573 5414
rect 26741 5437 26791 5462
rect 26741 5417 26754 5437
rect 26774 5417 26791 5437
rect 26741 5385 26791 5417
rect 26949 5435 26999 5462
rect 26949 5415 26972 5435
rect 26992 5415 26999 5435
rect 26949 5385 26999 5415
rect 31784 5566 31834 5582
rect 32002 5566 32052 5582
rect 32210 5566 32260 5582
rect 33143 5562 33193 5592
rect 33143 5542 33150 5562
rect 33170 5542 33193 5562
rect 33143 5515 33193 5542
rect 33351 5560 33401 5592
rect 33351 5540 33368 5560
rect 33388 5540 33401 5560
rect 33351 5515 33401 5540
rect 33569 5563 33619 5592
rect 33569 5543 33586 5563
rect 33606 5543 33619 5563
rect 33569 5515 33619 5543
rect 29577 5437 29627 5453
rect 29785 5437 29835 5453
rect 30003 5437 30053 5453
rect 25626 5306 25676 5334
rect 27321 5378 27371 5391
rect 27539 5378 27589 5391
rect 27747 5378 27797 5391
rect 28779 5389 28829 5402
rect 28987 5389 29037 5402
rect 29205 5389 29255 5402
rect 30887 5447 30937 5475
rect 26523 5327 26573 5343
rect 26741 5327 26791 5343
rect 26949 5327 26999 5343
rect 22944 5238 22994 5266
rect 15894 5097 15944 5125
rect 17783 5125 17833 5138
rect 18001 5125 18051 5138
rect 18209 5125 18259 5138
rect 20836 5180 20886 5193
rect 21044 5180 21094 5193
rect 21262 5180 21312 5193
rect 22944 5218 22957 5238
rect 22977 5218 22994 5238
rect 22944 5189 22994 5218
rect 23162 5241 23212 5266
rect 23162 5221 23175 5241
rect 23195 5221 23212 5241
rect 23162 5189 23212 5221
rect 23370 5239 23420 5266
rect 23370 5219 23393 5239
rect 23413 5219 23420 5239
rect 23370 5189 23420 5219
rect 24098 5203 24148 5219
rect 24306 5203 24356 5219
rect 24524 5203 24574 5219
rect 29577 5365 29627 5395
rect 29577 5345 29584 5365
rect 29604 5345 29627 5365
rect 29577 5318 29627 5345
rect 29785 5363 29835 5395
rect 29785 5343 29802 5363
rect 29822 5343 29835 5363
rect 29785 5318 29835 5343
rect 30003 5366 30053 5395
rect 30003 5346 30020 5366
rect 30040 5346 30053 5366
rect 30887 5427 30900 5447
rect 30920 5427 30937 5447
rect 30887 5398 30937 5427
rect 31105 5450 31155 5475
rect 31105 5430 31118 5450
rect 31138 5430 31155 5450
rect 31105 5398 31155 5430
rect 31313 5448 31363 5475
rect 31313 5428 31336 5448
rect 31356 5428 31363 5448
rect 31313 5398 31363 5428
rect 33941 5450 33991 5466
rect 34149 5450 34199 5466
rect 34367 5450 34417 5466
rect 30003 5318 30053 5346
rect 31685 5391 31735 5404
rect 31903 5391 31953 5404
rect 32111 5391 32161 5404
rect 33143 5402 33193 5415
rect 33351 5402 33401 5415
rect 33569 5402 33619 5415
rect 30887 5340 30937 5356
rect 31105 5340 31155 5356
rect 31313 5340 31363 5356
rect 27321 5250 27371 5278
rect 13517 5023 13567 5051
rect 11104 4971 11154 4984
rect 11312 4971 11362 4984
rect 11530 4971 11580 4984
rect 13517 5003 13530 5023
rect 13550 5003 13567 5023
rect 13517 4974 13567 5003
rect 13735 5026 13785 5051
rect 13735 5006 13748 5026
rect 13768 5006 13785 5026
rect 13735 4974 13785 5006
rect 13943 5024 13993 5051
rect 13943 5004 13966 5024
rect 13986 5004 13993 5024
rect 13943 4974 13993 5004
rect 18580 5118 18630 5134
rect 18798 5118 18848 5134
rect 19006 5118 19056 5134
rect 19734 5118 19784 5148
rect 19734 5098 19741 5118
rect 19761 5098 19784 5118
rect 19734 5071 19784 5098
rect 19942 5116 19992 5148
rect 19942 5096 19959 5116
rect 19979 5096 19992 5116
rect 19942 5071 19992 5096
rect 20160 5119 20210 5148
rect 22147 5138 22197 5151
rect 22365 5138 22415 5151
rect 22573 5138 22623 5151
rect 25200 5193 25250 5206
rect 25408 5193 25458 5206
rect 25626 5193 25676 5206
rect 27321 5230 27334 5250
rect 27354 5230 27371 5250
rect 27321 5201 27371 5230
rect 27539 5253 27589 5278
rect 27539 5233 27552 5253
rect 27572 5233 27589 5253
rect 27539 5201 27589 5233
rect 27747 5251 27797 5278
rect 27747 5231 27770 5251
rect 27790 5231 27797 5251
rect 27747 5201 27797 5231
rect 28475 5215 28525 5231
rect 28683 5215 28733 5231
rect 28901 5215 28951 5231
rect 33941 5378 33991 5408
rect 33941 5358 33948 5378
rect 33968 5358 33991 5378
rect 33941 5331 33991 5358
rect 34149 5376 34199 5408
rect 34149 5356 34166 5376
rect 34186 5356 34199 5376
rect 34149 5331 34199 5356
rect 34367 5379 34417 5408
rect 34367 5359 34384 5379
rect 34404 5359 34417 5379
rect 34367 5331 34417 5359
rect 31685 5263 31735 5291
rect 20160 5099 20177 5119
rect 20197 5099 20210 5119
rect 20160 5071 20210 5099
rect 15468 4984 15518 4997
rect 15676 4984 15726 4997
rect 15894 4984 15944 4997
rect 17783 4997 17833 5025
rect 17783 4977 17796 4997
rect 17816 4977 17833 4997
rect 412 4878 462 4894
rect 630 4878 680 4894
rect 838 4878 888 4894
rect 4776 4891 4826 4907
rect 4994 4891 5044 4907
rect 5202 4891 5252 4907
rect 9153 4903 9203 4919
rect 9371 4903 9421 4919
rect 9579 4903 9629 4919
rect 13517 4916 13567 4932
rect 13735 4916 13785 4932
rect 13943 4916 13993 4932
rect 17783 4948 17833 4977
rect 18001 5000 18051 5025
rect 18001 4980 18014 5000
rect 18034 4980 18051 5000
rect 18001 4948 18051 4980
rect 18209 4998 18259 5025
rect 18209 4978 18232 4998
rect 18252 4978 18259 4998
rect 18209 4948 18259 4978
rect 22944 5131 22994 5147
rect 23162 5131 23212 5147
rect 23370 5131 23420 5147
rect 24098 5131 24148 5161
rect 24098 5111 24105 5131
rect 24125 5111 24148 5131
rect 24098 5084 24148 5111
rect 24306 5129 24356 5161
rect 24306 5109 24323 5129
rect 24343 5109 24356 5129
rect 24306 5084 24356 5109
rect 24524 5132 24574 5161
rect 26524 5150 26574 5163
rect 26742 5150 26792 5163
rect 26950 5150 27000 5163
rect 29577 5205 29627 5218
rect 29785 5205 29835 5218
rect 30003 5205 30053 5218
rect 31685 5243 31698 5263
rect 31718 5243 31735 5263
rect 31685 5214 31735 5243
rect 31903 5266 31953 5291
rect 31903 5246 31916 5266
rect 31936 5246 31953 5266
rect 31903 5214 31953 5246
rect 32111 5264 32161 5291
rect 32111 5244 32134 5264
rect 32154 5244 32161 5264
rect 32111 5214 32161 5244
rect 32839 5228 32889 5244
rect 33047 5228 33097 5244
rect 33265 5228 33315 5244
rect 24524 5112 24541 5132
rect 24561 5112 24574 5132
rect 24524 5084 24574 5112
rect 22147 5010 22197 5038
rect 19734 4958 19784 4971
rect 19942 4958 19992 4971
rect 20160 4958 20210 4971
rect 22147 4990 22160 5010
rect 22180 4990 22197 5010
rect 22147 4961 22197 4990
rect 22365 5013 22415 5038
rect 22365 4993 22378 5013
rect 22398 4993 22415 5013
rect 22365 4961 22415 4993
rect 22573 5011 22623 5038
rect 22573 4991 22596 5011
rect 22616 4991 22623 5011
rect 22573 4961 22623 4991
rect 27321 5143 27371 5159
rect 27539 5143 27589 5159
rect 27747 5143 27797 5159
rect 28475 5143 28525 5173
rect 28475 5123 28482 5143
rect 28502 5123 28525 5143
rect 28475 5096 28525 5123
rect 28683 5141 28733 5173
rect 28683 5121 28700 5141
rect 28720 5121 28733 5141
rect 28683 5096 28733 5121
rect 28901 5144 28951 5173
rect 30888 5163 30938 5176
rect 31106 5163 31156 5176
rect 31314 5163 31364 5176
rect 33941 5218 33991 5231
rect 34149 5218 34199 5231
rect 34367 5218 34417 5231
rect 28901 5124 28918 5144
rect 28938 5124 28951 5144
rect 28901 5096 28951 5124
rect 26524 5022 26574 5050
rect 24098 4971 24148 4984
rect 24306 4971 24356 4984
rect 24524 4971 24574 4984
rect 26524 5002 26537 5022
rect 26557 5002 26574 5022
rect 26524 4973 26574 5002
rect 26742 5025 26792 5050
rect 26742 5005 26755 5025
rect 26775 5005 26792 5025
rect 26742 4973 26792 5005
rect 26950 5023 27000 5050
rect 26950 5003 26973 5023
rect 26993 5003 27000 5023
rect 26950 4973 27000 5003
rect 31685 5156 31735 5172
rect 31903 5156 31953 5172
rect 32111 5156 32161 5172
rect 32839 5156 32889 5186
rect 32839 5136 32846 5156
rect 32866 5136 32889 5156
rect 32839 5109 32889 5136
rect 33047 5154 33097 5186
rect 33047 5134 33064 5154
rect 33084 5134 33097 5154
rect 33047 5109 33097 5134
rect 33265 5157 33315 5186
rect 33265 5137 33282 5157
rect 33302 5137 33315 5157
rect 33265 5109 33315 5137
rect 30888 5035 30938 5063
rect 28475 4983 28525 4996
rect 28683 4983 28733 4996
rect 28901 4983 28951 4996
rect 30888 5015 30901 5035
rect 30921 5015 30938 5035
rect 30888 4986 30938 5015
rect 31106 5038 31156 5063
rect 31106 5018 31119 5038
rect 31139 5018 31156 5038
rect 31106 4986 31156 5018
rect 31314 5036 31364 5063
rect 31314 5016 31337 5036
rect 31357 5016 31364 5036
rect 31314 4986 31364 5016
rect 32839 4996 32889 5009
rect 33047 4996 33097 5009
rect 33265 4996 33315 5009
rect 17783 4890 17833 4906
rect 18001 4890 18051 4906
rect 18209 4890 18259 4906
rect 22147 4903 22197 4919
rect 22365 4903 22415 4919
rect 22573 4903 22623 4919
rect 26524 4915 26574 4931
rect 26742 4915 26792 4931
rect 26950 4915 27000 4931
rect 30888 4928 30938 4944
rect 31106 4928 31156 4944
rect 31314 4928 31364 4944
rect 3445 4794 3495 4810
rect 3653 4794 3703 4810
rect 3871 4794 3921 4810
rect 7809 4807 7859 4823
rect 8017 4807 8067 4823
rect 8235 4807 8285 4823
rect 12186 4819 12236 4835
rect 12394 4819 12444 4835
rect 12612 4819 12662 4835
rect 16550 4832 16600 4848
rect 16758 4832 16808 4848
rect 16976 4832 17026 4848
rect 1494 4729 1544 4742
rect 1712 4729 1762 4742
rect 1920 4729 1970 4742
rect 3445 4722 3495 4752
rect 3445 4702 3452 4722
rect 3472 4702 3495 4722
rect 3445 4675 3495 4702
rect 3653 4720 3703 4752
rect 3653 4700 3670 4720
rect 3690 4700 3703 4720
rect 3653 4675 3703 4700
rect 3871 4723 3921 4752
rect 3871 4703 3888 4723
rect 3908 4703 3921 4723
rect 5858 4742 5908 4755
rect 6076 4742 6126 4755
rect 6284 4742 6334 4755
rect 3871 4675 3921 4703
rect 1494 4601 1544 4629
rect 1494 4581 1507 4601
rect 1527 4581 1544 4601
rect 1494 4552 1544 4581
rect 1712 4604 1762 4629
rect 1712 4584 1725 4604
rect 1745 4584 1762 4604
rect 1712 4552 1762 4584
rect 1920 4602 1970 4629
rect 1920 4582 1943 4602
rect 1963 4582 1970 4602
rect 1920 4552 1970 4582
rect 2648 4566 2698 4582
rect 2856 4566 2906 4582
rect 3074 4566 3124 4582
rect 7809 4735 7859 4765
rect 7809 4715 7816 4735
rect 7836 4715 7859 4735
rect 7809 4688 7859 4715
rect 8017 4733 8067 4765
rect 8017 4713 8034 4733
rect 8054 4713 8067 4733
rect 8017 4688 8067 4713
rect 8235 4736 8285 4765
rect 8235 4716 8252 4736
rect 8272 4716 8285 4736
rect 10235 4754 10285 4767
rect 10453 4754 10503 4767
rect 10661 4754 10711 4767
rect 8235 4688 8285 4716
rect 5858 4614 5908 4642
rect 5858 4594 5871 4614
rect 5891 4594 5908 4614
rect 392 4507 442 4520
rect 610 4507 660 4520
rect 818 4507 868 4520
rect 3445 4562 3495 4575
rect 3653 4562 3703 4575
rect 3871 4562 3921 4575
rect 5858 4565 5908 4594
rect 6076 4617 6126 4642
rect 6076 4597 6089 4617
rect 6109 4597 6126 4617
rect 6076 4565 6126 4597
rect 6284 4615 6334 4642
rect 6284 4595 6307 4615
rect 6327 4595 6334 4615
rect 6284 4565 6334 4595
rect 7012 4579 7062 4595
rect 7220 4579 7270 4595
rect 7438 4579 7488 4595
rect 12186 4747 12236 4777
rect 12186 4727 12193 4747
rect 12213 4727 12236 4747
rect 12186 4700 12236 4727
rect 12394 4745 12444 4777
rect 12394 4725 12411 4745
rect 12431 4725 12444 4745
rect 12394 4700 12444 4725
rect 12612 4748 12662 4777
rect 12612 4728 12629 4748
rect 12649 4728 12662 4748
rect 14599 4767 14649 4780
rect 14817 4767 14867 4780
rect 15025 4767 15075 4780
rect 12612 4700 12662 4728
rect 10235 4626 10285 4654
rect 10235 4606 10248 4626
rect 10268 4606 10285 4626
rect 1494 4494 1544 4510
rect 1712 4494 1762 4510
rect 1920 4494 1970 4510
rect 2648 4494 2698 4524
rect 2648 4474 2655 4494
rect 2675 4474 2698 4494
rect 2648 4447 2698 4474
rect 2856 4492 2906 4524
rect 2856 4472 2873 4492
rect 2893 4472 2906 4492
rect 2856 4447 2906 4472
rect 3074 4495 3124 4524
rect 3074 4475 3091 4495
rect 3111 4475 3124 4495
rect 4756 4520 4806 4533
rect 4974 4520 5024 4533
rect 5182 4520 5232 4533
rect 7809 4575 7859 4588
rect 8017 4575 8067 4588
rect 8235 4575 8285 4588
rect 10235 4577 10285 4606
rect 10453 4629 10503 4654
rect 10453 4609 10466 4629
rect 10486 4609 10503 4629
rect 10453 4577 10503 4609
rect 10661 4627 10711 4654
rect 10661 4607 10684 4627
rect 10704 4607 10711 4627
rect 10661 4577 10711 4607
rect 11389 4591 11439 4607
rect 11597 4591 11647 4607
rect 11815 4591 11865 4607
rect 16550 4760 16600 4790
rect 16550 4740 16557 4760
rect 16577 4740 16600 4760
rect 16550 4713 16600 4740
rect 16758 4758 16808 4790
rect 16758 4738 16775 4758
rect 16795 4738 16808 4758
rect 16758 4713 16808 4738
rect 16976 4761 17026 4790
rect 20816 4806 20866 4822
rect 21024 4806 21074 4822
rect 21242 4806 21292 4822
rect 25180 4819 25230 4835
rect 25388 4819 25438 4835
rect 25606 4819 25656 4835
rect 29557 4831 29607 4847
rect 29765 4831 29815 4847
rect 29983 4831 30033 4847
rect 33921 4844 33971 4860
rect 34129 4844 34179 4860
rect 34347 4844 34397 4860
rect 16976 4741 16993 4761
rect 17013 4741 17026 4761
rect 16976 4713 17026 4741
rect 18865 4741 18915 4754
rect 19083 4741 19133 4754
rect 19291 4741 19341 4754
rect 14599 4639 14649 4667
rect 14599 4619 14612 4639
rect 14632 4619 14649 4639
rect 3074 4447 3124 4475
rect 392 4379 442 4407
rect 392 4359 405 4379
rect 425 4359 442 4379
rect 392 4330 442 4359
rect 610 4382 660 4407
rect 610 4362 623 4382
rect 643 4362 660 4382
rect 610 4330 660 4362
rect 818 4380 868 4407
rect 818 4360 841 4380
rect 861 4360 868 4380
rect 818 4330 868 4360
rect 5858 4507 5908 4523
rect 6076 4507 6126 4523
rect 6284 4507 6334 4523
rect 7012 4507 7062 4537
rect 7012 4487 7019 4507
rect 7039 4487 7062 4507
rect 7012 4460 7062 4487
rect 7220 4505 7270 4537
rect 7220 4485 7237 4505
rect 7257 4485 7270 4505
rect 7220 4460 7270 4485
rect 7438 4508 7488 4537
rect 7438 4488 7455 4508
rect 7475 4488 7488 4508
rect 9133 4532 9183 4545
rect 9351 4532 9401 4545
rect 9559 4532 9609 4545
rect 12186 4587 12236 4600
rect 12394 4587 12444 4600
rect 12612 4587 12662 4600
rect 14599 4590 14649 4619
rect 14817 4642 14867 4667
rect 14817 4622 14830 4642
rect 14850 4622 14867 4642
rect 14817 4590 14867 4622
rect 15025 4640 15075 4667
rect 15025 4620 15048 4640
rect 15068 4620 15075 4640
rect 15025 4590 15075 4620
rect 15753 4604 15803 4620
rect 15961 4604 16011 4620
rect 16179 4604 16229 4620
rect 20816 4734 20866 4764
rect 20816 4714 20823 4734
rect 20843 4714 20866 4734
rect 20816 4687 20866 4714
rect 21024 4732 21074 4764
rect 21024 4712 21041 4732
rect 21061 4712 21074 4732
rect 21024 4687 21074 4712
rect 21242 4735 21292 4764
rect 21242 4715 21259 4735
rect 21279 4715 21292 4735
rect 23229 4754 23279 4767
rect 23447 4754 23497 4767
rect 23655 4754 23705 4767
rect 21242 4687 21292 4715
rect 7438 4460 7488 4488
rect 3446 4382 3496 4398
rect 3654 4382 3704 4398
rect 3872 4382 3922 4398
rect 1190 4323 1240 4336
rect 1408 4323 1458 4336
rect 1616 4323 1666 4336
rect 2648 4334 2698 4347
rect 2856 4334 2906 4347
rect 3074 4334 3124 4347
rect 4756 4392 4806 4420
rect 392 4272 442 4288
rect 610 4272 660 4288
rect 818 4272 868 4288
rect 3446 4310 3496 4340
rect 3446 4290 3453 4310
rect 3473 4290 3496 4310
rect 3446 4263 3496 4290
rect 3654 4308 3704 4340
rect 3654 4288 3671 4308
rect 3691 4288 3704 4308
rect 3654 4263 3704 4288
rect 3872 4311 3922 4340
rect 3872 4291 3889 4311
rect 3909 4291 3922 4311
rect 4756 4372 4769 4392
rect 4789 4372 4806 4392
rect 4756 4343 4806 4372
rect 4974 4395 5024 4420
rect 4974 4375 4987 4395
rect 5007 4375 5024 4395
rect 4974 4343 5024 4375
rect 5182 4393 5232 4420
rect 5182 4373 5205 4393
rect 5225 4373 5232 4393
rect 5182 4343 5232 4373
rect 10235 4519 10285 4535
rect 10453 4519 10503 4535
rect 10661 4519 10711 4535
rect 11389 4519 11439 4549
rect 11389 4499 11396 4519
rect 11416 4499 11439 4519
rect 11389 4472 11439 4499
rect 11597 4517 11647 4549
rect 11597 4497 11614 4517
rect 11634 4497 11647 4517
rect 11597 4472 11647 4497
rect 11815 4520 11865 4549
rect 11815 4500 11832 4520
rect 11852 4500 11865 4520
rect 13497 4545 13547 4558
rect 13715 4545 13765 4558
rect 13923 4545 13973 4558
rect 16550 4600 16600 4613
rect 16758 4600 16808 4613
rect 16976 4600 17026 4613
rect 18865 4613 18915 4641
rect 11815 4472 11865 4500
rect 7810 4395 7860 4411
rect 8018 4395 8068 4411
rect 8236 4395 8286 4411
rect 3872 4263 3922 4291
rect 5554 4336 5604 4349
rect 5772 4336 5822 4349
rect 5980 4336 6030 4349
rect 7012 4347 7062 4360
rect 7220 4347 7270 4360
rect 7438 4347 7488 4360
rect 9133 4404 9183 4432
rect 4756 4285 4806 4301
rect 4974 4285 5024 4301
rect 5182 4285 5232 4301
rect 1190 4195 1240 4223
rect 1190 4175 1203 4195
rect 1223 4175 1240 4195
rect 1190 4146 1240 4175
rect 1408 4198 1458 4223
rect 1408 4178 1421 4198
rect 1441 4178 1458 4198
rect 1408 4146 1458 4178
rect 1616 4196 1666 4223
rect 1616 4176 1639 4196
rect 1659 4176 1666 4196
rect 1616 4146 1666 4176
rect 2549 4156 2599 4172
rect 2757 4156 2807 4172
rect 2975 4156 3025 4172
rect 7810 4323 7860 4353
rect 7810 4303 7817 4323
rect 7837 4303 7860 4323
rect 7810 4276 7860 4303
rect 8018 4321 8068 4353
rect 8018 4301 8035 4321
rect 8055 4301 8068 4321
rect 8018 4276 8068 4301
rect 8236 4324 8286 4353
rect 8236 4304 8253 4324
rect 8273 4304 8286 4324
rect 9133 4384 9146 4404
rect 9166 4384 9183 4404
rect 9133 4355 9183 4384
rect 9351 4407 9401 4432
rect 9351 4387 9364 4407
rect 9384 4387 9401 4407
rect 9351 4355 9401 4387
rect 9559 4405 9609 4432
rect 9559 4385 9582 4405
rect 9602 4385 9609 4405
rect 9559 4355 9609 4385
rect 14599 4532 14649 4548
rect 14817 4532 14867 4548
rect 15025 4532 15075 4548
rect 15753 4532 15803 4562
rect 15753 4512 15760 4532
rect 15780 4512 15803 4532
rect 15753 4485 15803 4512
rect 15961 4530 16011 4562
rect 15961 4510 15978 4530
rect 15998 4510 16011 4530
rect 15961 4485 16011 4510
rect 16179 4533 16229 4562
rect 16179 4513 16196 4533
rect 16216 4513 16229 4533
rect 18865 4593 18878 4613
rect 18898 4593 18915 4613
rect 18865 4564 18915 4593
rect 19083 4616 19133 4641
rect 19083 4596 19096 4616
rect 19116 4596 19133 4616
rect 19083 4564 19133 4596
rect 19291 4614 19341 4641
rect 19291 4594 19314 4614
rect 19334 4594 19341 4614
rect 19291 4564 19341 4594
rect 20019 4578 20069 4594
rect 20227 4578 20277 4594
rect 20445 4578 20495 4594
rect 25180 4747 25230 4777
rect 25180 4727 25187 4747
rect 25207 4727 25230 4747
rect 25180 4700 25230 4727
rect 25388 4745 25438 4777
rect 25388 4725 25405 4745
rect 25425 4725 25438 4745
rect 25388 4700 25438 4725
rect 25606 4748 25656 4777
rect 25606 4728 25623 4748
rect 25643 4728 25656 4748
rect 27606 4766 27656 4779
rect 27824 4766 27874 4779
rect 28032 4766 28082 4779
rect 25606 4700 25656 4728
rect 23229 4626 23279 4654
rect 23229 4606 23242 4626
rect 23262 4606 23279 4626
rect 16179 4485 16229 4513
rect 17763 4519 17813 4532
rect 17981 4519 18031 4532
rect 18189 4519 18239 4532
rect 20816 4574 20866 4587
rect 21024 4574 21074 4587
rect 21242 4574 21292 4587
rect 23229 4577 23279 4606
rect 23447 4629 23497 4654
rect 23447 4609 23460 4629
rect 23480 4609 23497 4629
rect 23447 4577 23497 4609
rect 23655 4627 23705 4654
rect 23655 4607 23678 4627
rect 23698 4607 23705 4627
rect 23655 4577 23705 4607
rect 24383 4591 24433 4607
rect 24591 4591 24641 4607
rect 24809 4591 24859 4607
rect 29557 4759 29607 4789
rect 29557 4739 29564 4759
rect 29584 4739 29607 4759
rect 29557 4712 29607 4739
rect 29765 4757 29815 4789
rect 29765 4737 29782 4757
rect 29802 4737 29815 4757
rect 29765 4712 29815 4737
rect 29983 4760 30033 4789
rect 29983 4740 30000 4760
rect 30020 4740 30033 4760
rect 31970 4779 32020 4792
rect 32188 4779 32238 4792
rect 32396 4779 32446 4792
rect 29983 4712 30033 4740
rect 27606 4638 27656 4666
rect 27606 4618 27619 4638
rect 27639 4618 27656 4638
rect 12187 4407 12237 4423
rect 12395 4407 12445 4423
rect 12613 4407 12663 4423
rect 8236 4276 8286 4304
rect 9931 4348 9981 4361
rect 10149 4348 10199 4361
rect 10357 4348 10407 4361
rect 11389 4359 11439 4372
rect 11597 4359 11647 4372
rect 11815 4359 11865 4372
rect 13497 4417 13547 4445
rect 9133 4297 9183 4313
rect 9351 4297 9401 4313
rect 9559 4297 9609 4313
rect 5554 4208 5604 4236
rect 393 4095 443 4108
rect 611 4095 661 4108
rect 819 4095 869 4108
rect 3446 4150 3496 4163
rect 3654 4150 3704 4163
rect 3872 4150 3922 4163
rect 5554 4188 5567 4208
rect 5587 4188 5604 4208
rect 5554 4159 5604 4188
rect 5772 4211 5822 4236
rect 5772 4191 5785 4211
rect 5805 4191 5822 4211
rect 5772 4159 5822 4191
rect 5980 4209 6030 4236
rect 5980 4189 6003 4209
rect 6023 4189 6030 4209
rect 5980 4159 6030 4189
rect 6913 4169 6963 4185
rect 7121 4169 7171 4185
rect 7339 4169 7389 4185
rect 12187 4335 12237 4365
rect 12187 4315 12194 4335
rect 12214 4315 12237 4335
rect 12187 4288 12237 4315
rect 12395 4333 12445 4365
rect 12395 4313 12412 4333
rect 12432 4313 12445 4333
rect 12395 4288 12445 4313
rect 12613 4336 12663 4365
rect 12613 4316 12630 4336
rect 12650 4316 12663 4336
rect 13497 4397 13510 4417
rect 13530 4397 13547 4417
rect 13497 4368 13547 4397
rect 13715 4420 13765 4445
rect 13715 4400 13728 4420
rect 13748 4400 13765 4420
rect 13715 4368 13765 4400
rect 13923 4418 13973 4445
rect 13923 4398 13946 4418
rect 13966 4398 13973 4418
rect 13923 4368 13973 4398
rect 16551 4420 16601 4436
rect 16759 4420 16809 4436
rect 16977 4420 17027 4436
rect 12613 4288 12663 4316
rect 14295 4361 14345 4374
rect 14513 4361 14563 4374
rect 14721 4361 14771 4374
rect 15753 4372 15803 4385
rect 15961 4372 16011 4385
rect 16179 4372 16229 4385
rect 18865 4506 18915 4522
rect 19083 4506 19133 4522
rect 19291 4506 19341 4522
rect 20019 4506 20069 4536
rect 20019 4486 20026 4506
rect 20046 4486 20069 4506
rect 20019 4459 20069 4486
rect 20227 4504 20277 4536
rect 20227 4484 20244 4504
rect 20264 4484 20277 4504
rect 20227 4459 20277 4484
rect 20445 4507 20495 4536
rect 20445 4487 20462 4507
rect 20482 4487 20495 4507
rect 22127 4532 22177 4545
rect 22345 4532 22395 4545
rect 22553 4532 22603 4545
rect 25180 4587 25230 4600
rect 25388 4587 25438 4600
rect 25606 4587 25656 4600
rect 27606 4589 27656 4618
rect 27824 4641 27874 4666
rect 27824 4621 27837 4641
rect 27857 4621 27874 4641
rect 27824 4589 27874 4621
rect 28032 4639 28082 4666
rect 28032 4619 28055 4639
rect 28075 4619 28082 4639
rect 28032 4589 28082 4619
rect 28760 4603 28810 4619
rect 28968 4603 29018 4619
rect 29186 4603 29236 4619
rect 33921 4772 33971 4802
rect 33921 4752 33928 4772
rect 33948 4752 33971 4772
rect 33921 4725 33971 4752
rect 34129 4770 34179 4802
rect 34129 4750 34146 4770
rect 34166 4750 34179 4770
rect 34129 4725 34179 4750
rect 34347 4773 34397 4802
rect 34347 4753 34364 4773
rect 34384 4753 34397 4773
rect 34347 4725 34397 4753
rect 31970 4651 32020 4679
rect 31970 4631 31983 4651
rect 32003 4631 32020 4651
rect 20445 4459 20495 4487
rect 13497 4310 13547 4326
rect 13715 4310 13765 4326
rect 13923 4310 13973 4326
rect 9931 4220 9981 4248
rect 1190 4088 1240 4104
rect 1408 4088 1458 4104
rect 1616 4088 1666 4104
rect 2549 4084 2599 4114
rect 2549 4064 2556 4084
rect 2576 4064 2599 4084
rect 2549 4037 2599 4064
rect 2757 4082 2807 4114
rect 2757 4062 2774 4082
rect 2794 4062 2807 4082
rect 2757 4037 2807 4062
rect 2975 4085 3025 4114
rect 4757 4108 4807 4121
rect 4975 4108 5025 4121
rect 5183 4108 5233 4121
rect 7810 4163 7860 4176
rect 8018 4163 8068 4176
rect 8236 4163 8286 4176
rect 9931 4200 9944 4220
rect 9964 4200 9981 4220
rect 9931 4171 9981 4200
rect 10149 4223 10199 4248
rect 10149 4203 10162 4223
rect 10182 4203 10199 4223
rect 10149 4171 10199 4203
rect 10357 4221 10407 4248
rect 10357 4201 10380 4221
rect 10400 4201 10407 4221
rect 10357 4171 10407 4201
rect 11290 4181 11340 4197
rect 11498 4181 11548 4197
rect 11716 4181 11766 4197
rect 16551 4348 16601 4378
rect 16551 4328 16558 4348
rect 16578 4328 16601 4348
rect 16551 4301 16601 4328
rect 16759 4346 16809 4378
rect 16759 4326 16776 4346
rect 16796 4326 16809 4346
rect 16759 4301 16809 4326
rect 16977 4349 17027 4378
rect 16977 4329 16994 4349
rect 17014 4329 17027 4349
rect 17763 4391 17813 4419
rect 16977 4301 17027 4329
rect 17763 4371 17776 4391
rect 17796 4371 17813 4391
rect 17763 4342 17813 4371
rect 17981 4394 18031 4419
rect 17981 4374 17994 4394
rect 18014 4374 18031 4394
rect 17981 4342 18031 4374
rect 18189 4392 18239 4419
rect 18189 4372 18212 4392
rect 18232 4372 18239 4392
rect 18189 4342 18239 4372
rect 23229 4519 23279 4535
rect 23447 4519 23497 4535
rect 23655 4519 23705 4535
rect 24383 4519 24433 4549
rect 24383 4499 24390 4519
rect 24410 4499 24433 4519
rect 24383 4472 24433 4499
rect 24591 4517 24641 4549
rect 24591 4497 24608 4517
rect 24628 4497 24641 4517
rect 24591 4472 24641 4497
rect 24809 4520 24859 4549
rect 24809 4500 24826 4520
rect 24846 4500 24859 4520
rect 26504 4544 26554 4557
rect 26722 4544 26772 4557
rect 26930 4544 26980 4557
rect 29557 4599 29607 4612
rect 29765 4599 29815 4612
rect 29983 4599 30033 4612
rect 31970 4602 32020 4631
rect 32188 4654 32238 4679
rect 32188 4634 32201 4654
rect 32221 4634 32238 4654
rect 32188 4602 32238 4634
rect 32396 4652 32446 4679
rect 32396 4632 32419 4652
rect 32439 4632 32446 4652
rect 32396 4602 32446 4632
rect 33124 4616 33174 4632
rect 33332 4616 33382 4632
rect 33550 4616 33600 4632
rect 24809 4472 24859 4500
rect 20817 4394 20867 4410
rect 21025 4394 21075 4410
rect 21243 4394 21293 4410
rect 14295 4233 14345 4261
rect 2975 4065 2992 4085
rect 3012 4065 3025 4085
rect 2975 4037 3025 4065
rect 393 3967 443 3995
rect 393 3947 406 3967
rect 426 3947 443 3967
rect 393 3918 443 3947
rect 611 3970 661 3995
rect 611 3950 624 3970
rect 644 3950 661 3970
rect 611 3918 661 3950
rect 819 3968 869 3995
rect 819 3948 842 3968
rect 862 3948 869 3968
rect 819 3918 869 3948
rect 5554 4101 5604 4117
rect 5772 4101 5822 4117
rect 5980 4101 6030 4117
rect 6913 4097 6963 4127
rect 6913 4077 6920 4097
rect 6940 4077 6963 4097
rect 6913 4050 6963 4077
rect 7121 4095 7171 4127
rect 7121 4075 7138 4095
rect 7158 4075 7171 4095
rect 7121 4050 7171 4075
rect 7339 4098 7389 4127
rect 9134 4120 9184 4133
rect 9352 4120 9402 4133
rect 9560 4120 9610 4133
rect 12187 4175 12237 4188
rect 12395 4175 12445 4188
rect 12613 4175 12663 4188
rect 14295 4213 14308 4233
rect 14328 4213 14345 4233
rect 14295 4184 14345 4213
rect 14513 4236 14563 4261
rect 14513 4216 14526 4236
rect 14546 4216 14563 4236
rect 14513 4184 14563 4216
rect 14721 4234 14771 4261
rect 14721 4214 14744 4234
rect 14764 4214 14771 4234
rect 14721 4184 14771 4214
rect 15654 4194 15704 4210
rect 15862 4194 15912 4210
rect 16080 4194 16130 4210
rect 18561 4335 18611 4348
rect 18779 4335 18829 4348
rect 18987 4335 19037 4348
rect 20019 4346 20069 4359
rect 20227 4346 20277 4359
rect 20445 4346 20495 4359
rect 22127 4404 22177 4432
rect 17763 4284 17813 4300
rect 17981 4284 18031 4300
rect 18189 4284 18239 4300
rect 20817 4322 20867 4352
rect 20817 4302 20824 4322
rect 20844 4302 20867 4322
rect 20817 4275 20867 4302
rect 21025 4320 21075 4352
rect 21025 4300 21042 4320
rect 21062 4300 21075 4320
rect 21025 4275 21075 4300
rect 21243 4323 21293 4352
rect 21243 4303 21260 4323
rect 21280 4303 21293 4323
rect 22127 4384 22140 4404
rect 22160 4384 22177 4404
rect 22127 4355 22177 4384
rect 22345 4407 22395 4432
rect 22345 4387 22358 4407
rect 22378 4387 22395 4407
rect 22345 4355 22395 4387
rect 22553 4405 22603 4432
rect 22553 4385 22576 4405
rect 22596 4385 22603 4405
rect 22553 4355 22603 4385
rect 27606 4531 27656 4547
rect 27824 4531 27874 4547
rect 28032 4531 28082 4547
rect 28760 4531 28810 4561
rect 28760 4511 28767 4531
rect 28787 4511 28810 4531
rect 28760 4484 28810 4511
rect 28968 4529 29018 4561
rect 28968 4509 28985 4529
rect 29005 4509 29018 4529
rect 28968 4484 29018 4509
rect 29186 4532 29236 4561
rect 29186 4512 29203 4532
rect 29223 4512 29236 4532
rect 30868 4557 30918 4570
rect 31086 4557 31136 4570
rect 31294 4557 31344 4570
rect 33921 4612 33971 4625
rect 34129 4612 34179 4625
rect 34347 4612 34397 4625
rect 29186 4484 29236 4512
rect 25181 4407 25231 4423
rect 25389 4407 25439 4423
rect 25607 4407 25657 4423
rect 21243 4275 21293 4303
rect 22925 4348 22975 4361
rect 23143 4348 23193 4361
rect 23351 4348 23401 4361
rect 24383 4359 24433 4372
rect 24591 4359 24641 4372
rect 24809 4359 24859 4372
rect 26504 4416 26554 4444
rect 22127 4297 22177 4313
rect 22345 4297 22395 4313
rect 22553 4297 22603 4313
rect 7339 4078 7356 4098
rect 7376 4078 7389 4098
rect 7339 4050 7389 4078
rect 4757 3980 4807 4008
rect 2549 3924 2599 3937
rect 2757 3924 2807 3937
rect 2975 3924 3025 3937
rect 4757 3960 4770 3980
rect 4790 3960 4807 3980
rect 4757 3931 4807 3960
rect 4975 3983 5025 4008
rect 4975 3963 4988 3983
rect 5008 3963 5025 3983
rect 4975 3931 5025 3963
rect 5183 3981 5233 4008
rect 5183 3961 5206 3981
rect 5226 3961 5233 3981
rect 5183 3931 5233 3961
rect 9931 4113 9981 4129
rect 10149 4113 10199 4129
rect 10357 4113 10407 4129
rect 11290 4109 11340 4139
rect 11290 4089 11297 4109
rect 11317 4089 11340 4109
rect 11290 4062 11340 4089
rect 11498 4107 11548 4139
rect 11498 4087 11515 4107
rect 11535 4087 11548 4107
rect 11498 4062 11548 4087
rect 11716 4110 11766 4139
rect 13498 4133 13548 4146
rect 13716 4133 13766 4146
rect 13924 4133 13974 4146
rect 16551 4188 16601 4201
rect 16759 4188 16809 4201
rect 16977 4188 17027 4201
rect 18561 4207 18611 4235
rect 18561 4187 18574 4207
rect 18594 4187 18611 4207
rect 18561 4158 18611 4187
rect 18779 4210 18829 4235
rect 18779 4190 18792 4210
rect 18812 4190 18829 4210
rect 18779 4158 18829 4190
rect 18987 4208 19037 4235
rect 18987 4188 19010 4208
rect 19030 4188 19037 4208
rect 18987 4158 19037 4188
rect 19920 4168 19970 4184
rect 20128 4168 20178 4184
rect 20346 4168 20396 4184
rect 25181 4335 25231 4365
rect 25181 4315 25188 4335
rect 25208 4315 25231 4335
rect 25181 4288 25231 4315
rect 25389 4333 25439 4365
rect 25389 4313 25406 4333
rect 25426 4313 25439 4333
rect 25389 4288 25439 4313
rect 25607 4336 25657 4365
rect 25607 4316 25624 4336
rect 25644 4316 25657 4336
rect 26504 4396 26517 4416
rect 26537 4396 26554 4416
rect 26504 4367 26554 4396
rect 26722 4419 26772 4444
rect 26722 4399 26735 4419
rect 26755 4399 26772 4419
rect 26722 4367 26772 4399
rect 26930 4417 26980 4444
rect 26930 4397 26953 4417
rect 26973 4397 26980 4417
rect 26930 4367 26980 4397
rect 31970 4544 32020 4560
rect 32188 4544 32238 4560
rect 32396 4544 32446 4560
rect 33124 4544 33174 4574
rect 33124 4524 33131 4544
rect 33151 4524 33174 4544
rect 33124 4497 33174 4524
rect 33332 4542 33382 4574
rect 33332 4522 33349 4542
rect 33369 4522 33382 4542
rect 33332 4497 33382 4522
rect 33550 4545 33600 4574
rect 33550 4525 33567 4545
rect 33587 4525 33600 4545
rect 33550 4497 33600 4525
rect 29558 4419 29608 4435
rect 29766 4419 29816 4435
rect 29984 4419 30034 4435
rect 25607 4288 25657 4316
rect 27302 4360 27352 4373
rect 27520 4360 27570 4373
rect 27728 4360 27778 4373
rect 28760 4371 28810 4384
rect 28968 4371 29018 4384
rect 29186 4371 29236 4384
rect 30868 4429 30918 4457
rect 26504 4309 26554 4325
rect 26722 4309 26772 4325
rect 26930 4309 26980 4325
rect 22925 4220 22975 4248
rect 11716 4090 11733 4110
rect 11753 4090 11766 4110
rect 11716 4062 11766 4090
rect 9134 3992 9184 4020
rect 6913 3937 6963 3950
rect 7121 3937 7171 3950
rect 7339 3937 7389 3950
rect 9134 3972 9147 3992
rect 9167 3972 9184 3992
rect 9134 3943 9184 3972
rect 9352 3995 9402 4020
rect 9352 3975 9365 3995
rect 9385 3975 9402 3995
rect 9352 3943 9402 3975
rect 9560 3993 9610 4020
rect 9560 3973 9583 3993
rect 9603 3973 9610 3993
rect 9560 3943 9610 3973
rect 14295 4126 14345 4142
rect 14513 4126 14563 4142
rect 14721 4126 14771 4142
rect 15654 4122 15704 4152
rect 15654 4102 15661 4122
rect 15681 4102 15704 4122
rect 15654 4075 15704 4102
rect 15862 4120 15912 4152
rect 15862 4100 15879 4120
rect 15899 4100 15912 4120
rect 15862 4075 15912 4100
rect 16080 4123 16130 4152
rect 16080 4103 16097 4123
rect 16117 4103 16130 4123
rect 16080 4075 16130 4103
rect 17764 4107 17814 4120
rect 17982 4107 18032 4120
rect 18190 4107 18240 4120
rect 20817 4162 20867 4175
rect 21025 4162 21075 4175
rect 21243 4162 21293 4175
rect 22925 4200 22938 4220
rect 22958 4200 22975 4220
rect 22925 4171 22975 4200
rect 23143 4223 23193 4248
rect 23143 4203 23156 4223
rect 23176 4203 23193 4223
rect 23143 4171 23193 4203
rect 23351 4221 23401 4248
rect 23351 4201 23374 4221
rect 23394 4201 23401 4221
rect 23351 4171 23401 4201
rect 24284 4181 24334 4197
rect 24492 4181 24542 4197
rect 24710 4181 24760 4197
rect 29558 4347 29608 4377
rect 29558 4327 29565 4347
rect 29585 4327 29608 4347
rect 29558 4300 29608 4327
rect 29766 4345 29816 4377
rect 29766 4325 29783 4345
rect 29803 4325 29816 4345
rect 29766 4300 29816 4325
rect 29984 4348 30034 4377
rect 29984 4328 30001 4348
rect 30021 4328 30034 4348
rect 30868 4409 30881 4429
rect 30901 4409 30918 4429
rect 30868 4380 30918 4409
rect 31086 4432 31136 4457
rect 31086 4412 31099 4432
rect 31119 4412 31136 4432
rect 31086 4380 31136 4412
rect 31294 4430 31344 4457
rect 31294 4410 31317 4430
rect 31337 4410 31344 4430
rect 31294 4380 31344 4410
rect 33922 4432 33972 4448
rect 34130 4432 34180 4448
rect 34348 4432 34398 4448
rect 29984 4300 30034 4328
rect 31666 4373 31716 4386
rect 31884 4373 31934 4386
rect 32092 4373 32142 4386
rect 33124 4384 33174 4397
rect 33332 4384 33382 4397
rect 33550 4384 33600 4397
rect 30868 4322 30918 4338
rect 31086 4322 31136 4338
rect 31294 4322 31344 4338
rect 27302 4232 27352 4260
rect 13498 4005 13548 4033
rect 11290 3949 11340 3962
rect 11498 3949 11548 3962
rect 11716 3949 11766 3962
rect 13498 3985 13511 4005
rect 13531 3985 13548 4005
rect 13498 3956 13548 3985
rect 13716 4008 13766 4033
rect 13716 3988 13729 4008
rect 13749 3988 13766 4008
rect 13716 3956 13766 3988
rect 13924 4006 13974 4033
rect 13924 3986 13947 4006
rect 13967 3986 13974 4006
rect 13924 3956 13974 3986
rect 18561 4100 18611 4116
rect 18779 4100 18829 4116
rect 18987 4100 19037 4116
rect 19920 4096 19970 4126
rect 19920 4076 19927 4096
rect 19947 4076 19970 4096
rect 19920 4049 19970 4076
rect 20128 4094 20178 4126
rect 20128 4074 20145 4094
rect 20165 4074 20178 4094
rect 20128 4049 20178 4074
rect 20346 4097 20396 4126
rect 22128 4120 22178 4133
rect 22346 4120 22396 4133
rect 22554 4120 22604 4133
rect 25181 4175 25231 4188
rect 25389 4175 25439 4188
rect 25607 4175 25657 4188
rect 27302 4212 27315 4232
rect 27335 4212 27352 4232
rect 27302 4183 27352 4212
rect 27520 4235 27570 4260
rect 27520 4215 27533 4235
rect 27553 4215 27570 4235
rect 27520 4183 27570 4215
rect 27728 4233 27778 4260
rect 27728 4213 27751 4233
rect 27771 4213 27778 4233
rect 27728 4183 27778 4213
rect 28661 4193 28711 4209
rect 28869 4193 28919 4209
rect 29087 4193 29137 4209
rect 33922 4360 33972 4390
rect 33922 4340 33929 4360
rect 33949 4340 33972 4360
rect 33922 4313 33972 4340
rect 34130 4358 34180 4390
rect 34130 4338 34147 4358
rect 34167 4338 34180 4358
rect 34130 4313 34180 4338
rect 34348 4361 34398 4390
rect 34348 4341 34365 4361
rect 34385 4341 34398 4361
rect 34348 4313 34398 4341
rect 31666 4245 31716 4273
rect 20346 4077 20363 4097
rect 20383 4077 20396 4097
rect 20346 4049 20396 4077
rect 15654 3962 15704 3975
rect 15862 3962 15912 3975
rect 16080 3962 16130 3975
rect 17764 3979 17814 4007
rect 17764 3959 17777 3979
rect 17797 3959 17814 3979
rect 393 3860 443 3876
rect 611 3860 661 3876
rect 819 3860 869 3876
rect 4757 3873 4807 3889
rect 4975 3873 5025 3889
rect 5183 3873 5233 3889
rect 9134 3885 9184 3901
rect 9352 3885 9402 3901
rect 9560 3885 9610 3901
rect 13498 3898 13548 3914
rect 13716 3898 13766 3914
rect 13924 3898 13974 3914
rect 17764 3930 17814 3959
rect 17982 3982 18032 4007
rect 17982 3962 17995 3982
rect 18015 3962 18032 3982
rect 17982 3930 18032 3962
rect 18190 3980 18240 4007
rect 18190 3960 18213 3980
rect 18233 3960 18240 3980
rect 18190 3930 18240 3960
rect 22925 4113 22975 4129
rect 23143 4113 23193 4129
rect 23351 4113 23401 4129
rect 24284 4109 24334 4139
rect 24284 4089 24291 4109
rect 24311 4089 24334 4109
rect 24284 4062 24334 4089
rect 24492 4107 24542 4139
rect 24492 4087 24509 4107
rect 24529 4087 24542 4107
rect 24492 4062 24542 4087
rect 24710 4110 24760 4139
rect 26505 4132 26555 4145
rect 26723 4132 26773 4145
rect 26931 4132 26981 4145
rect 29558 4187 29608 4200
rect 29766 4187 29816 4200
rect 29984 4187 30034 4200
rect 31666 4225 31679 4245
rect 31699 4225 31716 4245
rect 31666 4196 31716 4225
rect 31884 4248 31934 4273
rect 31884 4228 31897 4248
rect 31917 4228 31934 4248
rect 31884 4196 31934 4228
rect 32092 4246 32142 4273
rect 32092 4226 32115 4246
rect 32135 4226 32142 4246
rect 32092 4196 32142 4226
rect 33025 4206 33075 4222
rect 33233 4206 33283 4222
rect 33451 4206 33501 4222
rect 24710 4090 24727 4110
rect 24747 4090 24760 4110
rect 24710 4062 24760 4090
rect 22128 3992 22178 4020
rect 19920 3936 19970 3949
rect 20128 3936 20178 3949
rect 20346 3936 20396 3949
rect 22128 3972 22141 3992
rect 22161 3972 22178 3992
rect 22128 3943 22178 3972
rect 22346 3995 22396 4020
rect 22346 3975 22359 3995
rect 22379 3975 22396 3995
rect 22346 3943 22396 3975
rect 22554 3993 22604 4020
rect 22554 3973 22577 3993
rect 22597 3973 22604 3993
rect 22554 3943 22604 3973
rect 27302 4125 27352 4141
rect 27520 4125 27570 4141
rect 27728 4125 27778 4141
rect 28661 4121 28711 4151
rect 28661 4101 28668 4121
rect 28688 4101 28711 4121
rect 28661 4074 28711 4101
rect 28869 4119 28919 4151
rect 28869 4099 28886 4119
rect 28906 4099 28919 4119
rect 28869 4074 28919 4099
rect 29087 4122 29137 4151
rect 30869 4145 30919 4158
rect 31087 4145 31137 4158
rect 31295 4145 31345 4158
rect 33922 4200 33972 4213
rect 34130 4200 34180 4213
rect 34348 4200 34398 4213
rect 29087 4102 29104 4122
rect 29124 4102 29137 4122
rect 29087 4074 29137 4102
rect 26505 4004 26555 4032
rect 24284 3949 24334 3962
rect 24492 3949 24542 3962
rect 24710 3949 24760 3962
rect 26505 3984 26518 4004
rect 26538 3984 26555 4004
rect 26505 3955 26555 3984
rect 26723 4007 26773 4032
rect 26723 3987 26736 4007
rect 26756 3987 26773 4007
rect 26723 3955 26773 3987
rect 26931 4005 26981 4032
rect 26931 3985 26954 4005
rect 26974 3985 26981 4005
rect 26931 3955 26981 3985
rect 31666 4138 31716 4154
rect 31884 4138 31934 4154
rect 32092 4138 32142 4154
rect 33025 4134 33075 4164
rect 33025 4114 33032 4134
rect 33052 4114 33075 4134
rect 33025 4087 33075 4114
rect 33233 4132 33283 4164
rect 33233 4112 33250 4132
rect 33270 4112 33283 4132
rect 33233 4087 33283 4112
rect 33451 4135 33501 4164
rect 33451 4115 33468 4135
rect 33488 4115 33501 4135
rect 33451 4087 33501 4115
rect 30869 4017 30919 4045
rect 28661 3961 28711 3974
rect 28869 3961 28919 3974
rect 29087 3961 29137 3974
rect 30869 3997 30882 4017
rect 30902 3997 30919 4017
rect 30869 3968 30919 3997
rect 31087 4020 31137 4045
rect 31087 4000 31100 4020
rect 31120 4000 31137 4020
rect 31087 3968 31137 4000
rect 31295 4018 31345 4045
rect 31295 3998 31318 4018
rect 31338 3998 31345 4018
rect 31295 3968 31345 3998
rect 33025 3974 33075 3987
rect 33233 3974 33283 3987
rect 33451 3974 33501 3987
rect 17764 3872 17814 3888
rect 17982 3872 18032 3888
rect 18190 3872 18240 3888
rect 22128 3885 22178 3901
rect 22346 3885 22396 3901
rect 22554 3885 22604 3901
rect 26505 3897 26555 3913
rect 26723 3897 26773 3913
rect 26931 3897 26981 3913
rect 30869 3910 30919 3926
rect 31087 3910 31137 3926
rect 31295 3910 31345 3926
rect 3428 3776 3478 3792
rect 3636 3776 3686 3792
rect 3854 3776 3904 3792
rect 7792 3789 7842 3805
rect 8000 3789 8050 3805
rect 8218 3789 8268 3805
rect 12169 3801 12219 3817
rect 12377 3801 12427 3817
rect 12595 3801 12645 3817
rect 16533 3814 16583 3830
rect 16741 3814 16791 3830
rect 16959 3814 17009 3830
rect 1272 3715 1322 3728
rect 1490 3715 1540 3728
rect 1698 3715 1748 3728
rect 3428 3704 3478 3734
rect 3428 3684 3435 3704
rect 3455 3684 3478 3704
rect 3428 3657 3478 3684
rect 3636 3702 3686 3734
rect 3636 3682 3653 3702
rect 3673 3682 3686 3702
rect 3636 3657 3686 3682
rect 3854 3705 3904 3734
rect 3854 3685 3871 3705
rect 3891 3685 3904 3705
rect 5636 3728 5686 3741
rect 5854 3728 5904 3741
rect 6062 3728 6112 3741
rect 3854 3657 3904 3685
rect 1272 3587 1322 3615
rect 1272 3567 1285 3587
rect 1305 3567 1322 3587
rect 1272 3538 1322 3567
rect 1490 3590 1540 3615
rect 1490 3570 1503 3590
rect 1523 3570 1540 3590
rect 1490 3538 1540 3570
rect 1698 3588 1748 3615
rect 1698 3568 1721 3588
rect 1741 3568 1748 3588
rect 1698 3538 1748 3568
rect 2631 3548 2681 3564
rect 2839 3548 2889 3564
rect 3057 3548 3107 3564
rect 7792 3717 7842 3747
rect 7792 3697 7799 3717
rect 7819 3697 7842 3717
rect 7792 3670 7842 3697
rect 8000 3715 8050 3747
rect 8000 3695 8017 3715
rect 8037 3695 8050 3715
rect 8000 3670 8050 3695
rect 8218 3718 8268 3747
rect 8218 3698 8235 3718
rect 8255 3698 8268 3718
rect 10013 3740 10063 3753
rect 10231 3740 10281 3753
rect 10439 3740 10489 3753
rect 8218 3670 8268 3698
rect 5636 3600 5686 3628
rect 5636 3580 5649 3600
rect 5669 3580 5686 3600
rect 375 3489 425 3502
rect 593 3489 643 3502
rect 801 3489 851 3502
rect 3428 3544 3478 3557
rect 3636 3544 3686 3557
rect 3854 3544 3904 3557
rect 5636 3551 5686 3580
rect 5854 3603 5904 3628
rect 5854 3583 5867 3603
rect 5887 3583 5904 3603
rect 5854 3551 5904 3583
rect 6062 3601 6112 3628
rect 6062 3581 6085 3601
rect 6105 3581 6112 3601
rect 6062 3551 6112 3581
rect 6995 3561 7045 3577
rect 7203 3561 7253 3577
rect 7421 3561 7471 3577
rect 12169 3729 12219 3759
rect 12169 3709 12176 3729
rect 12196 3709 12219 3729
rect 12169 3682 12219 3709
rect 12377 3727 12427 3759
rect 12377 3707 12394 3727
rect 12414 3707 12427 3727
rect 12377 3682 12427 3707
rect 12595 3730 12645 3759
rect 12595 3710 12612 3730
rect 12632 3710 12645 3730
rect 14377 3753 14427 3766
rect 14595 3753 14645 3766
rect 14803 3753 14853 3766
rect 12595 3682 12645 3710
rect 10013 3612 10063 3640
rect 10013 3592 10026 3612
rect 10046 3592 10063 3612
rect 1272 3480 1322 3496
rect 1490 3480 1540 3496
rect 1698 3480 1748 3496
rect 2631 3476 2681 3506
rect 2631 3456 2638 3476
rect 2658 3456 2681 3476
rect 2631 3429 2681 3456
rect 2839 3474 2889 3506
rect 2839 3454 2856 3474
rect 2876 3454 2889 3474
rect 2839 3429 2889 3454
rect 3057 3477 3107 3506
rect 3057 3457 3074 3477
rect 3094 3457 3107 3477
rect 4739 3502 4789 3515
rect 4957 3502 5007 3515
rect 5165 3502 5215 3515
rect 7792 3557 7842 3570
rect 8000 3557 8050 3570
rect 8218 3557 8268 3570
rect 10013 3563 10063 3592
rect 10231 3615 10281 3640
rect 10231 3595 10244 3615
rect 10264 3595 10281 3615
rect 10231 3563 10281 3595
rect 10439 3613 10489 3640
rect 10439 3593 10462 3613
rect 10482 3593 10489 3613
rect 10439 3563 10489 3593
rect 11372 3573 11422 3589
rect 11580 3573 11630 3589
rect 11798 3573 11848 3589
rect 16533 3742 16583 3772
rect 16533 3722 16540 3742
rect 16560 3722 16583 3742
rect 16533 3695 16583 3722
rect 16741 3740 16791 3772
rect 16741 3720 16758 3740
rect 16778 3720 16791 3740
rect 16741 3695 16791 3720
rect 16959 3743 17009 3772
rect 20799 3788 20849 3804
rect 21007 3788 21057 3804
rect 21225 3788 21275 3804
rect 25163 3801 25213 3817
rect 25371 3801 25421 3817
rect 25589 3801 25639 3817
rect 29540 3813 29590 3829
rect 29748 3813 29798 3829
rect 29966 3813 30016 3829
rect 33904 3826 33954 3842
rect 34112 3826 34162 3842
rect 34330 3826 34380 3842
rect 16959 3723 16976 3743
rect 16996 3723 17009 3743
rect 16959 3695 17009 3723
rect 18643 3727 18693 3740
rect 18861 3727 18911 3740
rect 19069 3727 19119 3740
rect 14377 3625 14427 3653
rect 14377 3605 14390 3625
rect 14410 3605 14427 3625
rect 3057 3429 3107 3457
rect 375 3361 425 3389
rect 375 3341 388 3361
rect 408 3341 425 3361
rect 375 3312 425 3341
rect 593 3364 643 3389
rect 593 3344 606 3364
rect 626 3344 643 3364
rect 593 3312 643 3344
rect 801 3362 851 3389
rect 801 3342 824 3362
rect 844 3342 851 3362
rect 801 3312 851 3342
rect 5636 3493 5686 3509
rect 5854 3493 5904 3509
rect 6062 3493 6112 3509
rect 6995 3489 7045 3519
rect 6995 3469 7002 3489
rect 7022 3469 7045 3489
rect 6995 3442 7045 3469
rect 7203 3487 7253 3519
rect 7203 3467 7220 3487
rect 7240 3467 7253 3487
rect 7203 3442 7253 3467
rect 7421 3490 7471 3519
rect 7421 3470 7438 3490
rect 7458 3470 7471 3490
rect 9116 3514 9166 3527
rect 9334 3514 9384 3527
rect 9542 3514 9592 3527
rect 12169 3569 12219 3582
rect 12377 3569 12427 3582
rect 12595 3569 12645 3582
rect 14377 3576 14427 3605
rect 14595 3628 14645 3653
rect 14595 3608 14608 3628
rect 14628 3608 14645 3628
rect 14595 3576 14645 3608
rect 14803 3626 14853 3653
rect 14803 3606 14826 3626
rect 14846 3606 14853 3626
rect 14803 3576 14853 3606
rect 15736 3586 15786 3602
rect 15944 3586 15994 3602
rect 16162 3586 16212 3602
rect 20799 3716 20849 3746
rect 20799 3696 20806 3716
rect 20826 3696 20849 3716
rect 20799 3669 20849 3696
rect 21007 3714 21057 3746
rect 21007 3694 21024 3714
rect 21044 3694 21057 3714
rect 21007 3669 21057 3694
rect 21225 3717 21275 3746
rect 21225 3697 21242 3717
rect 21262 3697 21275 3717
rect 23007 3740 23057 3753
rect 23225 3740 23275 3753
rect 23433 3740 23483 3753
rect 21225 3669 21275 3697
rect 7421 3442 7471 3470
rect 3429 3364 3479 3380
rect 3637 3364 3687 3380
rect 3855 3364 3905 3380
rect 1173 3305 1223 3318
rect 1391 3305 1441 3318
rect 1599 3305 1649 3318
rect 2631 3316 2681 3329
rect 2839 3316 2889 3329
rect 3057 3316 3107 3329
rect 4739 3374 4789 3402
rect 375 3254 425 3270
rect 593 3254 643 3270
rect 801 3254 851 3270
rect 3429 3292 3479 3322
rect 3429 3272 3436 3292
rect 3456 3272 3479 3292
rect 3429 3245 3479 3272
rect 3637 3290 3687 3322
rect 3637 3270 3654 3290
rect 3674 3270 3687 3290
rect 3637 3245 3687 3270
rect 3855 3293 3905 3322
rect 3855 3273 3872 3293
rect 3892 3273 3905 3293
rect 4739 3354 4752 3374
rect 4772 3354 4789 3374
rect 4739 3325 4789 3354
rect 4957 3377 5007 3402
rect 4957 3357 4970 3377
rect 4990 3357 5007 3377
rect 4957 3325 5007 3357
rect 5165 3375 5215 3402
rect 5165 3355 5188 3375
rect 5208 3355 5215 3375
rect 5165 3325 5215 3355
rect 10013 3505 10063 3521
rect 10231 3505 10281 3521
rect 10439 3505 10489 3521
rect 11372 3501 11422 3531
rect 11372 3481 11379 3501
rect 11399 3481 11422 3501
rect 11372 3454 11422 3481
rect 11580 3499 11630 3531
rect 11580 3479 11597 3499
rect 11617 3479 11630 3499
rect 11580 3454 11630 3479
rect 11798 3502 11848 3531
rect 11798 3482 11815 3502
rect 11835 3482 11848 3502
rect 13480 3527 13530 3540
rect 13698 3527 13748 3540
rect 13906 3527 13956 3540
rect 16533 3582 16583 3595
rect 16741 3582 16791 3595
rect 16959 3582 17009 3595
rect 18643 3599 18693 3627
rect 18643 3579 18656 3599
rect 18676 3579 18693 3599
rect 18643 3550 18693 3579
rect 18861 3602 18911 3627
rect 18861 3582 18874 3602
rect 18894 3582 18911 3602
rect 18861 3550 18911 3582
rect 19069 3600 19119 3627
rect 19069 3580 19092 3600
rect 19112 3580 19119 3600
rect 19069 3550 19119 3580
rect 20002 3560 20052 3576
rect 20210 3560 20260 3576
rect 20428 3560 20478 3576
rect 25163 3729 25213 3759
rect 25163 3709 25170 3729
rect 25190 3709 25213 3729
rect 25163 3682 25213 3709
rect 25371 3727 25421 3759
rect 25371 3707 25388 3727
rect 25408 3707 25421 3727
rect 25371 3682 25421 3707
rect 25589 3730 25639 3759
rect 25589 3710 25606 3730
rect 25626 3710 25639 3730
rect 27384 3752 27434 3765
rect 27602 3752 27652 3765
rect 27810 3752 27860 3765
rect 25589 3682 25639 3710
rect 23007 3612 23057 3640
rect 23007 3592 23020 3612
rect 23040 3592 23057 3612
rect 11798 3454 11848 3482
rect 7793 3377 7843 3393
rect 8001 3377 8051 3393
rect 8219 3377 8269 3393
rect 3855 3245 3905 3273
rect 5537 3318 5587 3331
rect 5755 3318 5805 3331
rect 5963 3318 6013 3331
rect 6995 3329 7045 3342
rect 7203 3329 7253 3342
rect 7421 3329 7471 3342
rect 9116 3386 9166 3414
rect 4739 3267 4789 3283
rect 4957 3267 5007 3283
rect 5165 3267 5215 3283
rect 1173 3177 1223 3205
rect 1173 3157 1186 3177
rect 1206 3157 1223 3177
rect 1173 3128 1223 3157
rect 1391 3180 1441 3205
rect 1391 3160 1404 3180
rect 1424 3160 1441 3180
rect 1391 3128 1441 3160
rect 1599 3178 1649 3205
rect 1599 3158 1622 3178
rect 1642 3158 1649 3178
rect 1599 3128 1649 3158
rect 2466 3140 2516 3156
rect 2674 3140 2724 3156
rect 2892 3140 2942 3156
rect 7793 3305 7843 3335
rect 7793 3285 7800 3305
rect 7820 3285 7843 3305
rect 7793 3258 7843 3285
rect 8001 3303 8051 3335
rect 8001 3283 8018 3303
rect 8038 3283 8051 3303
rect 8001 3258 8051 3283
rect 8219 3306 8269 3335
rect 8219 3286 8236 3306
rect 8256 3286 8269 3306
rect 9116 3366 9129 3386
rect 9149 3366 9166 3386
rect 9116 3337 9166 3366
rect 9334 3389 9384 3414
rect 9334 3369 9347 3389
rect 9367 3369 9384 3389
rect 9334 3337 9384 3369
rect 9542 3387 9592 3414
rect 9542 3367 9565 3387
rect 9585 3367 9592 3387
rect 9542 3337 9592 3367
rect 14377 3518 14427 3534
rect 14595 3518 14645 3534
rect 14803 3518 14853 3534
rect 15736 3514 15786 3544
rect 15736 3494 15743 3514
rect 15763 3494 15786 3514
rect 15736 3467 15786 3494
rect 15944 3512 15994 3544
rect 15944 3492 15961 3512
rect 15981 3492 15994 3512
rect 15944 3467 15994 3492
rect 16162 3515 16212 3544
rect 16162 3495 16179 3515
rect 16199 3495 16212 3515
rect 16162 3467 16212 3495
rect 17746 3501 17796 3514
rect 17964 3501 18014 3514
rect 18172 3501 18222 3514
rect 20799 3556 20849 3569
rect 21007 3556 21057 3569
rect 21225 3556 21275 3569
rect 23007 3563 23057 3592
rect 23225 3615 23275 3640
rect 23225 3595 23238 3615
rect 23258 3595 23275 3615
rect 23225 3563 23275 3595
rect 23433 3613 23483 3640
rect 23433 3593 23456 3613
rect 23476 3593 23483 3613
rect 23433 3563 23483 3593
rect 24366 3573 24416 3589
rect 24574 3573 24624 3589
rect 24792 3573 24842 3589
rect 29540 3741 29590 3771
rect 29540 3721 29547 3741
rect 29567 3721 29590 3741
rect 29540 3694 29590 3721
rect 29748 3739 29798 3771
rect 29748 3719 29765 3739
rect 29785 3719 29798 3739
rect 29748 3694 29798 3719
rect 29966 3742 30016 3771
rect 29966 3722 29983 3742
rect 30003 3722 30016 3742
rect 31748 3765 31798 3778
rect 31966 3765 32016 3778
rect 32174 3765 32224 3778
rect 29966 3694 30016 3722
rect 27384 3624 27434 3652
rect 27384 3604 27397 3624
rect 27417 3604 27434 3624
rect 12170 3389 12220 3405
rect 12378 3389 12428 3405
rect 12596 3389 12646 3405
rect 8219 3258 8269 3286
rect 9914 3330 9964 3343
rect 10132 3330 10182 3343
rect 10340 3330 10390 3343
rect 11372 3341 11422 3354
rect 11580 3341 11630 3354
rect 11798 3341 11848 3354
rect 13480 3399 13530 3427
rect 9116 3279 9166 3295
rect 9334 3279 9384 3295
rect 9542 3279 9592 3295
rect 5537 3190 5587 3218
rect 376 3077 426 3090
rect 594 3077 644 3090
rect 802 3077 852 3090
rect 3429 3132 3479 3145
rect 3637 3132 3687 3145
rect 3855 3132 3905 3145
rect 5537 3170 5550 3190
rect 5570 3170 5587 3190
rect 5537 3141 5587 3170
rect 5755 3193 5805 3218
rect 5755 3173 5768 3193
rect 5788 3173 5805 3193
rect 5755 3141 5805 3173
rect 5963 3191 6013 3218
rect 5963 3171 5986 3191
rect 6006 3171 6013 3191
rect 5963 3141 6013 3171
rect 6830 3153 6880 3169
rect 7038 3153 7088 3169
rect 7256 3153 7306 3169
rect 12170 3317 12220 3347
rect 12170 3297 12177 3317
rect 12197 3297 12220 3317
rect 12170 3270 12220 3297
rect 12378 3315 12428 3347
rect 12378 3295 12395 3315
rect 12415 3295 12428 3315
rect 12378 3270 12428 3295
rect 12596 3318 12646 3347
rect 12596 3298 12613 3318
rect 12633 3298 12646 3318
rect 13480 3379 13493 3399
rect 13513 3379 13530 3399
rect 13480 3350 13530 3379
rect 13698 3402 13748 3427
rect 13698 3382 13711 3402
rect 13731 3382 13748 3402
rect 13698 3350 13748 3382
rect 13906 3400 13956 3427
rect 13906 3380 13929 3400
rect 13949 3380 13956 3400
rect 13906 3350 13956 3380
rect 16534 3402 16584 3418
rect 16742 3402 16792 3418
rect 16960 3402 17010 3418
rect 12596 3270 12646 3298
rect 14278 3343 14328 3356
rect 14496 3343 14546 3356
rect 14704 3343 14754 3356
rect 15736 3354 15786 3367
rect 15944 3354 15994 3367
rect 16162 3354 16212 3367
rect 18643 3492 18693 3508
rect 18861 3492 18911 3508
rect 19069 3492 19119 3508
rect 20002 3488 20052 3518
rect 20002 3468 20009 3488
rect 20029 3468 20052 3488
rect 20002 3441 20052 3468
rect 20210 3486 20260 3518
rect 20210 3466 20227 3486
rect 20247 3466 20260 3486
rect 20210 3441 20260 3466
rect 20428 3489 20478 3518
rect 20428 3469 20445 3489
rect 20465 3469 20478 3489
rect 22110 3514 22160 3527
rect 22328 3514 22378 3527
rect 22536 3514 22586 3527
rect 25163 3569 25213 3582
rect 25371 3569 25421 3582
rect 25589 3569 25639 3582
rect 27384 3575 27434 3604
rect 27602 3627 27652 3652
rect 27602 3607 27615 3627
rect 27635 3607 27652 3627
rect 27602 3575 27652 3607
rect 27810 3625 27860 3652
rect 27810 3605 27833 3625
rect 27853 3605 27860 3625
rect 27810 3575 27860 3605
rect 28743 3585 28793 3601
rect 28951 3585 29001 3601
rect 29169 3585 29219 3601
rect 33904 3754 33954 3784
rect 33904 3734 33911 3754
rect 33931 3734 33954 3754
rect 33904 3707 33954 3734
rect 34112 3752 34162 3784
rect 34112 3732 34129 3752
rect 34149 3732 34162 3752
rect 34112 3707 34162 3732
rect 34330 3755 34380 3784
rect 34330 3735 34347 3755
rect 34367 3735 34380 3755
rect 34330 3707 34380 3735
rect 31748 3637 31798 3665
rect 31748 3617 31761 3637
rect 31781 3617 31798 3637
rect 20428 3441 20478 3469
rect 13480 3292 13530 3308
rect 13698 3292 13748 3308
rect 13906 3292 13956 3308
rect 9914 3202 9964 3230
rect 1173 3070 1223 3086
rect 1391 3070 1441 3086
rect 1599 3070 1649 3086
rect 2466 3068 2516 3098
rect 2466 3048 2473 3068
rect 2493 3048 2516 3068
rect 2466 3021 2516 3048
rect 2674 3066 2724 3098
rect 2674 3046 2691 3066
rect 2711 3046 2724 3066
rect 2674 3021 2724 3046
rect 2892 3069 2942 3098
rect 4740 3090 4790 3103
rect 4958 3090 5008 3103
rect 5166 3090 5216 3103
rect 7793 3145 7843 3158
rect 8001 3145 8051 3158
rect 8219 3145 8269 3158
rect 9914 3182 9927 3202
rect 9947 3182 9964 3202
rect 9914 3153 9964 3182
rect 10132 3205 10182 3230
rect 10132 3185 10145 3205
rect 10165 3185 10182 3205
rect 10132 3153 10182 3185
rect 10340 3203 10390 3230
rect 10340 3183 10363 3203
rect 10383 3183 10390 3203
rect 10340 3153 10390 3183
rect 11207 3165 11257 3181
rect 11415 3165 11465 3181
rect 11633 3165 11683 3181
rect 16534 3330 16584 3360
rect 16534 3310 16541 3330
rect 16561 3310 16584 3330
rect 16534 3283 16584 3310
rect 16742 3328 16792 3360
rect 16742 3308 16759 3328
rect 16779 3308 16792 3328
rect 16742 3283 16792 3308
rect 16960 3331 17010 3360
rect 16960 3311 16977 3331
rect 16997 3311 17010 3331
rect 17746 3373 17796 3401
rect 16960 3283 17010 3311
rect 17746 3353 17759 3373
rect 17779 3353 17796 3373
rect 17746 3324 17796 3353
rect 17964 3376 18014 3401
rect 17964 3356 17977 3376
rect 17997 3356 18014 3376
rect 17964 3324 18014 3356
rect 18172 3374 18222 3401
rect 18172 3354 18195 3374
rect 18215 3354 18222 3374
rect 18172 3324 18222 3354
rect 23007 3505 23057 3521
rect 23225 3505 23275 3521
rect 23433 3505 23483 3521
rect 24366 3501 24416 3531
rect 24366 3481 24373 3501
rect 24393 3481 24416 3501
rect 24366 3454 24416 3481
rect 24574 3499 24624 3531
rect 24574 3479 24591 3499
rect 24611 3479 24624 3499
rect 24574 3454 24624 3479
rect 24792 3502 24842 3531
rect 24792 3482 24809 3502
rect 24829 3482 24842 3502
rect 26487 3526 26537 3539
rect 26705 3526 26755 3539
rect 26913 3526 26963 3539
rect 29540 3581 29590 3594
rect 29748 3581 29798 3594
rect 29966 3581 30016 3594
rect 31748 3588 31798 3617
rect 31966 3640 32016 3665
rect 31966 3620 31979 3640
rect 31999 3620 32016 3640
rect 31966 3588 32016 3620
rect 32174 3638 32224 3665
rect 32174 3618 32197 3638
rect 32217 3618 32224 3638
rect 32174 3588 32224 3618
rect 33107 3598 33157 3614
rect 33315 3598 33365 3614
rect 33533 3598 33583 3614
rect 24792 3454 24842 3482
rect 20800 3376 20850 3392
rect 21008 3376 21058 3392
rect 21226 3376 21276 3392
rect 14278 3215 14328 3243
rect 2892 3049 2909 3069
rect 2929 3049 2942 3069
rect 2892 3021 2942 3049
rect 376 2949 426 2977
rect 376 2929 389 2949
rect 409 2929 426 2949
rect 376 2900 426 2929
rect 594 2952 644 2977
rect 594 2932 607 2952
rect 627 2932 644 2952
rect 594 2900 644 2932
rect 802 2950 852 2977
rect 802 2930 825 2950
rect 845 2930 852 2950
rect 802 2900 852 2930
rect 5537 3083 5587 3099
rect 5755 3083 5805 3099
rect 5963 3083 6013 3099
rect 6830 3081 6880 3111
rect 6830 3061 6837 3081
rect 6857 3061 6880 3081
rect 6830 3034 6880 3061
rect 7038 3079 7088 3111
rect 7038 3059 7055 3079
rect 7075 3059 7088 3079
rect 7038 3034 7088 3059
rect 7256 3082 7306 3111
rect 9117 3102 9167 3115
rect 9335 3102 9385 3115
rect 9543 3102 9593 3115
rect 12170 3157 12220 3170
rect 12378 3157 12428 3170
rect 12596 3157 12646 3170
rect 14278 3195 14291 3215
rect 14311 3195 14328 3215
rect 14278 3166 14328 3195
rect 14496 3218 14546 3243
rect 14496 3198 14509 3218
rect 14529 3198 14546 3218
rect 14496 3166 14546 3198
rect 14704 3216 14754 3243
rect 14704 3196 14727 3216
rect 14747 3196 14754 3216
rect 14704 3166 14754 3196
rect 15571 3178 15621 3194
rect 15779 3178 15829 3194
rect 15997 3178 16047 3194
rect 18544 3317 18594 3330
rect 18762 3317 18812 3330
rect 18970 3317 19020 3330
rect 20002 3328 20052 3341
rect 20210 3328 20260 3341
rect 20428 3328 20478 3341
rect 22110 3386 22160 3414
rect 17746 3266 17796 3282
rect 17964 3266 18014 3282
rect 18172 3266 18222 3282
rect 20800 3304 20850 3334
rect 20800 3284 20807 3304
rect 20827 3284 20850 3304
rect 20800 3257 20850 3284
rect 21008 3302 21058 3334
rect 21008 3282 21025 3302
rect 21045 3282 21058 3302
rect 21008 3257 21058 3282
rect 21226 3305 21276 3334
rect 21226 3285 21243 3305
rect 21263 3285 21276 3305
rect 22110 3366 22123 3386
rect 22143 3366 22160 3386
rect 22110 3337 22160 3366
rect 22328 3389 22378 3414
rect 22328 3369 22341 3389
rect 22361 3369 22378 3389
rect 22328 3337 22378 3369
rect 22536 3387 22586 3414
rect 22536 3367 22559 3387
rect 22579 3367 22586 3387
rect 22536 3337 22586 3367
rect 27384 3517 27434 3533
rect 27602 3517 27652 3533
rect 27810 3517 27860 3533
rect 28743 3513 28793 3543
rect 28743 3493 28750 3513
rect 28770 3493 28793 3513
rect 28743 3466 28793 3493
rect 28951 3511 29001 3543
rect 28951 3491 28968 3511
rect 28988 3491 29001 3511
rect 28951 3466 29001 3491
rect 29169 3514 29219 3543
rect 29169 3494 29186 3514
rect 29206 3494 29219 3514
rect 30851 3539 30901 3552
rect 31069 3539 31119 3552
rect 31277 3539 31327 3552
rect 33904 3594 33954 3607
rect 34112 3594 34162 3607
rect 34330 3594 34380 3607
rect 29169 3466 29219 3494
rect 25164 3389 25214 3405
rect 25372 3389 25422 3405
rect 25590 3389 25640 3405
rect 21226 3257 21276 3285
rect 22908 3330 22958 3343
rect 23126 3330 23176 3343
rect 23334 3330 23384 3343
rect 24366 3341 24416 3354
rect 24574 3341 24624 3354
rect 24792 3341 24842 3354
rect 26487 3398 26537 3426
rect 22110 3279 22160 3295
rect 22328 3279 22378 3295
rect 22536 3279 22586 3295
rect 7256 3062 7273 3082
rect 7293 3062 7306 3082
rect 7256 3034 7306 3062
rect 4740 2962 4790 2990
rect 2466 2908 2516 2921
rect 2674 2908 2724 2921
rect 2892 2908 2942 2921
rect 4740 2942 4753 2962
rect 4773 2942 4790 2962
rect 4740 2913 4790 2942
rect 4958 2965 5008 2990
rect 4958 2945 4971 2965
rect 4991 2945 5008 2965
rect 4958 2913 5008 2945
rect 5166 2963 5216 2990
rect 5166 2943 5189 2963
rect 5209 2943 5216 2963
rect 5166 2913 5216 2943
rect 9914 3095 9964 3111
rect 10132 3095 10182 3111
rect 10340 3095 10390 3111
rect 11207 3093 11257 3123
rect 11207 3073 11214 3093
rect 11234 3073 11257 3093
rect 11207 3046 11257 3073
rect 11415 3091 11465 3123
rect 11415 3071 11432 3091
rect 11452 3071 11465 3091
rect 11415 3046 11465 3071
rect 11633 3094 11683 3123
rect 13481 3115 13531 3128
rect 13699 3115 13749 3128
rect 13907 3115 13957 3128
rect 16534 3170 16584 3183
rect 16742 3170 16792 3183
rect 16960 3170 17010 3183
rect 18544 3189 18594 3217
rect 18544 3169 18557 3189
rect 18577 3169 18594 3189
rect 18544 3140 18594 3169
rect 18762 3192 18812 3217
rect 18762 3172 18775 3192
rect 18795 3172 18812 3192
rect 18762 3140 18812 3172
rect 18970 3190 19020 3217
rect 18970 3170 18993 3190
rect 19013 3170 19020 3190
rect 18970 3140 19020 3170
rect 19837 3152 19887 3168
rect 20045 3152 20095 3168
rect 20263 3152 20313 3168
rect 25164 3317 25214 3347
rect 25164 3297 25171 3317
rect 25191 3297 25214 3317
rect 25164 3270 25214 3297
rect 25372 3315 25422 3347
rect 25372 3295 25389 3315
rect 25409 3295 25422 3315
rect 25372 3270 25422 3295
rect 25590 3318 25640 3347
rect 25590 3298 25607 3318
rect 25627 3298 25640 3318
rect 26487 3378 26500 3398
rect 26520 3378 26537 3398
rect 26487 3349 26537 3378
rect 26705 3401 26755 3426
rect 26705 3381 26718 3401
rect 26738 3381 26755 3401
rect 26705 3349 26755 3381
rect 26913 3399 26963 3426
rect 26913 3379 26936 3399
rect 26956 3379 26963 3399
rect 26913 3349 26963 3379
rect 31748 3530 31798 3546
rect 31966 3530 32016 3546
rect 32174 3530 32224 3546
rect 33107 3526 33157 3556
rect 33107 3506 33114 3526
rect 33134 3506 33157 3526
rect 33107 3479 33157 3506
rect 33315 3524 33365 3556
rect 33315 3504 33332 3524
rect 33352 3504 33365 3524
rect 33315 3479 33365 3504
rect 33533 3527 33583 3556
rect 33533 3507 33550 3527
rect 33570 3507 33583 3527
rect 33533 3479 33583 3507
rect 29541 3401 29591 3417
rect 29749 3401 29799 3417
rect 29967 3401 30017 3417
rect 25590 3270 25640 3298
rect 27285 3342 27335 3355
rect 27503 3342 27553 3355
rect 27711 3342 27761 3355
rect 28743 3353 28793 3366
rect 28951 3353 29001 3366
rect 29169 3353 29219 3366
rect 30851 3411 30901 3439
rect 26487 3291 26537 3307
rect 26705 3291 26755 3307
rect 26913 3291 26963 3307
rect 22908 3202 22958 3230
rect 11633 3074 11650 3094
rect 11670 3074 11683 3094
rect 11633 3046 11683 3074
rect 9117 2974 9167 3002
rect 6830 2921 6880 2934
rect 7038 2921 7088 2934
rect 7256 2921 7306 2934
rect 9117 2954 9130 2974
rect 9150 2954 9167 2974
rect 9117 2925 9167 2954
rect 9335 2977 9385 3002
rect 9335 2957 9348 2977
rect 9368 2957 9385 2977
rect 9335 2925 9385 2957
rect 9543 2975 9593 3002
rect 9543 2955 9566 2975
rect 9586 2955 9593 2975
rect 9543 2925 9593 2955
rect 14278 3108 14328 3124
rect 14496 3108 14546 3124
rect 14704 3108 14754 3124
rect 15571 3106 15621 3136
rect 15571 3086 15578 3106
rect 15598 3086 15621 3106
rect 15571 3059 15621 3086
rect 15779 3104 15829 3136
rect 15779 3084 15796 3104
rect 15816 3084 15829 3104
rect 15779 3059 15829 3084
rect 15997 3107 16047 3136
rect 15997 3087 16014 3107
rect 16034 3087 16047 3107
rect 15997 3059 16047 3087
rect 17747 3089 17797 3102
rect 17965 3089 18015 3102
rect 18173 3089 18223 3102
rect 20800 3144 20850 3157
rect 21008 3144 21058 3157
rect 21226 3144 21276 3157
rect 22908 3182 22921 3202
rect 22941 3182 22958 3202
rect 22908 3153 22958 3182
rect 23126 3205 23176 3230
rect 23126 3185 23139 3205
rect 23159 3185 23176 3205
rect 23126 3153 23176 3185
rect 23334 3203 23384 3230
rect 23334 3183 23357 3203
rect 23377 3183 23384 3203
rect 23334 3153 23384 3183
rect 24201 3165 24251 3181
rect 24409 3165 24459 3181
rect 24627 3165 24677 3181
rect 29541 3329 29591 3359
rect 29541 3309 29548 3329
rect 29568 3309 29591 3329
rect 29541 3282 29591 3309
rect 29749 3327 29799 3359
rect 29749 3307 29766 3327
rect 29786 3307 29799 3327
rect 29749 3282 29799 3307
rect 29967 3330 30017 3359
rect 29967 3310 29984 3330
rect 30004 3310 30017 3330
rect 30851 3391 30864 3411
rect 30884 3391 30901 3411
rect 30851 3362 30901 3391
rect 31069 3414 31119 3439
rect 31069 3394 31082 3414
rect 31102 3394 31119 3414
rect 31069 3362 31119 3394
rect 31277 3412 31327 3439
rect 31277 3392 31300 3412
rect 31320 3392 31327 3412
rect 31277 3362 31327 3392
rect 33905 3414 33955 3430
rect 34113 3414 34163 3430
rect 34331 3414 34381 3430
rect 29967 3282 30017 3310
rect 31649 3355 31699 3368
rect 31867 3355 31917 3368
rect 32075 3355 32125 3368
rect 33107 3366 33157 3379
rect 33315 3366 33365 3379
rect 33533 3366 33583 3379
rect 30851 3304 30901 3320
rect 31069 3304 31119 3320
rect 31277 3304 31327 3320
rect 27285 3214 27335 3242
rect 13481 2987 13531 3015
rect 11207 2933 11257 2946
rect 11415 2933 11465 2946
rect 11633 2933 11683 2946
rect 13481 2967 13494 2987
rect 13514 2967 13531 2987
rect 13481 2938 13531 2967
rect 13699 2990 13749 3015
rect 13699 2970 13712 2990
rect 13732 2970 13749 2990
rect 13699 2938 13749 2970
rect 13907 2988 13957 3015
rect 13907 2968 13930 2988
rect 13950 2968 13957 2988
rect 13907 2938 13957 2968
rect 18544 3082 18594 3098
rect 18762 3082 18812 3098
rect 18970 3082 19020 3098
rect 19837 3080 19887 3110
rect 19837 3060 19844 3080
rect 19864 3060 19887 3080
rect 19837 3033 19887 3060
rect 20045 3078 20095 3110
rect 20045 3058 20062 3078
rect 20082 3058 20095 3078
rect 20045 3033 20095 3058
rect 20263 3081 20313 3110
rect 22111 3102 22161 3115
rect 22329 3102 22379 3115
rect 22537 3102 22587 3115
rect 25164 3157 25214 3170
rect 25372 3157 25422 3170
rect 25590 3157 25640 3170
rect 27285 3194 27298 3214
rect 27318 3194 27335 3214
rect 27285 3165 27335 3194
rect 27503 3217 27553 3242
rect 27503 3197 27516 3217
rect 27536 3197 27553 3217
rect 27503 3165 27553 3197
rect 27711 3215 27761 3242
rect 27711 3195 27734 3215
rect 27754 3195 27761 3215
rect 27711 3165 27761 3195
rect 28578 3177 28628 3193
rect 28786 3177 28836 3193
rect 29004 3177 29054 3193
rect 33905 3342 33955 3372
rect 33905 3322 33912 3342
rect 33932 3322 33955 3342
rect 33905 3295 33955 3322
rect 34113 3340 34163 3372
rect 34113 3320 34130 3340
rect 34150 3320 34163 3340
rect 34113 3295 34163 3320
rect 34331 3343 34381 3372
rect 34331 3323 34348 3343
rect 34368 3323 34381 3343
rect 34331 3295 34381 3323
rect 31649 3227 31699 3255
rect 20263 3061 20280 3081
rect 20300 3061 20313 3081
rect 20263 3033 20313 3061
rect 15571 2946 15621 2959
rect 15779 2946 15829 2959
rect 15997 2946 16047 2959
rect 17747 2961 17797 2989
rect 17747 2941 17760 2961
rect 17780 2941 17797 2961
rect 376 2842 426 2858
rect 594 2842 644 2858
rect 802 2842 852 2858
rect 4740 2855 4790 2871
rect 4958 2855 5008 2871
rect 5166 2855 5216 2871
rect 9117 2867 9167 2883
rect 9335 2867 9385 2883
rect 9543 2867 9593 2883
rect 13481 2880 13531 2896
rect 13699 2880 13749 2896
rect 13907 2880 13957 2896
rect 17747 2912 17797 2941
rect 17965 2964 18015 2989
rect 17965 2944 17978 2964
rect 17998 2944 18015 2964
rect 17965 2912 18015 2944
rect 18173 2962 18223 2989
rect 18173 2942 18196 2962
rect 18216 2942 18223 2962
rect 18173 2912 18223 2942
rect 22908 3095 22958 3111
rect 23126 3095 23176 3111
rect 23334 3095 23384 3111
rect 24201 3093 24251 3123
rect 24201 3073 24208 3093
rect 24228 3073 24251 3093
rect 24201 3046 24251 3073
rect 24409 3091 24459 3123
rect 24409 3071 24426 3091
rect 24446 3071 24459 3091
rect 24409 3046 24459 3071
rect 24627 3094 24677 3123
rect 26488 3114 26538 3127
rect 26706 3114 26756 3127
rect 26914 3114 26964 3127
rect 29541 3169 29591 3182
rect 29749 3169 29799 3182
rect 29967 3169 30017 3182
rect 31649 3207 31662 3227
rect 31682 3207 31699 3227
rect 31649 3178 31699 3207
rect 31867 3230 31917 3255
rect 31867 3210 31880 3230
rect 31900 3210 31917 3230
rect 31867 3178 31917 3210
rect 32075 3228 32125 3255
rect 32075 3208 32098 3228
rect 32118 3208 32125 3228
rect 32075 3178 32125 3208
rect 32942 3190 32992 3206
rect 33150 3190 33200 3206
rect 33368 3190 33418 3206
rect 24627 3074 24644 3094
rect 24664 3074 24677 3094
rect 24627 3046 24677 3074
rect 22111 2974 22161 3002
rect 19837 2920 19887 2933
rect 20045 2920 20095 2933
rect 20263 2920 20313 2933
rect 22111 2954 22124 2974
rect 22144 2954 22161 2974
rect 22111 2925 22161 2954
rect 22329 2977 22379 3002
rect 22329 2957 22342 2977
rect 22362 2957 22379 2977
rect 22329 2925 22379 2957
rect 22537 2975 22587 3002
rect 22537 2955 22560 2975
rect 22580 2955 22587 2975
rect 22537 2925 22587 2955
rect 27285 3107 27335 3123
rect 27503 3107 27553 3123
rect 27711 3107 27761 3123
rect 28578 3105 28628 3135
rect 28578 3085 28585 3105
rect 28605 3085 28628 3105
rect 28578 3058 28628 3085
rect 28786 3103 28836 3135
rect 28786 3083 28803 3103
rect 28823 3083 28836 3103
rect 28786 3058 28836 3083
rect 29004 3106 29054 3135
rect 30852 3127 30902 3140
rect 31070 3127 31120 3140
rect 31278 3127 31328 3140
rect 33905 3182 33955 3195
rect 34113 3182 34163 3195
rect 34331 3182 34381 3195
rect 29004 3086 29021 3106
rect 29041 3086 29054 3106
rect 29004 3058 29054 3086
rect 26488 2986 26538 3014
rect 24201 2933 24251 2946
rect 24409 2933 24459 2946
rect 24627 2933 24677 2946
rect 26488 2966 26501 2986
rect 26521 2966 26538 2986
rect 26488 2937 26538 2966
rect 26706 2989 26756 3014
rect 26706 2969 26719 2989
rect 26739 2969 26756 2989
rect 26706 2937 26756 2969
rect 26914 2987 26964 3014
rect 26914 2967 26937 2987
rect 26957 2967 26964 2987
rect 26914 2937 26964 2967
rect 31649 3120 31699 3136
rect 31867 3120 31917 3136
rect 32075 3120 32125 3136
rect 32942 3118 32992 3148
rect 32942 3098 32949 3118
rect 32969 3098 32992 3118
rect 32942 3071 32992 3098
rect 33150 3116 33200 3148
rect 33150 3096 33167 3116
rect 33187 3096 33200 3116
rect 33150 3071 33200 3096
rect 33368 3119 33418 3148
rect 33368 3099 33385 3119
rect 33405 3099 33418 3119
rect 33368 3071 33418 3099
rect 30852 2999 30902 3027
rect 28578 2945 28628 2958
rect 28786 2945 28836 2958
rect 29004 2945 29054 2958
rect 30852 2979 30865 2999
rect 30885 2979 30902 2999
rect 30852 2950 30902 2979
rect 31070 3002 31120 3027
rect 31070 2982 31083 3002
rect 31103 2982 31120 3002
rect 31070 2950 31120 2982
rect 31278 3000 31328 3027
rect 31278 2980 31301 3000
rect 31321 2980 31328 3000
rect 31278 2950 31328 2980
rect 32942 2958 32992 2971
rect 33150 2958 33200 2971
rect 33368 2958 33418 2971
rect 17747 2854 17797 2870
rect 17965 2854 18015 2870
rect 18173 2854 18223 2870
rect 22111 2867 22161 2883
rect 22329 2867 22379 2883
rect 22537 2867 22587 2883
rect 26488 2879 26538 2895
rect 26706 2879 26756 2895
rect 26914 2879 26964 2895
rect 30852 2892 30902 2908
rect 31070 2892 31120 2908
rect 31278 2892 31328 2908
rect 3408 2758 3458 2774
rect 3616 2758 3666 2774
rect 3834 2758 3884 2774
rect 7772 2771 7822 2787
rect 7980 2771 8030 2787
rect 8198 2771 8248 2787
rect 12149 2783 12199 2799
rect 12357 2783 12407 2799
rect 12575 2783 12625 2799
rect 16513 2796 16563 2812
rect 16721 2796 16771 2812
rect 16939 2796 16989 2812
rect 1318 2695 1368 2708
rect 1536 2695 1586 2708
rect 1744 2695 1794 2708
rect 3408 2686 3458 2716
rect 3408 2666 3415 2686
rect 3435 2666 3458 2686
rect 3408 2639 3458 2666
rect 3616 2684 3666 2716
rect 3616 2664 3633 2684
rect 3653 2664 3666 2684
rect 3616 2639 3666 2664
rect 3834 2687 3884 2716
rect 3834 2667 3851 2687
rect 3871 2667 3884 2687
rect 5682 2708 5732 2721
rect 5900 2708 5950 2721
rect 6108 2708 6158 2721
rect 3834 2639 3884 2667
rect 1318 2567 1368 2595
rect 1318 2547 1331 2567
rect 1351 2547 1368 2567
rect 1318 2518 1368 2547
rect 1536 2570 1586 2595
rect 1536 2550 1549 2570
rect 1569 2550 1586 2570
rect 1536 2518 1586 2550
rect 1744 2568 1794 2595
rect 1744 2548 1767 2568
rect 1787 2548 1794 2568
rect 1744 2518 1794 2548
rect 2611 2530 2661 2546
rect 2819 2530 2869 2546
rect 3037 2530 3087 2546
rect 7772 2699 7822 2729
rect 7772 2679 7779 2699
rect 7799 2679 7822 2699
rect 7772 2652 7822 2679
rect 7980 2697 8030 2729
rect 7980 2677 7997 2697
rect 8017 2677 8030 2697
rect 7980 2652 8030 2677
rect 8198 2700 8248 2729
rect 8198 2680 8215 2700
rect 8235 2680 8248 2700
rect 10059 2720 10109 2733
rect 10277 2720 10327 2733
rect 10485 2720 10535 2733
rect 8198 2652 8248 2680
rect 5682 2580 5732 2608
rect 5682 2560 5695 2580
rect 5715 2560 5732 2580
rect 355 2471 405 2484
rect 573 2471 623 2484
rect 781 2471 831 2484
rect 3408 2526 3458 2539
rect 3616 2526 3666 2539
rect 3834 2526 3884 2539
rect 5682 2531 5732 2560
rect 5900 2583 5950 2608
rect 5900 2563 5913 2583
rect 5933 2563 5950 2583
rect 5900 2531 5950 2563
rect 6108 2581 6158 2608
rect 6108 2561 6131 2581
rect 6151 2561 6158 2581
rect 6108 2531 6158 2561
rect 6975 2543 7025 2559
rect 7183 2543 7233 2559
rect 7401 2543 7451 2559
rect 12149 2711 12199 2741
rect 12149 2691 12156 2711
rect 12176 2691 12199 2711
rect 12149 2664 12199 2691
rect 12357 2709 12407 2741
rect 12357 2689 12374 2709
rect 12394 2689 12407 2709
rect 12357 2664 12407 2689
rect 12575 2712 12625 2741
rect 12575 2692 12592 2712
rect 12612 2692 12625 2712
rect 14423 2733 14473 2746
rect 14641 2733 14691 2746
rect 14849 2733 14899 2746
rect 12575 2664 12625 2692
rect 10059 2592 10109 2620
rect 10059 2572 10072 2592
rect 10092 2572 10109 2592
rect 1318 2460 1368 2476
rect 1536 2460 1586 2476
rect 1744 2460 1794 2476
rect 2611 2458 2661 2488
rect 2611 2438 2618 2458
rect 2638 2438 2661 2458
rect 2611 2411 2661 2438
rect 2819 2456 2869 2488
rect 2819 2436 2836 2456
rect 2856 2436 2869 2456
rect 2819 2411 2869 2436
rect 3037 2459 3087 2488
rect 3037 2439 3054 2459
rect 3074 2439 3087 2459
rect 4719 2484 4769 2497
rect 4937 2484 4987 2497
rect 5145 2484 5195 2497
rect 7772 2539 7822 2552
rect 7980 2539 8030 2552
rect 8198 2539 8248 2552
rect 10059 2543 10109 2572
rect 10277 2595 10327 2620
rect 10277 2575 10290 2595
rect 10310 2575 10327 2595
rect 10277 2543 10327 2575
rect 10485 2593 10535 2620
rect 10485 2573 10508 2593
rect 10528 2573 10535 2593
rect 10485 2543 10535 2573
rect 11352 2555 11402 2571
rect 11560 2555 11610 2571
rect 11778 2555 11828 2571
rect 16513 2724 16563 2754
rect 16513 2704 16520 2724
rect 16540 2704 16563 2724
rect 16513 2677 16563 2704
rect 16721 2722 16771 2754
rect 16721 2702 16738 2722
rect 16758 2702 16771 2722
rect 16721 2677 16771 2702
rect 16939 2725 16989 2754
rect 20779 2770 20829 2786
rect 20987 2770 21037 2786
rect 21205 2770 21255 2786
rect 25143 2783 25193 2799
rect 25351 2783 25401 2799
rect 25569 2783 25619 2799
rect 29520 2795 29570 2811
rect 29728 2795 29778 2811
rect 29946 2795 29996 2811
rect 33884 2808 33934 2824
rect 34092 2808 34142 2824
rect 34310 2808 34360 2824
rect 16939 2705 16956 2725
rect 16976 2705 16989 2725
rect 16939 2677 16989 2705
rect 18689 2707 18739 2720
rect 18907 2707 18957 2720
rect 19115 2707 19165 2720
rect 14423 2605 14473 2633
rect 14423 2585 14436 2605
rect 14456 2585 14473 2605
rect 3037 2411 3087 2439
rect 355 2343 405 2371
rect 355 2323 368 2343
rect 388 2323 405 2343
rect 355 2294 405 2323
rect 573 2346 623 2371
rect 573 2326 586 2346
rect 606 2326 623 2346
rect 573 2294 623 2326
rect 781 2344 831 2371
rect 781 2324 804 2344
rect 824 2324 831 2344
rect 781 2294 831 2324
rect 5682 2473 5732 2489
rect 5900 2473 5950 2489
rect 6108 2473 6158 2489
rect 6975 2471 7025 2501
rect 6975 2451 6982 2471
rect 7002 2451 7025 2471
rect 6975 2424 7025 2451
rect 7183 2469 7233 2501
rect 7183 2449 7200 2469
rect 7220 2449 7233 2469
rect 7183 2424 7233 2449
rect 7401 2472 7451 2501
rect 7401 2452 7418 2472
rect 7438 2452 7451 2472
rect 9096 2496 9146 2509
rect 9314 2496 9364 2509
rect 9522 2496 9572 2509
rect 12149 2551 12199 2564
rect 12357 2551 12407 2564
rect 12575 2551 12625 2564
rect 14423 2556 14473 2585
rect 14641 2608 14691 2633
rect 14641 2588 14654 2608
rect 14674 2588 14691 2608
rect 14641 2556 14691 2588
rect 14849 2606 14899 2633
rect 14849 2586 14872 2606
rect 14892 2586 14899 2606
rect 14849 2556 14899 2586
rect 15716 2568 15766 2584
rect 15924 2568 15974 2584
rect 16142 2568 16192 2584
rect 20779 2698 20829 2728
rect 20779 2678 20786 2698
rect 20806 2678 20829 2698
rect 20779 2651 20829 2678
rect 20987 2696 21037 2728
rect 20987 2676 21004 2696
rect 21024 2676 21037 2696
rect 20987 2651 21037 2676
rect 21205 2699 21255 2728
rect 21205 2679 21222 2699
rect 21242 2679 21255 2699
rect 23053 2720 23103 2733
rect 23271 2720 23321 2733
rect 23479 2720 23529 2733
rect 21205 2651 21255 2679
rect 7401 2424 7451 2452
rect 3409 2346 3459 2362
rect 3617 2346 3667 2362
rect 3835 2346 3885 2362
rect 1153 2287 1203 2300
rect 1371 2287 1421 2300
rect 1579 2287 1629 2300
rect 2611 2298 2661 2311
rect 2819 2298 2869 2311
rect 3037 2298 3087 2311
rect 4719 2356 4769 2384
rect 355 2236 405 2252
rect 573 2236 623 2252
rect 781 2236 831 2252
rect 3409 2274 3459 2304
rect 3409 2254 3416 2274
rect 3436 2254 3459 2274
rect 3409 2227 3459 2254
rect 3617 2272 3667 2304
rect 3617 2252 3634 2272
rect 3654 2252 3667 2272
rect 3617 2227 3667 2252
rect 3835 2275 3885 2304
rect 3835 2255 3852 2275
rect 3872 2255 3885 2275
rect 4719 2336 4732 2356
rect 4752 2336 4769 2356
rect 4719 2307 4769 2336
rect 4937 2359 4987 2384
rect 4937 2339 4950 2359
rect 4970 2339 4987 2359
rect 4937 2307 4987 2339
rect 5145 2357 5195 2384
rect 5145 2337 5168 2357
rect 5188 2337 5195 2357
rect 5145 2307 5195 2337
rect 10059 2485 10109 2501
rect 10277 2485 10327 2501
rect 10485 2485 10535 2501
rect 11352 2483 11402 2513
rect 11352 2463 11359 2483
rect 11379 2463 11402 2483
rect 11352 2436 11402 2463
rect 11560 2481 11610 2513
rect 11560 2461 11577 2481
rect 11597 2461 11610 2481
rect 11560 2436 11610 2461
rect 11778 2484 11828 2513
rect 11778 2464 11795 2484
rect 11815 2464 11828 2484
rect 13460 2509 13510 2522
rect 13678 2509 13728 2522
rect 13886 2509 13936 2522
rect 16513 2564 16563 2577
rect 16721 2564 16771 2577
rect 16939 2564 16989 2577
rect 18689 2579 18739 2607
rect 18689 2559 18702 2579
rect 18722 2559 18739 2579
rect 18689 2530 18739 2559
rect 18907 2582 18957 2607
rect 18907 2562 18920 2582
rect 18940 2562 18957 2582
rect 18907 2530 18957 2562
rect 19115 2580 19165 2607
rect 19115 2560 19138 2580
rect 19158 2560 19165 2580
rect 19115 2530 19165 2560
rect 19982 2542 20032 2558
rect 20190 2542 20240 2558
rect 20408 2542 20458 2558
rect 25143 2711 25193 2741
rect 25143 2691 25150 2711
rect 25170 2691 25193 2711
rect 25143 2664 25193 2691
rect 25351 2709 25401 2741
rect 25351 2689 25368 2709
rect 25388 2689 25401 2709
rect 25351 2664 25401 2689
rect 25569 2712 25619 2741
rect 25569 2692 25586 2712
rect 25606 2692 25619 2712
rect 27430 2732 27480 2745
rect 27648 2732 27698 2745
rect 27856 2732 27906 2745
rect 25569 2664 25619 2692
rect 23053 2592 23103 2620
rect 23053 2572 23066 2592
rect 23086 2572 23103 2592
rect 11778 2436 11828 2464
rect 7773 2359 7823 2375
rect 7981 2359 8031 2375
rect 8199 2359 8249 2375
rect 3835 2227 3885 2255
rect 5517 2300 5567 2313
rect 5735 2300 5785 2313
rect 5943 2300 5993 2313
rect 6975 2311 7025 2324
rect 7183 2311 7233 2324
rect 7401 2311 7451 2324
rect 9096 2368 9146 2396
rect 4719 2249 4769 2265
rect 4937 2249 4987 2265
rect 5145 2249 5195 2265
rect 1153 2159 1203 2187
rect 1153 2139 1166 2159
rect 1186 2139 1203 2159
rect 1153 2110 1203 2139
rect 1371 2162 1421 2187
rect 1371 2142 1384 2162
rect 1404 2142 1421 2162
rect 1371 2110 1421 2142
rect 1579 2160 1629 2187
rect 1579 2140 1602 2160
rect 1622 2140 1629 2160
rect 1579 2110 1629 2140
rect 2512 2120 2562 2136
rect 2720 2120 2770 2136
rect 2938 2120 2988 2136
rect 7773 2287 7823 2317
rect 7773 2267 7780 2287
rect 7800 2267 7823 2287
rect 7773 2240 7823 2267
rect 7981 2285 8031 2317
rect 7981 2265 7998 2285
rect 8018 2265 8031 2285
rect 7981 2240 8031 2265
rect 8199 2288 8249 2317
rect 8199 2268 8216 2288
rect 8236 2268 8249 2288
rect 9096 2348 9109 2368
rect 9129 2348 9146 2368
rect 9096 2319 9146 2348
rect 9314 2371 9364 2396
rect 9314 2351 9327 2371
rect 9347 2351 9364 2371
rect 9314 2319 9364 2351
rect 9522 2369 9572 2396
rect 9522 2349 9545 2369
rect 9565 2349 9572 2369
rect 9522 2319 9572 2349
rect 14423 2498 14473 2514
rect 14641 2498 14691 2514
rect 14849 2498 14899 2514
rect 15716 2496 15766 2526
rect 15716 2476 15723 2496
rect 15743 2476 15766 2496
rect 15716 2449 15766 2476
rect 15924 2494 15974 2526
rect 15924 2474 15941 2494
rect 15961 2474 15974 2494
rect 15924 2449 15974 2474
rect 16142 2497 16192 2526
rect 16142 2477 16159 2497
rect 16179 2477 16192 2497
rect 16142 2449 16192 2477
rect 17726 2483 17776 2496
rect 17944 2483 17994 2496
rect 18152 2483 18202 2496
rect 20779 2538 20829 2551
rect 20987 2538 21037 2551
rect 21205 2538 21255 2551
rect 23053 2543 23103 2572
rect 23271 2595 23321 2620
rect 23271 2575 23284 2595
rect 23304 2575 23321 2595
rect 23271 2543 23321 2575
rect 23479 2593 23529 2620
rect 23479 2573 23502 2593
rect 23522 2573 23529 2593
rect 23479 2543 23529 2573
rect 24346 2555 24396 2571
rect 24554 2555 24604 2571
rect 24772 2555 24822 2571
rect 29520 2723 29570 2753
rect 29520 2703 29527 2723
rect 29547 2703 29570 2723
rect 29520 2676 29570 2703
rect 29728 2721 29778 2753
rect 29728 2701 29745 2721
rect 29765 2701 29778 2721
rect 29728 2676 29778 2701
rect 29946 2724 29996 2753
rect 29946 2704 29963 2724
rect 29983 2704 29996 2724
rect 31794 2745 31844 2758
rect 32012 2745 32062 2758
rect 32220 2745 32270 2758
rect 29946 2676 29996 2704
rect 27430 2604 27480 2632
rect 27430 2584 27443 2604
rect 27463 2584 27480 2604
rect 12150 2371 12200 2387
rect 12358 2371 12408 2387
rect 12576 2371 12626 2387
rect 8199 2240 8249 2268
rect 9894 2312 9944 2325
rect 10112 2312 10162 2325
rect 10320 2312 10370 2325
rect 11352 2323 11402 2336
rect 11560 2323 11610 2336
rect 11778 2323 11828 2336
rect 13460 2381 13510 2409
rect 9096 2261 9146 2277
rect 9314 2261 9364 2277
rect 9522 2261 9572 2277
rect 5517 2172 5567 2200
rect 356 2059 406 2072
rect 574 2059 624 2072
rect 782 2059 832 2072
rect 3409 2114 3459 2127
rect 3617 2114 3667 2127
rect 3835 2114 3885 2127
rect 5517 2152 5530 2172
rect 5550 2152 5567 2172
rect 5517 2123 5567 2152
rect 5735 2175 5785 2200
rect 5735 2155 5748 2175
rect 5768 2155 5785 2175
rect 5735 2123 5785 2155
rect 5943 2173 5993 2200
rect 5943 2153 5966 2173
rect 5986 2153 5993 2173
rect 5943 2123 5993 2153
rect 6876 2133 6926 2149
rect 7084 2133 7134 2149
rect 7302 2133 7352 2149
rect 12150 2299 12200 2329
rect 12150 2279 12157 2299
rect 12177 2279 12200 2299
rect 12150 2252 12200 2279
rect 12358 2297 12408 2329
rect 12358 2277 12375 2297
rect 12395 2277 12408 2297
rect 12358 2252 12408 2277
rect 12576 2300 12626 2329
rect 12576 2280 12593 2300
rect 12613 2280 12626 2300
rect 13460 2361 13473 2381
rect 13493 2361 13510 2381
rect 13460 2332 13510 2361
rect 13678 2384 13728 2409
rect 13678 2364 13691 2384
rect 13711 2364 13728 2384
rect 13678 2332 13728 2364
rect 13886 2382 13936 2409
rect 13886 2362 13909 2382
rect 13929 2362 13936 2382
rect 13886 2332 13936 2362
rect 16514 2384 16564 2400
rect 16722 2384 16772 2400
rect 16940 2384 16990 2400
rect 12576 2252 12626 2280
rect 14258 2325 14308 2338
rect 14476 2325 14526 2338
rect 14684 2325 14734 2338
rect 15716 2336 15766 2349
rect 15924 2336 15974 2349
rect 16142 2336 16192 2349
rect 18689 2472 18739 2488
rect 18907 2472 18957 2488
rect 19115 2472 19165 2488
rect 19982 2470 20032 2500
rect 19982 2450 19989 2470
rect 20009 2450 20032 2470
rect 19982 2423 20032 2450
rect 20190 2468 20240 2500
rect 20190 2448 20207 2468
rect 20227 2448 20240 2468
rect 20190 2423 20240 2448
rect 20408 2471 20458 2500
rect 20408 2451 20425 2471
rect 20445 2451 20458 2471
rect 22090 2496 22140 2509
rect 22308 2496 22358 2509
rect 22516 2496 22566 2509
rect 25143 2551 25193 2564
rect 25351 2551 25401 2564
rect 25569 2551 25619 2564
rect 27430 2555 27480 2584
rect 27648 2607 27698 2632
rect 27648 2587 27661 2607
rect 27681 2587 27698 2607
rect 27648 2555 27698 2587
rect 27856 2605 27906 2632
rect 27856 2585 27879 2605
rect 27899 2585 27906 2605
rect 27856 2555 27906 2585
rect 28723 2567 28773 2583
rect 28931 2567 28981 2583
rect 29149 2567 29199 2583
rect 33884 2736 33934 2766
rect 33884 2716 33891 2736
rect 33911 2716 33934 2736
rect 33884 2689 33934 2716
rect 34092 2734 34142 2766
rect 34092 2714 34109 2734
rect 34129 2714 34142 2734
rect 34092 2689 34142 2714
rect 34310 2737 34360 2766
rect 34310 2717 34327 2737
rect 34347 2717 34360 2737
rect 34310 2689 34360 2717
rect 31794 2617 31844 2645
rect 31794 2597 31807 2617
rect 31827 2597 31844 2617
rect 20408 2423 20458 2451
rect 13460 2274 13510 2290
rect 13678 2274 13728 2290
rect 13886 2274 13936 2290
rect 9894 2184 9944 2212
rect 1153 2052 1203 2068
rect 1371 2052 1421 2068
rect 1579 2052 1629 2068
rect 2512 2048 2562 2078
rect 2512 2028 2519 2048
rect 2539 2028 2562 2048
rect 2512 2001 2562 2028
rect 2720 2046 2770 2078
rect 2720 2026 2737 2046
rect 2757 2026 2770 2046
rect 2720 2001 2770 2026
rect 2938 2049 2988 2078
rect 4720 2072 4770 2085
rect 4938 2072 4988 2085
rect 5146 2072 5196 2085
rect 7773 2127 7823 2140
rect 7981 2127 8031 2140
rect 8199 2127 8249 2140
rect 9894 2164 9907 2184
rect 9927 2164 9944 2184
rect 9894 2135 9944 2164
rect 10112 2187 10162 2212
rect 10112 2167 10125 2187
rect 10145 2167 10162 2187
rect 10112 2135 10162 2167
rect 10320 2185 10370 2212
rect 10320 2165 10343 2185
rect 10363 2165 10370 2185
rect 10320 2135 10370 2165
rect 11253 2145 11303 2161
rect 11461 2145 11511 2161
rect 11679 2145 11729 2161
rect 16514 2312 16564 2342
rect 16514 2292 16521 2312
rect 16541 2292 16564 2312
rect 16514 2265 16564 2292
rect 16722 2310 16772 2342
rect 16722 2290 16739 2310
rect 16759 2290 16772 2310
rect 16722 2265 16772 2290
rect 16940 2313 16990 2342
rect 16940 2293 16957 2313
rect 16977 2293 16990 2313
rect 17726 2355 17776 2383
rect 16940 2265 16990 2293
rect 17726 2335 17739 2355
rect 17759 2335 17776 2355
rect 17726 2306 17776 2335
rect 17944 2358 17994 2383
rect 17944 2338 17957 2358
rect 17977 2338 17994 2358
rect 17944 2306 17994 2338
rect 18152 2356 18202 2383
rect 18152 2336 18175 2356
rect 18195 2336 18202 2356
rect 18152 2306 18202 2336
rect 23053 2485 23103 2501
rect 23271 2485 23321 2501
rect 23479 2485 23529 2501
rect 24346 2483 24396 2513
rect 24346 2463 24353 2483
rect 24373 2463 24396 2483
rect 24346 2436 24396 2463
rect 24554 2481 24604 2513
rect 24554 2461 24571 2481
rect 24591 2461 24604 2481
rect 24554 2436 24604 2461
rect 24772 2484 24822 2513
rect 24772 2464 24789 2484
rect 24809 2464 24822 2484
rect 26467 2508 26517 2521
rect 26685 2508 26735 2521
rect 26893 2508 26943 2521
rect 29520 2563 29570 2576
rect 29728 2563 29778 2576
rect 29946 2563 29996 2576
rect 31794 2568 31844 2597
rect 32012 2620 32062 2645
rect 32012 2600 32025 2620
rect 32045 2600 32062 2620
rect 32012 2568 32062 2600
rect 32220 2618 32270 2645
rect 32220 2598 32243 2618
rect 32263 2598 32270 2618
rect 32220 2568 32270 2598
rect 33087 2580 33137 2596
rect 33295 2580 33345 2596
rect 33513 2580 33563 2596
rect 24772 2436 24822 2464
rect 20780 2358 20830 2374
rect 20988 2358 21038 2374
rect 21206 2358 21256 2374
rect 14258 2197 14308 2225
rect 2938 2029 2955 2049
rect 2975 2029 2988 2049
rect 2938 2001 2988 2029
rect 356 1931 406 1959
rect 356 1911 369 1931
rect 389 1911 406 1931
rect 356 1882 406 1911
rect 574 1934 624 1959
rect 574 1914 587 1934
rect 607 1914 624 1934
rect 574 1882 624 1914
rect 782 1932 832 1959
rect 782 1912 805 1932
rect 825 1912 832 1932
rect 782 1882 832 1912
rect 5517 2065 5567 2081
rect 5735 2065 5785 2081
rect 5943 2065 5993 2081
rect 6876 2061 6926 2091
rect 6876 2041 6883 2061
rect 6903 2041 6926 2061
rect 6876 2014 6926 2041
rect 7084 2059 7134 2091
rect 7084 2039 7101 2059
rect 7121 2039 7134 2059
rect 7084 2014 7134 2039
rect 7302 2062 7352 2091
rect 9097 2084 9147 2097
rect 9315 2084 9365 2097
rect 9523 2084 9573 2097
rect 12150 2139 12200 2152
rect 12358 2139 12408 2152
rect 12576 2139 12626 2152
rect 14258 2177 14271 2197
rect 14291 2177 14308 2197
rect 14258 2148 14308 2177
rect 14476 2200 14526 2225
rect 14476 2180 14489 2200
rect 14509 2180 14526 2200
rect 14476 2148 14526 2180
rect 14684 2198 14734 2225
rect 14684 2178 14707 2198
rect 14727 2178 14734 2198
rect 14684 2148 14734 2178
rect 15617 2158 15667 2174
rect 15825 2158 15875 2174
rect 16043 2158 16093 2174
rect 18524 2299 18574 2312
rect 18742 2299 18792 2312
rect 18950 2299 19000 2312
rect 19982 2310 20032 2323
rect 20190 2310 20240 2323
rect 20408 2310 20458 2323
rect 22090 2368 22140 2396
rect 17726 2248 17776 2264
rect 17944 2248 17994 2264
rect 18152 2248 18202 2264
rect 20780 2286 20830 2316
rect 20780 2266 20787 2286
rect 20807 2266 20830 2286
rect 20780 2239 20830 2266
rect 20988 2284 21038 2316
rect 20988 2264 21005 2284
rect 21025 2264 21038 2284
rect 20988 2239 21038 2264
rect 21206 2287 21256 2316
rect 21206 2267 21223 2287
rect 21243 2267 21256 2287
rect 22090 2348 22103 2368
rect 22123 2348 22140 2368
rect 22090 2319 22140 2348
rect 22308 2371 22358 2396
rect 22308 2351 22321 2371
rect 22341 2351 22358 2371
rect 22308 2319 22358 2351
rect 22516 2369 22566 2396
rect 22516 2349 22539 2369
rect 22559 2349 22566 2369
rect 22516 2319 22566 2349
rect 27430 2497 27480 2513
rect 27648 2497 27698 2513
rect 27856 2497 27906 2513
rect 28723 2495 28773 2525
rect 28723 2475 28730 2495
rect 28750 2475 28773 2495
rect 28723 2448 28773 2475
rect 28931 2493 28981 2525
rect 28931 2473 28948 2493
rect 28968 2473 28981 2493
rect 28931 2448 28981 2473
rect 29149 2496 29199 2525
rect 29149 2476 29166 2496
rect 29186 2476 29199 2496
rect 30831 2521 30881 2534
rect 31049 2521 31099 2534
rect 31257 2521 31307 2534
rect 33884 2576 33934 2589
rect 34092 2576 34142 2589
rect 34310 2576 34360 2589
rect 29149 2448 29199 2476
rect 25144 2371 25194 2387
rect 25352 2371 25402 2387
rect 25570 2371 25620 2387
rect 21206 2239 21256 2267
rect 22888 2312 22938 2325
rect 23106 2312 23156 2325
rect 23314 2312 23364 2325
rect 24346 2323 24396 2336
rect 24554 2323 24604 2336
rect 24772 2323 24822 2336
rect 26467 2380 26517 2408
rect 22090 2261 22140 2277
rect 22308 2261 22358 2277
rect 22516 2261 22566 2277
rect 7302 2042 7319 2062
rect 7339 2042 7352 2062
rect 7302 2014 7352 2042
rect 4720 1944 4770 1972
rect 2512 1888 2562 1901
rect 2720 1888 2770 1901
rect 2938 1888 2988 1901
rect 4720 1924 4733 1944
rect 4753 1924 4770 1944
rect 4720 1895 4770 1924
rect 4938 1947 4988 1972
rect 4938 1927 4951 1947
rect 4971 1927 4988 1947
rect 4938 1895 4988 1927
rect 5146 1945 5196 1972
rect 5146 1925 5169 1945
rect 5189 1925 5196 1945
rect 5146 1895 5196 1925
rect 9894 2077 9944 2093
rect 10112 2077 10162 2093
rect 10320 2077 10370 2093
rect 11253 2073 11303 2103
rect 11253 2053 11260 2073
rect 11280 2053 11303 2073
rect 11253 2026 11303 2053
rect 11461 2071 11511 2103
rect 11461 2051 11478 2071
rect 11498 2051 11511 2071
rect 11461 2026 11511 2051
rect 11679 2074 11729 2103
rect 13461 2097 13511 2110
rect 13679 2097 13729 2110
rect 13887 2097 13937 2110
rect 16514 2152 16564 2165
rect 16722 2152 16772 2165
rect 16940 2152 16990 2165
rect 18524 2171 18574 2199
rect 18524 2151 18537 2171
rect 18557 2151 18574 2171
rect 18524 2122 18574 2151
rect 18742 2174 18792 2199
rect 18742 2154 18755 2174
rect 18775 2154 18792 2174
rect 18742 2122 18792 2154
rect 18950 2172 19000 2199
rect 18950 2152 18973 2172
rect 18993 2152 19000 2172
rect 18950 2122 19000 2152
rect 19883 2132 19933 2148
rect 20091 2132 20141 2148
rect 20309 2132 20359 2148
rect 25144 2299 25194 2329
rect 25144 2279 25151 2299
rect 25171 2279 25194 2299
rect 25144 2252 25194 2279
rect 25352 2297 25402 2329
rect 25352 2277 25369 2297
rect 25389 2277 25402 2297
rect 25352 2252 25402 2277
rect 25570 2300 25620 2329
rect 25570 2280 25587 2300
rect 25607 2280 25620 2300
rect 26467 2360 26480 2380
rect 26500 2360 26517 2380
rect 26467 2331 26517 2360
rect 26685 2383 26735 2408
rect 26685 2363 26698 2383
rect 26718 2363 26735 2383
rect 26685 2331 26735 2363
rect 26893 2381 26943 2408
rect 26893 2361 26916 2381
rect 26936 2361 26943 2381
rect 26893 2331 26943 2361
rect 31794 2510 31844 2526
rect 32012 2510 32062 2526
rect 32220 2510 32270 2526
rect 33087 2508 33137 2538
rect 33087 2488 33094 2508
rect 33114 2488 33137 2508
rect 33087 2461 33137 2488
rect 33295 2506 33345 2538
rect 33295 2486 33312 2506
rect 33332 2486 33345 2506
rect 33295 2461 33345 2486
rect 33513 2509 33563 2538
rect 33513 2489 33530 2509
rect 33550 2489 33563 2509
rect 33513 2461 33563 2489
rect 29521 2383 29571 2399
rect 29729 2383 29779 2399
rect 29947 2383 29997 2399
rect 25570 2252 25620 2280
rect 27265 2324 27315 2337
rect 27483 2324 27533 2337
rect 27691 2324 27741 2337
rect 28723 2335 28773 2348
rect 28931 2335 28981 2348
rect 29149 2335 29199 2348
rect 30831 2393 30881 2421
rect 26467 2273 26517 2289
rect 26685 2273 26735 2289
rect 26893 2273 26943 2289
rect 22888 2184 22938 2212
rect 11679 2054 11696 2074
rect 11716 2054 11729 2074
rect 11679 2026 11729 2054
rect 9097 1956 9147 1984
rect 6876 1901 6926 1914
rect 7084 1901 7134 1914
rect 7302 1901 7352 1914
rect 9097 1936 9110 1956
rect 9130 1936 9147 1956
rect 9097 1907 9147 1936
rect 9315 1959 9365 1984
rect 9315 1939 9328 1959
rect 9348 1939 9365 1959
rect 9315 1907 9365 1939
rect 9523 1957 9573 1984
rect 9523 1937 9546 1957
rect 9566 1937 9573 1957
rect 9523 1907 9573 1937
rect 14258 2090 14308 2106
rect 14476 2090 14526 2106
rect 14684 2090 14734 2106
rect 15617 2086 15667 2116
rect 15617 2066 15624 2086
rect 15644 2066 15667 2086
rect 15617 2039 15667 2066
rect 15825 2084 15875 2116
rect 15825 2064 15842 2084
rect 15862 2064 15875 2084
rect 15825 2039 15875 2064
rect 16043 2087 16093 2116
rect 16043 2067 16060 2087
rect 16080 2067 16093 2087
rect 16043 2039 16093 2067
rect 17727 2071 17777 2084
rect 17945 2071 17995 2084
rect 18153 2071 18203 2084
rect 20780 2126 20830 2139
rect 20988 2126 21038 2139
rect 21206 2126 21256 2139
rect 22888 2164 22901 2184
rect 22921 2164 22938 2184
rect 22888 2135 22938 2164
rect 23106 2187 23156 2212
rect 23106 2167 23119 2187
rect 23139 2167 23156 2187
rect 23106 2135 23156 2167
rect 23314 2185 23364 2212
rect 23314 2165 23337 2185
rect 23357 2165 23364 2185
rect 23314 2135 23364 2165
rect 24247 2145 24297 2161
rect 24455 2145 24505 2161
rect 24673 2145 24723 2161
rect 29521 2311 29571 2341
rect 29521 2291 29528 2311
rect 29548 2291 29571 2311
rect 29521 2264 29571 2291
rect 29729 2309 29779 2341
rect 29729 2289 29746 2309
rect 29766 2289 29779 2309
rect 29729 2264 29779 2289
rect 29947 2312 29997 2341
rect 29947 2292 29964 2312
rect 29984 2292 29997 2312
rect 30831 2373 30844 2393
rect 30864 2373 30881 2393
rect 30831 2344 30881 2373
rect 31049 2396 31099 2421
rect 31049 2376 31062 2396
rect 31082 2376 31099 2396
rect 31049 2344 31099 2376
rect 31257 2394 31307 2421
rect 31257 2374 31280 2394
rect 31300 2374 31307 2394
rect 31257 2344 31307 2374
rect 33885 2396 33935 2412
rect 34093 2396 34143 2412
rect 34311 2396 34361 2412
rect 29947 2264 29997 2292
rect 31629 2337 31679 2350
rect 31847 2337 31897 2350
rect 32055 2337 32105 2350
rect 33087 2348 33137 2361
rect 33295 2348 33345 2361
rect 33513 2348 33563 2361
rect 30831 2286 30881 2302
rect 31049 2286 31099 2302
rect 31257 2286 31307 2302
rect 27265 2196 27315 2224
rect 13461 1969 13511 1997
rect 11253 1913 11303 1926
rect 11461 1913 11511 1926
rect 11679 1913 11729 1926
rect 13461 1949 13474 1969
rect 13494 1949 13511 1969
rect 13461 1920 13511 1949
rect 13679 1972 13729 1997
rect 13679 1952 13692 1972
rect 13712 1952 13729 1972
rect 13679 1920 13729 1952
rect 13887 1970 13937 1997
rect 13887 1950 13910 1970
rect 13930 1950 13937 1970
rect 13887 1920 13937 1950
rect 18524 2064 18574 2080
rect 18742 2064 18792 2080
rect 18950 2064 19000 2080
rect 19883 2060 19933 2090
rect 19883 2040 19890 2060
rect 19910 2040 19933 2060
rect 19883 2013 19933 2040
rect 20091 2058 20141 2090
rect 20091 2038 20108 2058
rect 20128 2038 20141 2058
rect 20091 2013 20141 2038
rect 20309 2061 20359 2090
rect 22091 2084 22141 2097
rect 22309 2084 22359 2097
rect 22517 2084 22567 2097
rect 25144 2139 25194 2152
rect 25352 2139 25402 2152
rect 25570 2139 25620 2152
rect 27265 2176 27278 2196
rect 27298 2176 27315 2196
rect 27265 2147 27315 2176
rect 27483 2199 27533 2224
rect 27483 2179 27496 2199
rect 27516 2179 27533 2199
rect 27483 2147 27533 2179
rect 27691 2197 27741 2224
rect 27691 2177 27714 2197
rect 27734 2177 27741 2197
rect 27691 2147 27741 2177
rect 28624 2157 28674 2173
rect 28832 2157 28882 2173
rect 29050 2157 29100 2173
rect 33885 2324 33935 2354
rect 33885 2304 33892 2324
rect 33912 2304 33935 2324
rect 33885 2277 33935 2304
rect 34093 2322 34143 2354
rect 34093 2302 34110 2322
rect 34130 2302 34143 2322
rect 34093 2277 34143 2302
rect 34311 2325 34361 2354
rect 34311 2305 34328 2325
rect 34348 2305 34361 2325
rect 34311 2277 34361 2305
rect 31629 2209 31679 2237
rect 20309 2041 20326 2061
rect 20346 2041 20359 2061
rect 20309 2013 20359 2041
rect 15617 1926 15667 1939
rect 15825 1926 15875 1939
rect 16043 1926 16093 1939
rect 17727 1943 17777 1971
rect 17727 1923 17740 1943
rect 17760 1923 17777 1943
rect 356 1824 406 1840
rect 574 1824 624 1840
rect 782 1824 832 1840
rect 4720 1837 4770 1853
rect 4938 1837 4988 1853
rect 5146 1837 5196 1853
rect 9097 1849 9147 1865
rect 9315 1849 9365 1865
rect 9523 1849 9573 1865
rect 13461 1862 13511 1878
rect 13679 1862 13729 1878
rect 13887 1862 13937 1878
rect 17727 1894 17777 1923
rect 17945 1946 17995 1971
rect 17945 1926 17958 1946
rect 17978 1926 17995 1946
rect 17945 1894 17995 1926
rect 18153 1944 18203 1971
rect 18153 1924 18176 1944
rect 18196 1924 18203 1944
rect 18153 1894 18203 1924
rect 22888 2077 22938 2093
rect 23106 2077 23156 2093
rect 23314 2077 23364 2093
rect 24247 2073 24297 2103
rect 24247 2053 24254 2073
rect 24274 2053 24297 2073
rect 24247 2026 24297 2053
rect 24455 2071 24505 2103
rect 24455 2051 24472 2071
rect 24492 2051 24505 2071
rect 24455 2026 24505 2051
rect 24673 2074 24723 2103
rect 26468 2096 26518 2109
rect 26686 2096 26736 2109
rect 26894 2096 26944 2109
rect 29521 2151 29571 2164
rect 29729 2151 29779 2164
rect 29947 2151 29997 2164
rect 31629 2189 31642 2209
rect 31662 2189 31679 2209
rect 31629 2160 31679 2189
rect 31847 2212 31897 2237
rect 31847 2192 31860 2212
rect 31880 2192 31897 2212
rect 31847 2160 31897 2192
rect 32055 2210 32105 2237
rect 32055 2190 32078 2210
rect 32098 2190 32105 2210
rect 32055 2160 32105 2190
rect 32988 2170 33038 2186
rect 33196 2170 33246 2186
rect 33414 2170 33464 2186
rect 24673 2054 24690 2074
rect 24710 2054 24723 2074
rect 24673 2026 24723 2054
rect 22091 1956 22141 1984
rect 19883 1900 19933 1913
rect 20091 1900 20141 1913
rect 20309 1900 20359 1913
rect 22091 1936 22104 1956
rect 22124 1936 22141 1956
rect 22091 1907 22141 1936
rect 22309 1959 22359 1984
rect 22309 1939 22322 1959
rect 22342 1939 22359 1959
rect 22309 1907 22359 1939
rect 22517 1957 22567 1984
rect 22517 1937 22540 1957
rect 22560 1937 22567 1957
rect 22517 1907 22567 1937
rect 27265 2089 27315 2105
rect 27483 2089 27533 2105
rect 27691 2089 27741 2105
rect 28624 2085 28674 2115
rect 28624 2065 28631 2085
rect 28651 2065 28674 2085
rect 28624 2038 28674 2065
rect 28832 2083 28882 2115
rect 28832 2063 28849 2083
rect 28869 2063 28882 2083
rect 28832 2038 28882 2063
rect 29050 2086 29100 2115
rect 30832 2109 30882 2122
rect 31050 2109 31100 2122
rect 31258 2109 31308 2122
rect 33885 2164 33935 2177
rect 34093 2164 34143 2177
rect 34311 2164 34361 2177
rect 29050 2066 29067 2086
rect 29087 2066 29100 2086
rect 29050 2038 29100 2066
rect 26468 1968 26518 1996
rect 24247 1913 24297 1926
rect 24455 1913 24505 1926
rect 24673 1913 24723 1926
rect 26468 1948 26481 1968
rect 26501 1948 26518 1968
rect 26468 1919 26518 1948
rect 26686 1971 26736 1996
rect 26686 1951 26699 1971
rect 26719 1951 26736 1971
rect 26686 1919 26736 1951
rect 26894 1969 26944 1996
rect 26894 1949 26917 1969
rect 26937 1949 26944 1969
rect 26894 1919 26944 1949
rect 31629 2102 31679 2118
rect 31847 2102 31897 2118
rect 32055 2102 32105 2118
rect 32988 2098 33038 2128
rect 32988 2078 32995 2098
rect 33015 2078 33038 2098
rect 32988 2051 33038 2078
rect 33196 2096 33246 2128
rect 33196 2076 33213 2096
rect 33233 2076 33246 2096
rect 33196 2051 33246 2076
rect 33414 2099 33464 2128
rect 33414 2079 33431 2099
rect 33451 2079 33464 2099
rect 33414 2051 33464 2079
rect 30832 1981 30882 2009
rect 28624 1925 28674 1938
rect 28832 1925 28882 1938
rect 29050 1925 29100 1938
rect 30832 1961 30845 1981
rect 30865 1961 30882 1981
rect 30832 1932 30882 1961
rect 31050 1984 31100 2009
rect 31050 1964 31063 1984
rect 31083 1964 31100 1984
rect 31050 1932 31100 1964
rect 31258 1982 31308 2009
rect 31258 1962 31281 1982
rect 31301 1962 31308 1982
rect 31258 1932 31308 1962
rect 32988 1938 33038 1951
rect 33196 1938 33246 1951
rect 33414 1938 33464 1951
rect 17727 1836 17777 1852
rect 17945 1836 17995 1852
rect 18153 1836 18203 1852
rect 22091 1849 22141 1865
rect 22309 1849 22359 1865
rect 22517 1849 22567 1865
rect 26468 1861 26518 1877
rect 26686 1861 26736 1877
rect 26894 1861 26944 1877
rect 30832 1874 30882 1890
rect 31050 1874 31100 1890
rect 31258 1874 31308 1890
rect 3391 1740 3441 1756
rect 3599 1740 3649 1756
rect 3817 1740 3867 1756
rect 7755 1753 7805 1769
rect 7963 1753 8013 1769
rect 8181 1753 8231 1769
rect 12132 1765 12182 1781
rect 12340 1765 12390 1781
rect 12558 1765 12608 1781
rect 16496 1778 16546 1794
rect 16704 1778 16754 1794
rect 16922 1778 16972 1794
rect 1235 1679 1285 1692
rect 1453 1679 1503 1692
rect 1661 1679 1711 1692
rect 3391 1668 3441 1698
rect 3391 1648 3398 1668
rect 3418 1648 3441 1668
rect 3391 1621 3441 1648
rect 3599 1666 3649 1698
rect 3599 1646 3616 1666
rect 3636 1646 3649 1666
rect 3599 1621 3649 1646
rect 3817 1669 3867 1698
rect 3817 1649 3834 1669
rect 3854 1649 3867 1669
rect 5599 1692 5649 1705
rect 5817 1692 5867 1705
rect 6025 1692 6075 1705
rect 3817 1621 3867 1649
rect 1235 1551 1285 1579
rect 1235 1531 1248 1551
rect 1268 1531 1285 1551
rect 1235 1502 1285 1531
rect 1453 1554 1503 1579
rect 1453 1534 1466 1554
rect 1486 1534 1503 1554
rect 1453 1502 1503 1534
rect 1661 1552 1711 1579
rect 1661 1532 1684 1552
rect 1704 1532 1711 1552
rect 1661 1502 1711 1532
rect 2594 1512 2644 1528
rect 2802 1512 2852 1528
rect 3020 1512 3070 1528
rect 7755 1681 7805 1711
rect 7755 1661 7762 1681
rect 7782 1661 7805 1681
rect 7755 1634 7805 1661
rect 7963 1679 8013 1711
rect 7963 1659 7980 1679
rect 8000 1659 8013 1679
rect 7963 1634 8013 1659
rect 8181 1682 8231 1711
rect 8181 1662 8198 1682
rect 8218 1662 8231 1682
rect 9976 1704 10026 1717
rect 10194 1704 10244 1717
rect 10402 1704 10452 1717
rect 8181 1634 8231 1662
rect 5599 1564 5649 1592
rect 5599 1544 5612 1564
rect 5632 1544 5649 1564
rect 338 1453 388 1466
rect 556 1453 606 1466
rect 764 1453 814 1466
rect 3391 1508 3441 1521
rect 3599 1508 3649 1521
rect 3817 1508 3867 1521
rect 5599 1515 5649 1544
rect 5817 1567 5867 1592
rect 5817 1547 5830 1567
rect 5850 1547 5867 1567
rect 5817 1515 5867 1547
rect 6025 1565 6075 1592
rect 6025 1545 6048 1565
rect 6068 1545 6075 1565
rect 6025 1515 6075 1545
rect 6958 1525 7008 1541
rect 7166 1525 7216 1541
rect 7384 1525 7434 1541
rect 12132 1693 12182 1723
rect 12132 1673 12139 1693
rect 12159 1673 12182 1693
rect 12132 1646 12182 1673
rect 12340 1691 12390 1723
rect 12340 1671 12357 1691
rect 12377 1671 12390 1691
rect 12340 1646 12390 1671
rect 12558 1694 12608 1723
rect 12558 1674 12575 1694
rect 12595 1674 12608 1694
rect 14340 1717 14390 1730
rect 14558 1717 14608 1730
rect 14766 1717 14816 1730
rect 12558 1646 12608 1674
rect 9976 1576 10026 1604
rect 9976 1556 9989 1576
rect 10009 1556 10026 1576
rect 1235 1444 1285 1460
rect 1453 1444 1503 1460
rect 1661 1444 1711 1460
rect 2594 1440 2644 1470
rect 2594 1420 2601 1440
rect 2621 1420 2644 1440
rect 2594 1393 2644 1420
rect 2802 1438 2852 1470
rect 2802 1418 2819 1438
rect 2839 1418 2852 1438
rect 2802 1393 2852 1418
rect 3020 1441 3070 1470
rect 3020 1421 3037 1441
rect 3057 1421 3070 1441
rect 4702 1466 4752 1479
rect 4920 1466 4970 1479
rect 5128 1466 5178 1479
rect 7755 1521 7805 1534
rect 7963 1521 8013 1534
rect 8181 1521 8231 1534
rect 9976 1527 10026 1556
rect 10194 1579 10244 1604
rect 10194 1559 10207 1579
rect 10227 1559 10244 1579
rect 10194 1527 10244 1559
rect 10402 1577 10452 1604
rect 10402 1557 10425 1577
rect 10445 1557 10452 1577
rect 10402 1527 10452 1557
rect 11335 1537 11385 1553
rect 11543 1537 11593 1553
rect 11761 1537 11811 1553
rect 16496 1706 16546 1736
rect 16496 1686 16503 1706
rect 16523 1686 16546 1706
rect 16496 1659 16546 1686
rect 16704 1704 16754 1736
rect 16704 1684 16721 1704
rect 16741 1684 16754 1704
rect 16704 1659 16754 1684
rect 16922 1707 16972 1736
rect 20762 1752 20812 1768
rect 20970 1752 21020 1768
rect 21188 1752 21238 1768
rect 25126 1765 25176 1781
rect 25334 1765 25384 1781
rect 25552 1765 25602 1781
rect 29503 1777 29553 1793
rect 29711 1777 29761 1793
rect 29929 1777 29979 1793
rect 33867 1790 33917 1806
rect 34075 1790 34125 1806
rect 34293 1790 34343 1806
rect 16922 1687 16939 1707
rect 16959 1687 16972 1707
rect 16922 1659 16972 1687
rect 18606 1691 18656 1704
rect 18824 1691 18874 1704
rect 19032 1691 19082 1704
rect 14340 1589 14390 1617
rect 14340 1569 14353 1589
rect 14373 1569 14390 1589
rect 3020 1393 3070 1421
rect 338 1325 388 1353
rect 338 1305 351 1325
rect 371 1305 388 1325
rect 338 1276 388 1305
rect 556 1328 606 1353
rect 556 1308 569 1328
rect 589 1308 606 1328
rect 556 1276 606 1308
rect 764 1326 814 1353
rect 764 1306 787 1326
rect 807 1306 814 1326
rect 764 1276 814 1306
rect 5599 1457 5649 1473
rect 5817 1457 5867 1473
rect 6025 1457 6075 1473
rect 6958 1453 7008 1483
rect 6958 1433 6965 1453
rect 6985 1433 7008 1453
rect 6958 1406 7008 1433
rect 7166 1451 7216 1483
rect 7166 1431 7183 1451
rect 7203 1431 7216 1451
rect 7166 1406 7216 1431
rect 7384 1454 7434 1483
rect 7384 1434 7401 1454
rect 7421 1434 7434 1454
rect 9079 1478 9129 1491
rect 9297 1478 9347 1491
rect 9505 1478 9555 1491
rect 12132 1533 12182 1546
rect 12340 1533 12390 1546
rect 12558 1533 12608 1546
rect 14340 1540 14390 1569
rect 14558 1592 14608 1617
rect 14558 1572 14571 1592
rect 14591 1572 14608 1592
rect 14558 1540 14608 1572
rect 14766 1590 14816 1617
rect 14766 1570 14789 1590
rect 14809 1570 14816 1590
rect 14766 1540 14816 1570
rect 15699 1550 15749 1566
rect 15907 1550 15957 1566
rect 16125 1550 16175 1566
rect 20762 1680 20812 1710
rect 20762 1660 20769 1680
rect 20789 1660 20812 1680
rect 20762 1633 20812 1660
rect 20970 1678 21020 1710
rect 20970 1658 20987 1678
rect 21007 1658 21020 1678
rect 20970 1633 21020 1658
rect 21188 1681 21238 1710
rect 21188 1661 21205 1681
rect 21225 1661 21238 1681
rect 22970 1704 23020 1717
rect 23188 1704 23238 1717
rect 23396 1704 23446 1717
rect 21188 1633 21238 1661
rect 7384 1406 7434 1434
rect 3392 1328 3442 1344
rect 3600 1328 3650 1344
rect 3818 1328 3868 1344
rect 1136 1269 1186 1282
rect 1354 1269 1404 1282
rect 1562 1269 1612 1282
rect 2594 1280 2644 1293
rect 2802 1280 2852 1293
rect 3020 1280 3070 1293
rect 4702 1338 4752 1366
rect 338 1218 388 1234
rect 556 1218 606 1234
rect 764 1218 814 1234
rect 3392 1256 3442 1286
rect 3392 1236 3399 1256
rect 3419 1236 3442 1256
rect 3392 1209 3442 1236
rect 3600 1254 3650 1286
rect 3600 1234 3617 1254
rect 3637 1234 3650 1254
rect 3600 1209 3650 1234
rect 3818 1257 3868 1286
rect 3818 1237 3835 1257
rect 3855 1237 3868 1257
rect 4702 1318 4715 1338
rect 4735 1318 4752 1338
rect 4702 1289 4752 1318
rect 4920 1341 4970 1366
rect 4920 1321 4933 1341
rect 4953 1321 4970 1341
rect 4920 1289 4970 1321
rect 5128 1339 5178 1366
rect 5128 1319 5151 1339
rect 5171 1319 5178 1339
rect 5128 1289 5178 1319
rect 9976 1469 10026 1485
rect 10194 1469 10244 1485
rect 10402 1469 10452 1485
rect 11335 1465 11385 1495
rect 11335 1445 11342 1465
rect 11362 1445 11385 1465
rect 11335 1418 11385 1445
rect 11543 1463 11593 1495
rect 11543 1443 11560 1463
rect 11580 1443 11593 1463
rect 11543 1418 11593 1443
rect 11761 1466 11811 1495
rect 11761 1446 11778 1466
rect 11798 1446 11811 1466
rect 13443 1491 13493 1504
rect 13661 1491 13711 1504
rect 13869 1491 13919 1504
rect 16496 1546 16546 1559
rect 16704 1546 16754 1559
rect 16922 1546 16972 1559
rect 18606 1563 18656 1591
rect 18606 1543 18619 1563
rect 18639 1543 18656 1563
rect 18606 1514 18656 1543
rect 18824 1566 18874 1591
rect 18824 1546 18837 1566
rect 18857 1546 18874 1566
rect 18824 1514 18874 1546
rect 19032 1564 19082 1591
rect 19032 1544 19055 1564
rect 19075 1544 19082 1564
rect 19032 1514 19082 1544
rect 19965 1524 20015 1540
rect 20173 1524 20223 1540
rect 20391 1524 20441 1540
rect 25126 1693 25176 1723
rect 25126 1673 25133 1693
rect 25153 1673 25176 1693
rect 25126 1646 25176 1673
rect 25334 1691 25384 1723
rect 25334 1671 25351 1691
rect 25371 1671 25384 1691
rect 25334 1646 25384 1671
rect 25552 1694 25602 1723
rect 25552 1674 25569 1694
rect 25589 1674 25602 1694
rect 27347 1716 27397 1729
rect 27565 1716 27615 1729
rect 27773 1716 27823 1729
rect 25552 1646 25602 1674
rect 22970 1576 23020 1604
rect 22970 1556 22983 1576
rect 23003 1556 23020 1576
rect 11761 1418 11811 1446
rect 7756 1341 7806 1357
rect 7964 1341 8014 1357
rect 8182 1341 8232 1357
rect 3818 1209 3868 1237
rect 5500 1282 5550 1295
rect 5718 1282 5768 1295
rect 5926 1282 5976 1295
rect 6958 1293 7008 1306
rect 7166 1293 7216 1306
rect 7384 1293 7434 1306
rect 9079 1350 9129 1378
rect 4702 1231 4752 1247
rect 4920 1231 4970 1247
rect 5128 1231 5178 1247
rect 1136 1141 1186 1169
rect 1136 1121 1149 1141
rect 1169 1121 1186 1141
rect 1136 1092 1186 1121
rect 1354 1144 1404 1169
rect 1354 1124 1367 1144
rect 1387 1124 1404 1144
rect 1354 1092 1404 1124
rect 1562 1142 1612 1169
rect 1562 1122 1585 1142
rect 1605 1122 1612 1142
rect 1562 1092 1612 1122
rect 7756 1269 7806 1299
rect 7756 1249 7763 1269
rect 7783 1249 7806 1269
rect 7756 1222 7806 1249
rect 7964 1267 8014 1299
rect 7964 1247 7981 1267
rect 8001 1247 8014 1267
rect 7964 1222 8014 1247
rect 8182 1270 8232 1299
rect 8182 1250 8199 1270
rect 8219 1250 8232 1270
rect 9079 1330 9092 1350
rect 9112 1330 9129 1350
rect 9079 1301 9129 1330
rect 9297 1353 9347 1378
rect 9297 1333 9310 1353
rect 9330 1333 9347 1353
rect 9297 1301 9347 1333
rect 9505 1351 9555 1378
rect 9505 1331 9528 1351
rect 9548 1331 9555 1351
rect 9505 1301 9555 1331
rect 14340 1482 14390 1498
rect 14558 1482 14608 1498
rect 14766 1482 14816 1498
rect 15699 1478 15749 1508
rect 15699 1458 15706 1478
rect 15726 1458 15749 1478
rect 15699 1431 15749 1458
rect 15907 1476 15957 1508
rect 15907 1456 15924 1476
rect 15944 1456 15957 1476
rect 15907 1431 15957 1456
rect 16125 1479 16175 1508
rect 16125 1459 16142 1479
rect 16162 1459 16175 1479
rect 16125 1431 16175 1459
rect 17709 1465 17759 1478
rect 17927 1465 17977 1478
rect 18135 1465 18185 1478
rect 20762 1520 20812 1533
rect 20970 1520 21020 1533
rect 21188 1520 21238 1533
rect 22970 1527 23020 1556
rect 23188 1579 23238 1604
rect 23188 1559 23201 1579
rect 23221 1559 23238 1579
rect 23188 1527 23238 1559
rect 23396 1577 23446 1604
rect 23396 1557 23419 1577
rect 23439 1557 23446 1577
rect 23396 1527 23446 1557
rect 24329 1537 24379 1553
rect 24537 1537 24587 1553
rect 24755 1537 24805 1553
rect 29503 1705 29553 1735
rect 29503 1685 29510 1705
rect 29530 1685 29553 1705
rect 29503 1658 29553 1685
rect 29711 1703 29761 1735
rect 29711 1683 29728 1703
rect 29748 1683 29761 1703
rect 29711 1658 29761 1683
rect 29929 1706 29979 1735
rect 29929 1686 29946 1706
rect 29966 1686 29979 1706
rect 31711 1729 31761 1742
rect 31929 1729 31979 1742
rect 32137 1729 32187 1742
rect 29929 1658 29979 1686
rect 27347 1588 27397 1616
rect 27347 1568 27360 1588
rect 27380 1568 27397 1588
rect 12133 1353 12183 1369
rect 12341 1353 12391 1369
rect 12559 1353 12609 1369
rect 8182 1222 8232 1250
rect 9877 1294 9927 1307
rect 10095 1294 10145 1307
rect 10303 1294 10353 1307
rect 11335 1305 11385 1318
rect 11543 1305 11593 1318
rect 11761 1305 11811 1318
rect 13443 1363 13493 1391
rect 9079 1243 9129 1259
rect 9297 1243 9347 1259
rect 9505 1243 9555 1259
rect 5500 1154 5550 1182
rect 3392 1096 3442 1109
rect 3600 1096 3650 1109
rect 3818 1096 3868 1109
rect 5500 1134 5513 1154
rect 5533 1134 5550 1154
rect 5500 1105 5550 1134
rect 5718 1157 5768 1182
rect 5718 1137 5731 1157
rect 5751 1137 5768 1157
rect 5718 1105 5768 1137
rect 5926 1155 5976 1182
rect 5926 1135 5949 1155
rect 5969 1135 5976 1155
rect 5926 1105 5976 1135
rect 12133 1281 12183 1311
rect 12133 1261 12140 1281
rect 12160 1261 12183 1281
rect 12133 1234 12183 1261
rect 12341 1279 12391 1311
rect 12341 1259 12358 1279
rect 12378 1259 12391 1279
rect 12341 1234 12391 1259
rect 12559 1282 12609 1311
rect 12559 1262 12576 1282
rect 12596 1262 12609 1282
rect 13443 1343 13456 1363
rect 13476 1343 13493 1363
rect 13443 1314 13493 1343
rect 13661 1366 13711 1391
rect 13661 1346 13674 1366
rect 13694 1346 13711 1366
rect 13661 1314 13711 1346
rect 13869 1364 13919 1391
rect 13869 1344 13892 1364
rect 13912 1344 13919 1364
rect 13869 1314 13919 1344
rect 16497 1366 16547 1382
rect 16705 1366 16755 1382
rect 16923 1366 16973 1382
rect 12559 1234 12609 1262
rect 14241 1307 14291 1320
rect 14459 1307 14509 1320
rect 14667 1307 14717 1320
rect 15699 1318 15749 1331
rect 15907 1318 15957 1331
rect 16125 1318 16175 1331
rect 18606 1456 18656 1472
rect 18824 1456 18874 1472
rect 19032 1456 19082 1472
rect 19965 1452 20015 1482
rect 19965 1432 19972 1452
rect 19992 1432 20015 1452
rect 19965 1405 20015 1432
rect 20173 1450 20223 1482
rect 20173 1430 20190 1450
rect 20210 1430 20223 1450
rect 20173 1405 20223 1430
rect 20391 1453 20441 1482
rect 20391 1433 20408 1453
rect 20428 1433 20441 1453
rect 22073 1478 22123 1491
rect 22291 1478 22341 1491
rect 22499 1478 22549 1491
rect 25126 1533 25176 1546
rect 25334 1533 25384 1546
rect 25552 1533 25602 1546
rect 27347 1539 27397 1568
rect 27565 1591 27615 1616
rect 27565 1571 27578 1591
rect 27598 1571 27615 1591
rect 27565 1539 27615 1571
rect 27773 1589 27823 1616
rect 27773 1569 27796 1589
rect 27816 1569 27823 1589
rect 27773 1539 27823 1569
rect 28706 1549 28756 1565
rect 28914 1549 28964 1565
rect 29132 1549 29182 1565
rect 33867 1718 33917 1748
rect 33867 1698 33874 1718
rect 33894 1698 33917 1718
rect 33867 1671 33917 1698
rect 34075 1716 34125 1748
rect 34075 1696 34092 1716
rect 34112 1696 34125 1716
rect 34075 1671 34125 1696
rect 34293 1719 34343 1748
rect 34293 1699 34310 1719
rect 34330 1699 34343 1719
rect 34293 1671 34343 1699
rect 31711 1601 31761 1629
rect 31711 1581 31724 1601
rect 31744 1581 31761 1601
rect 20391 1405 20441 1433
rect 13443 1256 13493 1272
rect 13661 1256 13711 1272
rect 13869 1256 13919 1272
rect 9877 1166 9927 1194
rect 7756 1109 7806 1122
rect 7964 1109 8014 1122
rect 8182 1109 8232 1122
rect 9877 1146 9890 1166
rect 9910 1146 9927 1166
rect 9877 1117 9927 1146
rect 10095 1169 10145 1194
rect 10095 1149 10108 1169
rect 10128 1149 10145 1169
rect 10095 1117 10145 1149
rect 10303 1167 10353 1194
rect 10303 1147 10326 1167
rect 10346 1147 10353 1167
rect 10303 1117 10353 1147
rect 16497 1294 16547 1324
rect 16497 1274 16504 1294
rect 16524 1274 16547 1294
rect 16497 1247 16547 1274
rect 16705 1292 16755 1324
rect 16705 1272 16722 1292
rect 16742 1272 16755 1292
rect 16705 1247 16755 1272
rect 16923 1295 16973 1324
rect 16923 1275 16940 1295
rect 16960 1275 16973 1295
rect 17709 1337 17759 1365
rect 16923 1247 16973 1275
rect 17709 1317 17722 1337
rect 17742 1317 17759 1337
rect 17709 1288 17759 1317
rect 17927 1340 17977 1365
rect 17927 1320 17940 1340
rect 17960 1320 17977 1340
rect 17927 1288 17977 1320
rect 18135 1338 18185 1365
rect 18135 1318 18158 1338
rect 18178 1318 18185 1338
rect 18135 1288 18185 1318
rect 22970 1469 23020 1485
rect 23188 1469 23238 1485
rect 23396 1469 23446 1485
rect 24329 1465 24379 1495
rect 24329 1445 24336 1465
rect 24356 1445 24379 1465
rect 24329 1418 24379 1445
rect 24537 1463 24587 1495
rect 24537 1443 24554 1463
rect 24574 1443 24587 1463
rect 24537 1418 24587 1443
rect 24755 1466 24805 1495
rect 24755 1446 24772 1466
rect 24792 1446 24805 1466
rect 26450 1490 26500 1503
rect 26668 1490 26718 1503
rect 26876 1490 26926 1503
rect 29503 1545 29553 1558
rect 29711 1545 29761 1558
rect 29929 1545 29979 1558
rect 31711 1552 31761 1581
rect 31929 1604 31979 1629
rect 31929 1584 31942 1604
rect 31962 1584 31979 1604
rect 31929 1552 31979 1584
rect 32137 1602 32187 1629
rect 32137 1582 32160 1602
rect 32180 1582 32187 1602
rect 32137 1552 32187 1582
rect 33070 1562 33120 1578
rect 33278 1562 33328 1578
rect 33496 1562 33546 1578
rect 24755 1418 24805 1446
rect 20763 1340 20813 1356
rect 20971 1340 21021 1356
rect 21189 1340 21239 1356
rect 14241 1179 14291 1207
rect 12133 1121 12183 1134
rect 12341 1121 12391 1134
rect 12559 1121 12609 1134
rect 14241 1159 14254 1179
rect 14274 1159 14291 1179
rect 14241 1130 14291 1159
rect 14459 1182 14509 1207
rect 14459 1162 14472 1182
rect 14492 1162 14509 1182
rect 14459 1130 14509 1162
rect 14667 1180 14717 1207
rect 14667 1160 14690 1180
rect 14710 1160 14717 1180
rect 14667 1130 14717 1160
rect 18507 1281 18557 1294
rect 18725 1281 18775 1294
rect 18933 1281 18983 1294
rect 19965 1292 20015 1305
rect 20173 1292 20223 1305
rect 20391 1292 20441 1305
rect 22073 1350 22123 1378
rect 17709 1230 17759 1246
rect 17927 1230 17977 1246
rect 18135 1230 18185 1246
rect 20763 1268 20813 1298
rect 20763 1248 20770 1268
rect 20790 1248 20813 1268
rect 20763 1221 20813 1248
rect 20971 1266 21021 1298
rect 20971 1246 20988 1266
rect 21008 1246 21021 1266
rect 20971 1221 21021 1246
rect 21189 1269 21239 1298
rect 21189 1249 21206 1269
rect 21226 1249 21239 1269
rect 22073 1330 22086 1350
rect 22106 1330 22123 1350
rect 22073 1301 22123 1330
rect 22291 1353 22341 1378
rect 22291 1333 22304 1353
rect 22324 1333 22341 1353
rect 22291 1301 22341 1333
rect 22499 1351 22549 1378
rect 22499 1331 22522 1351
rect 22542 1331 22549 1351
rect 22499 1301 22549 1331
rect 27347 1481 27397 1497
rect 27565 1481 27615 1497
rect 27773 1481 27823 1497
rect 28706 1477 28756 1507
rect 28706 1457 28713 1477
rect 28733 1457 28756 1477
rect 28706 1430 28756 1457
rect 28914 1475 28964 1507
rect 28914 1455 28931 1475
rect 28951 1455 28964 1475
rect 28914 1430 28964 1455
rect 29132 1478 29182 1507
rect 29132 1458 29149 1478
rect 29169 1458 29182 1478
rect 30814 1503 30864 1516
rect 31032 1503 31082 1516
rect 31240 1503 31290 1516
rect 33867 1558 33917 1571
rect 34075 1558 34125 1571
rect 34293 1558 34343 1571
rect 29132 1430 29182 1458
rect 25127 1353 25177 1369
rect 25335 1353 25385 1369
rect 25553 1353 25603 1369
rect 21189 1221 21239 1249
rect 22871 1294 22921 1307
rect 23089 1294 23139 1307
rect 23297 1294 23347 1307
rect 24329 1305 24379 1318
rect 24537 1305 24587 1318
rect 24755 1305 24805 1318
rect 26450 1362 26500 1390
rect 22073 1243 22123 1259
rect 22291 1243 22341 1259
rect 22499 1243 22549 1259
rect 16497 1134 16547 1147
rect 16705 1134 16755 1147
rect 16923 1134 16973 1147
rect 18507 1153 18557 1181
rect 339 1041 389 1054
rect 557 1041 607 1054
rect 765 1041 815 1054
rect 1136 1034 1186 1050
rect 1354 1034 1404 1050
rect 1562 1034 1612 1050
rect 4703 1054 4753 1067
rect 4921 1054 4971 1067
rect 5129 1054 5179 1067
rect 339 913 389 941
rect 339 893 352 913
rect 372 893 389 913
rect 339 864 389 893
rect 557 916 607 941
rect 557 896 570 916
rect 590 896 607 916
rect 557 864 607 896
rect 765 914 815 941
rect 5500 1047 5550 1063
rect 5718 1047 5768 1063
rect 5926 1047 5976 1063
rect 9080 1066 9130 1079
rect 9298 1066 9348 1079
rect 9506 1066 9556 1079
rect 765 894 788 914
rect 808 894 815 914
rect 765 864 815 894
rect 4703 926 4753 954
rect 4703 906 4716 926
rect 4736 906 4753 926
rect 4703 877 4753 906
rect 4921 929 4971 954
rect 4921 909 4934 929
rect 4954 909 4971 929
rect 4921 877 4971 909
rect 5129 927 5179 954
rect 9877 1059 9927 1075
rect 10095 1059 10145 1075
rect 10303 1059 10353 1075
rect 13444 1079 13494 1092
rect 13662 1079 13712 1092
rect 13870 1079 13920 1092
rect 18507 1133 18520 1153
rect 18540 1133 18557 1153
rect 18507 1104 18557 1133
rect 18725 1156 18775 1181
rect 18725 1136 18738 1156
rect 18758 1136 18775 1156
rect 18725 1104 18775 1136
rect 18933 1154 18983 1181
rect 18933 1134 18956 1154
rect 18976 1134 18983 1154
rect 18933 1104 18983 1134
rect 25127 1281 25177 1311
rect 25127 1261 25134 1281
rect 25154 1261 25177 1281
rect 25127 1234 25177 1261
rect 25335 1279 25385 1311
rect 25335 1259 25352 1279
rect 25372 1259 25385 1279
rect 25335 1234 25385 1259
rect 25553 1282 25603 1311
rect 25553 1262 25570 1282
rect 25590 1262 25603 1282
rect 26450 1342 26463 1362
rect 26483 1342 26500 1362
rect 26450 1313 26500 1342
rect 26668 1365 26718 1390
rect 26668 1345 26681 1365
rect 26701 1345 26718 1365
rect 26668 1313 26718 1345
rect 26876 1363 26926 1390
rect 26876 1343 26899 1363
rect 26919 1343 26926 1363
rect 26876 1313 26926 1343
rect 31711 1494 31761 1510
rect 31929 1494 31979 1510
rect 32137 1494 32187 1510
rect 33070 1490 33120 1520
rect 33070 1470 33077 1490
rect 33097 1470 33120 1490
rect 33070 1443 33120 1470
rect 33278 1488 33328 1520
rect 33278 1468 33295 1488
rect 33315 1468 33328 1488
rect 33278 1443 33328 1468
rect 33496 1491 33546 1520
rect 33496 1471 33513 1491
rect 33533 1471 33546 1491
rect 33496 1443 33546 1471
rect 29504 1365 29554 1381
rect 29712 1365 29762 1381
rect 29930 1365 29980 1381
rect 25553 1234 25603 1262
rect 27248 1306 27298 1319
rect 27466 1306 27516 1319
rect 27674 1306 27724 1319
rect 28706 1317 28756 1330
rect 28914 1317 28964 1330
rect 29132 1317 29182 1330
rect 30814 1375 30864 1403
rect 26450 1255 26500 1271
rect 26668 1255 26718 1271
rect 26876 1255 26926 1271
rect 22871 1166 22921 1194
rect 20763 1108 20813 1121
rect 20971 1108 21021 1121
rect 21189 1108 21239 1121
rect 22871 1146 22884 1166
rect 22904 1146 22921 1166
rect 22871 1117 22921 1146
rect 23089 1169 23139 1194
rect 23089 1149 23102 1169
rect 23122 1149 23139 1169
rect 23089 1117 23139 1149
rect 23297 1167 23347 1194
rect 23297 1147 23320 1167
rect 23340 1147 23347 1167
rect 23297 1117 23347 1147
rect 29504 1293 29554 1323
rect 29504 1273 29511 1293
rect 29531 1273 29554 1293
rect 29504 1246 29554 1273
rect 29712 1291 29762 1323
rect 29712 1271 29729 1291
rect 29749 1271 29762 1291
rect 29712 1246 29762 1271
rect 29930 1294 29980 1323
rect 29930 1274 29947 1294
rect 29967 1274 29980 1294
rect 30814 1355 30827 1375
rect 30847 1355 30864 1375
rect 30814 1326 30864 1355
rect 31032 1378 31082 1403
rect 31032 1358 31045 1378
rect 31065 1358 31082 1378
rect 31032 1326 31082 1358
rect 31240 1376 31290 1403
rect 31240 1356 31263 1376
rect 31283 1356 31290 1376
rect 31240 1326 31290 1356
rect 33868 1378 33918 1394
rect 34076 1378 34126 1394
rect 34294 1378 34344 1394
rect 29930 1246 29980 1274
rect 31612 1319 31662 1332
rect 31830 1319 31880 1332
rect 32038 1319 32088 1332
rect 33070 1330 33120 1343
rect 33278 1330 33328 1343
rect 33496 1330 33546 1343
rect 30814 1268 30864 1284
rect 31032 1268 31082 1284
rect 31240 1268 31290 1284
rect 27248 1178 27298 1206
rect 25127 1121 25177 1134
rect 25335 1121 25385 1134
rect 25553 1121 25603 1134
rect 27248 1158 27261 1178
rect 27281 1158 27298 1178
rect 27248 1129 27298 1158
rect 27466 1181 27516 1206
rect 27466 1161 27479 1181
rect 27499 1161 27516 1181
rect 27466 1129 27516 1161
rect 27674 1179 27724 1206
rect 27674 1159 27697 1179
rect 27717 1159 27724 1179
rect 27674 1129 27724 1159
rect 33868 1306 33918 1336
rect 33868 1286 33875 1306
rect 33895 1286 33918 1306
rect 33868 1259 33918 1286
rect 34076 1304 34126 1336
rect 34076 1284 34093 1304
rect 34113 1284 34126 1304
rect 34076 1259 34126 1284
rect 34294 1307 34344 1336
rect 34294 1287 34311 1307
rect 34331 1287 34344 1307
rect 34294 1259 34344 1287
rect 31612 1191 31662 1219
rect 29504 1133 29554 1146
rect 29712 1133 29762 1146
rect 29930 1133 29980 1146
rect 31612 1171 31625 1191
rect 31645 1171 31662 1191
rect 31612 1142 31662 1171
rect 31830 1194 31880 1219
rect 31830 1174 31843 1194
rect 31863 1174 31880 1194
rect 31830 1142 31880 1174
rect 32038 1192 32088 1219
rect 32038 1172 32061 1192
rect 32081 1172 32088 1192
rect 32038 1142 32088 1172
rect 33868 1146 33918 1159
rect 34076 1146 34126 1159
rect 34294 1146 34344 1159
rect 5129 907 5152 927
rect 5172 907 5179 927
rect 5129 877 5179 907
rect 9080 938 9130 966
rect 9080 918 9093 938
rect 9113 918 9130 938
rect 9080 889 9130 918
rect 9298 941 9348 966
rect 9298 921 9311 941
rect 9331 921 9348 941
rect 9298 889 9348 921
rect 9506 939 9556 966
rect 14241 1072 14291 1088
rect 14459 1072 14509 1088
rect 14667 1072 14717 1088
rect 17710 1053 17760 1066
rect 17928 1053 17978 1066
rect 18136 1053 18186 1066
rect 9506 919 9529 939
rect 9549 919 9556 939
rect 9506 889 9556 919
rect 13444 951 13494 979
rect 13444 931 13457 951
rect 13477 931 13494 951
rect 13444 902 13494 931
rect 13662 954 13712 979
rect 13662 934 13675 954
rect 13695 934 13712 954
rect 13662 902 13712 934
rect 13870 952 13920 979
rect 13870 932 13893 952
rect 13913 932 13920 952
rect 13870 902 13920 932
rect 18507 1046 18557 1062
rect 18725 1046 18775 1062
rect 18933 1046 18983 1062
rect 22074 1066 22124 1079
rect 22292 1066 22342 1079
rect 22500 1066 22550 1079
rect 17710 925 17760 953
rect 17710 905 17723 925
rect 17743 905 17760 925
rect 339 806 389 822
rect 557 806 607 822
rect 765 806 815 822
rect 4703 819 4753 835
rect 4921 819 4971 835
rect 5129 819 5179 835
rect 9080 831 9130 847
rect 9298 831 9348 847
rect 9506 831 9556 847
rect 13444 844 13494 860
rect 13662 844 13712 860
rect 13870 844 13920 860
rect 17710 876 17760 905
rect 17928 928 17978 953
rect 17928 908 17941 928
rect 17961 908 17978 928
rect 17928 876 17978 908
rect 18136 926 18186 953
rect 22871 1059 22921 1075
rect 23089 1059 23139 1075
rect 23297 1059 23347 1075
rect 26451 1078 26501 1091
rect 26669 1078 26719 1091
rect 26877 1078 26927 1091
rect 18136 906 18159 926
rect 18179 906 18186 926
rect 18136 876 18186 906
rect 22074 938 22124 966
rect 22074 918 22087 938
rect 22107 918 22124 938
rect 22074 889 22124 918
rect 22292 941 22342 966
rect 22292 921 22305 941
rect 22325 921 22342 941
rect 22292 889 22342 921
rect 22500 939 22550 966
rect 27248 1071 27298 1087
rect 27466 1071 27516 1087
rect 27674 1071 27724 1087
rect 30815 1091 30865 1104
rect 31033 1091 31083 1104
rect 31241 1091 31291 1104
rect 22500 919 22523 939
rect 22543 919 22550 939
rect 22500 889 22550 919
rect 26451 950 26501 978
rect 26451 930 26464 950
rect 26484 930 26501 950
rect 26451 901 26501 930
rect 26669 953 26719 978
rect 26669 933 26682 953
rect 26702 933 26719 953
rect 26669 901 26719 933
rect 26877 951 26927 978
rect 31612 1084 31662 1100
rect 31830 1084 31880 1100
rect 32038 1084 32088 1100
rect 26877 931 26900 951
rect 26920 931 26927 951
rect 26877 901 26927 931
rect 30815 963 30865 991
rect 30815 943 30828 963
rect 30848 943 30865 963
rect 30815 914 30865 943
rect 31033 966 31083 991
rect 31033 946 31046 966
rect 31066 946 31083 966
rect 31033 914 31083 946
rect 31241 964 31291 991
rect 31241 944 31264 964
rect 31284 944 31291 964
rect 31241 914 31291 944
rect 17710 818 17760 834
rect 17928 818 17978 834
rect 18136 818 18186 834
rect 22074 831 22124 847
rect 22292 831 22342 847
rect 22500 831 22550 847
rect 26451 843 26501 859
rect 26669 843 26719 859
rect 26877 843 26927 859
rect 30815 856 30865 872
rect 31033 856 31083 872
rect 31241 856 31291 872
rect 14657 503 14707 516
rect 14875 503 14925 516
rect 15083 503 15133 516
rect 32028 515 32078 528
rect 32246 515 32296 528
rect 32454 515 32504 528
rect 5916 478 5966 491
rect 6134 478 6184 491
rect 6342 478 6392 491
rect 10293 490 10343 503
rect 10511 490 10561 503
rect 10719 490 10769 503
rect 1552 465 1602 478
rect 1770 465 1820 478
rect 1978 465 2028 478
rect 4041 391 4091 404
rect 4259 391 4309 404
rect 4467 391 4517 404
rect 1552 337 1602 365
rect 1552 317 1565 337
rect 1585 317 1602 337
rect 1552 288 1602 317
rect 1770 340 1820 365
rect 1770 320 1783 340
rect 1803 320 1820 340
rect 1770 288 1820 320
rect 1978 338 2028 365
rect 1978 318 2001 338
rect 2021 318 2028 338
rect 1978 288 2028 318
rect 8489 415 8539 428
rect 8707 415 8757 428
rect 8915 415 8965 428
rect 5916 350 5966 378
rect 5916 330 5929 350
rect 5949 330 5966 350
rect 5916 301 5966 330
rect 6134 353 6184 378
rect 6134 333 6147 353
rect 6167 333 6184 353
rect 6134 301 6184 333
rect 6342 351 6392 378
rect 6342 331 6365 351
rect 6385 331 6392 351
rect 6342 301 6392 331
rect 12782 416 12832 429
rect 13000 416 13050 429
rect 13208 416 13258 429
rect 10293 362 10343 390
rect 10293 342 10306 362
rect 10326 342 10343 362
rect 4041 263 4091 291
rect 1552 230 1602 246
rect 1770 230 1820 246
rect 1978 230 2028 246
rect 4041 243 4054 263
rect 4074 243 4091 263
rect 4041 214 4091 243
rect 4259 266 4309 291
rect 4259 246 4272 266
rect 4292 246 4309 266
rect 4259 214 4309 246
rect 4467 264 4517 291
rect 4467 244 4490 264
rect 4510 244 4517 264
rect 8489 287 8539 315
rect 8489 267 8502 287
rect 8522 267 8539 287
rect 4467 214 4517 244
rect 5916 243 5966 259
rect 6134 243 6184 259
rect 6342 243 6392 259
rect 8489 238 8539 267
rect 8707 290 8757 315
rect 8707 270 8720 290
rect 8740 270 8757 290
rect 8707 238 8757 270
rect 8915 288 8965 315
rect 10293 313 10343 342
rect 10511 365 10561 390
rect 10511 345 10524 365
rect 10544 345 10561 365
rect 10511 313 10561 345
rect 10719 363 10769 390
rect 10719 343 10742 363
rect 10762 343 10769 363
rect 10719 313 10769 343
rect 23287 490 23337 503
rect 23505 490 23555 503
rect 23713 490 23763 503
rect 27664 502 27714 515
rect 27882 502 27932 515
rect 28090 502 28140 515
rect 18923 477 18973 490
rect 19141 477 19191 490
rect 19349 477 19399 490
rect 14657 375 14707 403
rect 14657 355 14670 375
rect 14690 355 14707 375
rect 14657 326 14707 355
rect 14875 378 14925 403
rect 14875 358 14888 378
rect 14908 358 14925 378
rect 14875 326 14925 358
rect 15083 376 15133 403
rect 21412 403 21462 416
rect 21630 403 21680 416
rect 21838 403 21888 416
rect 15083 356 15106 376
rect 15126 356 15133 376
rect 15083 326 15133 356
rect 16979 352 17029 365
rect 17197 352 17247 365
rect 17405 352 17455 365
rect 8915 268 8938 288
rect 8958 268 8965 288
rect 12782 288 12832 316
rect 8915 238 8965 268
rect 10293 255 10343 271
rect 10511 255 10561 271
rect 10719 255 10769 271
rect 12782 268 12795 288
rect 12815 268 12832 288
rect 12782 239 12832 268
rect 13000 291 13050 316
rect 13000 271 13013 291
rect 13033 271 13050 291
rect 13000 239 13050 271
rect 13208 289 13258 316
rect 13208 269 13231 289
rect 13251 269 13258 289
rect 13208 239 13258 269
rect 14657 268 14707 284
rect 14875 268 14925 284
rect 15083 268 15133 284
rect 18923 349 18973 377
rect 18923 329 18936 349
rect 18956 329 18973 349
rect 18923 300 18973 329
rect 19141 352 19191 377
rect 19141 332 19154 352
rect 19174 332 19191 352
rect 19141 300 19191 332
rect 19349 350 19399 377
rect 19349 330 19372 350
rect 19392 330 19399 350
rect 19349 300 19399 330
rect 25860 427 25910 440
rect 26078 427 26128 440
rect 26286 427 26336 440
rect 23287 362 23337 390
rect 23287 342 23300 362
rect 23320 342 23337 362
rect 23287 313 23337 342
rect 23505 365 23555 390
rect 23505 345 23518 365
rect 23538 345 23555 365
rect 23505 313 23555 345
rect 23713 363 23763 390
rect 23713 343 23736 363
rect 23756 343 23763 363
rect 23713 313 23763 343
rect 30153 428 30203 441
rect 30371 428 30421 441
rect 30579 428 30629 441
rect 27664 374 27714 402
rect 27664 354 27677 374
rect 27697 354 27714 374
rect 21412 275 21462 303
rect 16979 224 17029 252
rect 16979 204 16992 224
rect 17012 204 17029 224
rect 8489 180 8539 196
rect 8707 180 8757 196
rect 8915 180 8965 196
rect 12782 181 12832 197
rect 13000 181 13050 197
rect 13208 181 13258 197
rect 16979 175 17029 204
rect 17197 227 17247 252
rect 17197 207 17210 227
rect 17230 207 17247 227
rect 17197 175 17247 207
rect 17405 225 17455 252
rect 18923 242 18973 258
rect 19141 242 19191 258
rect 19349 242 19399 258
rect 21412 255 21425 275
rect 21445 255 21462 275
rect 21412 226 21462 255
rect 21630 278 21680 303
rect 21630 258 21643 278
rect 21663 258 21680 278
rect 21630 226 21680 258
rect 21838 276 21888 303
rect 21838 256 21861 276
rect 21881 256 21888 276
rect 25860 299 25910 327
rect 25860 279 25873 299
rect 25893 279 25910 299
rect 21838 226 21888 256
rect 23287 255 23337 271
rect 23505 255 23555 271
rect 23713 255 23763 271
rect 25860 250 25910 279
rect 26078 302 26128 327
rect 26078 282 26091 302
rect 26111 282 26128 302
rect 26078 250 26128 282
rect 26286 300 26336 327
rect 27664 325 27714 354
rect 27882 377 27932 402
rect 27882 357 27895 377
rect 27915 357 27932 377
rect 27882 325 27932 357
rect 28090 375 28140 402
rect 28090 355 28113 375
rect 28133 355 28140 375
rect 28090 325 28140 355
rect 32028 387 32078 415
rect 32028 367 32041 387
rect 32061 367 32078 387
rect 32028 338 32078 367
rect 32246 390 32296 415
rect 32246 370 32259 390
rect 32279 370 32296 390
rect 32246 338 32296 370
rect 32454 388 32504 415
rect 32454 368 32477 388
rect 32497 368 32504 388
rect 32454 338 32504 368
rect 26286 280 26309 300
rect 26329 280 26336 300
rect 30153 300 30203 328
rect 26286 250 26336 280
rect 27664 267 27714 283
rect 27882 267 27932 283
rect 28090 267 28140 283
rect 30153 280 30166 300
rect 30186 280 30203 300
rect 30153 251 30203 280
rect 30371 303 30421 328
rect 30371 283 30384 303
rect 30404 283 30421 303
rect 30371 251 30421 283
rect 30579 301 30629 328
rect 30579 281 30602 301
rect 30622 281 30629 301
rect 30579 251 30629 281
rect 32028 280 32078 296
rect 32246 280 32296 296
rect 32454 280 32504 296
rect 17405 205 17428 225
rect 17448 205 17455 225
rect 17405 175 17455 205
rect 25860 192 25910 208
rect 26078 192 26128 208
rect 26286 192 26336 208
rect 30153 193 30203 209
rect 30371 193 30421 209
rect 30579 193 30629 209
rect 4041 156 4091 172
rect 4259 156 4309 172
rect 4467 156 4517 172
rect 21412 168 21462 184
rect 21630 168 21680 184
rect 21838 168 21888 184
rect 16979 117 17029 133
rect 17197 117 17247 133
rect 17405 117 17455 133
<< polycont >>
rect 3525 8774 3545 8794
rect 3743 8772 3763 8792
rect 3961 8775 3981 8795
rect 7889 8787 7909 8807
rect 8107 8785 8127 8805
rect 8325 8788 8345 8808
rect 12266 8799 12286 8819
rect 12484 8797 12504 8817
rect 12702 8800 12722 8820
rect 16630 8812 16650 8832
rect 16848 8810 16868 8830
rect 17066 8813 17086 8833
rect 20896 8786 20916 8806
rect 21114 8784 21134 8804
rect 21332 8787 21352 8807
rect 25260 8799 25280 8819
rect 25478 8797 25498 8817
rect 25696 8800 25716 8820
rect 29637 8811 29657 8831
rect 2728 8546 2748 8566
rect 2946 8544 2966 8564
rect 3164 8547 3184 8567
rect 478 8431 498 8451
rect 696 8434 716 8454
rect 914 8432 934 8452
rect 7092 8559 7112 8579
rect 7310 8557 7330 8577
rect 7528 8560 7548 8580
rect 3526 8362 3546 8382
rect 3744 8360 3764 8380
rect 3962 8363 3982 8383
rect 4842 8444 4862 8464
rect 5060 8447 5080 8467
rect 5278 8445 5298 8465
rect 11469 8571 11489 8591
rect 11687 8569 11707 8589
rect 11905 8572 11925 8592
rect 1276 8247 1296 8267
rect 1494 8250 1514 8270
rect 1712 8248 1732 8268
rect 7890 8375 7910 8395
rect 8108 8373 8128 8393
rect 8326 8376 8346 8396
rect 9219 8456 9239 8476
rect 9437 8459 9457 8479
rect 9655 8457 9675 8477
rect 15833 8584 15853 8604
rect 16051 8582 16071 8602
rect 16269 8585 16289 8605
rect 29855 8809 29875 8829
rect 30073 8812 30093 8832
rect 34001 8824 34021 8844
rect 34219 8822 34239 8842
rect 34437 8825 34457 8845
rect 5640 8260 5660 8280
rect 5858 8263 5878 8283
rect 6076 8261 6096 8281
rect 12267 8387 12287 8407
rect 12485 8385 12505 8405
rect 12703 8388 12723 8408
rect 13583 8469 13603 8489
rect 13801 8472 13821 8492
rect 14019 8470 14039 8490
rect 20099 8558 20119 8578
rect 20317 8556 20337 8576
rect 20535 8559 20555 8579
rect 2629 8136 2649 8156
rect 2847 8134 2867 8154
rect 10017 8272 10037 8292
rect 10235 8275 10255 8295
rect 10453 8273 10473 8293
rect 16631 8400 16651 8420
rect 16849 8398 16869 8418
rect 17067 8401 17087 8421
rect 17849 8443 17869 8463
rect 18067 8446 18087 8466
rect 18285 8444 18305 8464
rect 24463 8571 24483 8591
rect 24681 8569 24701 8589
rect 24899 8572 24919 8592
rect 3065 8137 3085 8157
rect 479 8019 499 8039
rect 697 8022 717 8042
rect 915 8020 935 8040
rect 6993 8149 7013 8169
rect 7211 8147 7231 8167
rect 14381 8285 14401 8305
rect 14599 8288 14619 8308
rect 14817 8286 14837 8306
rect 20897 8374 20917 8394
rect 21115 8372 21135 8392
rect 21333 8375 21353 8395
rect 22213 8456 22233 8476
rect 22431 8459 22451 8479
rect 22649 8457 22669 8477
rect 28840 8583 28860 8603
rect 29058 8581 29078 8601
rect 29276 8584 29296 8604
rect 7429 8150 7449 8170
rect 4843 8032 4863 8052
rect 5061 8035 5081 8055
rect 5279 8033 5299 8053
rect 11370 8161 11390 8181
rect 11588 8159 11608 8179
rect 18647 8259 18667 8279
rect 18865 8262 18885 8282
rect 19083 8260 19103 8280
rect 25261 8387 25281 8407
rect 25479 8385 25499 8405
rect 25697 8388 25717 8408
rect 26590 8468 26610 8488
rect 26808 8471 26828 8491
rect 27026 8469 27046 8489
rect 33204 8596 33224 8616
rect 33422 8594 33442 8614
rect 33640 8597 33660 8617
rect 11806 8162 11826 8182
rect 9220 8044 9240 8064
rect 9438 8047 9458 8067
rect 9656 8045 9676 8065
rect 15734 8174 15754 8194
rect 15952 8172 15972 8192
rect 16170 8175 16190 8195
rect 23011 8272 23031 8292
rect 23229 8275 23249 8295
rect 23447 8273 23467 8293
rect 29638 8399 29658 8419
rect 29856 8397 29876 8417
rect 30074 8400 30094 8420
rect 30954 8481 30974 8501
rect 31172 8484 31192 8504
rect 31390 8482 31410 8502
rect 13584 8057 13604 8077
rect 13802 8060 13822 8080
rect 14020 8058 14040 8078
rect 20000 8148 20020 8168
rect 20218 8146 20238 8166
rect 27388 8284 27408 8304
rect 27606 8287 27626 8307
rect 27824 8285 27844 8305
rect 34002 8412 34022 8432
rect 34220 8410 34240 8430
rect 34438 8413 34458 8433
rect 20436 8149 20456 8169
rect 17850 8031 17870 8051
rect 18068 8034 18088 8054
rect 18286 8032 18306 8052
rect 24364 8161 24384 8181
rect 24582 8159 24602 8179
rect 31752 8297 31772 8317
rect 31970 8300 31990 8320
rect 32188 8298 32208 8318
rect 24800 8162 24820 8182
rect 22214 8044 22234 8064
rect 22432 8047 22452 8067
rect 22650 8045 22670 8065
rect 28741 8173 28761 8193
rect 28959 8171 28979 8191
rect 29177 8174 29197 8194
rect 26591 8056 26611 8076
rect 26809 8059 26829 8079
rect 27027 8057 27047 8077
rect 33105 8186 33125 8206
rect 33323 8184 33343 8204
rect 33541 8187 33561 8207
rect 30955 8069 30975 8089
rect 31173 8072 31193 8092
rect 31391 8070 31411 8090
rect 3508 7756 3528 7776
rect 3726 7754 3746 7774
rect 3944 7757 3964 7777
rect 1358 7639 1378 7659
rect 1576 7642 1596 7662
rect 1794 7640 1814 7660
rect 7872 7769 7892 7789
rect 8090 7767 8110 7787
rect 8308 7770 8328 7790
rect 5722 7652 5742 7672
rect 5940 7655 5960 7675
rect 6158 7653 6178 7673
rect 12249 7781 12269 7801
rect 12467 7779 12487 7799
rect 12685 7782 12705 7802
rect 10099 7664 10119 7684
rect 2711 7528 2731 7548
rect 2929 7526 2949 7546
rect 3147 7529 3167 7549
rect 10317 7667 10337 7687
rect 10535 7665 10555 7685
rect 16613 7794 16633 7814
rect 16831 7792 16851 7812
rect 17049 7795 17069 7815
rect 14463 7677 14483 7697
rect 461 7413 481 7433
rect 679 7416 699 7436
rect 897 7414 917 7434
rect 7075 7541 7095 7561
rect 7293 7539 7313 7559
rect 7511 7542 7531 7562
rect 14681 7680 14701 7700
rect 14899 7678 14919 7698
rect 20879 7768 20899 7788
rect 21097 7766 21117 7786
rect 21315 7769 21335 7789
rect 3509 7344 3529 7364
rect 3727 7342 3747 7362
rect 3945 7345 3965 7365
rect 4825 7426 4845 7446
rect 5043 7429 5063 7449
rect 5261 7427 5281 7447
rect 11452 7553 11472 7573
rect 11670 7551 11690 7571
rect 11888 7554 11908 7574
rect 18729 7651 18749 7671
rect 18947 7654 18967 7674
rect 19165 7652 19185 7672
rect 25243 7781 25263 7801
rect 25461 7779 25481 7799
rect 25679 7782 25699 7802
rect 23093 7664 23113 7684
rect 1259 7229 1279 7249
rect 1477 7232 1497 7252
rect 1695 7230 1715 7250
rect 7873 7357 7893 7377
rect 8091 7355 8111 7375
rect 8309 7358 8329 7378
rect 9202 7438 9222 7458
rect 9420 7441 9440 7461
rect 9638 7439 9658 7459
rect 15816 7566 15836 7586
rect 16034 7564 16054 7584
rect 16252 7567 16272 7587
rect 23311 7667 23331 7687
rect 23529 7665 23549 7685
rect 29620 7793 29640 7813
rect 29838 7791 29858 7811
rect 30056 7794 30076 7814
rect 27470 7676 27490 7696
rect 5623 7242 5643 7262
rect 5841 7245 5861 7265
rect 6059 7243 6079 7263
rect 12250 7369 12270 7389
rect 12468 7367 12488 7387
rect 12686 7370 12706 7390
rect 13566 7451 13586 7471
rect 13784 7454 13804 7474
rect 14002 7452 14022 7472
rect 20082 7540 20102 7560
rect 20300 7538 20320 7558
rect 20518 7541 20538 7561
rect 27688 7679 27708 7699
rect 27906 7677 27926 7697
rect 33984 7806 34004 7826
rect 34202 7804 34222 7824
rect 34420 7807 34440 7827
rect 31834 7689 31854 7709
rect 2546 7120 2566 7140
rect 2764 7118 2784 7138
rect 10000 7254 10020 7274
rect 10218 7257 10238 7277
rect 10436 7255 10456 7275
rect 16614 7382 16634 7402
rect 16832 7380 16852 7400
rect 17050 7383 17070 7403
rect 17832 7425 17852 7445
rect 18050 7428 18070 7448
rect 18268 7426 18288 7446
rect 24446 7553 24466 7573
rect 24664 7551 24684 7571
rect 24882 7554 24902 7574
rect 32052 7692 32072 7712
rect 32270 7690 32290 7710
rect 2982 7121 3002 7141
rect 462 7001 482 7021
rect 680 7004 700 7024
rect 898 7002 918 7022
rect 6910 7133 6930 7153
rect 7128 7131 7148 7151
rect 14364 7267 14384 7287
rect 14582 7270 14602 7290
rect 14800 7268 14820 7288
rect 20880 7356 20900 7376
rect 21098 7354 21118 7374
rect 21316 7357 21336 7377
rect 22196 7438 22216 7458
rect 22414 7441 22434 7461
rect 22632 7439 22652 7459
rect 28823 7565 28843 7585
rect 29041 7563 29061 7583
rect 29259 7566 29279 7586
rect 7346 7134 7366 7154
rect 4826 7014 4846 7034
rect 5044 7017 5064 7037
rect 5262 7015 5282 7035
rect 11287 7145 11307 7165
rect 11505 7143 11525 7163
rect 18630 7241 18650 7261
rect 18848 7244 18868 7264
rect 19066 7242 19086 7262
rect 25244 7369 25264 7389
rect 25462 7367 25482 7387
rect 25680 7370 25700 7390
rect 26573 7450 26593 7470
rect 26791 7453 26811 7473
rect 27009 7451 27029 7471
rect 33187 7578 33207 7598
rect 33405 7576 33425 7596
rect 33623 7579 33643 7599
rect 11723 7146 11743 7166
rect 9203 7026 9223 7046
rect 9421 7029 9441 7049
rect 9639 7027 9659 7047
rect 15651 7158 15671 7178
rect 15869 7156 15889 7176
rect 16087 7159 16107 7179
rect 22994 7254 23014 7274
rect 23212 7257 23232 7277
rect 23430 7255 23450 7275
rect 29621 7381 29641 7401
rect 29839 7379 29859 7399
rect 30057 7382 30077 7402
rect 30937 7463 30957 7483
rect 31155 7466 31175 7486
rect 31373 7464 31393 7484
rect 13567 7039 13587 7059
rect 13785 7042 13805 7062
rect 14003 7040 14023 7060
rect 19917 7132 19937 7152
rect 20135 7130 20155 7150
rect 27371 7266 27391 7286
rect 27589 7269 27609 7289
rect 27807 7267 27827 7287
rect 33985 7394 34005 7414
rect 34203 7392 34223 7412
rect 34421 7395 34441 7415
rect 20353 7133 20373 7153
rect 17833 7013 17853 7033
rect 18051 7016 18071 7036
rect 18269 7014 18289 7034
rect 24281 7145 24301 7165
rect 24499 7143 24519 7163
rect 31735 7279 31755 7299
rect 31953 7282 31973 7302
rect 32171 7280 32191 7300
rect 24717 7146 24737 7166
rect 22197 7026 22217 7046
rect 22415 7029 22435 7049
rect 22633 7027 22653 7047
rect 28658 7157 28678 7177
rect 28876 7155 28896 7175
rect 29094 7158 29114 7178
rect 26574 7038 26594 7058
rect 26792 7041 26812 7061
rect 27010 7039 27030 7059
rect 33022 7170 33042 7190
rect 33240 7168 33260 7188
rect 33458 7171 33478 7191
rect 30938 7051 30958 7071
rect 31156 7054 31176 7074
rect 31374 7052 31394 7072
rect 3488 6738 3508 6758
rect 3706 6736 3726 6756
rect 3924 6739 3944 6759
rect 1404 6619 1424 6639
rect 1622 6622 1642 6642
rect 1840 6620 1860 6640
rect 7852 6751 7872 6771
rect 8070 6749 8090 6769
rect 8288 6752 8308 6772
rect 5768 6632 5788 6652
rect 5986 6635 6006 6655
rect 6204 6633 6224 6653
rect 12229 6763 12249 6783
rect 12447 6761 12467 6781
rect 12665 6764 12685 6784
rect 10145 6644 10165 6664
rect 2691 6510 2711 6530
rect 2909 6508 2929 6528
rect 3127 6511 3147 6531
rect 10363 6647 10383 6667
rect 10581 6645 10601 6665
rect 16593 6776 16613 6796
rect 16811 6774 16831 6794
rect 17029 6777 17049 6797
rect 14509 6657 14529 6677
rect 441 6395 461 6415
rect 659 6398 679 6418
rect 877 6396 897 6416
rect 7055 6523 7075 6543
rect 7273 6521 7293 6541
rect 7491 6524 7511 6544
rect 14727 6660 14747 6680
rect 14945 6658 14965 6678
rect 20859 6750 20879 6770
rect 21077 6748 21097 6768
rect 21295 6751 21315 6771
rect 3489 6326 3509 6346
rect 3707 6324 3727 6344
rect 3925 6327 3945 6347
rect 4805 6408 4825 6428
rect 5023 6411 5043 6431
rect 5241 6409 5261 6429
rect 11432 6535 11452 6555
rect 11650 6533 11670 6553
rect 11868 6536 11888 6556
rect 18775 6631 18795 6651
rect 18993 6634 19013 6654
rect 19211 6632 19231 6652
rect 25223 6763 25243 6783
rect 25441 6761 25461 6781
rect 25659 6764 25679 6784
rect 23139 6644 23159 6664
rect 1239 6211 1259 6231
rect 1457 6214 1477 6234
rect 1675 6212 1695 6232
rect 7853 6339 7873 6359
rect 8071 6337 8091 6357
rect 8289 6340 8309 6360
rect 9182 6420 9202 6440
rect 9400 6423 9420 6443
rect 9618 6421 9638 6441
rect 15796 6548 15816 6568
rect 16014 6546 16034 6566
rect 16232 6549 16252 6569
rect 23357 6647 23377 6667
rect 23575 6645 23595 6665
rect 29600 6775 29620 6795
rect 29818 6773 29838 6793
rect 30036 6776 30056 6796
rect 27516 6656 27536 6676
rect 5603 6224 5623 6244
rect 5821 6227 5841 6247
rect 6039 6225 6059 6245
rect 12230 6351 12250 6371
rect 12448 6349 12468 6369
rect 12666 6352 12686 6372
rect 13546 6433 13566 6453
rect 13764 6436 13784 6456
rect 13982 6434 14002 6454
rect 20062 6522 20082 6542
rect 20280 6520 20300 6540
rect 20498 6523 20518 6543
rect 27734 6659 27754 6679
rect 27952 6657 27972 6677
rect 33964 6788 33984 6808
rect 34182 6786 34202 6806
rect 34400 6789 34420 6809
rect 31880 6669 31900 6689
rect 2592 6100 2612 6120
rect 2810 6098 2830 6118
rect 9980 6236 10000 6256
rect 10198 6239 10218 6259
rect 10416 6237 10436 6257
rect 16594 6364 16614 6384
rect 16812 6362 16832 6382
rect 17030 6365 17050 6385
rect 17812 6407 17832 6427
rect 18030 6410 18050 6430
rect 18248 6408 18268 6428
rect 24426 6535 24446 6555
rect 24644 6533 24664 6553
rect 24862 6536 24882 6556
rect 32098 6672 32118 6692
rect 32316 6670 32336 6690
rect 3028 6101 3048 6121
rect 442 5983 462 6003
rect 660 5986 680 6006
rect 878 5984 898 6004
rect 6956 6113 6976 6133
rect 7174 6111 7194 6131
rect 14344 6249 14364 6269
rect 14562 6252 14582 6272
rect 14780 6250 14800 6270
rect 20860 6338 20880 6358
rect 21078 6336 21098 6356
rect 21296 6339 21316 6359
rect 22176 6420 22196 6440
rect 22394 6423 22414 6443
rect 22612 6421 22632 6441
rect 28803 6547 28823 6567
rect 29021 6545 29041 6565
rect 29239 6548 29259 6568
rect 7392 6114 7412 6134
rect 4806 5996 4826 6016
rect 5024 5999 5044 6019
rect 5242 5997 5262 6017
rect 11333 6125 11353 6145
rect 11551 6123 11571 6143
rect 18610 6223 18630 6243
rect 18828 6226 18848 6246
rect 19046 6224 19066 6244
rect 25224 6351 25244 6371
rect 25442 6349 25462 6369
rect 25660 6352 25680 6372
rect 26553 6432 26573 6452
rect 26771 6435 26791 6455
rect 26989 6433 27009 6453
rect 33167 6560 33187 6580
rect 33385 6558 33405 6578
rect 33603 6561 33623 6581
rect 11769 6126 11789 6146
rect 9183 6008 9203 6028
rect 9401 6011 9421 6031
rect 9619 6009 9639 6029
rect 15697 6138 15717 6158
rect 15915 6136 15935 6156
rect 16133 6139 16153 6159
rect 22974 6236 22994 6256
rect 23192 6239 23212 6259
rect 23410 6237 23430 6257
rect 29601 6363 29621 6383
rect 29819 6361 29839 6381
rect 30037 6364 30057 6384
rect 30917 6445 30937 6465
rect 31135 6448 31155 6468
rect 31353 6446 31373 6466
rect 13547 6021 13567 6041
rect 13765 6024 13785 6044
rect 13983 6022 14003 6042
rect 19963 6112 19983 6132
rect 20181 6110 20201 6130
rect 27351 6248 27371 6268
rect 27569 6251 27589 6271
rect 27787 6249 27807 6269
rect 33965 6376 33985 6396
rect 34183 6374 34203 6394
rect 34401 6377 34421 6397
rect 20399 6113 20419 6133
rect 17813 5995 17833 6015
rect 18031 5998 18051 6018
rect 18249 5996 18269 6016
rect 24327 6125 24347 6145
rect 24545 6123 24565 6143
rect 31715 6261 31735 6281
rect 31933 6264 31953 6284
rect 32151 6262 32171 6282
rect 24763 6126 24783 6146
rect 22177 6008 22197 6028
rect 22395 6011 22415 6031
rect 22613 6009 22633 6029
rect 28704 6137 28724 6157
rect 28922 6135 28942 6155
rect 29140 6138 29160 6158
rect 26554 6020 26574 6040
rect 26772 6023 26792 6043
rect 26990 6021 27010 6041
rect 33068 6150 33088 6170
rect 33286 6148 33306 6168
rect 33504 6151 33524 6171
rect 30918 6033 30938 6053
rect 31136 6036 31156 6056
rect 31354 6034 31374 6054
rect 3471 5720 3491 5740
rect 3689 5718 3709 5738
rect 3907 5721 3927 5741
rect 1321 5603 1341 5623
rect 1539 5606 1559 5626
rect 1757 5604 1777 5624
rect 7835 5733 7855 5753
rect 8053 5731 8073 5751
rect 8271 5734 8291 5754
rect 5685 5616 5705 5636
rect 5903 5619 5923 5639
rect 6121 5617 6141 5637
rect 12212 5745 12232 5765
rect 12430 5743 12450 5763
rect 12648 5746 12668 5766
rect 10062 5628 10082 5648
rect 2674 5492 2694 5512
rect 2892 5490 2912 5510
rect 3110 5493 3130 5513
rect 10280 5631 10300 5651
rect 10498 5629 10518 5649
rect 16576 5758 16596 5778
rect 16794 5756 16814 5776
rect 17012 5759 17032 5779
rect 14426 5641 14446 5661
rect 424 5377 444 5397
rect 642 5380 662 5400
rect 860 5378 880 5398
rect 7038 5505 7058 5525
rect 7256 5503 7276 5523
rect 7474 5506 7494 5526
rect 14644 5644 14664 5664
rect 14862 5642 14882 5662
rect 20842 5732 20862 5752
rect 21060 5730 21080 5750
rect 21278 5733 21298 5753
rect 3472 5308 3492 5328
rect 3690 5306 3710 5326
rect 3908 5309 3928 5329
rect 4788 5390 4808 5410
rect 5006 5393 5026 5413
rect 5224 5391 5244 5411
rect 11415 5517 11435 5537
rect 11633 5515 11653 5535
rect 11851 5518 11871 5538
rect 18692 5615 18712 5635
rect 18910 5618 18930 5638
rect 19128 5616 19148 5636
rect 25206 5745 25226 5765
rect 25424 5743 25444 5763
rect 25642 5746 25662 5766
rect 23056 5628 23076 5648
rect 1222 5193 1242 5213
rect 1440 5196 1460 5216
rect 1658 5194 1678 5214
rect 7836 5321 7856 5341
rect 8054 5319 8074 5339
rect 8272 5322 8292 5342
rect 9165 5402 9185 5422
rect 9383 5405 9403 5425
rect 9601 5403 9621 5423
rect 15779 5530 15799 5550
rect 15997 5528 16017 5548
rect 16215 5531 16235 5551
rect 23274 5631 23294 5651
rect 23492 5629 23512 5649
rect 29583 5757 29603 5777
rect 29801 5755 29821 5775
rect 30019 5758 30039 5778
rect 27433 5640 27453 5660
rect 5586 5206 5606 5226
rect 5804 5209 5824 5229
rect 6022 5207 6042 5227
rect 12213 5333 12233 5353
rect 12431 5331 12451 5351
rect 12649 5334 12669 5354
rect 13529 5415 13549 5435
rect 13747 5418 13767 5438
rect 13965 5416 13985 5436
rect 20045 5504 20065 5524
rect 20263 5502 20283 5522
rect 20481 5505 20501 5525
rect 27651 5643 27671 5663
rect 27869 5641 27889 5661
rect 33947 5770 33967 5790
rect 34165 5768 34185 5788
rect 34383 5771 34403 5791
rect 31797 5653 31817 5673
rect 2370 5086 2390 5106
rect 2588 5084 2608 5104
rect 9963 5218 9983 5238
rect 10181 5221 10201 5241
rect 10399 5219 10419 5239
rect 16577 5346 16597 5366
rect 16795 5344 16815 5364
rect 17013 5347 17033 5367
rect 17795 5389 17815 5409
rect 18013 5392 18033 5412
rect 18231 5390 18251 5410
rect 24409 5517 24429 5537
rect 24627 5515 24647 5535
rect 24845 5518 24865 5538
rect 32015 5656 32035 5676
rect 32233 5654 32253 5674
rect 2806 5087 2826 5107
rect 425 4965 445 4985
rect 643 4968 663 4988
rect 861 4966 881 4986
rect 6734 5099 6754 5119
rect 6952 5097 6972 5117
rect 14327 5231 14347 5251
rect 14545 5234 14565 5254
rect 14763 5232 14783 5252
rect 20843 5320 20863 5340
rect 21061 5318 21081 5338
rect 21279 5321 21299 5341
rect 22159 5402 22179 5422
rect 22377 5405 22397 5425
rect 22595 5403 22615 5423
rect 28786 5529 28806 5549
rect 29004 5527 29024 5547
rect 29222 5530 29242 5550
rect 7170 5100 7190 5120
rect 4789 4978 4809 4998
rect 5007 4981 5027 5001
rect 5225 4979 5245 4999
rect 11111 5111 11131 5131
rect 11329 5109 11349 5129
rect 11547 5112 11567 5132
rect 9166 4990 9186 5010
rect 9384 4993 9404 5013
rect 9602 4991 9622 5011
rect 15475 5124 15495 5144
rect 15693 5122 15713 5142
rect 15911 5125 15931 5145
rect 18593 5205 18613 5225
rect 18811 5208 18831 5228
rect 19029 5206 19049 5226
rect 25207 5333 25227 5353
rect 25425 5331 25445 5351
rect 25643 5334 25663 5354
rect 26536 5414 26556 5434
rect 26754 5417 26774 5437
rect 26972 5415 26992 5435
rect 33150 5542 33170 5562
rect 33368 5540 33388 5560
rect 33586 5543 33606 5563
rect 22957 5218 22977 5238
rect 23175 5221 23195 5241
rect 23393 5219 23413 5239
rect 29584 5345 29604 5365
rect 29802 5343 29822 5363
rect 30020 5346 30040 5366
rect 30900 5427 30920 5447
rect 31118 5430 31138 5450
rect 31336 5428 31356 5448
rect 13530 5003 13550 5023
rect 13748 5006 13768 5026
rect 13966 5004 13986 5024
rect 19741 5098 19761 5118
rect 19959 5096 19979 5116
rect 27334 5230 27354 5250
rect 27552 5233 27572 5253
rect 27770 5231 27790 5251
rect 33948 5358 33968 5378
rect 34166 5356 34186 5376
rect 34384 5359 34404 5379
rect 20177 5099 20197 5119
rect 17796 4977 17816 4997
rect 18014 4980 18034 5000
rect 18232 4978 18252 4998
rect 24105 5111 24125 5131
rect 24323 5109 24343 5129
rect 31698 5243 31718 5263
rect 31916 5246 31936 5266
rect 32134 5244 32154 5264
rect 24541 5112 24561 5132
rect 22160 4990 22180 5010
rect 22378 4993 22398 5013
rect 22596 4991 22616 5011
rect 28482 5123 28502 5143
rect 28700 5121 28720 5141
rect 28918 5124 28938 5144
rect 26537 5002 26557 5022
rect 26755 5005 26775 5025
rect 26973 5003 26993 5023
rect 32846 5136 32866 5156
rect 33064 5134 33084 5154
rect 33282 5137 33302 5157
rect 30901 5015 30921 5035
rect 31119 5018 31139 5038
rect 31337 5016 31357 5036
rect 3452 4702 3472 4722
rect 3670 4700 3690 4720
rect 3888 4703 3908 4723
rect 1507 4581 1527 4601
rect 1725 4584 1745 4604
rect 1943 4582 1963 4602
rect 7816 4715 7836 4735
rect 8034 4713 8054 4733
rect 8252 4716 8272 4736
rect 5871 4594 5891 4614
rect 6089 4597 6109 4617
rect 6307 4595 6327 4615
rect 12193 4727 12213 4747
rect 12411 4725 12431 4745
rect 12629 4728 12649 4748
rect 10248 4606 10268 4626
rect 2655 4474 2675 4494
rect 2873 4472 2893 4492
rect 3091 4475 3111 4495
rect 10466 4609 10486 4629
rect 10684 4607 10704 4627
rect 16557 4740 16577 4760
rect 16775 4738 16795 4758
rect 16993 4741 17013 4761
rect 14612 4619 14632 4639
rect 405 4359 425 4379
rect 623 4362 643 4382
rect 841 4360 861 4380
rect 7019 4487 7039 4507
rect 7237 4485 7257 4505
rect 7455 4488 7475 4508
rect 14830 4622 14850 4642
rect 15048 4620 15068 4640
rect 20823 4714 20843 4734
rect 21041 4712 21061 4732
rect 21259 4715 21279 4735
rect 3453 4290 3473 4310
rect 3671 4288 3691 4308
rect 3889 4291 3909 4311
rect 4769 4372 4789 4392
rect 4987 4375 5007 4395
rect 5205 4373 5225 4393
rect 11396 4499 11416 4519
rect 11614 4497 11634 4517
rect 11832 4500 11852 4520
rect 1203 4175 1223 4195
rect 1421 4178 1441 4198
rect 1639 4176 1659 4196
rect 7817 4303 7837 4323
rect 8035 4301 8055 4321
rect 8253 4304 8273 4324
rect 9146 4384 9166 4404
rect 9364 4387 9384 4407
rect 9582 4385 9602 4405
rect 15760 4512 15780 4532
rect 15978 4510 15998 4530
rect 16196 4513 16216 4533
rect 18878 4593 18898 4613
rect 19096 4596 19116 4616
rect 19314 4594 19334 4614
rect 25187 4727 25207 4747
rect 25405 4725 25425 4745
rect 25623 4728 25643 4748
rect 23242 4606 23262 4626
rect 23460 4609 23480 4629
rect 23678 4607 23698 4627
rect 29564 4739 29584 4759
rect 29782 4737 29802 4757
rect 30000 4740 30020 4760
rect 27619 4618 27639 4638
rect 5567 4188 5587 4208
rect 5785 4191 5805 4211
rect 6003 4189 6023 4209
rect 12194 4315 12214 4335
rect 12412 4313 12432 4333
rect 12630 4316 12650 4336
rect 13510 4397 13530 4417
rect 13728 4400 13748 4420
rect 13946 4398 13966 4418
rect 20026 4486 20046 4506
rect 20244 4484 20264 4504
rect 20462 4487 20482 4507
rect 27837 4621 27857 4641
rect 28055 4619 28075 4639
rect 33928 4752 33948 4772
rect 34146 4750 34166 4770
rect 34364 4753 34384 4773
rect 31983 4631 32003 4651
rect 2556 4064 2576 4084
rect 2774 4062 2794 4082
rect 9944 4200 9964 4220
rect 10162 4203 10182 4223
rect 10380 4201 10400 4221
rect 16558 4328 16578 4348
rect 16776 4326 16796 4346
rect 16994 4329 17014 4349
rect 17776 4371 17796 4391
rect 17994 4374 18014 4394
rect 18212 4372 18232 4392
rect 24390 4499 24410 4519
rect 24608 4497 24628 4517
rect 24826 4500 24846 4520
rect 32201 4634 32221 4654
rect 32419 4632 32439 4652
rect 2992 4065 3012 4085
rect 406 3947 426 3967
rect 624 3950 644 3970
rect 842 3948 862 3968
rect 6920 4077 6940 4097
rect 7138 4075 7158 4095
rect 14308 4213 14328 4233
rect 14526 4216 14546 4236
rect 14744 4214 14764 4234
rect 20824 4302 20844 4322
rect 21042 4300 21062 4320
rect 21260 4303 21280 4323
rect 22140 4384 22160 4404
rect 22358 4387 22378 4407
rect 22576 4385 22596 4405
rect 28767 4511 28787 4531
rect 28985 4509 29005 4529
rect 29203 4512 29223 4532
rect 7356 4078 7376 4098
rect 4770 3960 4790 3980
rect 4988 3963 5008 3983
rect 5206 3961 5226 3981
rect 11297 4089 11317 4109
rect 11515 4087 11535 4107
rect 18574 4187 18594 4207
rect 18792 4190 18812 4210
rect 19010 4188 19030 4208
rect 25188 4315 25208 4335
rect 25406 4313 25426 4333
rect 25624 4316 25644 4336
rect 26517 4396 26537 4416
rect 26735 4399 26755 4419
rect 26953 4397 26973 4417
rect 33131 4524 33151 4544
rect 33349 4522 33369 4542
rect 33567 4525 33587 4545
rect 11733 4090 11753 4110
rect 9147 3972 9167 3992
rect 9365 3975 9385 3995
rect 9583 3973 9603 3993
rect 15661 4102 15681 4122
rect 15879 4100 15899 4120
rect 16097 4103 16117 4123
rect 22938 4200 22958 4220
rect 23156 4203 23176 4223
rect 23374 4201 23394 4221
rect 29565 4327 29585 4347
rect 29783 4325 29803 4345
rect 30001 4328 30021 4348
rect 30881 4409 30901 4429
rect 31099 4412 31119 4432
rect 31317 4410 31337 4430
rect 13511 3985 13531 4005
rect 13729 3988 13749 4008
rect 13947 3986 13967 4006
rect 19927 4076 19947 4096
rect 20145 4074 20165 4094
rect 27315 4212 27335 4232
rect 27533 4215 27553 4235
rect 27751 4213 27771 4233
rect 33929 4340 33949 4360
rect 34147 4338 34167 4358
rect 34365 4341 34385 4361
rect 20363 4077 20383 4097
rect 17777 3959 17797 3979
rect 17995 3962 18015 3982
rect 18213 3960 18233 3980
rect 24291 4089 24311 4109
rect 24509 4087 24529 4107
rect 31679 4225 31699 4245
rect 31897 4228 31917 4248
rect 32115 4226 32135 4246
rect 24727 4090 24747 4110
rect 22141 3972 22161 3992
rect 22359 3975 22379 3995
rect 22577 3973 22597 3993
rect 28668 4101 28688 4121
rect 28886 4099 28906 4119
rect 29104 4102 29124 4122
rect 26518 3984 26538 4004
rect 26736 3987 26756 4007
rect 26954 3985 26974 4005
rect 33032 4114 33052 4134
rect 33250 4112 33270 4132
rect 33468 4115 33488 4135
rect 30882 3997 30902 4017
rect 31100 4000 31120 4020
rect 31318 3998 31338 4018
rect 3435 3684 3455 3704
rect 3653 3682 3673 3702
rect 3871 3685 3891 3705
rect 1285 3567 1305 3587
rect 1503 3570 1523 3590
rect 1721 3568 1741 3588
rect 7799 3697 7819 3717
rect 8017 3695 8037 3715
rect 8235 3698 8255 3718
rect 5649 3580 5669 3600
rect 5867 3583 5887 3603
rect 6085 3581 6105 3601
rect 12176 3709 12196 3729
rect 12394 3707 12414 3727
rect 12612 3710 12632 3730
rect 10026 3592 10046 3612
rect 2638 3456 2658 3476
rect 2856 3454 2876 3474
rect 3074 3457 3094 3477
rect 10244 3595 10264 3615
rect 10462 3593 10482 3613
rect 16540 3722 16560 3742
rect 16758 3720 16778 3740
rect 16976 3723 16996 3743
rect 14390 3605 14410 3625
rect 388 3341 408 3361
rect 606 3344 626 3364
rect 824 3342 844 3362
rect 7002 3469 7022 3489
rect 7220 3467 7240 3487
rect 7438 3470 7458 3490
rect 14608 3608 14628 3628
rect 14826 3606 14846 3626
rect 20806 3696 20826 3716
rect 21024 3694 21044 3714
rect 21242 3697 21262 3717
rect 3436 3272 3456 3292
rect 3654 3270 3674 3290
rect 3872 3273 3892 3293
rect 4752 3354 4772 3374
rect 4970 3357 4990 3377
rect 5188 3355 5208 3375
rect 11379 3481 11399 3501
rect 11597 3479 11617 3499
rect 11815 3482 11835 3502
rect 18656 3579 18676 3599
rect 18874 3582 18894 3602
rect 19092 3580 19112 3600
rect 25170 3709 25190 3729
rect 25388 3707 25408 3727
rect 25606 3710 25626 3730
rect 23020 3592 23040 3612
rect 1186 3157 1206 3177
rect 1404 3160 1424 3180
rect 1622 3158 1642 3178
rect 7800 3285 7820 3305
rect 8018 3283 8038 3303
rect 8236 3286 8256 3306
rect 9129 3366 9149 3386
rect 9347 3369 9367 3389
rect 9565 3367 9585 3387
rect 15743 3494 15763 3514
rect 15961 3492 15981 3512
rect 16179 3495 16199 3515
rect 23238 3595 23258 3615
rect 23456 3593 23476 3613
rect 29547 3721 29567 3741
rect 29765 3719 29785 3739
rect 29983 3722 30003 3742
rect 27397 3604 27417 3624
rect 5550 3170 5570 3190
rect 5768 3173 5788 3193
rect 5986 3171 6006 3191
rect 12177 3297 12197 3317
rect 12395 3295 12415 3315
rect 12613 3298 12633 3318
rect 13493 3379 13513 3399
rect 13711 3382 13731 3402
rect 13929 3380 13949 3400
rect 20009 3468 20029 3488
rect 20227 3466 20247 3486
rect 20445 3469 20465 3489
rect 27615 3607 27635 3627
rect 27833 3605 27853 3625
rect 33911 3734 33931 3754
rect 34129 3732 34149 3752
rect 34347 3735 34367 3755
rect 31761 3617 31781 3637
rect 2473 3048 2493 3068
rect 2691 3046 2711 3066
rect 9927 3182 9947 3202
rect 10145 3185 10165 3205
rect 10363 3183 10383 3203
rect 16541 3310 16561 3330
rect 16759 3308 16779 3328
rect 16977 3311 16997 3331
rect 17759 3353 17779 3373
rect 17977 3356 17997 3376
rect 18195 3354 18215 3374
rect 24373 3481 24393 3501
rect 24591 3479 24611 3499
rect 24809 3482 24829 3502
rect 31979 3620 31999 3640
rect 32197 3618 32217 3638
rect 2909 3049 2929 3069
rect 389 2929 409 2949
rect 607 2932 627 2952
rect 825 2930 845 2950
rect 6837 3061 6857 3081
rect 7055 3059 7075 3079
rect 14291 3195 14311 3215
rect 14509 3198 14529 3218
rect 14727 3196 14747 3216
rect 20807 3284 20827 3304
rect 21025 3282 21045 3302
rect 21243 3285 21263 3305
rect 22123 3366 22143 3386
rect 22341 3369 22361 3389
rect 22559 3367 22579 3387
rect 28750 3493 28770 3513
rect 28968 3491 28988 3511
rect 29186 3494 29206 3514
rect 7273 3062 7293 3082
rect 4753 2942 4773 2962
rect 4971 2945 4991 2965
rect 5189 2943 5209 2963
rect 11214 3073 11234 3093
rect 11432 3071 11452 3091
rect 18557 3169 18577 3189
rect 18775 3172 18795 3192
rect 18993 3170 19013 3190
rect 25171 3297 25191 3317
rect 25389 3295 25409 3315
rect 25607 3298 25627 3318
rect 26500 3378 26520 3398
rect 26718 3381 26738 3401
rect 26936 3379 26956 3399
rect 33114 3506 33134 3526
rect 33332 3504 33352 3524
rect 33550 3507 33570 3527
rect 11650 3074 11670 3094
rect 9130 2954 9150 2974
rect 9348 2957 9368 2977
rect 9566 2955 9586 2975
rect 15578 3086 15598 3106
rect 15796 3084 15816 3104
rect 16014 3087 16034 3107
rect 22921 3182 22941 3202
rect 23139 3185 23159 3205
rect 23357 3183 23377 3203
rect 29548 3309 29568 3329
rect 29766 3307 29786 3327
rect 29984 3310 30004 3330
rect 30864 3391 30884 3411
rect 31082 3394 31102 3414
rect 31300 3392 31320 3412
rect 13494 2967 13514 2987
rect 13712 2970 13732 2990
rect 13930 2968 13950 2988
rect 19844 3060 19864 3080
rect 20062 3058 20082 3078
rect 27298 3194 27318 3214
rect 27516 3197 27536 3217
rect 27734 3195 27754 3215
rect 33912 3322 33932 3342
rect 34130 3320 34150 3340
rect 34348 3323 34368 3343
rect 20280 3061 20300 3081
rect 17760 2941 17780 2961
rect 17978 2944 17998 2964
rect 18196 2942 18216 2962
rect 24208 3073 24228 3093
rect 24426 3071 24446 3091
rect 31662 3207 31682 3227
rect 31880 3210 31900 3230
rect 32098 3208 32118 3228
rect 24644 3074 24664 3094
rect 22124 2954 22144 2974
rect 22342 2957 22362 2977
rect 22560 2955 22580 2975
rect 28585 3085 28605 3105
rect 28803 3083 28823 3103
rect 29021 3086 29041 3106
rect 26501 2966 26521 2986
rect 26719 2969 26739 2989
rect 26937 2967 26957 2987
rect 32949 3098 32969 3118
rect 33167 3096 33187 3116
rect 33385 3099 33405 3119
rect 30865 2979 30885 2999
rect 31083 2982 31103 3002
rect 31301 2980 31321 3000
rect 3415 2666 3435 2686
rect 3633 2664 3653 2684
rect 3851 2667 3871 2687
rect 1331 2547 1351 2567
rect 1549 2550 1569 2570
rect 1767 2548 1787 2568
rect 7779 2679 7799 2699
rect 7997 2677 8017 2697
rect 8215 2680 8235 2700
rect 5695 2560 5715 2580
rect 5913 2563 5933 2583
rect 6131 2561 6151 2581
rect 12156 2691 12176 2711
rect 12374 2689 12394 2709
rect 12592 2692 12612 2712
rect 10072 2572 10092 2592
rect 2618 2438 2638 2458
rect 2836 2436 2856 2456
rect 3054 2439 3074 2459
rect 10290 2575 10310 2595
rect 10508 2573 10528 2593
rect 16520 2704 16540 2724
rect 16738 2702 16758 2722
rect 16956 2705 16976 2725
rect 14436 2585 14456 2605
rect 368 2323 388 2343
rect 586 2326 606 2346
rect 804 2324 824 2344
rect 6982 2451 7002 2471
rect 7200 2449 7220 2469
rect 7418 2452 7438 2472
rect 14654 2588 14674 2608
rect 14872 2586 14892 2606
rect 20786 2678 20806 2698
rect 21004 2676 21024 2696
rect 21222 2679 21242 2699
rect 3416 2254 3436 2274
rect 3634 2252 3654 2272
rect 3852 2255 3872 2275
rect 4732 2336 4752 2356
rect 4950 2339 4970 2359
rect 5168 2337 5188 2357
rect 11359 2463 11379 2483
rect 11577 2461 11597 2481
rect 11795 2464 11815 2484
rect 18702 2559 18722 2579
rect 18920 2562 18940 2582
rect 19138 2560 19158 2580
rect 25150 2691 25170 2711
rect 25368 2689 25388 2709
rect 25586 2692 25606 2712
rect 23066 2572 23086 2592
rect 1166 2139 1186 2159
rect 1384 2142 1404 2162
rect 1602 2140 1622 2160
rect 7780 2267 7800 2287
rect 7998 2265 8018 2285
rect 8216 2268 8236 2288
rect 9109 2348 9129 2368
rect 9327 2351 9347 2371
rect 9545 2349 9565 2369
rect 15723 2476 15743 2496
rect 15941 2474 15961 2494
rect 16159 2477 16179 2497
rect 23284 2575 23304 2595
rect 23502 2573 23522 2593
rect 29527 2703 29547 2723
rect 29745 2701 29765 2721
rect 29963 2704 29983 2724
rect 27443 2584 27463 2604
rect 5530 2152 5550 2172
rect 5748 2155 5768 2175
rect 5966 2153 5986 2173
rect 12157 2279 12177 2299
rect 12375 2277 12395 2297
rect 12593 2280 12613 2300
rect 13473 2361 13493 2381
rect 13691 2364 13711 2384
rect 13909 2362 13929 2382
rect 19989 2450 20009 2470
rect 20207 2448 20227 2468
rect 20425 2451 20445 2471
rect 27661 2587 27681 2607
rect 27879 2585 27899 2605
rect 33891 2716 33911 2736
rect 34109 2714 34129 2734
rect 34327 2717 34347 2737
rect 31807 2597 31827 2617
rect 2519 2028 2539 2048
rect 2737 2026 2757 2046
rect 9907 2164 9927 2184
rect 10125 2167 10145 2187
rect 10343 2165 10363 2185
rect 16521 2292 16541 2312
rect 16739 2290 16759 2310
rect 16957 2293 16977 2313
rect 17739 2335 17759 2355
rect 17957 2338 17977 2358
rect 18175 2336 18195 2356
rect 24353 2463 24373 2483
rect 24571 2461 24591 2481
rect 24789 2464 24809 2484
rect 32025 2600 32045 2620
rect 32243 2598 32263 2618
rect 2955 2029 2975 2049
rect 369 1911 389 1931
rect 587 1914 607 1934
rect 805 1912 825 1932
rect 6883 2041 6903 2061
rect 7101 2039 7121 2059
rect 14271 2177 14291 2197
rect 14489 2180 14509 2200
rect 14707 2178 14727 2198
rect 20787 2266 20807 2286
rect 21005 2264 21025 2284
rect 21223 2267 21243 2287
rect 22103 2348 22123 2368
rect 22321 2351 22341 2371
rect 22539 2349 22559 2369
rect 28730 2475 28750 2495
rect 28948 2473 28968 2493
rect 29166 2476 29186 2496
rect 7319 2042 7339 2062
rect 4733 1924 4753 1944
rect 4951 1927 4971 1947
rect 5169 1925 5189 1945
rect 11260 2053 11280 2073
rect 11478 2051 11498 2071
rect 18537 2151 18557 2171
rect 18755 2154 18775 2174
rect 18973 2152 18993 2172
rect 25151 2279 25171 2299
rect 25369 2277 25389 2297
rect 25587 2280 25607 2300
rect 26480 2360 26500 2380
rect 26698 2363 26718 2383
rect 26916 2361 26936 2381
rect 33094 2488 33114 2508
rect 33312 2486 33332 2506
rect 33530 2489 33550 2509
rect 11696 2054 11716 2074
rect 9110 1936 9130 1956
rect 9328 1939 9348 1959
rect 9546 1937 9566 1957
rect 15624 2066 15644 2086
rect 15842 2064 15862 2084
rect 16060 2067 16080 2087
rect 22901 2164 22921 2184
rect 23119 2167 23139 2187
rect 23337 2165 23357 2185
rect 29528 2291 29548 2311
rect 29746 2289 29766 2309
rect 29964 2292 29984 2312
rect 30844 2373 30864 2393
rect 31062 2376 31082 2396
rect 31280 2374 31300 2394
rect 13474 1949 13494 1969
rect 13692 1952 13712 1972
rect 13910 1950 13930 1970
rect 19890 2040 19910 2060
rect 20108 2038 20128 2058
rect 27278 2176 27298 2196
rect 27496 2179 27516 2199
rect 27714 2177 27734 2197
rect 33892 2304 33912 2324
rect 34110 2302 34130 2322
rect 34328 2305 34348 2325
rect 20326 2041 20346 2061
rect 17740 1923 17760 1943
rect 17958 1926 17978 1946
rect 18176 1924 18196 1944
rect 24254 2053 24274 2073
rect 24472 2051 24492 2071
rect 31642 2189 31662 2209
rect 31860 2192 31880 2212
rect 32078 2190 32098 2210
rect 24690 2054 24710 2074
rect 22104 1936 22124 1956
rect 22322 1939 22342 1959
rect 22540 1937 22560 1957
rect 28631 2065 28651 2085
rect 28849 2063 28869 2083
rect 29067 2066 29087 2086
rect 26481 1948 26501 1968
rect 26699 1951 26719 1971
rect 26917 1949 26937 1969
rect 32995 2078 33015 2098
rect 33213 2076 33233 2096
rect 33431 2079 33451 2099
rect 30845 1961 30865 1981
rect 31063 1964 31083 1984
rect 31281 1962 31301 1982
rect 3398 1648 3418 1668
rect 3616 1646 3636 1666
rect 3834 1649 3854 1669
rect 1248 1531 1268 1551
rect 1466 1534 1486 1554
rect 1684 1532 1704 1552
rect 7762 1661 7782 1681
rect 7980 1659 8000 1679
rect 8198 1662 8218 1682
rect 5612 1544 5632 1564
rect 5830 1547 5850 1567
rect 6048 1545 6068 1565
rect 12139 1673 12159 1693
rect 12357 1671 12377 1691
rect 12575 1674 12595 1694
rect 9989 1556 10009 1576
rect 2601 1420 2621 1440
rect 2819 1418 2839 1438
rect 3037 1421 3057 1441
rect 10207 1559 10227 1579
rect 10425 1557 10445 1577
rect 16503 1686 16523 1706
rect 16721 1684 16741 1704
rect 16939 1687 16959 1707
rect 14353 1569 14373 1589
rect 351 1305 371 1325
rect 569 1308 589 1328
rect 787 1306 807 1326
rect 6965 1433 6985 1453
rect 7183 1431 7203 1451
rect 7401 1434 7421 1454
rect 14571 1572 14591 1592
rect 14789 1570 14809 1590
rect 20769 1660 20789 1680
rect 20987 1658 21007 1678
rect 21205 1661 21225 1681
rect 3399 1236 3419 1256
rect 3617 1234 3637 1254
rect 3835 1237 3855 1257
rect 4715 1318 4735 1338
rect 4933 1321 4953 1341
rect 5151 1319 5171 1339
rect 11342 1445 11362 1465
rect 11560 1443 11580 1463
rect 11778 1446 11798 1466
rect 18619 1543 18639 1563
rect 18837 1546 18857 1566
rect 19055 1544 19075 1564
rect 25133 1673 25153 1693
rect 25351 1671 25371 1691
rect 25569 1674 25589 1694
rect 22983 1556 23003 1576
rect 1149 1121 1169 1141
rect 1367 1124 1387 1144
rect 1585 1122 1605 1142
rect 7763 1249 7783 1269
rect 7981 1247 8001 1267
rect 8199 1250 8219 1270
rect 9092 1330 9112 1350
rect 9310 1333 9330 1353
rect 9528 1331 9548 1351
rect 15706 1458 15726 1478
rect 15924 1456 15944 1476
rect 16142 1459 16162 1479
rect 23201 1559 23221 1579
rect 23419 1557 23439 1577
rect 29510 1685 29530 1705
rect 29728 1683 29748 1703
rect 29946 1686 29966 1706
rect 27360 1568 27380 1588
rect 5513 1134 5533 1154
rect 5731 1137 5751 1157
rect 5949 1135 5969 1155
rect 12140 1261 12160 1281
rect 12358 1259 12378 1279
rect 12576 1262 12596 1282
rect 13456 1343 13476 1363
rect 13674 1346 13694 1366
rect 13892 1344 13912 1364
rect 19972 1432 19992 1452
rect 20190 1430 20210 1450
rect 20408 1433 20428 1453
rect 27578 1571 27598 1591
rect 27796 1569 27816 1589
rect 33874 1698 33894 1718
rect 34092 1696 34112 1716
rect 34310 1699 34330 1719
rect 31724 1581 31744 1601
rect 9890 1146 9910 1166
rect 10108 1149 10128 1169
rect 10326 1147 10346 1167
rect 16504 1274 16524 1294
rect 16722 1272 16742 1292
rect 16940 1275 16960 1295
rect 17722 1317 17742 1337
rect 17940 1320 17960 1340
rect 18158 1318 18178 1338
rect 24336 1445 24356 1465
rect 24554 1443 24574 1463
rect 24772 1446 24792 1466
rect 31942 1584 31962 1604
rect 32160 1582 32180 1602
rect 14254 1159 14274 1179
rect 14472 1162 14492 1182
rect 14690 1160 14710 1180
rect 20770 1248 20790 1268
rect 20988 1246 21008 1266
rect 21206 1249 21226 1269
rect 22086 1330 22106 1350
rect 22304 1333 22324 1353
rect 22522 1331 22542 1351
rect 28713 1457 28733 1477
rect 28931 1455 28951 1475
rect 29149 1458 29169 1478
rect 352 893 372 913
rect 570 896 590 916
rect 788 894 808 914
rect 4716 906 4736 926
rect 4934 909 4954 929
rect 18520 1133 18540 1153
rect 18738 1136 18758 1156
rect 18956 1134 18976 1154
rect 25134 1261 25154 1281
rect 25352 1259 25372 1279
rect 25570 1262 25590 1282
rect 26463 1342 26483 1362
rect 26681 1345 26701 1365
rect 26899 1343 26919 1363
rect 33077 1470 33097 1490
rect 33295 1468 33315 1488
rect 33513 1471 33533 1491
rect 22884 1146 22904 1166
rect 23102 1149 23122 1169
rect 23320 1147 23340 1167
rect 29511 1273 29531 1293
rect 29729 1271 29749 1291
rect 29947 1274 29967 1294
rect 30827 1355 30847 1375
rect 31045 1358 31065 1378
rect 31263 1356 31283 1376
rect 27261 1158 27281 1178
rect 27479 1161 27499 1181
rect 27697 1159 27717 1179
rect 33875 1286 33895 1306
rect 34093 1284 34113 1304
rect 34311 1287 34331 1307
rect 31625 1171 31645 1191
rect 31843 1174 31863 1194
rect 32061 1172 32081 1192
rect 5152 907 5172 927
rect 9093 918 9113 938
rect 9311 921 9331 941
rect 9529 919 9549 939
rect 13457 931 13477 951
rect 13675 934 13695 954
rect 13893 932 13913 952
rect 17723 905 17743 925
rect 17941 908 17961 928
rect 18159 906 18179 926
rect 22087 918 22107 938
rect 22305 921 22325 941
rect 22523 919 22543 939
rect 26464 930 26484 950
rect 26682 933 26702 953
rect 26900 931 26920 951
rect 30828 943 30848 963
rect 31046 946 31066 966
rect 31264 944 31284 964
rect 1565 317 1585 337
rect 1783 320 1803 340
rect 2001 318 2021 338
rect 5929 330 5949 350
rect 6147 333 6167 353
rect 6365 331 6385 351
rect 10306 342 10326 362
rect 4054 243 4074 263
rect 4272 246 4292 266
rect 4490 244 4510 264
rect 8502 267 8522 287
rect 8720 270 8740 290
rect 10524 345 10544 365
rect 10742 343 10762 363
rect 14670 355 14690 375
rect 14888 358 14908 378
rect 15106 356 15126 376
rect 8938 268 8958 288
rect 12795 268 12815 288
rect 13013 271 13033 291
rect 13231 269 13251 289
rect 18936 329 18956 349
rect 19154 332 19174 352
rect 19372 330 19392 350
rect 23300 342 23320 362
rect 23518 345 23538 365
rect 23736 343 23756 363
rect 27677 354 27697 374
rect 16992 204 17012 224
rect 17210 207 17230 227
rect 21425 255 21445 275
rect 21643 258 21663 278
rect 21861 256 21881 276
rect 25873 279 25893 299
rect 26091 282 26111 302
rect 27895 357 27915 377
rect 28113 355 28133 375
rect 32041 367 32061 387
rect 32259 370 32279 390
rect 32477 368 32497 388
rect 26309 280 26329 300
rect 30166 280 30186 300
rect 30384 283 30404 303
rect 30602 281 30622 301
rect 17428 205 17448 225
<< ndiffres >>
rect 4181 8859 4238 8878
rect 4181 8841 4199 8859
rect 4217 8856 4238 8859
rect 4217 8841 4332 8856
rect 240 8801 301 8817
rect 145 8797 301 8801
rect 145 8779 263 8797
rect 281 8779 301 8797
rect 145 8758 301 8779
rect 145 8757 245 8758
rect 146 8721 188 8757
rect 4181 8818 4332 8841
rect 8545 8872 8602 8891
rect 8545 8854 8563 8872
rect 8581 8869 8602 8872
rect 8581 8854 8696 8869
rect 4290 8782 4332 8818
rect 4604 8814 4665 8830
rect 4509 8810 4665 8814
rect 4509 8792 4627 8810
rect 4645 8792 4665 8810
rect 4233 8781 4333 8782
rect 4177 8760 4333 8781
rect 4509 8771 4665 8792
rect 4509 8770 4609 8771
rect 146 8698 297 8721
rect 146 8683 261 8698
rect 240 8680 261 8683
rect 279 8680 297 8698
rect 240 8661 297 8680
rect 4177 8742 4197 8760
rect 4215 8742 4333 8760
rect 4177 8738 4333 8742
rect 4177 8722 4238 8738
rect 4510 8734 4552 8770
rect 8545 8831 8696 8854
rect 12922 8884 12979 8903
rect 12922 8866 12940 8884
rect 12958 8881 12979 8884
rect 12958 8866 13073 8881
rect 8654 8795 8696 8831
rect 8981 8826 9042 8842
rect 8886 8822 9042 8826
rect 8886 8804 9004 8822
rect 9022 8804 9042 8822
rect 8597 8794 8697 8795
rect 8541 8773 8697 8794
rect 8886 8783 9042 8804
rect 8886 8782 8986 8783
rect 4510 8711 4661 8734
rect 4510 8696 4625 8711
rect 4604 8693 4625 8696
rect 4643 8693 4661 8711
rect 4604 8674 4661 8693
rect 4174 8641 4231 8660
rect 8541 8755 8561 8773
rect 8579 8755 8697 8773
rect 8541 8751 8697 8755
rect 8541 8735 8602 8751
rect 8887 8746 8929 8782
rect 12922 8843 13073 8866
rect 17286 8897 17343 8916
rect 17286 8879 17304 8897
rect 17322 8894 17343 8897
rect 17322 8879 17437 8894
rect 13031 8807 13073 8843
rect 13345 8839 13406 8855
rect 13250 8835 13406 8839
rect 13250 8817 13368 8835
rect 13386 8817 13406 8835
rect 12974 8806 13074 8807
rect 12918 8785 13074 8806
rect 13250 8796 13406 8817
rect 13250 8795 13350 8796
rect 8887 8723 9038 8746
rect 8887 8708 9002 8723
rect 8981 8705 9002 8708
rect 9020 8705 9038 8723
rect 8981 8686 9038 8705
rect 4174 8623 4192 8641
rect 4210 8638 4231 8641
rect 4210 8623 4325 8638
rect 4174 8600 4325 8623
rect 8538 8654 8595 8673
rect 12918 8767 12938 8785
rect 12956 8767 13074 8785
rect 12918 8763 13074 8767
rect 12918 8747 12979 8763
rect 13251 8759 13293 8795
rect 17286 8856 17437 8879
rect 17395 8820 17437 8856
rect 21552 8871 21609 8890
rect 21552 8853 21570 8871
rect 21588 8868 21609 8871
rect 21588 8853 21703 8868
rect 17338 8819 17438 8820
rect 17282 8798 17438 8819
rect 17611 8813 17672 8829
rect 13251 8736 13402 8759
rect 13251 8721 13366 8736
rect 13345 8718 13366 8721
rect 13384 8718 13402 8736
rect 13345 8699 13402 8718
rect 8538 8636 8556 8654
rect 8574 8651 8595 8654
rect 8574 8636 8689 8651
rect 8538 8613 8689 8636
rect 12915 8666 12972 8685
rect 17282 8780 17302 8798
rect 17320 8780 17438 8798
rect 17282 8776 17438 8780
rect 17516 8809 17672 8813
rect 17516 8791 17634 8809
rect 17652 8791 17672 8809
rect 17282 8760 17343 8776
rect 17516 8770 17672 8791
rect 17516 8769 17616 8770
rect 17517 8733 17559 8769
rect 21552 8830 21703 8853
rect 25916 8884 25973 8903
rect 25916 8866 25934 8884
rect 25952 8881 25973 8884
rect 25952 8866 26067 8881
rect 21661 8794 21703 8830
rect 21975 8826 22036 8842
rect 21880 8822 22036 8826
rect 21880 8804 21998 8822
rect 22016 8804 22036 8822
rect 21604 8793 21704 8794
rect 21548 8772 21704 8793
rect 21880 8783 22036 8804
rect 21880 8782 21980 8783
rect 17517 8710 17668 8733
rect 12915 8648 12933 8666
rect 12951 8663 12972 8666
rect 12951 8648 13066 8663
rect 12915 8625 13066 8648
rect 17279 8679 17336 8698
rect 17517 8695 17632 8710
rect 17279 8661 17297 8679
rect 17315 8676 17336 8679
rect 17611 8692 17632 8695
rect 17650 8692 17668 8710
rect 17315 8661 17430 8676
rect 17611 8673 17668 8692
rect 17279 8638 17430 8661
rect 21548 8754 21568 8772
rect 21586 8754 21704 8772
rect 21548 8750 21704 8754
rect 21548 8734 21609 8750
rect 21881 8746 21923 8782
rect 25916 8843 26067 8866
rect 30293 8896 30350 8915
rect 30293 8878 30311 8896
rect 30329 8893 30350 8896
rect 30329 8878 30444 8893
rect 26025 8807 26067 8843
rect 26352 8838 26413 8854
rect 26257 8834 26413 8838
rect 26257 8816 26375 8834
rect 26393 8816 26413 8834
rect 25968 8806 26068 8807
rect 25912 8785 26068 8806
rect 26257 8795 26413 8816
rect 26257 8794 26357 8795
rect 21881 8723 22032 8746
rect 21881 8708 21996 8723
rect 21975 8705 21996 8708
rect 22014 8705 22032 8723
rect 21975 8686 22032 8705
rect 235 8477 296 8493
rect 4283 8564 4325 8600
rect 4226 8563 4326 8564
rect 4170 8542 4326 8563
rect 4170 8524 4190 8542
rect 4208 8524 4326 8542
rect 4170 8520 4326 8524
rect 140 8473 296 8477
rect 140 8455 258 8473
rect 276 8455 296 8473
rect 140 8434 296 8455
rect 140 8433 240 8434
rect 141 8397 183 8433
rect 4170 8504 4231 8520
rect 4599 8490 4660 8506
rect 8647 8577 8689 8613
rect 8590 8576 8690 8577
rect 8534 8555 8690 8576
rect 8534 8537 8554 8555
rect 8572 8537 8690 8555
rect 8534 8533 8690 8537
rect 4504 8486 4660 8490
rect 4168 8458 4225 8477
rect 141 8374 292 8397
rect 141 8359 256 8374
rect 235 8356 256 8359
rect 274 8356 292 8374
rect 4168 8440 4186 8458
rect 4204 8455 4225 8458
rect 4504 8468 4622 8486
rect 4640 8468 4660 8486
rect 4204 8440 4319 8455
rect 4504 8447 4660 8468
rect 4504 8446 4604 8447
rect 4168 8417 4319 8440
rect 235 8337 292 8356
rect 229 8294 290 8310
rect 4277 8381 4319 8417
rect 4505 8410 4547 8446
rect 8534 8517 8595 8533
rect 8976 8502 9037 8518
rect 13024 8589 13066 8625
rect 12967 8588 13067 8589
rect 12911 8567 13067 8588
rect 12911 8549 12931 8567
rect 12949 8549 13067 8567
rect 12911 8545 13067 8549
rect 8881 8498 9037 8502
rect 8532 8471 8589 8490
rect 4505 8387 4656 8410
rect 4220 8380 4320 8381
rect 4164 8359 4320 8380
rect 4505 8372 4620 8387
rect 4164 8341 4184 8359
rect 4202 8341 4320 8359
rect 4599 8369 4620 8372
rect 4638 8369 4656 8387
rect 8532 8453 8550 8471
rect 8568 8468 8589 8471
rect 8881 8480 8999 8498
rect 9017 8480 9037 8498
rect 8568 8453 8683 8468
rect 8881 8459 9037 8480
rect 8881 8458 8981 8459
rect 8532 8430 8683 8453
rect 4599 8350 4656 8369
rect 4164 8337 4320 8341
rect 134 8290 290 8294
rect 134 8272 252 8290
rect 270 8272 290 8290
rect 134 8251 290 8272
rect 134 8250 234 8251
rect 135 8214 177 8250
rect 4164 8321 4225 8337
rect 4593 8307 4654 8323
rect 8641 8394 8683 8430
rect 8882 8422 8924 8458
rect 12911 8529 12972 8545
rect 13340 8515 13401 8531
rect 17388 8602 17430 8638
rect 21545 8653 21602 8672
rect 25912 8767 25932 8785
rect 25950 8767 26068 8785
rect 25912 8763 26068 8767
rect 25912 8747 25973 8763
rect 26258 8758 26300 8794
rect 30293 8855 30444 8878
rect 34657 8909 34714 8928
rect 34657 8891 34675 8909
rect 34693 8906 34714 8909
rect 34693 8891 34808 8906
rect 30402 8819 30444 8855
rect 30716 8851 30777 8867
rect 30621 8847 30777 8851
rect 30621 8829 30739 8847
rect 30757 8829 30777 8847
rect 30345 8818 30445 8819
rect 30289 8797 30445 8818
rect 30621 8808 30777 8829
rect 30621 8807 30721 8808
rect 26258 8735 26409 8758
rect 26258 8720 26373 8735
rect 26352 8717 26373 8720
rect 26391 8717 26409 8735
rect 26352 8698 26409 8717
rect 21545 8635 21563 8653
rect 21581 8650 21602 8653
rect 21581 8635 21696 8650
rect 21545 8612 21696 8635
rect 25909 8666 25966 8685
rect 30289 8779 30309 8797
rect 30327 8779 30445 8797
rect 30289 8775 30445 8779
rect 30289 8759 30350 8775
rect 30622 8771 30664 8807
rect 34657 8868 34808 8891
rect 34766 8832 34808 8868
rect 34709 8831 34809 8832
rect 34653 8810 34809 8831
rect 30622 8748 30773 8771
rect 30622 8733 30737 8748
rect 30716 8730 30737 8733
rect 30755 8730 30773 8748
rect 30716 8711 30773 8730
rect 25909 8648 25927 8666
rect 25945 8663 25966 8666
rect 25945 8648 26060 8663
rect 25909 8625 26060 8648
rect 30286 8678 30343 8697
rect 34653 8792 34673 8810
rect 34691 8792 34809 8810
rect 34653 8788 34809 8792
rect 34653 8772 34714 8788
rect 30286 8660 30304 8678
rect 30322 8675 30343 8678
rect 30322 8660 30437 8675
rect 30286 8637 30437 8660
rect 34650 8691 34707 8710
rect 34650 8673 34668 8691
rect 34686 8688 34707 8691
rect 34686 8673 34801 8688
rect 34650 8650 34801 8673
rect 17331 8601 17431 8602
rect 17275 8580 17431 8601
rect 17275 8562 17295 8580
rect 17313 8562 17431 8580
rect 17275 8558 17431 8562
rect 13245 8511 13401 8515
rect 12909 8483 12966 8502
rect 8882 8399 9033 8422
rect 8584 8393 8684 8394
rect 8528 8372 8684 8393
rect 8882 8384 8997 8399
rect 8528 8354 8548 8372
rect 8566 8354 8684 8372
rect 8976 8381 8997 8384
rect 9015 8381 9033 8399
rect 12909 8465 12927 8483
rect 12945 8480 12966 8483
rect 13245 8493 13363 8511
rect 13381 8493 13401 8511
rect 12945 8465 13060 8480
rect 13245 8472 13401 8493
rect 13245 8471 13345 8472
rect 12909 8442 13060 8465
rect 8976 8362 9033 8381
rect 8528 8350 8684 8354
rect 4498 8303 4654 8307
rect 4498 8285 4616 8303
rect 4634 8285 4654 8303
rect 4498 8264 4654 8285
rect 4498 8263 4598 8264
rect 135 8191 286 8214
rect 135 8176 250 8191
rect 229 8173 250 8176
rect 268 8173 286 8191
rect 229 8154 286 8173
rect 4499 8227 4541 8263
rect 8528 8334 8589 8350
rect 8970 8319 9031 8335
rect 13018 8406 13060 8442
rect 13246 8435 13288 8471
rect 17275 8542 17336 8558
rect 17273 8496 17330 8515
rect 13246 8412 13397 8435
rect 12961 8405 13061 8406
rect 12905 8384 13061 8405
rect 13246 8397 13361 8412
rect 12905 8366 12925 8384
rect 12943 8366 13061 8384
rect 13340 8394 13361 8397
rect 13379 8394 13397 8412
rect 17273 8478 17291 8496
rect 17309 8493 17330 8496
rect 17309 8478 17424 8493
rect 17606 8489 17667 8505
rect 21654 8576 21696 8612
rect 21597 8575 21697 8576
rect 21541 8554 21697 8575
rect 21541 8536 21561 8554
rect 21579 8536 21697 8554
rect 21541 8532 21697 8536
rect 17273 8455 17424 8478
rect 13340 8375 13397 8394
rect 12905 8362 13061 8366
rect 8875 8315 9031 8319
rect 8875 8297 8993 8315
rect 9011 8297 9031 8315
rect 8875 8276 9031 8297
rect 8875 8275 8975 8276
rect 4499 8204 4650 8227
rect 4499 8189 4614 8204
rect 4593 8186 4614 8189
rect 4632 8186 4650 8204
rect 222 8076 283 8092
rect 127 8072 283 8076
rect 127 8054 245 8072
rect 263 8054 283 8072
rect 4593 8167 4650 8186
rect 8876 8239 8918 8275
rect 12905 8346 12966 8362
rect 13334 8332 13395 8348
rect 17382 8419 17424 8455
rect 17511 8485 17667 8489
rect 17511 8467 17629 8485
rect 17647 8467 17667 8485
rect 17511 8446 17667 8467
rect 17511 8445 17611 8446
rect 17325 8418 17425 8419
rect 17269 8397 17425 8418
rect 17269 8379 17289 8397
rect 17307 8379 17425 8397
rect 17269 8375 17425 8379
rect 17512 8409 17554 8445
rect 21541 8516 21602 8532
rect 21970 8502 22031 8518
rect 26018 8589 26060 8625
rect 25961 8588 26061 8589
rect 25905 8567 26061 8588
rect 25905 8549 25925 8567
rect 25943 8549 26061 8567
rect 25905 8545 26061 8549
rect 21875 8498 22031 8502
rect 21539 8470 21596 8489
rect 17512 8386 17663 8409
rect 13239 8328 13395 8332
rect 13239 8310 13357 8328
rect 13375 8310 13395 8328
rect 13239 8289 13395 8310
rect 13239 8288 13339 8289
rect 8876 8216 9027 8239
rect 8876 8201 8991 8216
rect 4163 8134 4220 8153
rect 4163 8116 4181 8134
rect 4199 8131 4220 8134
rect 4199 8116 4314 8131
rect 127 8033 283 8054
rect 127 8032 227 8033
rect 128 7996 170 8032
rect 128 7973 279 7996
rect 4163 8093 4314 8116
rect 4272 8057 4314 8093
rect 4586 8089 4647 8105
rect 4491 8085 4647 8089
rect 4491 8067 4609 8085
rect 4627 8067 4647 8085
rect 8970 8198 8991 8201
rect 9009 8198 9027 8216
rect 8970 8179 9027 8198
rect 13240 8252 13282 8288
rect 17269 8359 17330 8375
rect 17512 8371 17627 8386
rect 17606 8368 17627 8371
rect 17645 8368 17663 8386
rect 21539 8452 21557 8470
rect 21575 8467 21596 8470
rect 21875 8480 21993 8498
rect 22011 8480 22031 8498
rect 21575 8452 21690 8467
rect 21875 8459 22031 8480
rect 21875 8458 21975 8459
rect 21539 8429 21690 8452
rect 17606 8349 17663 8368
rect 17600 8306 17661 8322
rect 21648 8393 21690 8429
rect 21876 8422 21918 8458
rect 25905 8529 25966 8545
rect 26347 8514 26408 8530
rect 30395 8601 30437 8637
rect 30338 8600 30438 8601
rect 30282 8579 30438 8600
rect 30282 8561 30302 8579
rect 30320 8561 30438 8579
rect 30282 8557 30438 8561
rect 26252 8510 26408 8514
rect 25903 8483 25960 8502
rect 21876 8399 22027 8422
rect 21591 8392 21691 8393
rect 21535 8371 21691 8392
rect 21876 8384 21991 8399
rect 21535 8353 21555 8371
rect 21573 8353 21691 8371
rect 21970 8381 21991 8384
rect 22009 8381 22027 8399
rect 25903 8465 25921 8483
rect 25939 8480 25960 8483
rect 26252 8492 26370 8510
rect 26388 8492 26408 8510
rect 25939 8465 26054 8480
rect 26252 8471 26408 8492
rect 26252 8470 26352 8471
rect 25903 8442 26054 8465
rect 21970 8362 22027 8381
rect 21535 8349 21691 8353
rect 17505 8302 17661 8306
rect 17505 8284 17623 8302
rect 17641 8284 17661 8302
rect 13240 8229 13391 8252
rect 13240 8214 13355 8229
rect 13334 8211 13355 8214
rect 13373 8211 13391 8229
rect 8527 8147 8584 8166
rect 8527 8129 8545 8147
rect 8563 8144 8584 8147
rect 8563 8129 8678 8144
rect 4215 8056 4315 8057
rect 4159 8035 4315 8056
rect 4491 8046 4647 8067
rect 4491 8045 4591 8046
rect 4159 8017 4179 8035
rect 4197 8017 4315 8035
rect 4159 8013 4315 8017
rect 4159 7997 4220 8013
rect 4492 8009 4534 8045
rect 128 7958 243 7973
rect 222 7955 243 7958
rect 261 7955 279 7973
rect 222 7936 279 7955
rect 4492 7986 4643 8009
rect 8527 8106 8678 8129
rect 8636 8070 8678 8106
rect 8963 8101 9024 8117
rect 8868 8097 9024 8101
rect 8868 8079 8986 8097
rect 9004 8079 9024 8097
rect 13334 8192 13391 8211
rect 17505 8263 17661 8284
rect 17505 8262 17605 8263
rect 17506 8226 17548 8262
rect 21535 8333 21596 8349
rect 21964 8319 22025 8335
rect 26012 8406 26054 8442
rect 26253 8434 26295 8470
rect 30282 8541 30343 8557
rect 30711 8527 30772 8543
rect 34759 8614 34801 8650
rect 34702 8613 34802 8614
rect 34646 8592 34802 8613
rect 34646 8574 34666 8592
rect 34684 8574 34802 8592
rect 34646 8570 34802 8574
rect 30616 8523 30772 8527
rect 30280 8495 30337 8514
rect 26253 8411 26404 8434
rect 25955 8405 26055 8406
rect 25899 8384 26055 8405
rect 26253 8396 26368 8411
rect 25899 8366 25919 8384
rect 25937 8366 26055 8384
rect 26347 8393 26368 8396
rect 26386 8393 26404 8411
rect 30280 8477 30298 8495
rect 30316 8492 30337 8495
rect 30616 8505 30734 8523
rect 30752 8505 30772 8523
rect 30316 8477 30431 8492
rect 30616 8484 30772 8505
rect 30616 8483 30716 8484
rect 30280 8454 30431 8477
rect 26347 8374 26404 8393
rect 25899 8362 26055 8366
rect 21869 8315 22025 8319
rect 21869 8297 21987 8315
rect 22005 8297 22025 8315
rect 21869 8276 22025 8297
rect 21869 8275 21969 8276
rect 12904 8159 12961 8178
rect 12904 8141 12922 8159
rect 12940 8156 12961 8159
rect 12940 8141 13055 8156
rect 8579 8069 8679 8070
rect 8523 8048 8679 8069
rect 8868 8058 9024 8079
rect 8868 8057 8968 8058
rect 8523 8030 8543 8048
rect 8561 8030 8679 8048
rect 8523 8026 8679 8030
rect 8523 8010 8584 8026
rect 8869 8021 8911 8057
rect 4492 7971 4607 7986
rect 4586 7968 4607 7971
rect 4625 7968 4643 7986
rect 4586 7949 4643 7968
rect 8869 7998 9020 8021
rect 12904 8118 13055 8141
rect 13013 8082 13055 8118
rect 13327 8114 13388 8130
rect 13232 8110 13388 8114
rect 13232 8092 13350 8110
rect 13368 8092 13388 8110
rect 17506 8203 17657 8226
rect 17268 8172 17325 8191
rect 17506 8188 17621 8203
rect 17268 8154 17286 8172
rect 17304 8169 17325 8172
rect 17600 8185 17621 8188
rect 17639 8185 17657 8203
rect 17304 8154 17419 8169
rect 17600 8166 17657 8185
rect 21870 8239 21912 8275
rect 25899 8346 25960 8362
rect 26341 8331 26402 8347
rect 30389 8418 30431 8454
rect 30617 8447 30659 8483
rect 34646 8554 34707 8570
rect 34644 8508 34701 8527
rect 30617 8424 30768 8447
rect 30332 8417 30432 8418
rect 30276 8396 30432 8417
rect 30617 8409 30732 8424
rect 30276 8378 30296 8396
rect 30314 8378 30432 8396
rect 30711 8406 30732 8409
rect 30750 8406 30768 8424
rect 34644 8490 34662 8508
rect 34680 8505 34701 8508
rect 34680 8490 34795 8505
rect 34644 8467 34795 8490
rect 30711 8387 30768 8406
rect 30276 8374 30432 8378
rect 26246 8327 26402 8331
rect 26246 8309 26364 8327
rect 26382 8309 26402 8327
rect 26246 8288 26402 8309
rect 26246 8287 26346 8288
rect 21870 8216 22021 8239
rect 21870 8201 21985 8216
rect 21964 8198 21985 8201
rect 22003 8198 22021 8216
rect 12956 8081 13056 8082
rect 12900 8060 13056 8081
rect 13232 8071 13388 8092
rect 13232 8070 13332 8071
rect 12900 8042 12920 8060
rect 12938 8042 13056 8060
rect 12900 8038 13056 8042
rect 12900 8022 12961 8038
rect 13233 8034 13275 8070
rect 8869 7983 8984 7998
rect 8963 7980 8984 7983
rect 9002 7980 9020 7998
rect 8963 7961 9020 7980
rect 13233 8011 13384 8034
rect 17268 8131 17419 8154
rect 17377 8095 17419 8131
rect 17320 8094 17420 8095
rect 17264 8073 17420 8094
rect 17593 8088 17654 8104
rect 17264 8055 17284 8073
rect 17302 8055 17420 8073
rect 17264 8051 17420 8055
rect 17498 8084 17654 8088
rect 17498 8066 17616 8084
rect 17634 8066 17654 8084
rect 21964 8179 22021 8198
rect 26247 8251 26289 8287
rect 30276 8358 30337 8374
rect 30705 8344 30766 8360
rect 34753 8431 34795 8467
rect 34696 8430 34796 8431
rect 34640 8409 34796 8430
rect 34640 8391 34660 8409
rect 34678 8391 34796 8409
rect 34640 8387 34796 8391
rect 30610 8340 30766 8344
rect 30610 8322 30728 8340
rect 30746 8322 30766 8340
rect 30610 8301 30766 8322
rect 30610 8300 30710 8301
rect 26247 8228 26398 8251
rect 26247 8213 26362 8228
rect 21534 8146 21591 8165
rect 21534 8128 21552 8146
rect 21570 8143 21591 8146
rect 21570 8128 21685 8143
rect 17264 8035 17325 8051
rect 17498 8045 17654 8066
rect 17498 8044 17598 8045
rect 13233 7996 13348 8011
rect 13327 7993 13348 7996
rect 13366 7993 13384 8011
rect 13327 7974 13384 7993
rect 17499 8008 17541 8044
rect 17499 7985 17650 8008
rect 21534 8105 21685 8128
rect 21643 8069 21685 8105
rect 21957 8101 22018 8117
rect 21862 8097 22018 8101
rect 21862 8079 21980 8097
rect 21998 8079 22018 8097
rect 26341 8210 26362 8213
rect 26380 8210 26398 8228
rect 26341 8191 26398 8210
rect 30611 8264 30653 8300
rect 34640 8371 34701 8387
rect 30611 8241 30762 8264
rect 30611 8226 30726 8241
rect 30705 8223 30726 8226
rect 30744 8223 30762 8241
rect 25898 8159 25955 8178
rect 25898 8141 25916 8159
rect 25934 8156 25955 8159
rect 25934 8141 26049 8156
rect 21586 8068 21686 8069
rect 21530 8047 21686 8068
rect 21862 8058 22018 8079
rect 21862 8057 21962 8058
rect 21530 8029 21550 8047
rect 21568 8029 21686 8047
rect 21530 8025 21686 8029
rect 21530 8009 21591 8025
rect 21863 8021 21905 8057
rect 17499 7970 17614 7985
rect 17593 7967 17614 7970
rect 17632 7967 17650 7985
rect 17593 7948 17650 7967
rect 21863 7998 22014 8021
rect 25898 8118 26049 8141
rect 26007 8082 26049 8118
rect 26334 8113 26395 8129
rect 26239 8109 26395 8113
rect 26239 8091 26357 8109
rect 26375 8091 26395 8109
rect 30705 8204 30762 8223
rect 30275 8171 30332 8190
rect 30275 8153 30293 8171
rect 30311 8168 30332 8171
rect 30311 8153 30426 8168
rect 25950 8081 26050 8082
rect 25894 8060 26050 8081
rect 26239 8070 26395 8091
rect 26239 8069 26339 8070
rect 25894 8042 25914 8060
rect 25932 8042 26050 8060
rect 25894 8038 26050 8042
rect 25894 8022 25955 8038
rect 26240 8033 26282 8069
rect 21863 7983 21978 7998
rect 21957 7980 21978 7983
rect 21996 7980 22014 7998
rect 21957 7961 22014 7980
rect 26240 8010 26391 8033
rect 30275 8130 30426 8153
rect 30384 8094 30426 8130
rect 30698 8126 30759 8142
rect 30603 8122 30759 8126
rect 30603 8104 30721 8122
rect 30739 8104 30759 8122
rect 34639 8184 34696 8203
rect 34639 8166 34657 8184
rect 34675 8181 34696 8184
rect 34675 8166 34790 8181
rect 30327 8093 30427 8094
rect 30271 8072 30427 8093
rect 30603 8083 30759 8104
rect 30603 8082 30703 8083
rect 30271 8054 30291 8072
rect 30309 8054 30427 8072
rect 30271 8050 30427 8054
rect 30271 8034 30332 8050
rect 30604 8046 30646 8082
rect 26240 7995 26355 8010
rect 26334 7992 26355 7995
rect 26373 7992 26391 8010
rect 26334 7973 26391 7992
rect 30604 8023 30755 8046
rect 34639 8143 34790 8166
rect 34748 8107 34790 8143
rect 34691 8106 34791 8107
rect 34635 8085 34791 8106
rect 34635 8067 34655 8085
rect 34673 8067 34791 8085
rect 34635 8063 34791 8067
rect 34635 8047 34696 8063
rect 30604 8008 30719 8023
rect 30698 8005 30719 8008
rect 30737 8005 30755 8023
rect 30698 7986 30755 8005
rect 4164 7841 4221 7860
rect 4164 7823 4182 7841
rect 4200 7838 4221 7841
rect 4200 7823 4315 7838
rect 223 7783 284 7799
rect 128 7779 284 7783
rect 128 7761 246 7779
rect 264 7761 284 7779
rect 128 7740 284 7761
rect 128 7739 228 7740
rect 129 7703 171 7739
rect 129 7680 280 7703
rect 4164 7800 4315 7823
rect 8528 7854 8585 7873
rect 8528 7836 8546 7854
rect 8564 7851 8585 7854
rect 8564 7836 8679 7851
rect 4273 7764 4315 7800
rect 4587 7796 4648 7812
rect 4492 7792 4648 7796
rect 4492 7774 4610 7792
rect 4628 7774 4648 7792
rect 4216 7763 4316 7764
rect 4160 7742 4316 7763
rect 4492 7753 4648 7774
rect 4492 7752 4592 7753
rect 129 7665 244 7680
rect 223 7662 244 7665
rect 262 7662 280 7680
rect 223 7643 280 7662
rect 4160 7724 4180 7742
rect 4198 7724 4316 7742
rect 4160 7720 4316 7724
rect 4160 7704 4221 7720
rect 4493 7716 4535 7752
rect 4493 7693 4644 7716
rect 8528 7813 8679 7836
rect 12905 7866 12962 7885
rect 12905 7848 12923 7866
rect 12941 7863 12962 7866
rect 12941 7848 13056 7863
rect 8637 7777 8679 7813
rect 8964 7808 9025 7824
rect 8869 7804 9025 7808
rect 8869 7786 8987 7804
rect 9005 7786 9025 7804
rect 8580 7776 8680 7777
rect 8524 7755 8680 7776
rect 8869 7765 9025 7786
rect 8869 7764 8969 7765
rect 4493 7678 4608 7693
rect 4587 7675 4608 7678
rect 4626 7675 4644 7693
rect 4587 7656 4644 7675
rect 4157 7623 4214 7642
rect 8524 7737 8544 7755
rect 8562 7737 8680 7755
rect 8524 7733 8680 7737
rect 8524 7717 8585 7733
rect 8870 7728 8912 7764
rect 8870 7705 9021 7728
rect 12905 7825 13056 7848
rect 17269 7879 17326 7898
rect 17269 7861 17287 7879
rect 17305 7876 17326 7879
rect 17305 7861 17420 7876
rect 13014 7789 13056 7825
rect 13328 7821 13389 7837
rect 13233 7817 13389 7821
rect 13233 7799 13351 7817
rect 13369 7799 13389 7817
rect 12957 7788 13057 7789
rect 12901 7767 13057 7788
rect 13233 7778 13389 7799
rect 13233 7777 13333 7778
rect 8870 7690 8985 7705
rect 8964 7687 8985 7690
rect 9003 7687 9021 7705
rect 8964 7668 9021 7687
rect 4157 7605 4175 7623
rect 4193 7620 4214 7623
rect 4193 7605 4308 7620
rect 4157 7582 4308 7605
rect 218 7459 279 7475
rect 4266 7546 4308 7582
rect 8521 7636 8578 7655
rect 8521 7618 8539 7636
rect 8557 7633 8578 7636
rect 12901 7749 12921 7767
rect 12939 7749 13057 7767
rect 12901 7745 13057 7749
rect 12901 7729 12962 7745
rect 13234 7741 13276 7777
rect 13234 7718 13385 7741
rect 17269 7838 17420 7861
rect 17378 7802 17420 7838
rect 21535 7853 21592 7872
rect 21535 7835 21553 7853
rect 21571 7850 21592 7853
rect 21571 7835 21686 7850
rect 17321 7801 17421 7802
rect 17265 7780 17421 7801
rect 17594 7795 17655 7811
rect 13234 7703 13349 7718
rect 13328 7700 13349 7703
rect 13367 7700 13385 7718
rect 13328 7681 13385 7700
rect 8557 7618 8672 7633
rect 8521 7595 8672 7618
rect 4209 7545 4309 7546
rect 4153 7524 4309 7545
rect 4153 7506 4173 7524
rect 4191 7506 4309 7524
rect 4153 7502 4309 7506
rect 123 7455 279 7459
rect 123 7437 241 7455
rect 259 7437 279 7455
rect 123 7416 279 7437
rect 123 7415 223 7416
rect 124 7379 166 7415
rect 4153 7486 4214 7502
rect 4582 7472 4643 7488
rect 8630 7559 8672 7595
rect 12898 7648 12955 7667
rect 17265 7762 17285 7780
rect 17303 7762 17421 7780
rect 17265 7758 17421 7762
rect 17499 7791 17655 7795
rect 17499 7773 17617 7791
rect 17635 7773 17655 7791
rect 17265 7742 17326 7758
rect 17499 7752 17655 7773
rect 17499 7751 17599 7752
rect 17500 7715 17542 7751
rect 17500 7692 17651 7715
rect 21535 7812 21686 7835
rect 25899 7866 25956 7885
rect 25899 7848 25917 7866
rect 25935 7863 25956 7866
rect 25935 7848 26050 7863
rect 21644 7776 21686 7812
rect 21958 7808 22019 7824
rect 21863 7804 22019 7808
rect 21863 7786 21981 7804
rect 21999 7786 22019 7804
rect 21587 7775 21687 7776
rect 21531 7754 21687 7775
rect 21863 7765 22019 7786
rect 21863 7764 21963 7765
rect 12898 7630 12916 7648
rect 12934 7645 12955 7648
rect 12934 7630 13049 7645
rect 12898 7607 13049 7630
rect 8573 7558 8673 7559
rect 8517 7537 8673 7558
rect 8517 7519 8537 7537
rect 8555 7519 8673 7537
rect 8517 7515 8673 7519
rect 4487 7468 4643 7472
rect 4151 7440 4208 7459
rect 124 7356 275 7379
rect 124 7341 239 7356
rect 218 7338 239 7341
rect 257 7338 275 7356
rect 4151 7422 4169 7440
rect 4187 7437 4208 7440
rect 4487 7450 4605 7468
rect 4623 7450 4643 7468
rect 4187 7422 4302 7437
rect 4487 7429 4643 7450
rect 4487 7428 4587 7429
rect 4151 7399 4302 7422
rect 218 7319 275 7338
rect 212 7276 273 7292
rect 4260 7363 4302 7399
rect 4488 7392 4530 7428
rect 8517 7499 8578 7515
rect 8959 7484 9020 7500
rect 13007 7571 13049 7607
rect 17262 7661 17319 7680
rect 17500 7677 17615 7692
rect 17262 7643 17280 7661
rect 17298 7658 17319 7661
rect 17594 7674 17615 7677
rect 17633 7674 17651 7692
rect 17298 7643 17413 7658
rect 17594 7655 17651 7674
rect 17262 7620 17413 7643
rect 21531 7736 21551 7754
rect 21569 7736 21687 7754
rect 21531 7732 21687 7736
rect 21531 7716 21592 7732
rect 21864 7728 21906 7764
rect 21864 7705 22015 7728
rect 25899 7825 26050 7848
rect 30276 7878 30333 7897
rect 30276 7860 30294 7878
rect 30312 7875 30333 7878
rect 30312 7860 30427 7875
rect 26008 7789 26050 7825
rect 26335 7820 26396 7836
rect 26240 7816 26396 7820
rect 26240 7798 26358 7816
rect 26376 7798 26396 7816
rect 25951 7788 26051 7789
rect 25895 7767 26051 7788
rect 26240 7777 26396 7798
rect 26240 7776 26340 7777
rect 21864 7690 21979 7705
rect 21958 7687 21979 7690
rect 21997 7687 22015 7705
rect 21958 7668 22015 7687
rect 12950 7570 13050 7571
rect 12894 7549 13050 7570
rect 12894 7531 12914 7549
rect 12932 7531 13050 7549
rect 12894 7527 13050 7531
rect 8864 7480 9020 7484
rect 8515 7453 8572 7472
rect 4488 7369 4639 7392
rect 4203 7362 4303 7363
rect 4147 7341 4303 7362
rect 4488 7354 4603 7369
rect 4147 7323 4167 7341
rect 4185 7323 4303 7341
rect 4582 7351 4603 7354
rect 4621 7351 4639 7369
rect 8515 7435 8533 7453
rect 8551 7450 8572 7453
rect 8864 7462 8982 7480
rect 9000 7462 9020 7480
rect 8551 7435 8666 7450
rect 8864 7441 9020 7462
rect 8864 7440 8964 7441
rect 8515 7412 8666 7435
rect 4582 7332 4639 7351
rect 4147 7319 4303 7323
rect 117 7272 273 7276
rect 117 7254 235 7272
rect 253 7254 273 7272
rect 117 7233 273 7254
rect 117 7232 217 7233
rect 118 7196 160 7232
rect 4147 7303 4208 7319
rect 4576 7289 4637 7305
rect 8624 7376 8666 7412
rect 8865 7404 8907 7440
rect 12894 7511 12955 7527
rect 13323 7497 13384 7513
rect 17371 7584 17413 7620
rect 17314 7583 17414 7584
rect 17258 7562 17414 7583
rect 21528 7635 21585 7654
rect 25895 7749 25915 7767
rect 25933 7749 26051 7767
rect 25895 7745 26051 7749
rect 25895 7729 25956 7745
rect 26241 7740 26283 7776
rect 26241 7717 26392 7740
rect 30276 7837 30427 7860
rect 34640 7891 34697 7910
rect 34640 7873 34658 7891
rect 34676 7888 34697 7891
rect 34676 7873 34791 7888
rect 30385 7801 30427 7837
rect 30699 7833 30760 7849
rect 30604 7829 30760 7833
rect 30604 7811 30722 7829
rect 30740 7811 30760 7829
rect 30328 7800 30428 7801
rect 30272 7779 30428 7800
rect 30604 7790 30760 7811
rect 30604 7789 30704 7790
rect 26241 7702 26356 7717
rect 26335 7699 26356 7702
rect 26374 7699 26392 7717
rect 26335 7680 26392 7699
rect 21528 7617 21546 7635
rect 21564 7632 21585 7635
rect 21564 7617 21679 7632
rect 21528 7594 21679 7617
rect 17258 7544 17278 7562
rect 17296 7544 17414 7562
rect 17258 7540 17414 7544
rect 13228 7493 13384 7497
rect 12892 7465 12949 7484
rect 8865 7381 9016 7404
rect 8567 7375 8667 7376
rect 8511 7354 8667 7375
rect 8865 7366 8980 7381
rect 8511 7336 8531 7354
rect 8549 7336 8667 7354
rect 8959 7363 8980 7366
rect 8998 7363 9016 7381
rect 12892 7447 12910 7465
rect 12928 7462 12949 7465
rect 13228 7475 13346 7493
rect 13364 7475 13384 7493
rect 12928 7447 13043 7462
rect 13228 7454 13384 7475
rect 13228 7453 13328 7454
rect 12892 7424 13043 7447
rect 8959 7344 9016 7363
rect 8511 7332 8667 7336
rect 4481 7285 4637 7289
rect 4481 7267 4599 7285
rect 4617 7267 4637 7285
rect 4481 7246 4637 7267
rect 4481 7245 4581 7246
rect 118 7173 269 7196
rect 118 7158 233 7173
rect 212 7155 233 7158
rect 251 7155 269 7173
rect 212 7136 269 7155
rect 4482 7209 4524 7245
rect 8511 7316 8572 7332
rect 8953 7301 9014 7317
rect 13001 7388 13043 7424
rect 13229 7417 13271 7453
rect 17258 7524 17319 7540
rect 17256 7478 17313 7497
rect 13229 7394 13380 7417
rect 12944 7387 13044 7388
rect 12888 7366 13044 7387
rect 13229 7379 13344 7394
rect 12888 7348 12908 7366
rect 12926 7348 13044 7366
rect 13323 7376 13344 7379
rect 13362 7376 13380 7394
rect 17256 7460 17274 7478
rect 17292 7475 17313 7478
rect 17292 7460 17407 7475
rect 17589 7471 17650 7487
rect 21637 7558 21679 7594
rect 25892 7648 25949 7667
rect 25892 7630 25910 7648
rect 25928 7645 25949 7648
rect 30272 7761 30292 7779
rect 30310 7761 30428 7779
rect 30272 7757 30428 7761
rect 30272 7741 30333 7757
rect 30605 7753 30647 7789
rect 30605 7730 30756 7753
rect 34640 7850 34791 7873
rect 34749 7814 34791 7850
rect 34692 7813 34792 7814
rect 34636 7792 34792 7813
rect 30605 7715 30720 7730
rect 30699 7712 30720 7715
rect 30738 7712 30756 7730
rect 30699 7693 30756 7712
rect 25928 7630 26043 7645
rect 25892 7607 26043 7630
rect 21580 7557 21680 7558
rect 21524 7536 21680 7557
rect 21524 7518 21544 7536
rect 21562 7518 21680 7536
rect 21524 7514 21680 7518
rect 17256 7437 17407 7460
rect 13323 7357 13380 7376
rect 12888 7344 13044 7348
rect 8858 7297 9014 7301
rect 8858 7279 8976 7297
rect 8994 7279 9014 7297
rect 8858 7258 9014 7279
rect 8858 7257 8958 7258
rect 4482 7186 4633 7209
rect 4482 7171 4597 7186
rect 205 7058 266 7074
rect 110 7054 266 7058
rect 110 7036 228 7054
rect 246 7036 266 7054
rect 4576 7168 4597 7171
rect 4615 7168 4633 7186
rect 4576 7149 4633 7168
rect 8859 7221 8901 7257
rect 12888 7328 12949 7344
rect 13317 7314 13378 7330
rect 17365 7401 17407 7437
rect 17494 7467 17650 7471
rect 17494 7449 17612 7467
rect 17630 7449 17650 7467
rect 17494 7428 17650 7449
rect 17494 7427 17594 7428
rect 17308 7400 17408 7401
rect 17252 7379 17408 7400
rect 17252 7361 17272 7379
rect 17290 7361 17408 7379
rect 17252 7357 17408 7361
rect 17495 7391 17537 7427
rect 21524 7498 21585 7514
rect 21953 7484 22014 7500
rect 26001 7571 26043 7607
rect 30269 7660 30326 7679
rect 34636 7774 34656 7792
rect 34674 7774 34792 7792
rect 34636 7770 34792 7774
rect 34636 7754 34697 7770
rect 30269 7642 30287 7660
rect 30305 7657 30326 7660
rect 30305 7642 30420 7657
rect 30269 7619 30420 7642
rect 25944 7570 26044 7571
rect 25888 7549 26044 7570
rect 25888 7531 25908 7549
rect 25926 7531 26044 7549
rect 25888 7527 26044 7531
rect 21858 7480 22014 7484
rect 21522 7452 21579 7471
rect 17495 7368 17646 7391
rect 13222 7310 13378 7314
rect 13222 7292 13340 7310
rect 13358 7292 13378 7310
rect 13222 7271 13378 7292
rect 13222 7270 13322 7271
rect 8859 7198 9010 7221
rect 8859 7183 8974 7198
rect 4146 7116 4203 7135
rect 4146 7098 4164 7116
rect 4182 7113 4203 7116
rect 4182 7098 4297 7113
rect 110 7015 266 7036
rect 110 7014 210 7015
rect 111 6978 153 7014
rect 111 6955 262 6978
rect 4146 7075 4297 7098
rect 4255 7039 4297 7075
rect 4569 7071 4630 7087
rect 4474 7067 4630 7071
rect 4474 7049 4592 7067
rect 4610 7049 4630 7067
rect 8953 7180 8974 7183
rect 8992 7180 9010 7198
rect 8953 7161 9010 7180
rect 13223 7234 13265 7270
rect 17252 7341 17313 7357
rect 17495 7353 17610 7368
rect 17589 7350 17610 7353
rect 17628 7350 17646 7368
rect 21522 7434 21540 7452
rect 21558 7449 21579 7452
rect 21858 7462 21976 7480
rect 21994 7462 22014 7480
rect 21558 7434 21673 7449
rect 21858 7441 22014 7462
rect 21858 7440 21958 7441
rect 21522 7411 21673 7434
rect 17589 7331 17646 7350
rect 17583 7288 17644 7304
rect 21631 7375 21673 7411
rect 21859 7404 21901 7440
rect 25888 7511 25949 7527
rect 26330 7496 26391 7512
rect 30378 7583 30420 7619
rect 34633 7673 34690 7692
rect 34633 7655 34651 7673
rect 34669 7670 34690 7673
rect 34669 7655 34784 7670
rect 34633 7632 34784 7655
rect 30321 7582 30421 7583
rect 30265 7561 30421 7582
rect 30265 7543 30285 7561
rect 30303 7543 30421 7561
rect 30265 7539 30421 7543
rect 26235 7492 26391 7496
rect 25886 7465 25943 7484
rect 21859 7381 22010 7404
rect 21574 7374 21674 7375
rect 21518 7353 21674 7374
rect 21859 7366 21974 7381
rect 21518 7335 21538 7353
rect 21556 7335 21674 7353
rect 21953 7363 21974 7366
rect 21992 7363 22010 7381
rect 25886 7447 25904 7465
rect 25922 7462 25943 7465
rect 26235 7474 26353 7492
rect 26371 7474 26391 7492
rect 25922 7447 26037 7462
rect 26235 7453 26391 7474
rect 26235 7452 26335 7453
rect 25886 7424 26037 7447
rect 21953 7344 22010 7363
rect 21518 7331 21674 7335
rect 17488 7284 17644 7288
rect 17488 7266 17606 7284
rect 17624 7266 17644 7284
rect 13223 7211 13374 7234
rect 13223 7196 13338 7211
rect 8510 7129 8567 7148
rect 8510 7111 8528 7129
rect 8546 7126 8567 7129
rect 8546 7111 8661 7126
rect 4198 7038 4298 7039
rect 4142 7017 4298 7038
rect 4474 7028 4630 7049
rect 4474 7027 4574 7028
rect 4142 6999 4162 7017
rect 4180 6999 4298 7017
rect 4142 6995 4298 6999
rect 4142 6979 4203 6995
rect 4475 6991 4517 7027
rect 111 6940 226 6955
rect 205 6937 226 6940
rect 244 6937 262 6955
rect 205 6918 262 6937
rect 4475 6968 4626 6991
rect 8510 7088 8661 7111
rect 8619 7052 8661 7088
rect 8946 7083 9007 7099
rect 8851 7079 9007 7083
rect 8851 7061 8969 7079
rect 8987 7061 9007 7079
rect 13317 7193 13338 7196
rect 13356 7193 13374 7211
rect 13317 7174 13374 7193
rect 17488 7245 17644 7266
rect 17488 7244 17588 7245
rect 17489 7208 17531 7244
rect 21518 7315 21579 7331
rect 21947 7301 22008 7317
rect 25995 7388 26037 7424
rect 26236 7416 26278 7452
rect 30265 7523 30326 7539
rect 30694 7509 30755 7525
rect 34742 7596 34784 7632
rect 34685 7595 34785 7596
rect 34629 7574 34785 7595
rect 34629 7556 34649 7574
rect 34667 7556 34785 7574
rect 34629 7552 34785 7556
rect 30599 7505 30755 7509
rect 30263 7477 30320 7496
rect 26236 7393 26387 7416
rect 25938 7387 26038 7388
rect 25882 7366 26038 7387
rect 26236 7378 26351 7393
rect 25882 7348 25902 7366
rect 25920 7348 26038 7366
rect 26330 7375 26351 7378
rect 26369 7375 26387 7393
rect 30263 7459 30281 7477
rect 30299 7474 30320 7477
rect 30599 7487 30717 7505
rect 30735 7487 30755 7505
rect 30299 7459 30414 7474
rect 30599 7466 30755 7487
rect 30599 7465 30699 7466
rect 30263 7436 30414 7459
rect 26330 7356 26387 7375
rect 25882 7344 26038 7348
rect 21852 7297 22008 7301
rect 21852 7279 21970 7297
rect 21988 7279 22008 7297
rect 21852 7258 22008 7279
rect 21852 7257 21952 7258
rect 12887 7141 12944 7160
rect 12887 7123 12905 7141
rect 12923 7138 12944 7141
rect 12923 7123 13038 7138
rect 8562 7051 8662 7052
rect 8506 7030 8662 7051
rect 8851 7040 9007 7061
rect 8851 7039 8951 7040
rect 8506 7012 8526 7030
rect 8544 7012 8662 7030
rect 8506 7008 8662 7012
rect 8506 6992 8567 7008
rect 8852 7003 8894 7039
rect 4475 6953 4590 6968
rect 4569 6950 4590 6953
rect 4608 6950 4626 6968
rect 4569 6931 4626 6950
rect 8852 6980 9003 7003
rect 12887 7100 13038 7123
rect 12996 7064 13038 7100
rect 13310 7096 13371 7112
rect 13215 7092 13371 7096
rect 13215 7074 13333 7092
rect 13351 7074 13371 7092
rect 17489 7185 17640 7208
rect 17251 7154 17308 7173
rect 17489 7170 17604 7185
rect 17251 7136 17269 7154
rect 17287 7151 17308 7154
rect 17583 7167 17604 7170
rect 17622 7167 17640 7185
rect 17287 7136 17402 7151
rect 17583 7148 17640 7167
rect 21853 7221 21895 7257
rect 25882 7328 25943 7344
rect 26324 7313 26385 7329
rect 30372 7400 30414 7436
rect 30600 7429 30642 7465
rect 34629 7536 34690 7552
rect 34627 7490 34684 7509
rect 30600 7406 30751 7429
rect 30315 7399 30415 7400
rect 30259 7378 30415 7399
rect 30600 7391 30715 7406
rect 30259 7360 30279 7378
rect 30297 7360 30415 7378
rect 30694 7388 30715 7391
rect 30733 7388 30751 7406
rect 34627 7472 34645 7490
rect 34663 7487 34684 7490
rect 34663 7472 34778 7487
rect 34627 7449 34778 7472
rect 30694 7369 30751 7388
rect 30259 7356 30415 7360
rect 26229 7309 26385 7313
rect 26229 7291 26347 7309
rect 26365 7291 26385 7309
rect 26229 7270 26385 7291
rect 26229 7269 26329 7270
rect 21853 7198 22004 7221
rect 21853 7183 21968 7198
rect 12939 7063 13039 7064
rect 12883 7042 13039 7063
rect 13215 7053 13371 7074
rect 13215 7052 13315 7053
rect 12883 7024 12903 7042
rect 12921 7024 13039 7042
rect 12883 7020 13039 7024
rect 12883 7004 12944 7020
rect 13216 7016 13258 7052
rect 8852 6965 8967 6980
rect 8946 6962 8967 6965
rect 8985 6962 9003 6980
rect 8946 6943 9003 6962
rect 13216 6993 13367 7016
rect 17251 7113 17402 7136
rect 17360 7077 17402 7113
rect 17303 7076 17403 7077
rect 17247 7055 17403 7076
rect 17576 7070 17637 7086
rect 17247 7037 17267 7055
rect 17285 7037 17403 7055
rect 17247 7033 17403 7037
rect 17481 7066 17637 7070
rect 17481 7048 17599 7066
rect 17617 7048 17637 7066
rect 21947 7180 21968 7183
rect 21986 7180 22004 7198
rect 21947 7161 22004 7180
rect 26230 7233 26272 7269
rect 30259 7340 30320 7356
rect 30688 7326 30749 7342
rect 34736 7413 34778 7449
rect 34679 7412 34779 7413
rect 34623 7391 34779 7412
rect 34623 7373 34643 7391
rect 34661 7373 34779 7391
rect 34623 7369 34779 7373
rect 30593 7322 30749 7326
rect 30593 7304 30711 7322
rect 30729 7304 30749 7322
rect 30593 7283 30749 7304
rect 30593 7282 30693 7283
rect 26230 7210 26381 7233
rect 26230 7195 26345 7210
rect 21517 7128 21574 7147
rect 21517 7110 21535 7128
rect 21553 7125 21574 7128
rect 21553 7110 21668 7125
rect 17247 7017 17308 7033
rect 17481 7027 17637 7048
rect 17481 7026 17581 7027
rect 13216 6978 13331 6993
rect 13310 6975 13331 6978
rect 13349 6975 13367 6993
rect 13310 6956 13367 6975
rect 17482 6990 17524 7026
rect 17482 6967 17633 6990
rect 21517 7087 21668 7110
rect 21626 7051 21668 7087
rect 21940 7083 22001 7099
rect 21845 7079 22001 7083
rect 21845 7061 21963 7079
rect 21981 7061 22001 7079
rect 26324 7192 26345 7195
rect 26363 7192 26381 7210
rect 26324 7173 26381 7192
rect 30594 7246 30636 7282
rect 34623 7353 34684 7369
rect 30594 7223 30745 7246
rect 30594 7208 30709 7223
rect 25881 7141 25938 7160
rect 25881 7123 25899 7141
rect 25917 7138 25938 7141
rect 25917 7123 26032 7138
rect 21569 7050 21669 7051
rect 21513 7029 21669 7050
rect 21845 7040 22001 7061
rect 21845 7039 21945 7040
rect 21513 7011 21533 7029
rect 21551 7011 21669 7029
rect 21513 7007 21669 7011
rect 21513 6991 21574 7007
rect 21846 7003 21888 7039
rect 17482 6952 17597 6967
rect 17576 6949 17597 6952
rect 17615 6949 17633 6967
rect 17576 6930 17633 6949
rect 21846 6980 21997 7003
rect 25881 7100 26032 7123
rect 25990 7064 26032 7100
rect 26317 7095 26378 7111
rect 26222 7091 26378 7095
rect 26222 7073 26340 7091
rect 26358 7073 26378 7091
rect 30688 7205 30709 7208
rect 30727 7205 30745 7223
rect 30688 7186 30745 7205
rect 30258 7153 30315 7172
rect 30258 7135 30276 7153
rect 30294 7150 30315 7153
rect 30294 7135 30409 7150
rect 25933 7063 26033 7064
rect 25877 7042 26033 7063
rect 26222 7052 26378 7073
rect 26222 7051 26322 7052
rect 25877 7024 25897 7042
rect 25915 7024 26033 7042
rect 25877 7020 26033 7024
rect 25877 7004 25938 7020
rect 26223 7015 26265 7051
rect 21846 6965 21961 6980
rect 21940 6962 21961 6965
rect 21979 6962 21997 6980
rect 21940 6943 21997 6962
rect 26223 6992 26374 7015
rect 30258 7112 30409 7135
rect 30367 7076 30409 7112
rect 30681 7108 30742 7124
rect 30586 7104 30742 7108
rect 30586 7086 30704 7104
rect 30722 7086 30742 7104
rect 34622 7166 34679 7185
rect 34622 7148 34640 7166
rect 34658 7163 34679 7166
rect 34658 7148 34773 7163
rect 30310 7075 30410 7076
rect 30254 7054 30410 7075
rect 30586 7065 30742 7086
rect 30586 7064 30686 7065
rect 30254 7036 30274 7054
rect 30292 7036 30410 7054
rect 30254 7032 30410 7036
rect 30254 7016 30315 7032
rect 30587 7028 30629 7064
rect 26223 6977 26338 6992
rect 26317 6974 26338 6977
rect 26356 6974 26374 6992
rect 26317 6955 26374 6974
rect 30587 7005 30738 7028
rect 34622 7125 34773 7148
rect 34731 7089 34773 7125
rect 34674 7088 34774 7089
rect 34618 7067 34774 7088
rect 34618 7049 34638 7067
rect 34656 7049 34774 7067
rect 34618 7045 34774 7049
rect 34618 7029 34679 7045
rect 30587 6990 30702 7005
rect 30681 6987 30702 6990
rect 30720 6987 30738 7005
rect 30681 6968 30738 6987
rect 4144 6823 4201 6842
rect 4144 6805 4162 6823
rect 4180 6820 4201 6823
rect 4180 6805 4295 6820
rect 203 6765 264 6781
rect 108 6761 264 6765
rect 108 6743 226 6761
rect 244 6743 264 6761
rect 108 6722 264 6743
rect 108 6721 208 6722
rect 109 6685 151 6721
rect 109 6662 260 6685
rect 4144 6782 4295 6805
rect 8508 6836 8565 6855
rect 8508 6818 8526 6836
rect 8544 6833 8565 6836
rect 8544 6818 8659 6833
rect 4253 6746 4295 6782
rect 4567 6778 4628 6794
rect 4472 6774 4628 6778
rect 4472 6756 4590 6774
rect 4608 6756 4628 6774
rect 4196 6745 4296 6746
rect 4140 6724 4296 6745
rect 4472 6735 4628 6756
rect 4472 6734 4572 6735
rect 109 6647 224 6662
rect 203 6644 224 6647
rect 242 6644 260 6662
rect 203 6625 260 6644
rect 4140 6706 4160 6724
rect 4178 6706 4296 6724
rect 4140 6702 4296 6706
rect 4140 6686 4201 6702
rect 4473 6698 4515 6734
rect 4473 6675 4624 6698
rect 8508 6795 8659 6818
rect 12885 6848 12942 6867
rect 12885 6830 12903 6848
rect 12921 6845 12942 6848
rect 12921 6830 13036 6845
rect 8617 6759 8659 6795
rect 8944 6790 9005 6806
rect 8849 6786 9005 6790
rect 8849 6768 8967 6786
rect 8985 6768 9005 6786
rect 8560 6758 8660 6759
rect 8504 6737 8660 6758
rect 8849 6747 9005 6768
rect 8849 6746 8949 6747
rect 4473 6660 4588 6675
rect 4567 6657 4588 6660
rect 4606 6657 4624 6675
rect 4567 6638 4624 6657
rect 4137 6605 4194 6624
rect 4137 6587 4155 6605
rect 4173 6602 4194 6605
rect 8504 6719 8524 6737
rect 8542 6719 8660 6737
rect 8504 6715 8660 6719
rect 8504 6699 8565 6715
rect 8850 6710 8892 6746
rect 8850 6687 9001 6710
rect 12885 6807 13036 6830
rect 17249 6861 17306 6880
rect 17249 6843 17267 6861
rect 17285 6858 17306 6861
rect 17285 6843 17400 6858
rect 12994 6771 13036 6807
rect 13308 6803 13369 6819
rect 13213 6799 13369 6803
rect 13213 6781 13331 6799
rect 13349 6781 13369 6799
rect 12937 6770 13037 6771
rect 12881 6749 13037 6770
rect 13213 6760 13369 6781
rect 13213 6759 13313 6760
rect 8850 6672 8965 6687
rect 8944 6669 8965 6672
rect 8983 6669 9001 6687
rect 8944 6650 9001 6669
rect 4173 6587 4288 6602
rect 4137 6564 4288 6587
rect 198 6441 259 6457
rect 4246 6528 4288 6564
rect 8501 6618 8558 6637
rect 8501 6600 8519 6618
rect 8537 6615 8558 6618
rect 12881 6731 12901 6749
rect 12919 6731 13037 6749
rect 12881 6727 13037 6731
rect 12881 6711 12942 6727
rect 13214 6723 13256 6759
rect 13214 6700 13365 6723
rect 17249 6820 17400 6843
rect 17358 6784 17400 6820
rect 21515 6835 21572 6854
rect 21515 6817 21533 6835
rect 21551 6832 21572 6835
rect 21551 6817 21666 6832
rect 17301 6783 17401 6784
rect 17245 6762 17401 6783
rect 17574 6777 17635 6793
rect 13214 6685 13329 6700
rect 13308 6682 13329 6685
rect 13347 6682 13365 6700
rect 13308 6663 13365 6682
rect 8537 6600 8652 6615
rect 8501 6577 8652 6600
rect 4189 6527 4289 6528
rect 4133 6506 4289 6527
rect 4133 6488 4153 6506
rect 4171 6488 4289 6506
rect 4133 6484 4289 6488
rect 103 6437 259 6441
rect 103 6419 221 6437
rect 239 6419 259 6437
rect 103 6398 259 6419
rect 103 6397 203 6398
rect 104 6361 146 6397
rect 4133 6468 4194 6484
rect 4562 6454 4623 6470
rect 8610 6541 8652 6577
rect 12878 6630 12935 6649
rect 12878 6612 12896 6630
rect 12914 6627 12935 6630
rect 17245 6744 17265 6762
rect 17283 6744 17401 6762
rect 17245 6740 17401 6744
rect 17479 6773 17635 6777
rect 17479 6755 17597 6773
rect 17615 6755 17635 6773
rect 17245 6724 17306 6740
rect 17479 6734 17635 6755
rect 17479 6733 17579 6734
rect 17480 6697 17522 6733
rect 17480 6674 17631 6697
rect 21515 6794 21666 6817
rect 25879 6848 25936 6867
rect 25879 6830 25897 6848
rect 25915 6845 25936 6848
rect 25915 6830 26030 6845
rect 21624 6758 21666 6794
rect 21938 6790 21999 6806
rect 21843 6786 21999 6790
rect 21843 6768 21961 6786
rect 21979 6768 21999 6786
rect 21567 6757 21667 6758
rect 21511 6736 21667 6757
rect 21843 6747 21999 6768
rect 21843 6746 21943 6747
rect 12914 6612 13029 6627
rect 12878 6589 13029 6612
rect 8553 6540 8653 6541
rect 8497 6519 8653 6540
rect 8497 6501 8517 6519
rect 8535 6501 8653 6519
rect 8497 6497 8653 6501
rect 4467 6450 4623 6454
rect 4131 6422 4188 6441
rect 104 6338 255 6361
rect 104 6323 219 6338
rect 198 6320 219 6323
rect 237 6320 255 6338
rect 4131 6404 4149 6422
rect 4167 6419 4188 6422
rect 4467 6432 4585 6450
rect 4603 6432 4623 6450
rect 4167 6404 4282 6419
rect 4467 6411 4623 6432
rect 4467 6410 4567 6411
rect 4131 6381 4282 6404
rect 198 6301 255 6320
rect 192 6258 253 6274
rect 4240 6345 4282 6381
rect 4468 6374 4510 6410
rect 8497 6481 8558 6497
rect 8939 6466 9000 6482
rect 12987 6553 13029 6589
rect 17242 6643 17299 6662
rect 17480 6659 17595 6674
rect 17242 6625 17260 6643
rect 17278 6640 17299 6643
rect 17574 6656 17595 6659
rect 17613 6656 17631 6674
rect 17278 6625 17393 6640
rect 17574 6637 17631 6656
rect 17242 6602 17393 6625
rect 21511 6718 21531 6736
rect 21549 6718 21667 6736
rect 21511 6714 21667 6718
rect 21511 6698 21572 6714
rect 21844 6710 21886 6746
rect 21844 6687 21995 6710
rect 25879 6807 26030 6830
rect 30256 6860 30313 6879
rect 30256 6842 30274 6860
rect 30292 6857 30313 6860
rect 30292 6842 30407 6857
rect 25988 6771 26030 6807
rect 26315 6802 26376 6818
rect 26220 6798 26376 6802
rect 26220 6780 26338 6798
rect 26356 6780 26376 6798
rect 25931 6770 26031 6771
rect 25875 6749 26031 6770
rect 26220 6759 26376 6780
rect 26220 6758 26320 6759
rect 21844 6672 21959 6687
rect 21938 6669 21959 6672
rect 21977 6669 21995 6687
rect 21938 6650 21995 6669
rect 12930 6552 13030 6553
rect 12874 6531 13030 6552
rect 12874 6513 12894 6531
rect 12912 6513 13030 6531
rect 12874 6509 13030 6513
rect 8844 6462 9000 6466
rect 8495 6435 8552 6454
rect 4468 6351 4619 6374
rect 4183 6344 4283 6345
rect 4127 6323 4283 6344
rect 4468 6336 4583 6351
rect 4127 6305 4147 6323
rect 4165 6305 4283 6323
rect 4562 6333 4583 6336
rect 4601 6333 4619 6351
rect 8495 6417 8513 6435
rect 8531 6432 8552 6435
rect 8844 6444 8962 6462
rect 8980 6444 9000 6462
rect 8531 6417 8646 6432
rect 8844 6423 9000 6444
rect 8844 6422 8944 6423
rect 8495 6394 8646 6417
rect 4562 6314 4619 6333
rect 4127 6301 4283 6305
rect 97 6254 253 6258
rect 97 6236 215 6254
rect 233 6236 253 6254
rect 97 6215 253 6236
rect 97 6214 197 6215
rect 98 6178 140 6214
rect 4127 6285 4188 6301
rect 4556 6271 4617 6287
rect 8604 6358 8646 6394
rect 8845 6386 8887 6422
rect 12874 6493 12935 6509
rect 13303 6479 13364 6495
rect 17351 6566 17393 6602
rect 17294 6565 17394 6566
rect 17238 6544 17394 6565
rect 21508 6617 21565 6636
rect 21508 6599 21526 6617
rect 21544 6614 21565 6617
rect 25875 6731 25895 6749
rect 25913 6731 26031 6749
rect 25875 6727 26031 6731
rect 25875 6711 25936 6727
rect 26221 6722 26263 6758
rect 26221 6699 26372 6722
rect 30256 6819 30407 6842
rect 34620 6873 34677 6892
rect 34620 6855 34638 6873
rect 34656 6870 34677 6873
rect 34656 6855 34771 6870
rect 30365 6783 30407 6819
rect 30679 6815 30740 6831
rect 30584 6811 30740 6815
rect 30584 6793 30702 6811
rect 30720 6793 30740 6811
rect 30308 6782 30408 6783
rect 30252 6761 30408 6782
rect 30584 6772 30740 6793
rect 30584 6771 30684 6772
rect 26221 6684 26336 6699
rect 26315 6681 26336 6684
rect 26354 6681 26372 6699
rect 26315 6662 26372 6681
rect 21544 6599 21659 6614
rect 21508 6576 21659 6599
rect 17238 6526 17258 6544
rect 17276 6526 17394 6544
rect 17238 6522 17394 6526
rect 13208 6475 13364 6479
rect 12872 6447 12929 6466
rect 8845 6363 8996 6386
rect 8547 6357 8647 6358
rect 8491 6336 8647 6357
rect 8845 6348 8960 6363
rect 8491 6318 8511 6336
rect 8529 6318 8647 6336
rect 8939 6345 8960 6348
rect 8978 6345 8996 6363
rect 12872 6429 12890 6447
rect 12908 6444 12929 6447
rect 13208 6457 13326 6475
rect 13344 6457 13364 6475
rect 12908 6429 13023 6444
rect 13208 6436 13364 6457
rect 13208 6435 13308 6436
rect 12872 6406 13023 6429
rect 8939 6326 8996 6345
rect 8491 6314 8647 6318
rect 4461 6267 4617 6271
rect 4461 6249 4579 6267
rect 4597 6249 4617 6267
rect 4461 6228 4617 6249
rect 4461 6227 4561 6228
rect 98 6155 249 6178
rect 98 6140 213 6155
rect 192 6137 213 6140
rect 231 6137 249 6155
rect 192 6118 249 6137
rect 4462 6191 4504 6227
rect 8491 6298 8552 6314
rect 8933 6283 8994 6299
rect 12981 6370 13023 6406
rect 13209 6399 13251 6435
rect 17238 6506 17299 6522
rect 17236 6460 17293 6479
rect 13209 6376 13360 6399
rect 12924 6369 13024 6370
rect 12868 6348 13024 6369
rect 13209 6361 13324 6376
rect 12868 6330 12888 6348
rect 12906 6330 13024 6348
rect 13303 6358 13324 6361
rect 13342 6358 13360 6376
rect 17236 6442 17254 6460
rect 17272 6457 17293 6460
rect 17272 6442 17387 6457
rect 17569 6453 17630 6469
rect 21617 6540 21659 6576
rect 25872 6630 25929 6649
rect 25872 6612 25890 6630
rect 25908 6627 25929 6630
rect 30252 6743 30272 6761
rect 30290 6743 30408 6761
rect 30252 6739 30408 6743
rect 30252 6723 30313 6739
rect 30585 6735 30627 6771
rect 30585 6712 30736 6735
rect 34620 6832 34771 6855
rect 34729 6796 34771 6832
rect 34672 6795 34772 6796
rect 34616 6774 34772 6795
rect 30585 6697 30700 6712
rect 30679 6694 30700 6697
rect 30718 6694 30736 6712
rect 30679 6675 30736 6694
rect 25908 6612 26023 6627
rect 25872 6589 26023 6612
rect 21560 6539 21660 6540
rect 21504 6518 21660 6539
rect 21504 6500 21524 6518
rect 21542 6500 21660 6518
rect 21504 6496 21660 6500
rect 17236 6419 17387 6442
rect 13303 6339 13360 6358
rect 12868 6326 13024 6330
rect 8838 6279 8994 6283
rect 8838 6261 8956 6279
rect 8974 6261 8994 6279
rect 8838 6240 8994 6261
rect 8838 6239 8938 6240
rect 4462 6168 4613 6191
rect 4462 6153 4577 6168
rect 4556 6150 4577 6153
rect 4595 6150 4613 6168
rect 185 6040 246 6056
rect 90 6036 246 6040
rect 90 6018 208 6036
rect 226 6018 246 6036
rect 4556 6131 4613 6150
rect 8839 6203 8881 6239
rect 12868 6310 12929 6326
rect 13297 6296 13358 6312
rect 17345 6383 17387 6419
rect 17474 6449 17630 6453
rect 17474 6431 17592 6449
rect 17610 6431 17630 6449
rect 17474 6410 17630 6431
rect 17474 6409 17574 6410
rect 17288 6382 17388 6383
rect 17232 6361 17388 6382
rect 17232 6343 17252 6361
rect 17270 6343 17388 6361
rect 17232 6339 17388 6343
rect 17475 6373 17517 6409
rect 21504 6480 21565 6496
rect 21933 6466 21994 6482
rect 25981 6553 26023 6589
rect 30249 6642 30306 6661
rect 30249 6624 30267 6642
rect 30285 6639 30306 6642
rect 34616 6756 34636 6774
rect 34654 6756 34772 6774
rect 34616 6752 34772 6756
rect 34616 6736 34677 6752
rect 30285 6624 30400 6639
rect 30249 6601 30400 6624
rect 25924 6552 26024 6553
rect 25868 6531 26024 6552
rect 25868 6513 25888 6531
rect 25906 6513 26024 6531
rect 25868 6509 26024 6513
rect 21838 6462 21994 6466
rect 21502 6434 21559 6453
rect 17475 6350 17626 6373
rect 13202 6292 13358 6296
rect 13202 6274 13320 6292
rect 13338 6274 13358 6292
rect 13202 6253 13358 6274
rect 13202 6252 13302 6253
rect 8839 6180 8990 6203
rect 8839 6165 8954 6180
rect 4126 6098 4183 6117
rect 4126 6080 4144 6098
rect 4162 6095 4183 6098
rect 4162 6080 4277 6095
rect 90 5997 246 6018
rect 90 5996 190 5997
rect 91 5960 133 5996
rect 91 5937 242 5960
rect 4126 6057 4277 6080
rect 4235 6021 4277 6057
rect 4549 6053 4610 6069
rect 4454 6049 4610 6053
rect 4454 6031 4572 6049
rect 4590 6031 4610 6049
rect 8933 6162 8954 6165
rect 8972 6162 8990 6180
rect 8933 6143 8990 6162
rect 13203 6216 13245 6252
rect 17232 6323 17293 6339
rect 17475 6335 17590 6350
rect 17569 6332 17590 6335
rect 17608 6332 17626 6350
rect 21502 6416 21520 6434
rect 21538 6431 21559 6434
rect 21838 6444 21956 6462
rect 21974 6444 21994 6462
rect 21538 6416 21653 6431
rect 21838 6423 21994 6444
rect 21838 6422 21938 6423
rect 21502 6393 21653 6416
rect 17569 6313 17626 6332
rect 17563 6270 17624 6286
rect 21611 6357 21653 6393
rect 21839 6386 21881 6422
rect 25868 6493 25929 6509
rect 26310 6478 26371 6494
rect 30358 6565 30400 6601
rect 34613 6655 34670 6674
rect 34613 6637 34631 6655
rect 34649 6652 34670 6655
rect 34649 6637 34764 6652
rect 34613 6614 34764 6637
rect 30301 6564 30401 6565
rect 30245 6543 30401 6564
rect 30245 6525 30265 6543
rect 30283 6525 30401 6543
rect 30245 6521 30401 6525
rect 26215 6474 26371 6478
rect 25866 6447 25923 6466
rect 21839 6363 21990 6386
rect 21554 6356 21654 6357
rect 21498 6335 21654 6356
rect 21839 6348 21954 6363
rect 21498 6317 21518 6335
rect 21536 6317 21654 6335
rect 21933 6345 21954 6348
rect 21972 6345 21990 6363
rect 25866 6429 25884 6447
rect 25902 6444 25923 6447
rect 26215 6456 26333 6474
rect 26351 6456 26371 6474
rect 25902 6429 26017 6444
rect 26215 6435 26371 6456
rect 26215 6434 26315 6435
rect 25866 6406 26017 6429
rect 21933 6326 21990 6345
rect 21498 6313 21654 6317
rect 17468 6266 17624 6270
rect 17468 6248 17586 6266
rect 17604 6248 17624 6266
rect 13203 6193 13354 6216
rect 13203 6178 13318 6193
rect 13297 6175 13318 6178
rect 13336 6175 13354 6193
rect 8490 6111 8547 6130
rect 8490 6093 8508 6111
rect 8526 6108 8547 6111
rect 8526 6093 8641 6108
rect 4178 6020 4278 6021
rect 4122 5999 4278 6020
rect 4454 6010 4610 6031
rect 4454 6009 4554 6010
rect 4122 5981 4142 5999
rect 4160 5981 4278 5999
rect 4122 5977 4278 5981
rect 4122 5961 4183 5977
rect 4455 5973 4497 6009
rect 91 5922 206 5937
rect 185 5919 206 5922
rect 224 5919 242 5937
rect 185 5900 242 5919
rect 4455 5950 4606 5973
rect 8490 6070 8641 6093
rect 8599 6034 8641 6070
rect 8926 6065 8987 6081
rect 8831 6061 8987 6065
rect 8831 6043 8949 6061
rect 8967 6043 8987 6061
rect 13297 6156 13354 6175
rect 17468 6227 17624 6248
rect 17468 6226 17568 6227
rect 17469 6190 17511 6226
rect 21498 6297 21559 6313
rect 21927 6283 21988 6299
rect 25975 6370 26017 6406
rect 26216 6398 26258 6434
rect 30245 6505 30306 6521
rect 30674 6491 30735 6507
rect 34722 6578 34764 6614
rect 34665 6577 34765 6578
rect 34609 6556 34765 6577
rect 34609 6538 34629 6556
rect 34647 6538 34765 6556
rect 34609 6534 34765 6538
rect 30579 6487 30735 6491
rect 30243 6459 30300 6478
rect 26216 6375 26367 6398
rect 25918 6369 26018 6370
rect 25862 6348 26018 6369
rect 26216 6360 26331 6375
rect 25862 6330 25882 6348
rect 25900 6330 26018 6348
rect 26310 6357 26331 6360
rect 26349 6357 26367 6375
rect 30243 6441 30261 6459
rect 30279 6456 30300 6459
rect 30579 6469 30697 6487
rect 30715 6469 30735 6487
rect 30279 6441 30394 6456
rect 30579 6448 30735 6469
rect 30579 6447 30679 6448
rect 30243 6418 30394 6441
rect 26310 6338 26367 6357
rect 25862 6326 26018 6330
rect 21832 6279 21988 6283
rect 21832 6261 21950 6279
rect 21968 6261 21988 6279
rect 21832 6240 21988 6261
rect 21832 6239 21932 6240
rect 12867 6123 12924 6142
rect 12867 6105 12885 6123
rect 12903 6120 12924 6123
rect 12903 6105 13018 6120
rect 8542 6033 8642 6034
rect 8486 6012 8642 6033
rect 8831 6022 8987 6043
rect 8831 6021 8931 6022
rect 8486 5994 8506 6012
rect 8524 5994 8642 6012
rect 8486 5990 8642 5994
rect 8486 5974 8547 5990
rect 8832 5985 8874 6021
rect 4455 5935 4570 5950
rect 4549 5932 4570 5935
rect 4588 5932 4606 5950
rect 4549 5913 4606 5932
rect 8832 5962 8983 5985
rect 12867 6082 13018 6105
rect 12976 6046 13018 6082
rect 13290 6078 13351 6094
rect 13195 6074 13351 6078
rect 13195 6056 13313 6074
rect 13331 6056 13351 6074
rect 17469 6167 17620 6190
rect 17231 6136 17288 6155
rect 17469 6152 17584 6167
rect 17231 6118 17249 6136
rect 17267 6133 17288 6136
rect 17563 6149 17584 6152
rect 17602 6149 17620 6167
rect 17267 6118 17382 6133
rect 17563 6130 17620 6149
rect 21833 6203 21875 6239
rect 25862 6310 25923 6326
rect 26304 6295 26365 6311
rect 30352 6382 30394 6418
rect 30580 6411 30622 6447
rect 34609 6518 34670 6534
rect 34607 6472 34664 6491
rect 30580 6388 30731 6411
rect 30295 6381 30395 6382
rect 30239 6360 30395 6381
rect 30580 6373 30695 6388
rect 30239 6342 30259 6360
rect 30277 6342 30395 6360
rect 30674 6370 30695 6373
rect 30713 6370 30731 6388
rect 34607 6454 34625 6472
rect 34643 6469 34664 6472
rect 34643 6454 34758 6469
rect 34607 6431 34758 6454
rect 30674 6351 30731 6370
rect 30239 6338 30395 6342
rect 26209 6291 26365 6295
rect 26209 6273 26327 6291
rect 26345 6273 26365 6291
rect 26209 6252 26365 6273
rect 26209 6251 26309 6252
rect 21833 6180 21984 6203
rect 21833 6165 21948 6180
rect 21927 6162 21948 6165
rect 21966 6162 21984 6180
rect 12919 6045 13019 6046
rect 12863 6024 13019 6045
rect 13195 6035 13351 6056
rect 13195 6034 13295 6035
rect 12863 6006 12883 6024
rect 12901 6006 13019 6024
rect 12863 6002 13019 6006
rect 12863 5986 12924 6002
rect 13196 5998 13238 6034
rect 8832 5947 8947 5962
rect 8926 5944 8947 5947
rect 8965 5944 8983 5962
rect 8926 5925 8983 5944
rect 13196 5975 13347 5998
rect 17231 6095 17382 6118
rect 17340 6059 17382 6095
rect 17283 6058 17383 6059
rect 17227 6037 17383 6058
rect 17556 6052 17617 6068
rect 17227 6019 17247 6037
rect 17265 6019 17383 6037
rect 17227 6015 17383 6019
rect 17461 6048 17617 6052
rect 17461 6030 17579 6048
rect 17597 6030 17617 6048
rect 21927 6143 21984 6162
rect 26210 6215 26252 6251
rect 30239 6322 30300 6338
rect 30668 6308 30729 6324
rect 34716 6395 34758 6431
rect 34659 6394 34759 6395
rect 34603 6373 34759 6394
rect 34603 6355 34623 6373
rect 34641 6355 34759 6373
rect 34603 6351 34759 6355
rect 30573 6304 30729 6308
rect 30573 6286 30691 6304
rect 30709 6286 30729 6304
rect 30573 6265 30729 6286
rect 30573 6264 30673 6265
rect 26210 6192 26361 6215
rect 26210 6177 26325 6192
rect 21497 6110 21554 6129
rect 21497 6092 21515 6110
rect 21533 6107 21554 6110
rect 21533 6092 21648 6107
rect 17227 5999 17288 6015
rect 17461 6009 17617 6030
rect 17461 6008 17561 6009
rect 13196 5960 13311 5975
rect 13290 5957 13311 5960
rect 13329 5957 13347 5975
rect 13290 5938 13347 5957
rect 17462 5972 17504 6008
rect 17462 5949 17613 5972
rect 21497 6069 21648 6092
rect 21606 6033 21648 6069
rect 21920 6065 21981 6081
rect 21825 6061 21981 6065
rect 21825 6043 21943 6061
rect 21961 6043 21981 6061
rect 26304 6174 26325 6177
rect 26343 6174 26361 6192
rect 26304 6155 26361 6174
rect 30574 6228 30616 6264
rect 34603 6335 34664 6351
rect 30574 6205 30725 6228
rect 30574 6190 30689 6205
rect 30668 6187 30689 6190
rect 30707 6187 30725 6205
rect 25861 6123 25918 6142
rect 25861 6105 25879 6123
rect 25897 6120 25918 6123
rect 25897 6105 26012 6120
rect 21549 6032 21649 6033
rect 21493 6011 21649 6032
rect 21825 6022 21981 6043
rect 21825 6021 21925 6022
rect 21493 5993 21513 6011
rect 21531 5993 21649 6011
rect 21493 5989 21649 5993
rect 21493 5973 21554 5989
rect 21826 5985 21868 6021
rect 17462 5934 17577 5949
rect 17556 5931 17577 5934
rect 17595 5931 17613 5949
rect 17556 5912 17613 5931
rect 21826 5962 21977 5985
rect 25861 6082 26012 6105
rect 25970 6046 26012 6082
rect 26297 6077 26358 6093
rect 26202 6073 26358 6077
rect 26202 6055 26320 6073
rect 26338 6055 26358 6073
rect 30668 6168 30725 6187
rect 30238 6135 30295 6154
rect 30238 6117 30256 6135
rect 30274 6132 30295 6135
rect 30274 6117 30389 6132
rect 25913 6045 26013 6046
rect 25857 6024 26013 6045
rect 26202 6034 26358 6055
rect 26202 6033 26302 6034
rect 25857 6006 25877 6024
rect 25895 6006 26013 6024
rect 25857 6002 26013 6006
rect 25857 5986 25918 6002
rect 26203 5997 26245 6033
rect 21826 5947 21941 5962
rect 21920 5944 21941 5947
rect 21959 5944 21977 5962
rect 21920 5925 21977 5944
rect 26203 5974 26354 5997
rect 30238 6094 30389 6117
rect 30347 6058 30389 6094
rect 30661 6090 30722 6106
rect 30566 6086 30722 6090
rect 30566 6068 30684 6086
rect 30702 6068 30722 6086
rect 34602 6148 34659 6167
rect 34602 6130 34620 6148
rect 34638 6145 34659 6148
rect 34638 6130 34753 6145
rect 30290 6057 30390 6058
rect 30234 6036 30390 6057
rect 30566 6047 30722 6068
rect 30566 6046 30666 6047
rect 30234 6018 30254 6036
rect 30272 6018 30390 6036
rect 30234 6014 30390 6018
rect 30234 5998 30295 6014
rect 30567 6010 30609 6046
rect 26203 5959 26318 5974
rect 26297 5956 26318 5959
rect 26336 5956 26354 5974
rect 26297 5937 26354 5956
rect 30567 5987 30718 6010
rect 34602 6107 34753 6130
rect 34711 6071 34753 6107
rect 34654 6070 34754 6071
rect 34598 6049 34754 6070
rect 34598 6031 34618 6049
rect 34636 6031 34754 6049
rect 34598 6027 34754 6031
rect 34598 6011 34659 6027
rect 30567 5972 30682 5987
rect 30661 5969 30682 5972
rect 30700 5969 30718 5987
rect 30661 5950 30718 5969
rect 4127 5805 4184 5824
rect 4127 5787 4145 5805
rect 4163 5802 4184 5805
rect 4163 5787 4278 5802
rect 186 5747 247 5763
rect 91 5743 247 5747
rect 91 5725 209 5743
rect 227 5725 247 5743
rect 91 5704 247 5725
rect 91 5703 191 5704
rect 92 5667 134 5703
rect 92 5644 243 5667
rect 4127 5764 4278 5787
rect 8491 5818 8548 5837
rect 8491 5800 8509 5818
rect 8527 5815 8548 5818
rect 8527 5800 8642 5815
rect 4236 5728 4278 5764
rect 4550 5760 4611 5776
rect 4455 5756 4611 5760
rect 4455 5738 4573 5756
rect 4591 5738 4611 5756
rect 4179 5727 4279 5728
rect 4123 5706 4279 5727
rect 4455 5717 4611 5738
rect 4455 5716 4555 5717
rect 92 5629 207 5644
rect 186 5626 207 5629
rect 225 5626 243 5644
rect 186 5607 243 5626
rect 4123 5688 4143 5706
rect 4161 5688 4279 5706
rect 4123 5684 4279 5688
rect 4123 5668 4184 5684
rect 4456 5680 4498 5716
rect 4456 5657 4607 5680
rect 8491 5777 8642 5800
rect 12868 5830 12925 5849
rect 12868 5812 12886 5830
rect 12904 5827 12925 5830
rect 12904 5812 13019 5827
rect 8600 5741 8642 5777
rect 8927 5772 8988 5788
rect 8832 5768 8988 5772
rect 8832 5750 8950 5768
rect 8968 5750 8988 5768
rect 8543 5740 8643 5741
rect 8487 5719 8643 5740
rect 8832 5729 8988 5750
rect 8832 5728 8932 5729
rect 4456 5642 4571 5657
rect 4550 5639 4571 5642
rect 4589 5639 4607 5657
rect 4550 5620 4607 5639
rect 4120 5587 4177 5606
rect 8487 5701 8507 5719
rect 8525 5701 8643 5719
rect 8487 5697 8643 5701
rect 8487 5681 8548 5697
rect 8833 5692 8875 5728
rect 8833 5669 8984 5692
rect 12868 5789 13019 5812
rect 17232 5843 17289 5862
rect 17232 5825 17250 5843
rect 17268 5840 17289 5843
rect 17268 5825 17383 5840
rect 12977 5753 13019 5789
rect 13291 5785 13352 5801
rect 13196 5781 13352 5785
rect 13196 5763 13314 5781
rect 13332 5763 13352 5781
rect 12920 5752 13020 5753
rect 12864 5731 13020 5752
rect 13196 5742 13352 5763
rect 13196 5741 13296 5742
rect 8833 5654 8948 5669
rect 8927 5651 8948 5654
rect 8966 5651 8984 5669
rect 8927 5632 8984 5651
rect 4120 5569 4138 5587
rect 4156 5584 4177 5587
rect 4156 5569 4271 5584
rect 4120 5546 4271 5569
rect 181 5423 242 5439
rect 4229 5510 4271 5546
rect 8484 5600 8541 5619
rect 8484 5582 8502 5600
rect 8520 5597 8541 5600
rect 12864 5713 12884 5731
rect 12902 5713 13020 5731
rect 12864 5709 13020 5713
rect 12864 5693 12925 5709
rect 13197 5705 13239 5741
rect 13197 5682 13348 5705
rect 17232 5802 17383 5825
rect 17341 5766 17383 5802
rect 21498 5817 21555 5836
rect 21498 5799 21516 5817
rect 21534 5814 21555 5817
rect 21534 5799 21649 5814
rect 17284 5765 17384 5766
rect 17228 5744 17384 5765
rect 17557 5759 17618 5775
rect 13197 5667 13312 5682
rect 13291 5664 13312 5667
rect 13330 5664 13348 5682
rect 13291 5645 13348 5664
rect 8520 5582 8635 5597
rect 8484 5559 8635 5582
rect 4172 5509 4272 5510
rect 4116 5488 4272 5509
rect 4116 5470 4136 5488
rect 4154 5470 4272 5488
rect 4116 5466 4272 5470
rect 86 5419 242 5423
rect 86 5401 204 5419
rect 222 5401 242 5419
rect 86 5380 242 5401
rect 86 5379 186 5380
rect 87 5343 129 5379
rect 4116 5450 4177 5466
rect 4545 5436 4606 5452
rect 8593 5523 8635 5559
rect 12861 5612 12918 5631
rect 17228 5726 17248 5744
rect 17266 5726 17384 5744
rect 17228 5722 17384 5726
rect 17462 5755 17618 5759
rect 17462 5737 17580 5755
rect 17598 5737 17618 5755
rect 17228 5706 17289 5722
rect 17462 5716 17618 5737
rect 17462 5715 17562 5716
rect 17463 5679 17505 5715
rect 17463 5656 17614 5679
rect 21498 5776 21649 5799
rect 25862 5830 25919 5849
rect 25862 5812 25880 5830
rect 25898 5827 25919 5830
rect 25898 5812 26013 5827
rect 21607 5740 21649 5776
rect 21921 5772 21982 5788
rect 21826 5768 21982 5772
rect 21826 5750 21944 5768
rect 21962 5750 21982 5768
rect 21550 5739 21650 5740
rect 21494 5718 21650 5739
rect 21826 5729 21982 5750
rect 21826 5728 21926 5729
rect 12861 5594 12879 5612
rect 12897 5609 12918 5612
rect 12897 5594 13012 5609
rect 12861 5571 13012 5594
rect 8536 5522 8636 5523
rect 8480 5501 8636 5522
rect 8480 5483 8500 5501
rect 8518 5483 8636 5501
rect 8480 5479 8636 5483
rect 4450 5432 4606 5436
rect 4114 5404 4171 5423
rect 87 5320 238 5343
rect 87 5305 202 5320
rect 181 5302 202 5305
rect 220 5302 238 5320
rect 4114 5386 4132 5404
rect 4150 5401 4171 5404
rect 4450 5414 4568 5432
rect 4586 5414 4606 5432
rect 4150 5386 4265 5401
rect 4450 5393 4606 5414
rect 4450 5392 4550 5393
rect 4114 5363 4265 5386
rect 181 5283 238 5302
rect 175 5240 236 5256
rect 4223 5327 4265 5363
rect 4451 5356 4493 5392
rect 8480 5463 8541 5479
rect 8922 5448 8983 5464
rect 12970 5535 13012 5571
rect 17225 5625 17282 5644
rect 17463 5641 17578 5656
rect 17225 5607 17243 5625
rect 17261 5622 17282 5625
rect 17557 5638 17578 5641
rect 17596 5638 17614 5656
rect 17261 5607 17376 5622
rect 17557 5619 17614 5638
rect 17225 5584 17376 5607
rect 21494 5700 21514 5718
rect 21532 5700 21650 5718
rect 21494 5696 21650 5700
rect 21494 5680 21555 5696
rect 21827 5692 21869 5728
rect 21827 5669 21978 5692
rect 25862 5789 26013 5812
rect 30239 5842 30296 5861
rect 30239 5824 30257 5842
rect 30275 5839 30296 5842
rect 30275 5824 30390 5839
rect 25971 5753 26013 5789
rect 26298 5784 26359 5800
rect 26203 5780 26359 5784
rect 26203 5762 26321 5780
rect 26339 5762 26359 5780
rect 25914 5752 26014 5753
rect 25858 5731 26014 5752
rect 26203 5741 26359 5762
rect 26203 5740 26303 5741
rect 21827 5654 21942 5669
rect 21921 5651 21942 5654
rect 21960 5651 21978 5669
rect 21921 5632 21978 5651
rect 12913 5534 13013 5535
rect 12857 5513 13013 5534
rect 12857 5495 12877 5513
rect 12895 5495 13013 5513
rect 12857 5491 13013 5495
rect 8827 5444 8983 5448
rect 8478 5417 8535 5436
rect 4451 5333 4602 5356
rect 4166 5326 4266 5327
rect 4110 5305 4266 5326
rect 4451 5318 4566 5333
rect 4110 5287 4130 5305
rect 4148 5287 4266 5305
rect 4545 5315 4566 5318
rect 4584 5315 4602 5333
rect 8478 5399 8496 5417
rect 8514 5414 8535 5417
rect 8827 5426 8945 5444
rect 8963 5426 8983 5444
rect 8514 5399 8629 5414
rect 8827 5405 8983 5426
rect 8827 5404 8927 5405
rect 8478 5376 8629 5399
rect 4545 5296 4602 5315
rect 4110 5283 4266 5287
rect 80 5236 236 5240
rect 80 5218 198 5236
rect 216 5218 236 5236
rect 80 5197 236 5218
rect 80 5196 180 5197
rect 81 5160 123 5196
rect 4110 5267 4171 5283
rect 4539 5253 4600 5269
rect 8587 5340 8629 5376
rect 8828 5368 8870 5404
rect 12857 5475 12918 5491
rect 13286 5461 13347 5477
rect 17334 5548 17376 5584
rect 17277 5547 17377 5548
rect 17221 5526 17377 5547
rect 21491 5599 21548 5618
rect 25858 5713 25878 5731
rect 25896 5713 26014 5731
rect 25858 5709 26014 5713
rect 25858 5693 25919 5709
rect 26204 5704 26246 5740
rect 26204 5681 26355 5704
rect 30239 5801 30390 5824
rect 34603 5855 34660 5874
rect 34603 5837 34621 5855
rect 34639 5852 34660 5855
rect 34639 5837 34754 5852
rect 30348 5765 30390 5801
rect 30662 5797 30723 5813
rect 30567 5793 30723 5797
rect 30567 5775 30685 5793
rect 30703 5775 30723 5793
rect 30291 5764 30391 5765
rect 30235 5743 30391 5764
rect 30567 5754 30723 5775
rect 30567 5753 30667 5754
rect 26204 5666 26319 5681
rect 26298 5663 26319 5666
rect 26337 5663 26355 5681
rect 26298 5644 26355 5663
rect 21491 5581 21509 5599
rect 21527 5596 21548 5599
rect 21527 5581 21642 5596
rect 21491 5558 21642 5581
rect 17221 5508 17241 5526
rect 17259 5508 17377 5526
rect 17221 5504 17377 5508
rect 13191 5457 13347 5461
rect 12855 5429 12912 5448
rect 8828 5345 8979 5368
rect 8530 5339 8630 5340
rect 8474 5318 8630 5339
rect 8828 5330 8943 5345
rect 8474 5300 8494 5318
rect 8512 5300 8630 5318
rect 8922 5327 8943 5330
rect 8961 5327 8979 5345
rect 12855 5411 12873 5429
rect 12891 5426 12912 5429
rect 13191 5439 13309 5457
rect 13327 5439 13347 5457
rect 12891 5411 13006 5426
rect 13191 5418 13347 5439
rect 13191 5417 13291 5418
rect 12855 5388 13006 5411
rect 8922 5308 8979 5327
rect 8474 5296 8630 5300
rect 4444 5249 4600 5253
rect 4444 5231 4562 5249
rect 4580 5231 4600 5249
rect 4444 5210 4600 5231
rect 4444 5209 4544 5210
rect 81 5137 232 5160
rect 81 5122 196 5137
rect 175 5119 196 5122
rect 214 5119 232 5137
rect 175 5100 232 5119
rect 4445 5173 4487 5209
rect 8474 5280 8535 5296
rect 8916 5265 8977 5281
rect 12964 5352 13006 5388
rect 13192 5381 13234 5417
rect 17221 5488 17282 5504
rect 17219 5442 17276 5461
rect 13192 5358 13343 5381
rect 12907 5351 13007 5352
rect 12851 5330 13007 5351
rect 13192 5343 13307 5358
rect 12851 5312 12871 5330
rect 12889 5312 13007 5330
rect 13286 5340 13307 5343
rect 13325 5340 13343 5358
rect 17219 5424 17237 5442
rect 17255 5439 17276 5442
rect 17255 5424 17370 5439
rect 17552 5435 17613 5451
rect 21600 5522 21642 5558
rect 25855 5612 25912 5631
rect 25855 5594 25873 5612
rect 25891 5609 25912 5612
rect 30235 5725 30255 5743
rect 30273 5725 30391 5743
rect 30235 5721 30391 5725
rect 30235 5705 30296 5721
rect 30568 5717 30610 5753
rect 30568 5694 30719 5717
rect 34603 5814 34754 5837
rect 34712 5778 34754 5814
rect 34655 5777 34755 5778
rect 34599 5756 34755 5777
rect 30568 5679 30683 5694
rect 30662 5676 30683 5679
rect 30701 5676 30719 5694
rect 30662 5657 30719 5676
rect 25891 5594 26006 5609
rect 25855 5571 26006 5594
rect 21543 5521 21643 5522
rect 21487 5500 21643 5521
rect 21487 5482 21507 5500
rect 21525 5482 21643 5500
rect 21487 5478 21643 5482
rect 17219 5401 17370 5424
rect 13286 5321 13343 5340
rect 12851 5308 13007 5312
rect 8821 5261 8977 5265
rect 8821 5243 8939 5261
rect 8957 5243 8977 5261
rect 8821 5222 8977 5243
rect 8821 5221 8921 5222
rect 4445 5150 4596 5173
rect 168 5022 229 5038
rect 73 5018 229 5022
rect 73 5000 191 5018
rect 209 5000 229 5018
rect 4445 5135 4560 5150
rect 4539 5132 4560 5135
rect 4578 5132 4596 5150
rect 4539 5113 4596 5132
rect 8822 5185 8864 5221
rect 12851 5292 12912 5308
rect 13280 5278 13341 5294
rect 17328 5365 17370 5401
rect 17457 5431 17613 5435
rect 17457 5413 17575 5431
rect 17593 5413 17613 5431
rect 17457 5392 17613 5413
rect 17457 5391 17557 5392
rect 17271 5364 17371 5365
rect 17215 5343 17371 5364
rect 17215 5325 17235 5343
rect 17253 5325 17371 5343
rect 17215 5321 17371 5325
rect 17458 5355 17500 5391
rect 21487 5462 21548 5478
rect 21916 5448 21977 5464
rect 25964 5535 26006 5571
rect 30232 5624 30289 5643
rect 34599 5738 34619 5756
rect 34637 5738 34755 5756
rect 34599 5734 34755 5738
rect 34599 5718 34660 5734
rect 30232 5606 30250 5624
rect 30268 5621 30289 5624
rect 30268 5606 30383 5621
rect 30232 5583 30383 5606
rect 25907 5534 26007 5535
rect 25851 5513 26007 5534
rect 25851 5495 25871 5513
rect 25889 5495 26007 5513
rect 25851 5491 26007 5495
rect 21821 5444 21977 5448
rect 21485 5416 21542 5435
rect 17458 5332 17609 5355
rect 13185 5274 13341 5278
rect 13185 5256 13303 5274
rect 13321 5256 13341 5274
rect 13185 5235 13341 5256
rect 13185 5234 13285 5235
rect 8822 5162 8973 5185
rect 4109 5080 4166 5099
rect 4109 5062 4127 5080
rect 4145 5077 4166 5080
rect 4145 5062 4260 5077
rect 73 4979 229 5000
rect 73 4978 173 4979
rect 74 4942 116 4978
rect 74 4919 225 4942
rect 4109 5039 4260 5062
rect 4218 5003 4260 5039
rect 4532 5035 4593 5051
rect 4437 5031 4593 5035
rect 4437 5013 4555 5031
rect 4573 5013 4593 5031
rect 8822 5147 8937 5162
rect 8916 5144 8937 5147
rect 8955 5144 8973 5162
rect 8916 5125 8973 5144
rect 13186 5198 13228 5234
rect 17215 5305 17276 5321
rect 17458 5317 17573 5332
rect 17552 5314 17573 5317
rect 17591 5314 17609 5332
rect 21485 5398 21503 5416
rect 21521 5413 21542 5416
rect 21821 5426 21939 5444
rect 21957 5426 21977 5444
rect 21521 5398 21636 5413
rect 21821 5405 21977 5426
rect 21821 5404 21921 5405
rect 21485 5375 21636 5398
rect 17552 5295 17609 5314
rect 17546 5252 17607 5268
rect 21594 5339 21636 5375
rect 21822 5368 21864 5404
rect 25851 5475 25912 5491
rect 26293 5460 26354 5476
rect 30341 5547 30383 5583
rect 34596 5637 34653 5656
rect 34596 5619 34614 5637
rect 34632 5634 34653 5637
rect 34632 5619 34747 5634
rect 34596 5596 34747 5619
rect 30284 5546 30384 5547
rect 30228 5525 30384 5546
rect 30228 5507 30248 5525
rect 30266 5507 30384 5525
rect 30228 5503 30384 5507
rect 26198 5456 26354 5460
rect 25849 5429 25906 5448
rect 21822 5345 21973 5368
rect 21537 5338 21637 5339
rect 21481 5317 21637 5338
rect 21822 5330 21937 5345
rect 21481 5299 21501 5317
rect 21519 5299 21637 5317
rect 21916 5327 21937 5330
rect 21955 5327 21973 5345
rect 25849 5411 25867 5429
rect 25885 5426 25906 5429
rect 26198 5438 26316 5456
rect 26334 5438 26354 5456
rect 25885 5411 26000 5426
rect 26198 5417 26354 5438
rect 26198 5416 26298 5417
rect 25849 5388 26000 5411
rect 21916 5308 21973 5327
rect 21481 5295 21637 5299
rect 17451 5248 17607 5252
rect 17451 5230 17569 5248
rect 17587 5230 17607 5248
rect 13186 5175 13337 5198
rect 8473 5093 8530 5112
rect 8473 5075 8491 5093
rect 8509 5090 8530 5093
rect 8509 5075 8624 5090
rect 4161 5002 4261 5003
rect 4105 4981 4261 5002
rect 4437 4992 4593 5013
rect 4437 4991 4537 4992
rect 4105 4963 4125 4981
rect 4143 4963 4261 4981
rect 4105 4959 4261 4963
rect 4105 4943 4166 4959
rect 4438 4955 4480 4991
rect 74 4904 189 4919
rect 168 4901 189 4904
rect 207 4901 225 4919
rect 168 4882 225 4901
rect 4438 4932 4589 4955
rect 8473 5052 8624 5075
rect 8582 5016 8624 5052
rect 8909 5047 8970 5063
rect 8814 5043 8970 5047
rect 8814 5025 8932 5043
rect 8950 5025 8970 5043
rect 13186 5160 13301 5175
rect 13280 5157 13301 5160
rect 13319 5157 13337 5175
rect 13280 5138 13337 5157
rect 17451 5209 17607 5230
rect 17451 5208 17551 5209
rect 12850 5105 12907 5124
rect 12850 5087 12868 5105
rect 12886 5102 12907 5105
rect 12886 5087 13001 5102
rect 8525 5015 8625 5016
rect 8469 4994 8625 5015
rect 8814 5004 8970 5025
rect 8814 5003 8914 5004
rect 8469 4976 8489 4994
rect 8507 4976 8625 4994
rect 8469 4972 8625 4976
rect 8469 4956 8530 4972
rect 8815 4967 8857 5003
rect 4438 4917 4553 4932
rect 4532 4914 4553 4917
rect 4571 4914 4589 4932
rect 4532 4895 4589 4914
rect 8815 4944 8966 4967
rect 12850 5064 13001 5087
rect 12959 5028 13001 5064
rect 13273 5060 13334 5076
rect 13178 5056 13334 5060
rect 13178 5038 13296 5056
rect 13314 5038 13334 5056
rect 17452 5172 17494 5208
rect 21481 5279 21542 5295
rect 21910 5265 21971 5281
rect 25958 5352 26000 5388
rect 26199 5380 26241 5416
rect 30228 5487 30289 5503
rect 30657 5473 30718 5489
rect 34705 5560 34747 5596
rect 34648 5559 34748 5560
rect 34592 5538 34748 5559
rect 34592 5520 34612 5538
rect 34630 5520 34748 5538
rect 34592 5516 34748 5520
rect 30562 5469 30718 5473
rect 30226 5441 30283 5460
rect 26199 5357 26350 5380
rect 25901 5351 26001 5352
rect 25845 5330 26001 5351
rect 26199 5342 26314 5357
rect 25845 5312 25865 5330
rect 25883 5312 26001 5330
rect 26293 5339 26314 5342
rect 26332 5339 26350 5357
rect 30226 5423 30244 5441
rect 30262 5438 30283 5441
rect 30562 5451 30680 5469
rect 30698 5451 30718 5469
rect 30262 5423 30377 5438
rect 30562 5430 30718 5451
rect 30562 5429 30662 5430
rect 30226 5400 30377 5423
rect 26293 5320 26350 5339
rect 25845 5308 26001 5312
rect 21815 5261 21971 5265
rect 21815 5243 21933 5261
rect 21951 5243 21971 5261
rect 21815 5222 21971 5243
rect 21815 5221 21915 5222
rect 17452 5149 17603 5172
rect 17214 5118 17271 5137
rect 17452 5134 17567 5149
rect 17214 5100 17232 5118
rect 17250 5115 17271 5118
rect 17546 5131 17567 5134
rect 17585 5131 17603 5149
rect 17250 5100 17365 5115
rect 17546 5112 17603 5131
rect 21816 5185 21858 5221
rect 25845 5292 25906 5308
rect 26287 5277 26348 5293
rect 30335 5364 30377 5400
rect 30563 5393 30605 5429
rect 34592 5500 34653 5516
rect 34590 5454 34647 5473
rect 30563 5370 30714 5393
rect 30278 5363 30378 5364
rect 30222 5342 30378 5363
rect 30563 5355 30678 5370
rect 30222 5324 30242 5342
rect 30260 5324 30378 5342
rect 30657 5352 30678 5355
rect 30696 5352 30714 5370
rect 34590 5436 34608 5454
rect 34626 5451 34647 5454
rect 34626 5436 34741 5451
rect 34590 5413 34741 5436
rect 30657 5333 30714 5352
rect 30222 5320 30378 5324
rect 26192 5273 26348 5277
rect 26192 5255 26310 5273
rect 26328 5255 26348 5273
rect 26192 5234 26348 5255
rect 26192 5233 26292 5234
rect 21816 5162 21967 5185
rect 12902 5027 13002 5028
rect 12846 5006 13002 5027
rect 13178 5017 13334 5038
rect 13178 5016 13278 5017
rect 12846 4988 12866 5006
rect 12884 4988 13002 5006
rect 12846 4984 13002 4988
rect 12846 4968 12907 4984
rect 13179 4980 13221 5016
rect 8815 4929 8930 4944
rect 8909 4926 8930 4929
rect 8948 4926 8966 4944
rect 8909 4907 8966 4926
rect 13179 4957 13330 4980
rect 17214 5077 17365 5100
rect 17323 5041 17365 5077
rect 17266 5040 17366 5041
rect 17210 5019 17366 5040
rect 17539 5034 17600 5050
rect 17210 5001 17230 5019
rect 17248 5001 17366 5019
rect 17210 4997 17366 5001
rect 17444 5030 17600 5034
rect 17444 5012 17562 5030
rect 17580 5012 17600 5030
rect 21816 5147 21931 5162
rect 21910 5144 21931 5147
rect 21949 5144 21967 5162
rect 21910 5125 21967 5144
rect 26193 5197 26235 5233
rect 30222 5304 30283 5320
rect 30651 5290 30712 5306
rect 34699 5377 34741 5413
rect 34642 5376 34742 5377
rect 34586 5355 34742 5376
rect 34586 5337 34606 5355
rect 34624 5337 34742 5355
rect 34586 5333 34742 5337
rect 30556 5286 30712 5290
rect 30556 5268 30674 5286
rect 30692 5268 30712 5286
rect 30556 5247 30712 5268
rect 30556 5246 30656 5247
rect 26193 5174 26344 5197
rect 21480 5092 21537 5111
rect 21480 5074 21498 5092
rect 21516 5089 21537 5092
rect 21516 5074 21631 5089
rect 17210 4981 17271 4997
rect 17444 4991 17600 5012
rect 17444 4990 17544 4991
rect 13179 4942 13294 4957
rect 13273 4939 13294 4942
rect 13312 4939 13330 4957
rect 13273 4920 13330 4939
rect 17445 4954 17487 4990
rect 17445 4931 17596 4954
rect 21480 5051 21631 5074
rect 21589 5015 21631 5051
rect 21903 5047 21964 5063
rect 21808 5043 21964 5047
rect 21808 5025 21926 5043
rect 21944 5025 21964 5043
rect 26193 5159 26308 5174
rect 26287 5156 26308 5159
rect 26326 5156 26344 5174
rect 26287 5137 26344 5156
rect 30557 5210 30599 5246
rect 34586 5317 34647 5333
rect 30557 5187 30708 5210
rect 25844 5105 25901 5124
rect 25844 5087 25862 5105
rect 25880 5102 25901 5105
rect 25880 5087 25995 5102
rect 21532 5014 21632 5015
rect 21476 4993 21632 5014
rect 21808 5004 21964 5025
rect 21808 5003 21908 5004
rect 21476 4975 21496 4993
rect 21514 4975 21632 4993
rect 21476 4971 21632 4975
rect 21476 4955 21537 4971
rect 21809 4967 21851 5003
rect 17445 4916 17560 4931
rect 17539 4913 17560 4916
rect 17578 4913 17596 4931
rect 17539 4894 17596 4913
rect 21809 4944 21960 4967
rect 25844 5064 25995 5087
rect 25953 5028 25995 5064
rect 26280 5059 26341 5075
rect 26185 5055 26341 5059
rect 26185 5037 26303 5055
rect 26321 5037 26341 5055
rect 30557 5172 30672 5187
rect 30651 5169 30672 5172
rect 30690 5169 30708 5187
rect 30651 5150 30708 5169
rect 30221 5117 30278 5136
rect 30221 5099 30239 5117
rect 30257 5114 30278 5117
rect 30257 5099 30372 5114
rect 25896 5027 25996 5028
rect 25840 5006 25996 5027
rect 26185 5016 26341 5037
rect 26185 5015 26285 5016
rect 25840 4988 25860 5006
rect 25878 4988 25996 5006
rect 25840 4984 25996 4988
rect 25840 4968 25901 4984
rect 26186 4979 26228 5015
rect 21809 4929 21924 4944
rect 21903 4926 21924 4929
rect 21942 4926 21960 4944
rect 21903 4907 21960 4926
rect 26186 4956 26337 4979
rect 30221 5076 30372 5099
rect 30330 5040 30372 5076
rect 30644 5072 30705 5088
rect 30549 5068 30705 5072
rect 30549 5050 30667 5068
rect 30685 5050 30705 5068
rect 34585 5130 34642 5149
rect 34585 5112 34603 5130
rect 34621 5127 34642 5130
rect 34621 5112 34736 5127
rect 30273 5039 30373 5040
rect 30217 5018 30373 5039
rect 30549 5029 30705 5050
rect 30549 5028 30649 5029
rect 30217 5000 30237 5018
rect 30255 5000 30373 5018
rect 30217 4996 30373 5000
rect 30217 4980 30278 4996
rect 30550 4992 30592 5028
rect 26186 4941 26301 4956
rect 26280 4938 26301 4941
rect 26319 4938 26337 4956
rect 26280 4919 26337 4938
rect 30550 4969 30701 4992
rect 34585 5089 34736 5112
rect 34694 5053 34736 5089
rect 34637 5052 34737 5053
rect 34581 5031 34737 5052
rect 34581 5013 34601 5031
rect 34619 5013 34737 5031
rect 34581 5009 34737 5013
rect 34581 4993 34642 5009
rect 30550 4954 30665 4969
rect 30644 4951 30665 4954
rect 30683 4951 30701 4969
rect 30644 4932 30701 4951
rect 4108 4787 4165 4806
rect 4108 4769 4126 4787
rect 4144 4784 4165 4787
rect 4144 4769 4259 4784
rect 167 4729 228 4745
rect 72 4725 228 4729
rect 72 4707 190 4725
rect 208 4707 228 4725
rect 72 4686 228 4707
rect 72 4685 172 4686
rect 73 4649 115 4685
rect 73 4626 224 4649
rect 4108 4746 4259 4769
rect 8472 4800 8529 4819
rect 8472 4782 8490 4800
rect 8508 4797 8529 4800
rect 8508 4782 8623 4797
rect 4217 4710 4259 4746
rect 4531 4742 4592 4758
rect 4436 4738 4592 4742
rect 4436 4720 4554 4738
rect 4572 4720 4592 4738
rect 4160 4709 4260 4710
rect 4104 4688 4260 4709
rect 4436 4699 4592 4720
rect 4436 4698 4536 4699
rect 73 4611 188 4626
rect 167 4608 188 4611
rect 206 4608 224 4626
rect 167 4589 224 4608
rect 4104 4670 4124 4688
rect 4142 4670 4260 4688
rect 4104 4666 4260 4670
rect 4104 4650 4165 4666
rect 4437 4662 4479 4698
rect 4437 4639 4588 4662
rect 8472 4759 8623 4782
rect 12849 4812 12906 4831
rect 12849 4794 12867 4812
rect 12885 4809 12906 4812
rect 12885 4794 13000 4809
rect 8581 4723 8623 4759
rect 8908 4754 8969 4770
rect 8813 4750 8969 4754
rect 8813 4732 8931 4750
rect 8949 4732 8969 4750
rect 8524 4722 8624 4723
rect 8468 4701 8624 4722
rect 8813 4711 8969 4732
rect 8813 4710 8913 4711
rect 4437 4624 4552 4639
rect 4531 4621 4552 4624
rect 4570 4621 4588 4639
rect 4531 4602 4588 4621
rect 4101 4569 4158 4588
rect 4101 4551 4119 4569
rect 4137 4566 4158 4569
rect 4137 4551 4252 4566
rect 8468 4683 8488 4701
rect 8506 4683 8624 4701
rect 8468 4679 8624 4683
rect 8468 4663 8529 4679
rect 8814 4674 8856 4710
rect 8814 4651 8965 4674
rect 12849 4771 13000 4794
rect 17213 4825 17270 4844
rect 17213 4807 17231 4825
rect 17249 4822 17270 4825
rect 17249 4807 17364 4822
rect 12958 4735 13000 4771
rect 13272 4767 13333 4783
rect 13177 4763 13333 4767
rect 13177 4745 13295 4763
rect 13313 4745 13333 4763
rect 12901 4734 13001 4735
rect 12845 4713 13001 4734
rect 13177 4724 13333 4745
rect 13177 4723 13277 4724
rect 8814 4636 8929 4651
rect 8908 4633 8929 4636
rect 8947 4633 8965 4651
rect 8908 4614 8965 4633
rect 4101 4528 4252 4551
rect 162 4405 223 4421
rect 4210 4492 4252 4528
rect 8465 4582 8522 4601
rect 8465 4564 8483 4582
rect 8501 4579 8522 4582
rect 8501 4564 8616 4579
rect 12845 4695 12865 4713
rect 12883 4695 13001 4713
rect 12845 4691 13001 4695
rect 12845 4675 12906 4691
rect 13178 4687 13220 4723
rect 13178 4664 13329 4687
rect 17213 4784 17364 4807
rect 17322 4748 17364 4784
rect 21479 4799 21536 4818
rect 21479 4781 21497 4799
rect 21515 4796 21536 4799
rect 21515 4781 21630 4796
rect 17265 4747 17365 4748
rect 17209 4726 17365 4747
rect 17538 4741 17599 4757
rect 13178 4649 13293 4664
rect 13272 4646 13293 4649
rect 13311 4646 13329 4664
rect 13272 4627 13329 4646
rect 8465 4541 8616 4564
rect 4153 4491 4253 4492
rect 4097 4470 4253 4491
rect 4097 4452 4117 4470
rect 4135 4452 4253 4470
rect 4097 4448 4253 4452
rect 67 4401 223 4405
rect 67 4383 185 4401
rect 203 4383 223 4401
rect 67 4362 223 4383
rect 67 4361 167 4362
rect 68 4325 110 4361
rect 4097 4432 4158 4448
rect 4526 4418 4587 4434
rect 8574 4505 8616 4541
rect 12842 4594 12899 4613
rect 12842 4576 12860 4594
rect 12878 4591 12899 4594
rect 12878 4576 12993 4591
rect 17209 4708 17229 4726
rect 17247 4708 17365 4726
rect 17209 4704 17365 4708
rect 17443 4737 17599 4741
rect 17443 4719 17561 4737
rect 17579 4719 17599 4737
rect 17209 4688 17270 4704
rect 17443 4698 17599 4719
rect 17443 4697 17543 4698
rect 17444 4661 17486 4697
rect 17444 4638 17595 4661
rect 21479 4758 21630 4781
rect 25843 4812 25900 4831
rect 25843 4794 25861 4812
rect 25879 4809 25900 4812
rect 25879 4794 25994 4809
rect 21588 4722 21630 4758
rect 21902 4754 21963 4770
rect 21807 4750 21963 4754
rect 21807 4732 21925 4750
rect 21943 4732 21963 4750
rect 21531 4721 21631 4722
rect 21475 4700 21631 4721
rect 21807 4711 21963 4732
rect 21807 4710 21907 4711
rect 12842 4553 12993 4576
rect 8517 4504 8617 4505
rect 8461 4483 8617 4504
rect 8461 4465 8481 4483
rect 8499 4465 8617 4483
rect 8461 4461 8617 4465
rect 4431 4414 4587 4418
rect 4095 4386 4152 4405
rect 68 4302 219 4325
rect 68 4287 183 4302
rect 162 4284 183 4287
rect 201 4284 219 4302
rect 4095 4368 4113 4386
rect 4131 4383 4152 4386
rect 4431 4396 4549 4414
rect 4567 4396 4587 4414
rect 4131 4368 4246 4383
rect 4431 4375 4587 4396
rect 4431 4374 4531 4375
rect 4095 4345 4246 4368
rect 162 4265 219 4284
rect 156 4222 217 4238
rect 4204 4309 4246 4345
rect 4432 4338 4474 4374
rect 8461 4445 8522 4461
rect 8903 4430 8964 4446
rect 12951 4517 12993 4553
rect 17206 4607 17263 4626
rect 17444 4623 17559 4638
rect 17206 4589 17224 4607
rect 17242 4604 17263 4607
rect 17538 4620 17559 4623
rect 17577 4620 17595 4638
rect 17242 4589 17357 4604
rect 17538 4601 17595 4620
rect 17206 4566 17357 4589
rect 12894 4516 12994 4517
rect 12838 4495 12994 4516
rect 12838 4477 12858 4495
rect 12876 4477 12994 4495
rect 12838 4473 12994 4477
rect 8808 4426 8964 4430
rect 8459 4399 8516 4418
rect 4432 4315 4583 4338
rect 4147 4308 4247 4309
rect 4091 4287 4247 4308
rect 4432 4300 4547 4315
rect 4091 4269 4111 4287
rect 4129 4269 4247 4287
rect 4526 4297 4547 4300
rect 4565 4297 4583 4315
rect 8459 4381 8477 4399
rect 8495 4396 8516 4399
rect 8808 4408 8926 4426
rect 8944 4408 8964 4426
rect 8495 4381 8610 4396
rect 8808 4387 8964 4408
rect 8808 4386 8908 4387
rect 8459 4358 8610 4381
rect 4526 4278 4583 4297
rect 4091 4265 4247 4269
rect 61 4218 217 4222
rect 61 4200 179 4218
rect 197 4200 217 4218
rect 61 4179 217 4200
rect 61 4178 161 4179
rect 62 4142 104 4178
rect 4091 4249 4152 4265
rect 4520 4235 4581 4251
rect 8568 4322 8610 4358
rect 8809 4350 8851 4386
rect 12838 4457 12899 4473
rect 13267 4443 13328 4459
rect 17315 4530 17357 4566
rect 21475 4682 21495 4700
rect 21513 4682 21631 4700
rect 21475 4678 21631 4682
rect 21475 4662 21536 4678
rect 21808 4674 21850 4710
rect 21808 4651 21959 4674
rect 25843 4771 25994 4794
rect 30220 4824 30277 4843
rect 30220 4806 30238 4824
rect 30256 4821 30277 4824
rect 30256 4806 30371 4821
rect 25952 4735 25994 4771
rect 26279 4766 26340 4782
rect 26184 4762 26340 4766
rect 26184 4744 26302 4762
rect 26320 4744 26340 4762
rect 25895 4734 25995 4735
rect 25839 4713 25995 4734
rect 26184 4723 26340 4744
rect 26184 4722 26284 4723
rect 21808 4636 21923 4651
rect 21902 4633 21923 4636
rect 21941 4633 21959 4651
rect 21902 4614 21959 4633
rect 17258 4529 17358 4530
rect 17202 4508 17358 4529
rect 21472 4581 21529 4600
rect 21472 4563 21490 4581
rect 21508 4578 21529 4581
rect 21508 4563 21623 4578
rect 25839 4695 25859 4713
rect 25877 4695 25995 4713
rect 25839 4691 25995 4695
rect 25839 4675 25900 4691
rect 26185 4686 26227 4722
rect 26185 4663 26336 4686
rect 30220 4783 30371 4806
rect 34584 4837 34641 4856
rect 34584 4819 34602 4837
rect 34620 4834 34641 4837
rect 34620 4819 34735 4834
rect 30329 4747 30371 4783
rect 30643 4779 30704 4795
rect 30548 4775 30704 4779
rect 30548 4757 30666 4775
rect 30684 4757 30704 4775
rect 30272 4746 30372 4747
rect 30216 4725 30372 4746
rect 30548 4736 30704 4757
rect 30548 4735 30648 4736
rect 26185 4648 26300 4663
rect 26279 4645 26300 4648
rect 26318 4645 26336 4663
rect 26279 4626 26336 4645
rect 21472 4540 21623 4563
rect 17202 4490 17222 4508
rect 17240 4490 17358 4508
rect 17202 4486 17358 4490
rect 13172 4439 13328 4443
rect 12836 4411 12893 4430
rect 8809 4327 8960 4350
rect 8511 4321 8611 4322
rect 8455 4300 8611 4321
rect 8809 4312 8924 4327
rect 8455 4282 8475 4300
rect 8493 4282 8611 4300
rect 8903 4309 8924 4312
rect 8942 4309 8960 4327
rect 12836 4393 12854 4411
rect 12872 4408 12893 4411
rect 13172 4421 13290 4439
rect 13308 4421 13328 4439
rect 12872 4393 12987 4408
rect 13172 4400 13328 4421
rect 13172 4399 13272 4400
rect 12836 4370 12987 4393
rect 8903 4290 8960 4309
rect 8455 4278 8611 4282
rect 4425 4231 4581 4235
rect 4425 4213 4543 4231
rect 4561 4213 4581 4231
rect 4425 4192 4581 4213
rect 4425 4191 4525 4192
rect 62 4119 213 4142
rect 62 4104 177 4119
rect 156 4101 177 4104
rect 195 4101 213 4119
rect 156 4082 213 4101
rect 4426 4155 4468 4191
rect 8455 4262 8516 4278
rect 8897 4247 8958 4263
rect 12945 4334 12987 4370
rect 13173 4363 13215 4399
rect 17202 4470 17263 4486
rect 17200 4424 17257 4443
rect 13173 4340 13324 4363
rect 12888 4333 12988 4334
rect 12832 4312 12988 4333
rect 13173 4325 13288 4340
rect 12832 4294 12852 4312
rect 12870 4294 12988 4312
rect 13267 4322 13288 4325
rect 13306 4322 13324 4340
rect 17200 4406 17218 4424
rect 17236 4421 17257 4424
rect 17236 4406 17351 4421
rect 17533 4417 17594 4433
rect 21581 4504 21623 4540
rect 25836 4594 25893 4613
rect 25836 4576 25854 4594
rect 25872 4591 25893 4594
rect 25872 4576 25987 4591
rect 30216 4707 30236 4725
rect 30254 4707 30372 4725
rect 30216 4703 30372 4707
rect 30216 4687 30277 4703
rect 30549 4699 30591 4735
rect 30549 4676 30700 4699
rect 34584 4796 34735 4819
rect 34693 4760 34735 4796
rect 34636 4759 34736 4760
rect 34580 4738 34736 4759
rect 30549 4661 30664 4676
rect 30643 4658 30664 4661
rect 30682 4658 30700 4676
rect 30643 4639 30700 4658
rect 25836 4553 25987 4576
rect 21524 4503 21624 4504
rect 21468 4482 21624 4503
rect 21468 4464 21488 4482
rect 21506 4464 21624 4482
rect 21468 4460 21624 4464
rect 17200 4383 17351 4406
rect 13267 4303 13324 4322
rect 12832 4290 12988 4294
rect 8802 4243 8958 4247
rect 8802 4225 8920 4243
rect 8938 4225 8958 4243
rect 8802 4204 8958 4225
rect 8802 4203 8902 4204
rect 4426 4132 4577 4155
rect 4426 4117 4541 4132
rect 4520 4114 4541 4117
rect 4559 4114 4577 4132
rect 149 4004 210 4020
rect 54 4000 210 4004
rect 54 3982 172 4000
rect 190 3982 210 4000
rect 4520 4095 4577 4114
rect 8803 4167 8845 4203
rect 12832 4274 12893 4290
rect 13261 4260 13322 4276
rect 17309 4347 17351 4383
rect 17438 4413 17594 4417
rect 17438 4395 17556 4413
rect 17574 4395 17594 4413
rect 17438 4374 17594 4395
rect 17438 4373 17538 4374
rect 17252 4346 17352 4347
rect 17196 4325 17352 4346
rect 17196 4307 17216 4325
rect 17234 4307 17352 4325
rect 17196 4303 17352 4307
rect 17439 4337 17481 4373
rect 21468 4444 21529 4460
rect 21897 4430 21958 4446
rect 25945 4517 25987 4553
rect 30213 4606 30270 4625
rect 30213 4588 30231 4606
rect 30249 4603 30270 4606
rect 30249 4588 30364 4603
rect 34580 4720 34600 4738
rect 34618 4720 34736 4738
rect 34580 4716 34736 4720
rect 34580 4700 34641 4716
rect 30213 4565 30364 4588
rect 25888 4516 25988 4517
rect 25832 4495 25988 4516
rect 25832 4477 25852 4495
rect 25870 4477 25988 4495
rect 25832 4473 25988 4477
rect 21802 4426 21958 4430
rect 21466 4398 21523 4417
rect 17439 4314 17590 4337
rect 13166 4256 13322 4260
rect 13166 4238 13284 4256
rect 13302 4238 13322 4256
rect 13166 4217 13322 4238
rect 13166 4216 13266 4217
rect 8803 4144 8954 4167
rect 8803 4129 8918 4144
rect 4090 4062 4147 4081
rect 4090 4044 4108 4062
rect 4126 4059 4147 4062
rect 4126 4044 4241 4059
rect 54 3961 210 3982
rect 54 3960 154 3961
rect 55 3924 97 3960
rect 55 3901 206 3924
rect 4090 4021 4241 4044
rect 4199 3985 4241 4021
rect 4513 4017 4574 4033
rect 4418 4013 4574 4017
rect 4418 3995 4536 4013
rect 4554 3995 4574 4013
rect 8897 4126 8918 4129
rect 8936 4126 8954 4144
rect 8897 4107 8954 4126
rect 13167 4180 13209 4216
rect 17196 4287 17257 4303
rect 17439 4299 17554 4314
rect 17533 4296 17554 4299
rect 17572 4296 17590 4314
rect 21466 4380 21484 4398
rect 21502 4395 21523 4398
rect 21802 4408 21920 4426
rect 21938 4408 21958 4426
rect 21502 4380 21617 4395
rect 21802 4387 21958 4408
rect 21802 4386 21902 4387
rect 21466 4357 21617 4380
rect 17533 4277 17590 4296
rect 17527 4234 17588 4250
rect 21575 4321 21617 4357
rect 21803 4350 21845 4386
rect 25832 4457 25893 4473
rect 26274 4442 26335 4458
rect 30322 4529 30364 4565
rect 34577 4619 34634 4638
rect 34577 4601 34595 4619
rect 34613 4616 34634 4619
rect 34613 4601 34728 4616
rect 34577 4578 34728 4601
rect 30265 4528 30365 4529
rect 30209 4507 30365 4528
rect 30209 4489 30229 4507
rect 30247 4489 30365 4507
rect 30209 4485 30365 4489
rect 26179 4438 26335 4442
rect 25830 4411 25887 4430
rect 21803 4327 21954 4350
rect 21518 4320 21618 4321
rect 21462 4299 21618 4320
rect 21803 4312 21918 4327
rect 21462 4281 21482 4299
rect 21500 4281 21618 4299
rect 21897 4309 21918 4312
rect 21936 4309 21954 4327
rect 25830 4393 25848 4411
rect 25866 4408 25887 4411
rect 26179 4420 26297 4438
rect 26315 4420 26335 4438
rect 25866 4393 25981 4408
rect 26179 4399 26335 4420
rect 26179 4398 26279 4399
rect 25830 4370 25981 4393
rect 21897 4290 21954 4309
rect 21462 4277 21618 4281
rect 17432 4230 17588 4234
rect 17432 4212 17550 4230
rect 17568 4212 17588 4230
rect 13167 4157 13318 4180
rect 13167 4142 13282 4157
rect 13261 4139 13282 4142
rect 13300 4139 13318 4157
rect 8454 4075 8511 4094
rect 8454 4057 8472 4075
rect 8490 4072 8511 4075
rect 8490 4057 8605 4072
rect 4142 3984 4242 3985
rect 4086 3963 4242 3984
rect 4418 3974 4574 3995
rect 4418 3973 4518 3974
rect 4086 3945 4106 3963
rect 4124 3945 4242 3963
rect 4086 3941 4242 3945
rect 4086 3925 4147 3941
rect 4419 3937 4461 3973
rect 55 3886 170 3901
rect 149 3883 170 3886
rect 188 3883 206 3901
rect 149 3864 206 3883
rect 4419 3914 4570 3937
rect 8454 4034 8605 4057
rect 8563 3998 8605 4034
rect 8890 4029 8951 4045
rect 8795 4025 8951 4029
rect 8795 4007 8913 4025
rect 8931 4007 8951 4025
rect 13261 4120 13318 4139
rect 17432 4191 17588 4212
rect 17432 4190 17532 4191
rect 17433 4154 17475 4190
rect 21462 4261 21523 4277
rect 21891 4247 21952 4263
rect 25939 4334 25981 4370
rect 26180 4362 26222 4398
rect 30209 4469 30270 4485
rect 30638 4455 30699 4471
rect 34686 4542 34728 4578
rect 34629 4541 34729 4542
rect 34573 4520 34729 4541
rect 34573 4502 34593 4520
rect 34611 4502 34729 4520
rect 34573 4498 34729 4502
rect 30543 4451 30699 4455
rect 30207 4423 30264 4442
rect 26180 4339 26331 4362
rect 25882 4333 25982 4334
rect 25826 4312 25982 4333
rect 26180 4324 26295 4339
rect 25826 4294 25846 4312
rect 25864 4294 25982 4312
rect 26274 4321 26295 4324
rect 26313 4321 26331 4339
rect 30207 4405 30225 4423
rect 30243 4420 30264 4423
rect 30543 4433 30661 4451
rect 30679 4433 30699 4451
rect 30243 4405 30358 4420
rect 30543 4412 30699 4433
rect 30543 4411 30643 4412
rect 30207 4382 30358 4405
rect 26274 4302 26331 4321
rect 25826 4290 25982 4294
rect 21796 4243 21952 4247
rect 21796 4225 21914 4243
rect 21932 4225 21952 4243
rect 21796 4204 21952 4225
rect 21796 4203 21896 4204
rect 12831 4087 12888 4106
rect 12831 4069 12849 4087
rect 12867 4084 12888 4087
rect 12867 4069 12982 4084
rect 8506 3997 8606 3998
rect 8450 3976 8606 3997
rect 8795 3986 8951 4007
rect 8795 3985 8895 3986
rect 8450 3958 8470 3976
rect 8488 3958 8606 3976
rect 8450 3954 8606 3958
rect 8450 3938 8511 3954
rect 8796 3949 8838 3985
rect 4419 3899 4534 3914
rect 4513 3896 4534 3899
rect 4552 3896 4570 3914
rect 4513 3877 4570 3896
rect 8796 3926 8947 3949
rect 12831 4046 12982 4069
rect 12940 4010 12982 4046
rect 13254 4042 13315 4058
rect 13159 4038 13315 4042
rect 13159 4020 13277 4038
rect 13295 4020 13315 4038
rect 17433 4131 17584 4154
rect 17195 4100 17252 4119
rect 17433 4116 17548 4131
rect 17195 4082 17213 4100
rect 17231 4097 17252 4100
rect 17527 4113 17548 4116
rect 17566 4113 17584 4131
rect 17231 4082 17346 4097
rect 17527 4094 17584 4113
rect 21797 4167 21839 4203
rect 25826 4274 25887 4290
rect 26268 4259 26329 4275
rect 30316 4346 30358 4382
rect 30544 4375 30586 4411
rect 34573 4482 34634 4498
rect 34571 4436 34628 4455
rect 30544 4352 30695 4375
rect 30259 4345 30359 4346
rect 30203 4324 30359 4345
rect 30544 4337 30659 4352
rect 30203 4306 30223 4324
rect 30241 4306 30359 4324
rect 30638 4334 30659 4337
rect 30677 4334 30695 4352
rect 34571 4418 34589 4436
rect 34607 4433 34628 4436
rect 34607 4418 34722 4433
rect 34571 4395 34722 4418
rect 30638 4315 30695 4334
rect 30203 4302 30359 4306
rect 26173 4255 26329 4259
rect 26173 4237 26291 4255
rect 26309 4237 26329 4255
rect 26173 4216 26329 4237
rect 26173 4215 26273 4216
rect 21797 4144 21948 4167
rect 21797 4129 21912 4144
rect 21891 4126 21912 4129
rect 21930 4126 21948 4144
rect 12883 4009 12983 4010
rect 12827 3988 12983 4009
rect 13159 3999 13315 4020
rect 13159 3998 13259 3999
rect 12827 3970 12847 3988
rect 12865 3970 12983 3988
rect 12827 3966 12983 3970
rect 12827 3950 12888 3966
rect 13160 3962 13202 3998
rect 8796 3911 8911 3926
rect 8890 3908 8911 3911
rect 8929 3908 8947 3926
rect 8890 3889 8947 3908
rect 13160 3939 13311 3962
rect 17195 4059 17346 4082
rect 17304 4023 17346 4059
rect 17247 4022 17347 4023
rect 17191 4001 17347 4022
rect 17520 4016 17581 4032
rect 17191 3983 17211 4001
rect 17229 3983 17347 4001
rect 17191 3979 17347 3983
rect 17425 4012 17581 4016
rect 17425 3994 17543 4012
rect 17561 3994 17581 4012
rect 21891 4107 21948 4126
rect 26174 4179 26216 4215
rect 30203 4286 30264 4302
rect 30632 4272 30693 4288
rect 34680 4359 34722 4395
rect 34623 4358 34723 4359
rect 34567 4337 34723 4358
rect 34567 4319 34587 4337
rect 34605 4319 34723 4337
rect 34567 4315 34723 4319
rect 30537 4268 30693 4272
rect 30537 4250 30655 4268
rect 30673 4250 30693 4268
rect 30537 4229 30693 4250
rect 30537 4228 30637 4229
rect 26174 4156 26325 4179
rect 26174 4141 26289 4156
rect 21461 4074 21518 4093
rect 21461 4056 21479 4074
rect 21497 4071 21518 4074
rect 21497 4056 21612 4071
rect 17191 3963 17252 3979
rect 17425 3973 17581 3994
rect 17425 3972 17525 3973
rect 13160 3924 13275 3939
rect 13254 3921 13275 3924
rect 13293 3921 13311 3939
rect 13254 3902 13311 3921
rect 17426 3936 17468 3972
rect 17426 3913 17577 3936
rect 21461 4033 21612 4056
rect 21570 3997 21612 4033
rect 21884 4029 21945 4045
rect 21789 4025 21945 4029
rect 21789 4007 21907 4025
rect 21925 4007 21945 4025
rect 26268 4138 26289 4141
rect 26307 4138 26325 4156
rect 26268 4119 26325 4138
rect 30538 4192 30580 4228
rect 34567 4299 34628 4315
rect 30538 4169 30689 4192
rect 30538 4154 30653 4169
rect 30632 4151 30653 4154
rect 30671 4151 30689 4169
rect 25825 4087 25882 4106
rect 25825 4069 25843 4087
rect 25861 4084 25882 4087
rect 25861 4069 25976 4084
rect 21513 3996 21613 3997
rect 21457 3975 21613 3996
rect 21789 3986 21945 4007
rect 21789 3985 21889 3986
rect 21457 3957 21477 3975
rect 21495 3957 21613 3975
rect 21457 3953 21613 3957
rect 21457 3937 21518 3953
rect 21790 3949 21832 3985
rect 17426 3898 17541 3913
rect 17520 3895 17541 3898
rect 17559 3895 17577 3913
rect 17520 3876 17577 3895
rect 21790 3926 21941 3949
rect 25825 4046 25976 4069
rect 25934 4010 25976 4046
rect 26261 4041 26322 4057
rect 26166 4037 26322 4041
rect 26166 4019 26284 4037
rect 26302 4019 26322 4037
rect 30632 4132 30689 4151
rect 30202 4099 30259 4118
rect 30202 4081 30220 4099
rect 30238 4096 30259 4099
rect 30238 4081 30353 4096
rect 25877 4009 25977 4010
rect 25821 3988 25977 4009
rect 26166 3998 26322 4019
rect 26166 3997 26266 3998
rect 25821 3970 25841 3988
rect 25859 3970 25977 3988
rect 25821 3966 25977 3970
rect 25821 3950 25882 3966
rect 26167 3961 26209 3997
rect 21790 3911 21905 3926
rect 21884 3908 21905 3911
rect 21923 3908 21941 3926
rect 21884 3889 21941 3908
rect 26167 3938 26318 3961
rect 30202 4058 30353 4081
rect 30311 4022 30353 4058
rect 30625 4054 30686 4070
rect 30530 4050 30686 4054
rect 30530 4032 30648 4050
rect 30666 4032 30686 4050
rect 34566 4112 34623 4131
rect 34566 4094 34584 4112
rect 34602 4109 34623 4112
rect 34602 4094 34717 4109
rect 30254 4021 30354 4022
rect 30198 4000 30354 4021
rect 30530 4011 30686 4032
rect 30530 4010 30630 4011
rect 30198 3982 30218 4000
rect 30236 3982 30354 4000
rect 30198 3978 30354 3982
rect 30198 3962 30259 3978
rect 30531 3974 30573 4010
rect 26167 3923 26282 3938
rect 26261 3920 26282 3923
rect 26300 3920 26318 3938
rect 26261 3901 26318 3920
rect 30531 3951 30682 3974
rect 34566 4071 34717 4094
rect 34675 4035 34717 4071
rect 34618 4034 34718 4035
rect 34562 4013 34718 4034
rect 34562 3995 34582 4013
rect 34600 3995 34718 4013
rect 34562 3991 34718 3995
rect 34562 3975 34623 3991
rect 30531 3936 30646 3951
rect 30625 3933 30646 3936
rect 30664 3933 30682 3951
rect 30625 3914 30682 3933
rect 4091 3769 4148 3788
rect 4091 3751 4109 3769
rect 4127 3766 4148 3769
rect 4127 3751 4242 3766
rect 150 3711 211 3727
rect 55 3707 211 3711
rect 55 3689 173 3707
rect 191 3689 211 3707
rect 55 3668 211 3689
rect 55 3667 155 3668
rect 56 3631 98 3667
rect 56 3608 207 3631
rect 4091 3728 4242 3751
rect 8455 3782 8512 3801
rect 8455 3764 8473 3782
rect 8491 3779 8512 3782
rect 8491 3764 8606 3779
rect 4200 3692 4242 3728
rect 4514 3724 4575 3740
rect 4419 3720 4575 3724
rect 4419 3702 4537 3720
rect 4555 3702 4575 3720
rect 4143 3691 4243 3692
rect 4087 3670 4243 3691
rect 4419 3681 4575 3702
rect 4419 3680 4519 3681
rect 56 3593 171 3608
rect 150 3590 171 3593
rect 189 3590 207 3608
rect 150 3571 207 3590
rect 4087 3652 4107 3670
rect 4125 3652 4243 3670
rect 4087 3648 4243 3652
rect 4087 3632 4148 3648
rect 4420 3644 4462 3680
rect 4420 3621 4571 3644
rect 8455 3741 8606 3764
rect 12832 3794 12889 3813
rect 12832 3776 12850 3794
rect 12868 3791 12889 3794
rect 12868 3776 12983 3791
rect 8564 3705 8606 3741
rect 8891 3736 8952 3752
rect 8796 3732 8952 3736
rect 8796 3714 8914 3732
rect 8932 3714 8952 3732
rect 8507 3704 8607 3705
rect 8451 3683 8607 3704
rect 8796 3693 8952 3714
rect 8796 3692 8896 3693
rect 4420 3606 4535 3621
rect 4514 3603 4535 3606
rect 4553 3603 4571 3621
rect 4514 3584 4571 3603
rect 4084 3551 4141 3570
rect 8451 3665 8471 3683
rect 8489 3665 8607 3683
rect 8451 3661 8607 3665
rect 8451 3645 8512 3661
rect 8797 3656 8839 3692
rect 8797 3633 8948 3656
rect 12832 3753 12983 3776
rect 17196 3807 17253 3826
rect 17196 3789 17214 3807
rect 17232 3804 17253 3807
rect 17232 3789 17347 3804
rect 12941 3717 12983 3753
rect 13255 3749 13316 3765
rect 13160 3745 13316 3749
rect 13160 3727 13278 3745
rect 13296 3727 13316 3745
rect 12884 3716 12984 3717
rect 12828 3695 12984 3716
rect 13160 3706 13316 3727
rect 13160 3705 13260 3706
rect 8797 3618 8912 3633
rect 8891 3615 8912 3618
rect 8930 3615 8948 3633
rect 8891 3596 8948 3615
rect 4084 3533 4102 3551
rect 4120 3548 4141 3551
rect 4120 3533 4235 3548
rect 4084 3510 4235 3533
rect 145 3387 206 3403
rect 4193 3474 4235 3510
rect 8448 3564 8505 3583
rect 8448 3546 8466 3564
rect 8484 3561 8505 3564
rect 12828 3677 12848 3695
rect 12866 3677 12984 3695
rect 12828 3673 12984 3677
rect 12828 3657 12889 3673
rect 13161 3669 13203 3705
rect 13161 3646 13312 3669
rect 17196 3766 17347 3789
rect 17305 3730 17347 3766
rect 21462 3781 21519 3800
rect 21462 3763 21480 3781
rect 21498 3778 21519 3781
rect 21498 3763 21613 3778
rect 17248 3729 17348 3730
rect 17192 3708 17348 3729
rect 17521 3723 17582 3739
rect 13161 3631 13276 3646
rect 13255 3628 13276 3631
rect 13294 3628 13312 3646
rect 13255 3609 13312 3628
rect 8484 3546 8599 3561
rect 8448 3523 8599 3546
rect 4136 3473 4236 3474
rect 4080 3452 4236 3473
rect 4080 3434 4100 3452
rect 4118 3434 4236 3452
rect 4080 3430 4236 3434
rect 50 3383 206 3387
rect 50 3365 168 3383
rect 186 3365 206 3383
rect 50 3344 206 3365
rect 50 3343 150 3344
rect 51 3307 93 3343
rect 4080 3414 4141 3430
rect 4509 3400 4570 3416
rect 8557 3487 8599 3523
rect 12825 3576 12882 3595
rect 17192 3690 17212 3708
rect 17230 3690 17348 3708
rect 17192 3686 17348 3690
rect 17426 3719 17582 3723
rect 17426 3701 17544 3719
rect 17562 3701 17582 3719
rect 17192 3670 17253 3686
rect 17426 3680 17582 3701
rect 17426 3679 17526 3680
rect 17427 3643 17469 3679
rect 17427 3620 17578 3643
rect 21462 3740 21613 3763
rect 25826 3794 25883 3813
rect 25826 3776 25844 3794
rect 25862 3791 25883 3794
rect 25862 3776 25977 3791
rect 21571 3704 21613 3740
rect 21885 3736 21946 3752
rect 21790 3732 21946 3736
rect 21790 3714 21908 3732
rect 21926 3714 21946 3732
rect 21514 3703 21614 3704
rect 21458 3682 21614 3703
rect 21790 3693 21946 3714
rect 21790 3692 21890 3693
rect 12825 3558 12843 3576
rect 12861 3573 12882 3576
rect 12861 3558 12976 3573
rect 12825 3535 12976 3558
rect 8500 3486 8600 3487
rect 8444 3465 8600 3486
rect 8444 3447 8464 3465
rect 8482 3447 8600 3465
rect 8444 3443 8600 3447
rect 4414 3396 4570 3400
rect 4078 3368 4135 3387
rect 51 3284 202 3307
rect 51 3269 166 3284
rect 145 3266 166 3269
rect 184 3266 202 3284
rect 4078 3350 4096 3368
rect 4114 3365 4135 3368
rect 4414 3378 4532 3396
rect 4550 3378 4570 3396
rect 4114 3350 4229 3365
rect 4414 3357 4570 3378
rect 4414 3356 4514 3357
rect 4078 3327 4229 3350
rect 145 3247 202 3266
rect 139 3204 200 3220
rect 4187 3291 4229 3327
rect 4415 3320 4457 3356
rect 8444 3427 8505 3443
rect 8886 3412 8947 3428
rect 12934 3499 12976 3535
rect 17189 3589 17246 3608
rect 17427 3605 17542 3620
rect 17189 3571 17207 3589
rect 17225 3586 17246 3589
rect 17521 3602 17542 3605
rect 17560 3602 17578 3620
rect 17225 3571 17340 3586
rect 17521 3583 17578 3602
rect 17189 3548 17340 3571
rect 21458 3664 21478 3682
rect 21496 3664 21614 3682
rect 21458 3660 21614 3664
rect 21458 3644 21519 3660
rect 21791 3656 21833 3692
rect 21791 3633 21942 3656
rect 25826 3753 25977 3776
rect 30203 3806 30260 3825
rect 30203 3788 30221 3806
rect 30239 3803 30260 3806
rect 30239 3788 30354 3803
rect 25935 3717 25977 3753
rect 26262 3748 26323 3764
rect 26167 3744 26323 3748
rect 26167 3726 26285 3744
rect 26303 3726 26323 3744
rect 25878 3716 25978 3717
rect 25822 3695 25978 3716
rect 26167 3705 26323 3726
rect 26167 3704 26267 3705
rect 21791 3618 21906 3633
rect 21885 3615 21906 3618
rect 21924 3615 21942 3633
rect 21885 3596 21942 3615
rect 12877 3498 12977 3499
rect 12821 3477 12977 3498
rect 12821 3459 12841 3477
rect 12859 3459 12977 3477
rect 12821 3455 12977 3459
rect 8791 3408 8947 3412
rect 8442 3381 8499 3400
rect 4415 3297 4566 3320
rect 4130 3290 4230 3291
rect 4074 3269 4230 3290
rect 4415 3282 4530 3297
rect 4074 3251 4094 3269
rect 4112 3251 4230 3269
rect 4509 3279 4530 3282
rect 4548 3279 4566 3297
rect 8442 3363 8460 3381
rect 8478 3378 8499 3381
rect 8791 3390 8909 3408
rect 8927 3390 8947 3408
rect 8478 3363 8593 3378
rect 8791 3369 8947 3390
rect 8791 3368 8891 3369
rect 8442 3340 8593 3363
rect 4509 3260 4566 3279
rect 4074 3247 4230 3251
rect 44 3200 200 3204
rect 44 3182 162 3200
rect 180 3182 200 3200
rect 44 3161 200 3182
rect 44 3160 144 3161
rect 45 3124 87 3160
rect 4074 3231 4135 3247
rect 4503 3217 4564 3233
rect 8551 3304 8593 3340
rect 8792 3332 8834 3368
rect 12821 3439 12882 3455
rect 13250 3425 13311 3441
rect 17298 3512 17340 3548
rect 17241 3511 17341 3512
rect 17185 3490 17341 3511
rect 21455 3563 21512 3582
rect 25822 3677 25842 3695
rect 25860 3677 25978 3695
rect 25822 3673 25978 3677
rect 25822 3657 25883 3673
rect 26168 3668 26210 3704
rect 26168 3645 26319 3668
rect 30203 3765 30354 3788
rect 34567 3819 34624 3838
rect 34567 3801 34585 3819
rect 34603 3816 34624 3819
rect 34603 3801 34718 3816
rect 30312 3729 30354 3765
rect 30626 3761 30687 3777
rect 30531 3757 30687 3761
rect 30531 3739 30649 3757
rect 30667 3739 30687 3757
rect 30255 3728 30355 3729
rect 30199 3707 30355 3728
rect 30531 3718 30687 3739
rect 30531 3717 30631 3718
rect 26168 3630 26283 3645
rect 26262 3627 26283 3630
rect 26301 3627 26319 3645
rect 26262 3608 26319 3627
rect 21455 3545 21473 3563
rect 21491 3560 21512 3563
rect 21491 3545 21606 3560
rect 21455 3522 21606 3545
rect 17185 3472 17205 3490
rect 17223 3472 17341 3490
rect 17185 3468 17341 3472
rect 13155 3421 13311 3425
rect 12819 3393 12876 3412
rect 8792 3309 8943 3332
rect 8494 3303 8594 3304
rect 8438 3282 8594 3303
rect 8792 3294 8907 3309
rect 8438 3264 8458 3282
rect 8476 3264 8594 3282
rect 8886 3291 8907 3294
rect 8925 3291 8943 3309
rect 12819 3375 12837 3393
rect 12855 3390 12876 3393
rect 13155 3403 13273 3421
rect 13291 3403 13311 3421
rect 12855 3375 12970 3390
rect 13155 3382 13311 3403
rect 13155 3381 13255 3382
rect 12819 3352 12970 3375
rect 8886 3272 8943 3291
rect 8438 3260 8594 3264
rect 4408 3213 4564 3217
rect 4408 3195 4526 3213
rect 4544 3195 4564 3213
rect 4408 3174 4564 3195
rect 4408 3173 4508 3174
rect 45 3101 196 3124
rect 45 3086 160 3101
rect 139 3083 160 3086
rect 178 3083 196 3101
rect 139 3064 196 3083
rect 4409 3137 4451 3173
rect 8438 3244 8499 3260
rect 8880 3229 8941 3245
rect 12928 3316 12970 3352
rect 13156 3345 13198 3381
rect 17185 3452 17246 3468
rect 17183 3406 17240 3425
rect 13156 3322 13307 3345
rect 12871 3315 12971 3316
rect 12815 3294 12971 3315
rect 13156 3307 13271 3322
rect 12815 3276 12835 3294
rect 12853 3276 12971 3294
rect 13250 3304 13271 3307
rect 13289 3304 13307 3322
rect 17183 3388 17201 3406
rect 17219 3403 17240 3406
rect 17219 3388 17334 3403
rect 17516 3399 17577 3415
rect 21564 3486 21606 3522
rect 25819 3576 25876 3595
rect 25819 3558 25837 3576
rect 25855 3573 25876 3576
rect 30199 3689 30219 3707
rect 30237 3689 30355 3707
rect 30199 3685 30355 3689
rect 30199 3669 30260 3685
rect 30532 3681 30574 3717
rect 30532 3658 30683 3681
rect 34567 3778 34718 3801
rect 34676 3742 34718 3778
rect 34619 3741 34719 3742
rect 34563 3720 34719 3741
rect 30532 3643 30647 3658
rect 30626 3640 30647 3643
rect 30665 3640 30683 3658
rect 30626 3621 30683 3640
rect 25855 3558 25970 3573
rect 25819 3535 25970 3558
rect 21507 3485 21607 3486
rect 21451 3464 21607 3485
rect 21451 3446 21471 3464
rect 21489 3446 21607 3464
rect 21451 3442 21607 3446
rect 17183 3365 17334 3388
rect 13250 3285 13307 3304
rect 12815 3272 12971 3276
rect 8785 3225 8941 3229
rect 8785 3207 8903 3225
rect 8921 3207 8941 3225
rect 8785 3186 8941 3207
rect 8785 3185 8885 3186
rect 4409 3114 4560 3137
rect 4409 3099 4524 3114
rect 132 2986 193 3002
rect 37 2982 193 2986
rect 37 2964 155 2982
rect 173 2964 193 2982
rect 4503 3096 4524 3099
rect 4542 3096 4560 3114
rect 4503 3077 4560 3096
rect 8786 3149 8828 3185
rect 12815 3256 12876 3272
rect 13244 3242 13305 3258
rect 17292 3329 17334 3365
rect 17421 3395 17577 3399
rect 17421 3377 17539 3395
rect 17557 3377 17577 3395
rect 17421 3356 17577 3377
rect 17421 3355 17521 3356
rect 17235 3328 17335 3329
rect 17179 3307 17335 3328
rect 17179 3289 17199 3307
rect 17217 3289 17335 3307
rect 17179 3285 17335 3289
rect 17422 3319 17464 3355
rect 21451 3426 21512 3442
rect 21880 3412 21941 3428
rect 25928 3499 25970 3535
rect 30196 3588 30253 3607
rect 34563 3702 34583 3720
rect 34601 3702 34719 3720
rect 34563 3698 34719 3702
rect 34563 3682 34624 3698
rect 30196 3570 30214 3588
rect 30232 3585 30253 3588
rect 30232 3570 30347 3585
rect 30196 3547 30347 3570
rect 25871 3498 25971 3499
rect 25815 3477 25971 3498
rect 25815 3459 25835 3477
rect 25853 3459 25971 3477
rect 25815 3455 25971 3459
rect 21785 3408 21941 3412
rect 21449 3380 21506 3399
rect 17422 3296 17573 3319
rect 13149 3238 13305 3242
rect 13149 3220 13267 3238
rect 13285 3220 13305 3238
rect 13149 3199 13305 3220
rect 13149 3198 13249 3199
rect 8786 3126 8937 3149
rect 8786 3111 8901 3126
rect 4073 3044 4130 3063
rect 4073 3026 4091 3044
rect 4109 3041 4130 3044
rect 4109 3026 4224 3041
rect 37 2943 193 2964
rect 37 2942 137 2943
rect 38 2906 80 2942
rect 38 2883 189 2906
rect 4073 3003 4224 3026
rect 4182 2967 4224 3003
rect 4496 2999 4557 3015
rect 4401 2995 4557 2999
rect 4401 2977 4519 2995
rect 4537 2977 4557 2995
rect 8880 3108 8901 3111
rect 8919 3108 8937 3126
rect 8880 3089 8937 3108
rect 13150 3162 13192 3198
rect 17179 3269 17240 3285
rect 17422 3281 17537 3296
rect 17516 3278 17537 3281
rect 17555 3278 17573 3296
rect 21449 3362 21467 3380
rect 21485 3377 21506 3380
rect 21785 3390 21903 3408
rect 21921 3390 21941 3408
rect 21485 3362 21600 3377
rect 21785 3369 21941 3390
rect 21785 3368 21885 3369
rect 21449 3339 21600 3362
rect 17516 3259 17573 3278
rect 17510 3216 17571 3232
rect 21558 3303 21600 3339
rect 21786 3332 21828 3368
rect 25815 3439 25876 3455
rect 26257 3424 26318 3440
rect 30305 3511 30347 3547
rect 34560 3601 34617 3620
rect 34560 3583 34578 3601
rect 34596 3598 34617 3601
rect 34596 3583 34711 3598
rect 34560 3560 34711 3583
rect 30248 3510 30348 3511
rect 30192 3489 30348 3510
rect 30192 3471 30212 3489
rect 30230 3471 30348 3489
rect 30192 3467 30348 3471
rect 26162 3420 26318 3424
rect 25813 3393 25870 3412
rect 21786 3309 21937 3332
rect 21501 3302 21601 3303
rect 21445 3281 21601 3302
rect 21786 3294 21901 3309
rect 21445 3263 21465 3281
rect 21483 3263 21601 3281
rect 21880 3291 21901 3294
rect 21919 3291 21937 3309
rect 25813 3375 25831 3393
rect 25849 3390 25870 3393
rect 26162 3402 26280 3420
rect 26298 3402 26318 3420
rect 25849 3375 25964 3390
rect 26162 3381 26318 3402
rect 26162 3380 26262 3381
rect 25813 3352 25964 3375
rect 21880 3272 21937 3291
rect 21445 3259 21601 3263
rect 17415 3212 17571 3216
rect 17415 3194 17533 3212
rect 17551 3194 17571 3212
rect 13150 3139 13301 3162
rect 13150 3124 13265 3139
rect 8437 3057 8494 3076
rect 8437 3039 8455 3057
rect 8473 3054 8494 3057
rect 8473 3039 8588 3054
rect 4125 2966 4225 2967
rect 4069 2945 4225 2966
rect 4401 2956 4557 2977
rect 4401 2955 4501 2956
rect 4069 2927 4089 2945
rect 4107 2927 4225 2945
rect 4069 2923 4225 2927
rect 4069 2907 4130 2923
rect 4402 2919 4444 2955
rect 38 2868 153 2883
rect 132 2865 153 2868
rect 171 2865 189 2883
rect 132 2846 189 2865
rect 4402 2896 4553 2919
rect 8437 3016 8588 3039
rect 8546 2980 8588 3016
rect 8873 3011 8934 3027
rect 8778 3007 8934 3011
rect 8778 2989 8896 3007
rect 8914 2989 8934 3007
rect 13244 3121 13265 3124
rect 13283 3121 13301 3139
rect 13244 3102 13301 3121
rect 17415 3173 17571 3194
rect 17415 3172 17515 3173
rect 17416 3136 17458 3172
rect 21445 3243 21506 3259
rect 21874 3229 21935 3245
rect 25922 3316 25964 3352
rect 26163 3344 26205 3380
rect 30192 3451 30253 3467
rect 30621 3437 30682 3453
rect 34669 3524 34711 3560
rect 34612 3523 34712 3524
rect 34556 3502 34712 3523
rect 34556 3484 34576 3502
rect 34594 3484 34712 3502
rect 34556 3480 34712 3484
rect 30526 3433 30682 3437
rect 30190 3405 30247 3424
rect 26163 3321 26314 3344
rect 25865 3315 25965 3316
rect 25809 3294 25965 3315
rect 26163 3306 26278 3321
rect 25809 3276 25829 3294
rect 25847 3276 25965 3294
rect 26257 3303 26278 3306
rect 26296 3303 26314 3321
rect 30190 3387 30208 3405
rect 30226 3402 30247 3405
rect 30526 3415 30644 3433
rect 30662 3415 30682 3433
rect 30226 3387 30341 3402
rect 30526 3394 30682 3415
rect 30526 3393 30626 3394
rect 30190 3364 30341 3387
rect 26257 3284 26314 3303
rect 25809 3272 25965 3276
rect 21779 3225 21935 3229
rect 21779 3207 21897 3225
rect 21915 3207 21935 3225
rect 21779 3186 21935 3207
rect 21779 3185 21879 3186
rect 12814 3069 12871 3088
rect 12814 3051 12832 3069
rect 12850 3066 12871 3069
rect 12850 3051 12965 3066
rect 8489 2979 8589 2980
rect 8433 2958 8589 2979
rect 8778 2968 8934 2989
rect 8778 2967 8878 2968
rect 8433 2940 8453 2958
rect 8471 2940 8589 2958
rect 8433 2936 8589 2940
rect 8433 2920 8494 2936
rect 8779 2931 8821 2967
rect 4402 2881 4517 2896
rect 4496 2878 4517 2881
rect 4535 2878 4553 2896
rect 4496 2859 4553 2878
rect 8779 2908 8930 2931
rect 12814 3028 12965 3051
rect 12923 2992 12965 3028
rect 13237 3024 13298 3040
rect 13142 3020 13298 3024
rect 13142 3002 13260 3020
rect 13278 3002 13298 3020
rect 17416 3113 17567 3136
rect 17178 3082 17235 3101
rect 17416 3098 17531 3113
rect 17178 3064 17196 3082
rect 17214 3079 17235 3082
rect 17510 3095 17531 3098
rect 17549 3095 17567 3113
rect 17214 3064 17329 3079
rect 17510 3076 17567 3095
rect 21780 3149 21822 3185
rect 25809 3256 25870 3272
rect 26251 3241 26312 3257
rect 30299 3328 30341 3364
rect 30527 3357 30569 3393
rect 34556 3464 34617 3480
rect 34554 3418 34611 3437
rect 30527 3334 30678 3357
rect 30242 3327 30342 3328
rect 30186 3306 30342 3327
rect 30527 3319 30642 3334
rect 30186 3288 30206 3306
rect 30224 3288 30342 3306
rect 30621 3316 30642 3319
rect 30660 3316 30678 3334
rect 34554 3400 34572 3418
rect 34590 3415 34611 3418
rect 34590 3400 34705 3415
rect 34554 3377 34705 3400
rect 30621 3297 30678 3316
rect 30186 3284 30342 3288
rect 26156 3237 26312 3241
rect 26156 3219 26274 3237
rect 26292 3219 26312 3237
rect 26156 3198 26312 3219
rect 26156 3197 26256 3198
rect 21780 3126 21931 3149
rect 21780 3111 21895 3126
rect 12866 2991 12966 2992
rect 12810 2970 12966 2991
rect 13142 2981 13298 3002
rect 13142 2980 13242 2981
rect 12810 2952 12830 2970
rect 12848 2952 12966 2970
rect 12810 2948 12966 2952
rect 12810 2932 12871 2948
rect 13143 2944 13185 2980
rect 8779 2893 8894 2908
rect 8873 2890 8894 2893
rect 8912 2890 8930 2908
rect 8873 2871 8930 2890
rect 13143 2921 13294 2944
rect 17178 3041 17329 3064
rect 17287 3005 17329 3041
rect 17230 3004 17330 3005
rect 17174 2983 17330 3004
rect 17503 2998 17564 3014
rect 17174 2965 17194 2983
rect 17212 2965 17330 2983
rect 17174 2961 17330 2965
rect 17408 2994 17564 2998
rect 17408 2976 17526 2994
rect 17544 2976 17564 2994
rect 21874 3108 21895 3111
rect 21913 3108 21931 3126
rect 21874 3089 21931 3108
rect 26157 3161 26199 3197
rect 30186 3268 30247 3284
rect 30615 3254 30676 3270
rect 34663 3341 34705 3377
rect 34606 3340 34706 3341
rect 34550 3319 34706 3340
rect 34550 3301 34570 3319
rect 34588 3301 34706 3319
rect 34550 3297 34706 3301
rect 30520 3250 30676 3254
rect 30520 3232 30638 3250
rect 30656 3232 30676 3250
rect 30520 3211 30676 3232
rect 30520 3210 30620 3211
rect 26157 3138 26308 3161
rect 26157 3123 26272 3138
rect 21444 3056 21501 3075
rect 21444 3038 21462 3056
rect 21480 3053 21501 3056
rect 21480 3038 21595 3053
rect 17174 2945 17235 2961
rect 17408 2955 17564 2976
rect 17408 2954 17508 2955
rect 13143 2906 13258 2921
rect 13237 2903 13258 2906
rect 13276 2903 13294 2921
rect 13237 2884 13294 2903
rect 17409 2918 17451 2954
rect 17409 2895 17560 2918
rect 21444 3015 21595 3038
rect 21553 2979 21595 3015
rect 21867 3011 21928 3027
rect 21772 3007 21928 3011
rect 21772 2989 21890 3007
rect 21908 2989 21928 3007
rect 26251 3120 26272 3123
rect 26290 3120 26308 3138
rect 26251 3101 26308 3120
rect 30521 3174 30563 3210
rect 34550 3281 34611 3297
rect 30521 3151 30672 3174
rect 30521 3136 30636 3151
rect 25808 3069 25865 3088
rect 25808 3051 25826 3069
rect 25844 3066 25865 3069
rect 25844 3051 25959 3066
rect 21496 2978 21596 2979
rect 21440 2957 21596 2978
rect 21772 2968 21928 2989
rect 21772 2967 21872 2968
rect 21440 2939 21460 2957
rect 21478 2939 21596 2957
rect 21440 2935 21596 2939
rect 21440 2919 21501 2935
rect 21773 2931 21815 2967
rect 17409 2880 17524 2895
rect 17503 2877 17524 2880
rect 17542 2877 17560 2895
rect 17503 2858 17560 2877
rect 21773 2908 21924 2931
rect 25808 3028 25959 3051
rect 25917 2992 25959 3028
rect 26244 3023 26305 3039
rect 26149 3019 26305 3023
rect 26149 3001 26267 3019
rect 26285 3001 26305 3019
rect 30615 3133 30636 3136
rect 30654 3133 30672 3151
rect 30615 3114 30672 3133
rect 30185 3081 30242 3100
rect 30185 3063 30203 3081
rect 30221 3078 30242 3081
rect 30221 3063 30336 3078
rect 25860 2991 25960 2992
rect 25804 2970 25960 2991
rect 26149 2980 26305 3001
rect 26149 2979 26249 2980
rect 25804 2952 25824 2970
rect 25842 2952 25960 2970
rect 25804 2948 25960 2952
rect 25804 2932 25865 2948
rect 26150 2943 26192 2979
rect 21773 2893 21888 2908
rect 21867 2890 21888 2893
rect 21906 2890 21924 2908
rect 21867 2871 21924 2890
rect 26150 2920 26301 2943
rect 30185 3040 30336 3063
rect 30294 3004 30336 3040
rect 30608 3036 30669 3052
rect 30513 3032 30669 3036
rect 30513 3014 30631 3032
rect 30649 3014 30669 3032
rect 34549 3094 34606 3113
rect 34549 3076 34567 3094
rect 34585 3091 34606 3094
rect 34585 3076 34700 3091
rect 30237 3003 30337 3004
rect 30181 2982 30337 3003
rect 30513 2993 30669 3014
rect 30513 2992 30613 2993
rect 30181 2964 30201 2982
rect 30219 2964 30337 2982
rect 30181 2960 30337 2964
rect 30181 2944 30242 2960
rect 30514 2956 30556 2992
rect 26150 2905 26265 2920
rect 26244 2902 26265 2905
rect 26283 2902 26301 2920
rect 26244 2883 26301 2902
rect 30514 2933 30665 2956
rect 34549 3053 34700 3076
rect 34658 3017 34700 3053
rect 34601 3016 34701 3017
rect 34545 2995 34701 3016
rect 34545 2977 34565 2995
rect 34583 2977 34701 2995
rect 34545 2973 34701 2977
rect 34545 2957 34606 2973
rect 30514 2918 30629 2933
rect 30608 2915 30629 2918
rect 30647 2915 30665 2933
rect 30608 2896 30665 2915
rect 4071 2751 4128 2770
rect 4071 2733 4089 2751
rect 4107 2748 4128 2751
rect 4107 2733 4222 2748
rect 130 2693 191 2709
rect 35 2689 191 2693
rect 35 2671 153 2689
rect 171 2671 191 2689
rect 35 2650 191 2671
rect 35 2649 135 2650
rect 36 2613 78 2649
rect 36 2590 187 2613
rect 4071 2710 4222 2733
rect 8435 2764 8492 2783
rect 8435 2746 8453 2764
rect 8471 2761 8492 2764
rect 8471 2746 8586 2761
rect 4180 2674 4222 2710
rect 4494 2706 4555 2722
rect 4399 2702 4555 2706
rect 4399 2684 4517 2702
rect 4535 2684 4555 2702
rect 4123 2673 4223 2674
rect 4067 2652 4223 2673
rect 4399 2663 4555 2684
rect 4399 2662 4499 2663
rect 36 2575 151 2590
rect 130 2572 151 2575
rect 169 2572 187 2590
rect 130 2553 187 2572
rect 4067 2634 4087 2652
rect 4105 2634 4223 2652
rect 4067 2630 4223 2634
rect 4067 2614 4128 2630
rect 4400 2626 4442 2662
rect 4400 2603 4551 2626
rect 8435 2723 8586 2746
rect 12812 2776 12869 2795
rect 12812 2758 12830 2776
rect 12848 2773 12869 2776
rect 12848 2758 12963 2773
rect 8544 2687 8586 2723
rect 8871 2718 8932 2734
rect 8776 2714 8932 2718
rect 8776 2696 8894 2714
rect 8912 2696 8932 2714
rect 8487 2686 8587 2687
rect 8431 2665 8587 2686
rect 8776 2675 8932 2696
rect 8776 2674 8876 2675
rect 4400 2588 4515 2603
rect 4494 2585 4515 2588
rect 4533 2585 4551 2603
rect 4494 2566 4551 2585
rect 4064 2533 4121 2552
rect 4064 2515 4082 2533
rect 4100 2530 4121 2533
rect 8431 2647 8451 2665
rect 8469 2647 8587 2665
rect 8431 2643 8587 2647
rect 8431 2627 8492 2643
rect 8777 2638 8819 2674
rect 8777 2615 8928 2638
rect 12812 2735 12963 2758
rect 17176 2789 17233 2808
rect 17176 2771 17194 2789
rect 17212 2786 17233 2789
rect 17212 2771 17327 2786
rect 12921 2699 12963 2735
rect 13235 2731 13296 2747
rect 13140 2727 13296 2731
rect 13140 2709 13258 2727
rect 13276 2709 13296 2727
rect 12864 2698 12964 2699
rect 12808 2677 12964 2698
rect 13140 2688 13296 2709
rect 13140 2687 13240 2688
rect 8777 2600 8892 2615
rect 8871 2597 8892 2600
rect 8910 2597 8928 2615
rect 8871 2578 8928 2597
rect 4100 2515 4215 2530
rect 4064 2492 4215 2515
rect 125 2369 186 2385
rect 4173 2456 4215 2492
rect 8428 2546 8485 2565
rect 8428 2528 8446 2546
rect 8464 2543 8485 2546
rect 12808 2659 12828 2677
rect 12846 2659 12964 2677
rect 12808 2655 12964 2659
rect 12808 2639 12869 2655
rect 13141 2651 13183 2687
rect 13141 2628 13292 2651
rect 17176 2748 17327 2771
rect 17285 2712 17327 2748
rect 21442 2763 21499 2782
rect 21442 2745 21460 2763
rect 21478 2760 21499 2763
rect 21478 2745 21593 2760
rect 17228 2711 17328 2712
rect 17172 2690 17328 2711
rect 17501 2705 17562 2721
rect 13141 2613 13256 2628
rect 13235 2610 13256 2613
rect 13274 2610 13292 2628
rect 13235 2591 13292 2610
rect 8464 2528 8579 2543
rect 8428 2505 8579 2528
rect 4116 2455 4216 2456
rect 4060 2434 4216 2455
rect 4060 2416 4080 2434
rect 4098 2416 4216 2434
rect 4060 2412 4216 2416
rect 30 2365 186 2369
rect 30 2347 148 2365
rect 166 2347 186 2365
rect 30 2326 186 2347
rect 30 2325 130 2326
rect 31 2289 73 2325
rect 4060 2396 4121 2412
rect 4489 2382 4550 2398
rect 8537 2469 8579 2505
rect 12805 2558 12862 2577
rect 12805 2540 12823 2558
rect 12841 2555 12862 2558
rect 17172 2672 17192 2690
rect 17210 2672 17328 2690
rect 17172 2668 17328 2672
rect 17406 2701 17562 2705
rect 17406 2683 17524 2701
rect 17542 2683 17562 2701
rect 17172 2652 17233 2668
rect 17406 2662 17562 2683
rect 17406 2661 17506 2662
rect 17407 2625 17449 2661
rect 17407 2602 17558 2625
rect 21442 2722 21593 2745
rect 25806 2776 25863 2795
rect 25806 2758 25824 2776
rect 25842 2773 25863 2776
rect 25842 2758 25957 2773
rect 21551 2686 21593 2722
rect 21865 2718 21926 2734
rect 21770 2714 21926 2718
rect 21770 2696 21888 2714
rect 21906 2696 21926 2714
rect 21494 2685 21594 2686
rect 21438 2664 21594 2685
rect 21770 2675 21926 2696
rect 21770 2674 21870 2675
rect 12841 2540 12956 2555
rect 12805 2517 12956 2540
rect 8480 2468 8580 2469
rect 8424 2447 8580 2468
rect 8424 2429 8444 2447
rect 8462 2429 8580 2447
rect 8424 2425 8580 2429
rect 4394 2378 4550 2382
rect 4058 2350 4115 2369
rect 31 2266 182 2289
rect 31 2251 146 2266
rect 125 2248 146 2251
rect 164 2248 182 2266
rect 4058 2332 4076 2350
rect 4094 2347 4115 2350
rect 4394 2360 4512 2378
rect 4530 2360 4550 2378
rect 4094 2332 4209 2347
rect 4394 2339 4550 2360
rect 4394 2338 4494 2339
rect 4058 2309 4209 2332
rect 125 2229 182 2248
rect 119 2186 180 2202
rect 4167 2273 4209 2309
rect 4395 2302 4437 2338
rect 8424 2409 8485 2425
rect 8866 2394 8927 2410
rect 12914 2481 12956 2517
rect 17169 2571 17226 2590
rect 17407 2587 17522 2602
rect 17169 2553 17187 2571
rect 17205 2568 17226 2571
rect 17501 2584 17522 2587
rect 17540 2584 17558 2602
rect 17205 2553 17320 2568
rect 17501 2565 17558 2584
rect 17169 2530 17320 2553
rect 21438 2646 21458 2664
rect 21476 2646 21594 2664
rect 21438 2642 21594 2646
rect 21438 2626 21499 2642
rect 21771 2638 21813 2674
rect 21771 2615 21922 2638
rect 25806 2735 25957 2758
rect 30183 2788 30240 2807
rect 30183 2770 30201 2788
rect 30219 2785 30240 2788
rect 30219 2770 30334 2785
rect 25915 2699 25957 2735
rect 26242 2730 26303 2746
rect 26147 2726 26303 2730
rect 26147 2708 26265 2726
rect 26283 2708 26303 2726
rect 25858 2698 25958 2699
rect 25802 2677 25958 2698
rect 26147 2687 26303 2708
rect 26147 2686 26247 2687
rect 21771 2600 21886 2615
rect 21865 2597 21886 2600
rect 21904 2597 21922 2615
rect 21865 2578 21922 2597
rect 12857 2480 12957 2481
rect 12801 2459 12957 2480
rect 12801 2441 12821 2459
rect 12839 2441 12957 2459
rect 12801 2437 12957 2441
rect 8771 2390 8927 2394
rect 8422 2363 8479 2382
rect 4395 2279 4546 2302
rect 4110 2272 4210 2273
rect 4054 2251 4210 2272
rect 4395 2264 4510 2279
rect 4054 2233 4074 2251
rect 4092 2233 4210 2251
rect 4489 2261 4510 2264
rect 4528 2261 4546 2279
rect 8422 2345 8440 2363
rect 8458 2360 8479 2363
rect 8771 2372 8889 2390
rect 8907 2372 8927 2390
rect 8458 2345 8573 2360
rect 8771 2351 8927 2372
rect 8771 2350 8871 2351
rect 8422 2322 8573 2345
rect 4489 2242 4546 2261
rect 4054 2229 4210 2233
rect 24 2182 180 2186
rect 24 2164 142 2182
rect 160 2164 180 2182
rect 24 2143 180 2164
rect 24 2142 124 2143
rect 25 2106 67 2142
rect 4054 2213 4115 2229
rect 4483 2199 4544 2215
rect 8531 2286 8573 2322
rect 8772 2314 8814 2350
rect 12801 2421 12862 2437
rect 13230 2407 13291 2423
rect 17278 2494 17320 2530
rect 17221 2493 17321 2494
rect 17165 2472 17321 2493
rect 21435 2545 21492 2564
rect 21435 2527 21453 2545
rect 21471 2542 21492 2545
rect 25802 2659 25822 2677
rect 25840 2659 25958 2677
rect 25802 2655 25958 2659
rect 25802 2639 25863 2655
rect 26148 2650 26190 2686
rect 26148 2627 26299 2650
rect 30183 2747 30334 2770
rect 34547 2801 34604 2820
rect 34547 2783 34565 2801
rect 34583 2798 34604 2801
rect 34583 2783 34698 2798
rect 30292 2711 30334 2747
rect 30606 2743 30667 2759
rect 30511 2739 30667 2743
rect 30511 2721 30629 2739
rect 30647 2721 30667 2739
rect 30235 2710 30335 2711
rect 30179 2689 30335 2710
rect 30511 2700 30667 2721
rect 30511 2699 30611 2700
rect 26148 2612 26263 2627
rect 26242 2609 26263 2612
rect 26281 2609 26299 2627
rect 26242 2590 26299 2609
rect 21471 2527 21586 2542
rect 21435 2504 21586 2527
rect 17165 2454 17185 2472
rect 17203 2454 17321 2472
rect 17165 2450 17321 2454
rect 13135 2403 13291 2407
rect 12799 2375 12856 2394
rect 8772 2291 8923 2314
rect 8474 2285 8574 2286
rect 8418 2264 8574 2285
rect 8772 2276 8887 2291
rect 8418 2246 8438 2264
rect 8456 2246 8574 2264
rect 8866 2273 8887 2276
rect 8905 2273 8923 2291
rect 12799 2357 12817 2375
rect 12835 2372 12856 2375
rect 13135 2385 13253 2403
rect 13271 2385 13291 2403
rect 12835 2357 12950 2372
rect 13135 2364 13291 2385
rect 13135 2363 13235 2364
rect 12799 2334 12950 2357
rect 8866 2254 8923 2273
rect 8418 2242 8574 2246
rect 4388 2195 4544 2199
rect 4388 2177 4506 2195
rect 4524 2177 4544 2195
rect 4388 2156 4544 2177
rect 4388 2155 4488 2156
rect 25 2083 176 2106
rect 25 2068 140 2083
rect 119 2065 140 2068
rect 158 2065 176 2083
rect 119 2046 176 2065
rect 4389 2119 4431 2155
rect 8418 2226 8479 2242
rect 8860 2211 8921 2227
rect 12908 2298 12950 2334
rect 13136 2327 13178 2363
rect 17165 2434 17226 2450
rect 17163 2388 17220 2407
rect 13136 2304 13287 2327
rect 12851 2297 12951 2298
rect 12795 2276 12951 2297
rect 13136 2289 13251 2304
rect 12795 2258 12815 2276
rect 12833 2258 12951 2276
rect 13230 2286 13251 2289
rect 13269 2286 13287 2304
rect 17163 2370 17181 2388
rect 17199 2385 17220 2388
rect 17199 2370 17314 2385
rect 17496 2381 17557 2397
rect 21544 2468 21586 2504
rect 25799 2558 25856 2577
rect 25799 2540 25817 2558
rect 25835 2555 25856 2558
rect 30179 2671 30199 2689
rect 30217 2671 30335 2689
rect 30179 2667 30335 2671
rect 30179 2651 30240 2667
rect 30512 2663 30554 2699
rect 30512 2640 30663 2663
rect 34547 2760 34698 2783
rect 34656 2724 34698 2760
rect 34599 2723 34699 2724
rect 34543 2702 34699 2723
rect 30512 2625 30627 2640
rect 30606 2622 30627 2625
rect 30645 2622 30663 2640
rect 30606 2603 30663 2622
rect 25835 2540 25950 2555
rect 25799 2517 25950 2540
rect 21487 2467 21587 2468
rect 21431 2446 21587 2467
rect 21431 2428 21451 2446
rect 21469 2428 21587 2446
rect 21431 2424 21587 2428
rect 17163 2347 17314 2370
rect 13230 2267 13287 2286
rect 12795 2254 12951 2258
rect 8765 2207 8921 2211
rect 8765 2189 8883 2207
rect 8901 2189 8921 2207
rect 8765 2168 8921 2189
rect 8765 2167 8865 2168
rect 4389 2096 4540 2119
rect 4389 2081 4504 2096
rect 4483 2078 4504 2081
rect 4522 2078 4540 2096
rect 112 1968 173 1984
rect 17 1964 173 1968
rect 17 1946 135 1964
rect 153 1946 173 1964
rect 4483 2059 4540 2078
rect 8766 2131 8808 2167
rect 12795 2238 12856 2254
rect 13224 2224 13285 2240
rect 17272 2311 17314 2347
rect 17401 2377 17557 2381
rect 17401 2359 17519 2377
rect 17537 2359 17557 2377
rect 17401 2338 17557 2359
rect 17401 2337 17501 2338
rect 17215 2310 17315 2311
rect 17159 2289 17315 2310
rect 17159 2271 17179 2289
rect 17197 2271 17315 2289
rect 17159 2267 17315 2271
rect 17402 2301 17444 2337
rect 21431 2408 21492 2424
rect 21860 2394 21921 2410
rect 25908 2481 25950 2517
rect 30176 2570 30233 2589
rect 30176 2552 30194 2570
rect 30212 2567 30233 2570
rect 34543 2684 34563 2702
rect 34581 2684 34699 2702
rect 34543 2680 34699 2684
rect 34543 2664 34604 2680
rect 30212 2552 30327 2567
rect 30176 2529 30327 2552
rect 25851 2480 25951 2481
rect 25795 2459 25951 2480
rect 25795 2441 25815 2459
rect 25833 2441 25951 2459
rect 25795 2437 25951 2441
rect 21765 2390 21921 2394
rect 21429 2362 21486 2381
rect 17402 2278 17553 2301
rect 13129 2220 13285 2224
rect 13129 2202 13247 2220
rect 13265 2202 13285 2220
rect 13129 2181 13285 2202
rect 13129 2180 13229 2181
rect 8766 2108 8917 2131
rect 8766 2093 8881 2108
rect 4053 2026 4110 2045
rect 4053 2008 4071 2026
rect 4089 2023 4110 2026
rect 4089 2008 4204 2023
rect 17 1925 173 1946
rect 17 1924 117 1925
rect 18 1888 60 1924
rect 18 1865 169 1888
rect 4053 1985 4204 2008
rect 4162 1949 4204 1985
rect 4476 1981 4537 1997
rect 4381 1977 4537 1981
rect 4381 1959 4499 1977
rect 4517 1959 4537 1977
rect 8860 2090 8881 2093
rect 8899 2090 8917 2108
rect 8860 2071 8917 2090
rect 13130 2144 13172 2180
rect 17159 2251 17220 2267
rect 17402 2263 17517 2278
rect 17496 2260 17517 2263
rect 17535 2260 17553 2278
rect 21429 2344 21447 2362
rect 21465 2359 21486 2362
rect 21765 2372 21883 2390
rect 21901 2372 21921 2390
rect 21465 2344 21580 2359
rect 21765 2351 21921 2372
rect 21765 2350 21865 2351
rect 21429 2321 21580 2344
rect 17496 2241 17553 2260
rect 17490 2198 17551 2214
rect 21538 2285 21580 2321
rect 21766 2314 21808 2350
rect 25795 2421 25856 2437
rect 26237 2406 26298 2422
rect 30285 2493 30327 2529
rect 34540 2583 34597 2602
rect 34540 2565 34558 2583
rect 34576 2580 34597 2583
rect 34576 2565 34691 2580
rect 34540 2542 34691 2565
rect 30228 2492 30328 2493
rect 30172 2471 30328 2492
rect 30172 2453 30192 2471
rect 30210 2453 30328 2471
rect 30172 2449 30328 2453
rect 26142 2402 26298 2406
rect 25793 2375 25850 2394
rect 21766 2291 21917 2314
rect 21481 2284 21581 2285
rect 21425 2263 21581 2284
rect 21766 2276 21881 2291
rect 21425 2245 21445 2263
rect 21463 2245 21581 2263
rect 21860 2273 21881 2276
rect 21899 2273 21917 2291
rect 25793 2357 25811 2375
rect 25829 2372 25850 2375
rect 26142 2384 26260 2402
rect 26278 2384 26298 2402
rect 25829 2357 25944 2372
rect 26142 2363 26298 2384
rect 26142 2362 26242 2363
rect 25793 2334 25944 2357
rect 21860 2254 21917 2273
rect 21425 2241 21581 2245
rect 17395 2194 17551 2198
rect 17395 2176 17513 2194
rect 17531 2176 17551 2194
rect 13130 2121 13281 2144
rect 13130 2106 13245 2121
rect 13224 2103 13245 2106
rect 13263 2103 13281 2121
rect 8417 2039 8474 2058
rect 8417 2021 8435 2039
rect 8453 2036 8474 2039
rect 8453 2021 8568 2036
rect 4105 1948 4205 1949
rect 4049 1927 4205 1948
rect 4381 1938 4537 1959
rect 4381 1937 4481 1938
rect 4049 1909 4069 1927
rect 4087 1909 4205 1927
rect 4049 1905 4205 1909
rect 4049 1889 4110 1905
rect 4382 1901 4424 1937
rect 18 1850 133 1865
rect 112 1847 133 1850
rect 151 1847 169 1865
rect 112 1828 169 1847
rect 4382 1878 4533 1901
rect 8417 1998 8568 2021
rect 8526 1962 8568 1998
rect 8853 1993 8914 2009
rect 8758 1989 8914 1993
rect 8758 1971 8876 1989
rect 8894 1971 8914 1989
rect 13224 2084 13281 2103
rect 17395 2155 17551 2176
rect 17395 2154 17495 2155
rect 17396 2118 17438 2154
rect 21425 2225 21486 2241
rect 21854 2211 21915 2227
rect 25902 2298 25944 2334
rect 26143 2326 26185 2362
rect 30172 2433 30233 2449
rect 30601 2419 30662 2435
rect 34649 2506 34691 2542
rect 34592 2505 34692 2506
rect 34536 2484 34692 2505
rect 34536 2466 34556 2484
rect 34574 2466 34692 2484
rect 34536 2462 34692 2466
rect 30506 2415 30662 2419
rect 30170 2387 30227 2406
rect 26143 2303 26294 2326
rect 25845 2297 25945 2298
rect 25789 2276 25945 2297
rect 26143 2288 26258 2303
rect 25789 2258 25809 2276
rect 25827 2258 25945 2276
rect 26237 2285 26258 2288
rect 26276 2285 26294 2303
rect 30170 2369 30188 2387
rect 30206 2384 30227 2387
rect 30506 2397 30624 2415
rect 30642 2397 30662 2415
rect 30206 2369 30321 2384
rect 30506 2376 30662 2397
rect 30506 2375 30606 2376
rect 30170 2346 30321 2369
rect 26237 2266 26294 2285
rect 25789 2254 25945 2258
rect 21759 2207 21915 2211
rect 21759 2189 21877 2207
rect 21895 2189 21915 2207
rect 21759 2168 21915 2189
rect 21759 2167 21859 2168
rect 12794 2051 12851 2070
rect 12794 2033 12812 2051
rect 12830 2048 12851 2051
rect 12830 2033 12945 2048
rect 8469 1961 8569 1962
rect 8413 1940 8569 1961
rect 8758 1950 8914 1971
rect 8758 1949 8858 1950
rect 8413 1922 8433 1940
rect 8451 1922 8569 1940
rect 8413 1918 8569 1922
rect 8413 1902 8474 1918
rect 8759 1913 8801 1949
rect 4382 1863 4497 1878
rect 4476 1860 4497 1863
rect 4515 1860 4533 1878
rect 4476 1841 4533 1860
rect 8759 1890 8910 1913
rect 12794 2010 12945 2033
rect 12903 1974 12945 2010
rect 13217 2006 13278 2022
rect 13122 2002 13278 2006
rect 13122 1984 13240 2002
rect 13258 1984 13278 2002
rect 17396 2095 17547 2118
rect 17158 2064 17215 2083
rect 17396 2080 17511 2095
rect 17158 2046 17176 2064
rect 17194 2061 17215 2064
rect 17490 2077 17511 2080
rect 17529 2077 17547 2095
rect 17194 2046 17309 2061
rect 17490 2058 17547 2077
rect 21760 2131 21802 2167
rect 25789 2238 25850 2254
rect 26231 2223 26292 2239
rect 30279 2310 30321 2346
rect 30507 2339 30549 2375
rect 34536 2446 34597 2462
rect 34534 2400 34591 2419
rect 30507 2316 30658 2339
rect 30222 2309 30322 2310
rect 30166 2288 30322 2309
rect 30507 2301 30622 2316
rect 30166 2270 30186 2288
rect 30204 2270 30322 2288
rect 30601 2298 30622 2301
rect 30640 2298 30658 2316
rect 34534 2382 34552 2400
rect 34570 2397 34591 2400
rect 34570 2382 34685 2397
rect 34534 2359 34685 2382
rect 30601 2279 30658 2298
rect 30166 2266 30322 2270
rect 26136 2219 26292 2223
rect 26136 2201 26254 2219
rect 26272 2201 26292 2219
rect 26136 2180 26292 2201
rect 26136 2179 26236 2180
rect 21760 2108 21911 2131
rect 21760 2093 21875 2108
rect 21854 2090 21875 2093
rect 21893 2090 21911 2108
rect 12846 1973 12946 1974
rect 12790 1952 12946 1973
rect 13122 1963 13278 1984
rect 13122 1962 13222 1963
rect 12790 1934 12810 1952
rect 12828 1934 12946 1952
rect 12790 1930 12946 1934
rect 12790 1914 12851 1930
rect 13123 1926 13165 1962
rect 8759 1875 8874 1890
rect 8853 1872 8874 1875
rect 8892 1872 8910 1890
rect 8853 1853 8910 1872
rect 13123 1903 13274 1926
rect 17158 2023 17309 2046
rect 17267 1987 17309 2023
rect 17210 1986 17310 1987
rect 17154 1965 17310 1986
rect 17483 1980 17544 1996
rect 17154 1947 17174 1965
rect 17192 1947 17310 1965
rect 17154 1943 17310 1947
rect 17388 1976 17544 1980
rect 17388 1958 17506 1976
rect 17524 1958 17544 1976
rect 21854 2071 21911 2090
rect 26137 2143 26179 2179
rect 30166 2250 30227 2266
rect 30595 2236 30656 2252
rect 34643 2323 34685 2359
rect 34586 2322 34686 2323
rect 34530 2301 34686 2322
rect 34530 2283 34550 2301
rect 34568 2283 34686 2301
rect 34530 2279 34686 2283
rect 30500 2232 30656 2236
rect 30500 2214 30618 2232
rect 30636 2214 30656 2232
rect 30500 2193 30656 2214
rect 30500 2192 30600 2193
rect 26137 2120 26288 2143
rect 26137 2105 26252 2120
rect 21424 2038 21481 2057
rect 21424 2020 21442 2038
rect 21460 2035 21481 2038
rect 21460 2020 21575 2035
rect 17154 1927 17215 1943
rect 17388 1937 17544 1958
rect 17388 1936 17488 1937
rect 13123 1888 13238 1903
rect 13217 1885 13238 1888
rect 13256 1885 13274 1903
rect 13217 1866 13274 1885
rect 17389 1900 17431 1936
rect 17389 1877 17540 1900
rect 21424 1997 21575 2020
rect 21533 1961 21575 1997
rect 21847 1993 21908 2009
rect 21752 1989 21908 1993
rect 21752 1971 21870 1989
rect 21888 1971 21908 1989
rect 26231 2102 26252 2105
rect 26270 2102 26288 2120
rect 26231 2083 26288 2102
rect 30501 2156 30543 2192
rect 34530 2263 34591 2279
rect 30501 2133 30652 2156
rect 30501 2118 30616 2133
rect 30595 2115 30616 2118
rect 30634 2115 30652 2133
rect 25788 2051 25845 2070
rect 25788 2033 25806 2051
rect 25824 2048 25845 2051
rect 25824 2033 25939 2048
rect 21476 1960 21576 1961
rect 21420 1939 21576 1960
rect 21752 1950 21908 1971
rect 21752 1949 21852 1950
rect 21420 1921 21440 1939
rect 21458 1921 21576 1939
rect 21420 1917 21576 1921
rect 21420 1901 21481 1917
rect 21753 1913 21795 1949
rect 17389 1862 17504 1877
rect 17483 1859 17504 1862
rect 17522 1859 17540 1877
rect 17483 1840 17540 1859
rect 21753 1890 21904 1913
rect 25788 2010 25939 2033
rect 25897 1974 25939 2010
rect 26224 2005 26285 2021
rect 26129 2001 26285 2005
rect 26129 1983 26247 2001
rect 26265 1983 26285 2001
rect 30595 2096 30652 2115
rect 30165 2063 30222 2082
rect 30165 2045 30183 2063
rect 30201 2060 30222 2063
rect 30201 2045 30316 2060
rect 25840 1973 25940 1974
rect 25784 1952 25940 1973
rect 26129 1962 26285 1983
rect 26129 1961 26229 1962
rect 25784 1934 25804 1952
rect 25822 1934 25940 1952
rect 25784 1930 25940 1934
rect 25784 1914 25845 1930
rect 26130 1925 26172 1961
rect 21753 1875 21868 1890
rect 21847 1872 21868 1875
rect 21886 1872 21904 1890
rect 21847 1853 21904 1872
rect 26130 1902 26281 1925
rect 30165 2022 30316 2045
rect 30274 1986 30316 2022
rect 30588 2018 30649 2034
rect 30493 2014 30649 2018
rect 30493 1996 30611 2014
rect 30629 1996 30649 2014
rect 34529 2076 34586 2095
rect 34529 2058 34547 2076
rect 34565 2073 34586 2076
rect 34565 2058 34680 2073
rect 30217 1985 30317 1986
rect 30161 1964 30317 1985
rect 30493 1975 30649 1996
rect 30493 1974 30593 1975
rect 30161 1946 30181 1964
rect 30199 1946 30317 1964
rect 30161 1942 30317 1946
rect 30161 1926 30222 1942
rect 30494 1938 30536 1974
rect 26130 1887 26245 1902
rect 26224 1884 26245 1887
rect 26263 1884 26281 1902
rect 26224 1865 26281 1884
rect 30494 1915 30645 1938
rect 34529 2035 34680 2058
rect 34638 1999 34680 2035
rect 34581 1998 34681 1999
rect 34525 1977 34681 1998
rect 34525 1959 34545 1977
rect 34563 1959 34681 1977
rect 34525 1955 34681 1959
rect 34525 1939 34586 1955
rect 30494 1900 30609 1915
rect 30588 1897 30609 1900
rect 30627 1897 30645 1915
rect 30588 1878 30645 1897
rect 4054 1733 4111 1752
rect 4054 1715 4072 1733
rect 4090 1730 4111 1733
rect 4090 1715 4205 1730
rect 113 1675 174 1691
rect 18 1671 174 1675
rect 18 1653 136 1671
rect 154 1653 174 1671
rect 18 1632 174 1653
rect 18 1631 118 1632
rect 19 1595 61 1631
rect 19 1572 170 1595
rect 4054 1692 4205 1715
rect 8418 1746 8475 1765
rect 8418 1728 8436 1746
rect 8454 1743 8475 1746
rect 8454 1728 8569 1743
rect 4163 1656 4205 1692
rect 4477 1688 4538 1704
rect 4382 1684 4538 1688
rect 4382 1666 4500 1684
rect 4518 1666 4538 1684
rect 4106 1655 4206 1656
rect 4050 1634 4206 1655
rect 4382 1645 4538 1666
rect 4382 1644 4482 1645
rect 19 1557 134 1572
rect 113 1554 134 1557
rect 152 1554 170 1572
rect 113 1535 170 1554
rect 4050 1616 4070 1634
rect 4088 1616 4206 1634
rect 4050 1612 4206 1616
rect 4050 1596 4111 1612
rect 4383 1608 4425 1644
rect 4383 1585 4534 1608
rect 8418 1705 8569 1728
rect 12795 1758 12852 1777
rect 12795 1740 12813 1758
rect 12831 1755 12852 1758
rect 12831 1740 12946 1755
rect 8527 1669 8569 1705
rect 8854 1700 8915 1716
rect 8759 1696 8915 1700
rect 8759 1678 8877 1696
rect 8895 1678 8915 1696
rect 8470 1668 8570 1669
rect 8414 1647 8570 1668
rect 8759 1657 8915 1678
rect 8759 1656 8859 1657
rect 4383 1570 4498 1585
rect 4477 1567 4498 1570
rect 4516 1567 4534 1585
rect 4477 1548 4534 1567
rect 4047 1515 4104 1534
rect 8414 1629 8434 1647
rect 8452 1629 8570 1647
rect 8414 1625 8570 1629
rect 8414 1609 8475 1625
rect 8760 1620 8802 1656
rect 8760 1597 8911 1620
rect 12795 1717 12946 1740
rect 17159 1771 17216 1790
rect 17159 1753 17177 1771
rect 17195 1768 17216 1771
rect 17195 1753 17310 1768
rect 12904 1681 12946 1717
rect 13218 1713 13279 1729
rect 13123 1709 13279 1713
rect 13123 1691 13241 1709
rect 13259 1691 13279 1709
rect 12847 1680 12947 1681
rect 12791 1659 12947 1680
rect 13123 1670 13279 1691
rect 13123 1669 13223 1670
rect 8760 1582 8875 1597
rect 8854 1579 8875 1582
rect 8893 1579 8911 1597
rect 8854 1560 8911 1579
rect 4047 1497 4065 1515
rect 4083 1512 4104 1515
rect 4083 1497 4198 1512
rect 4047 1474 4198 1497
rect 108 1351 169 1367
rect 4156 1438 4198 1474
rect 8411 1528 8468 1547
rect 8411 1510 8429 1528
rect 8447 1525 8468 1528
rect 12791 1641 12811 1659
rect 12829 1641 12947 1659
rect 12791 1637 12947 1641
rect 12791 1621 12852 1637
rect 13124 1633 13166 1669
rect 13124 1610 13275 1633
rect 17159 1730 17310 1753
rect 17268 1694 17310 1730
rect 21425 1745 21482 1764
rect 21425 1727 21443 1745
rect 21461 1742 21482 1745
rect 21461 1727 21576 1742
rect 17211 1693 17311 1694
rect 17155 1672 17311 1693
rect 17484 1687 17545 1703
rect 13124 1595 13239 1610
rect 13218 1592 13239 1595
rect 13257 1592 13275 1610
rect 13218 1573 13275 1592
rect 8447 1510 8562 1525
rect 8411 1487 8562 1510
rect 4099 1437 4199 1438
rect 4043 1416 4199 1437
rect 4043 1398 4063 1416
rect 4081 1398 4199 1416
rect 4043 1394 4199 1398
rect 13 1347 169 1351
rect 13 1329 131 1347
rect 149 1329 169 1347
rect 13 1308 169 1329
rect 13 1307 113 1308
rect 14 1271 56 1307
rect 4043 1378 4104 1394
rect 4472 1364 4533 1380
rect 8520 1451 8562 1487
rect 12788 1540 12845 1559
rect 17155 1654 17175 1672
rect 17193 1654 17311 1672
rect 17155 1650 17311 1654
rect 17389 1683 17545 1687
rect 17389 1665 17507 1683
rect 17525 1665 17545 1683
rect 17155 1634 17216 1650
rect 17389 1644 17545 1665
rect 17389 1643 17489 1644
rect 17390 1607 17432 1643
rect 17390 1584 17541 1607
rect 21425 1704 21576 1727
rect 25789 1758 25846 1777
rect 25789 1740 25807 1758
rect 25825 1755 25846 1758
rect 25825 1740 25940 1755
rect 21534 1668 21576 1704
rect 21848 1700 21909 1716
rect 21753 1696 21909 1700
rect 21753 1678 21871 1696
rect 21889 1678 21909 1696
rect 21477 1667 21577 1668
rect 21421 1646 21577 1667
rect 21753 1657 21909 1678
rect 21753 1656 21853 1657
rect 12788 1522 12806 1540
rect 12824 1537 12845 1540
rect 12824 1522 12939 1537
rect 12788 1499 12939 1522
rect 8463 1450 8563 1451
rect 8407 1429 8563 1450
rect 8407 1411 8427 1429
rect 8445 1411 8563 1429
rect 8407 1407 8563 1411
rect 4377 1360 4533 1364
rect 4041 1332 4098 1351
rect 14 1248 165 1271
rect 14 1233 129 1248
rect 108 1230 129 1233
rect 147 1230 165 1248
rect 4041 1314 4059 1332
rect 4077 1329 4098 1332
rect 4377 1342 4495 1360
rect 4513 1342 4533 1360
rect 4077 1314 4192 1329
rect 4377 1321 4533 1342
rect 4377 1320 4477 1321
rect 4041 1291 4192 1314
rect 108 1211 165 1230
rect 102 1168 163 1184
rect 4150 1255 4192 1291
rect 4378 1284 4420 1320
rect 8407 1391 8468 1407
rect 8849 1376 8910 1392
rect 12897 1463 12939 1499
rect 17152 1553 17209 1572
rect 17390 1569 17505 1584
rect 17152 1535 17170 1553
rect 17188 1550 17209 1553
rect 17484 1566 17505 1569
rect 17523 1566 17541 1584
rect 17188 1535 17303 1550
rect 17484 1547 17541 1566
rect 17152 1512 17303 1535
rect 21421 1628 21441 1646
rect 21459 1628 21577 1646
rect 21421 1624 21577 1628
rect 21421 1608 21482 1624
rect 21754 1620 21796 1656
rect 21754 1597 21905 1620
rect 25789 1717 25940 1740
rect 30166 1770 30223 1789
rect 30166 1752 30184 1770
rect 30202 1767 30223 1770
rect 30202 1752 30317 1767
rect 25898 1681 25940 1717
rect 26225 1712 26286 1728
rect 26130 1708 26286 1712
rect 26130 1690 26248 1708
rect 26266 1690 26286 1708
rect 25841 1680 25941 1681
rect 25785 1659 25941 1680
rect 26130 1669 26286 1690
rect 26130 1668 26230 1669
rect 21754 1582 21869 1597
rect 21848 1579 21869 1582
rect 21887 1579 21905 1597
rect 21848 1560 21905 1579
rect 12840 1462 12940 1463
rect 12784 1441 12940 1462
rect 12784 1423 12804 1441
rect 12822 1423 12940 1441
rect 12784 1419 12940 1423
rect 8754 1372 8910 1376
rect 8405 1345 8462 1364
rect 4378 1261 4529 1284
rect 4093 1254 4193 1255
rect 4037 1233 4193 1254
rect 4378 1246 4493 1261
rect 4037 1215 4057 1233
rect 4075 1215 4193 1233
rect 4472 1243 4493 1246
rect 4511 1243 4529 1261
rect 8405 1327 8423 1345
rect 8441 1342 8462 1345
rect 8754 1354 8872 1372
rect 8890 1354 8910 1372
rect 8441 1327 8556 1342
rect 8754 1333 8910 1354
rect 8754 1332 8854 1333
rect 8405 1304 8556 1327
rect 4472 1224 4529 1243
rect 4037 1211 4193 1215
rect 7 1164 163 1168
rect 7 1146 125 1164
rect 143 1146 163 1164
rect 7 1125 163 1146
rect 7 1124 107 1125
rect 8 1088 50 1124
rect 4037 1195 4098 1211
rect 4466 1181 4527 1197
rect 8514 1268 8556 1304
rect 8755 1296 8797 1332
rect 12784 1403 12845 1419
rect 13213 1389 13274 1405
rect 17261 1476 17303 1512
rect 17204 1475 17304 1476
rect 17148 1454 17304 1475
rect 21418 1527 21475 1546
rect 25785 1641 25805 1659
rect 25823 1641 25941 1659
rect 25785 1637 25941 1641
rect 25785 1621 25846 1637
rect 26131 1632 26173 1668
rect 26131 1609 26282 1632
rect 30166 1729 30317 1752
rect 34530 1783 34587 1802
rect 34530 1765 34548 1783
rect 34566 1780 34587 1783
rect 34566 1765 34681 1780
rect 30275 1693 30317 1729
rect 30589 1725 30650 1741
rect 30494 1721 30650 1725
rect 30494 1703 30612 1721
rect 30630 1703 30650 1721
rect 30218 1692 30318 1693
rect 30162 1671 30318 1692
rect 30494 1682 30650 1703
rect 30494 1681 30594 1682
rect 26131 1594 26246 1609
rect 26225 1591 26246 1594
rect 26264 1591 26282 1609
rect 26225 1572 26282 1591
rect 21418 1509 21436 1527
rect 21454 1524 21475 1527
rect 21454 1509 21569 1524
rect 21418 1486 21569 1509
rect 17148 1436 17168 1454
rect 17186 1436 17304 1454
rect 17148 1432 17304 1436
rect 13118 1385 13274 1389
rect 12782 1357 12839 1376
rect 8755 1273 8906 1296
rect 8457 1267 8557 1268
rect 8401 1246 8557 1267
rect 8755 1258 8870 1273
rect 8401 1228 8421 1246
rect 8439 1228 8557 1246
rect 8849 1255 8870 1258
rect 8888 1255 8906 1273
rect 12782 1339 12800 1357
rect 12818 1354 12839 1357
rect 13118 1367 13236 1385
rect 13254 1367 13274 1385
rect 12818 1339 12933 1354
rect 13118 1346 13274 1367
rect 13118 1345 13218 1346
rect 12782 1316 12933 1339
rect 8849 1236 8906 1255
rect 8401 1224 8557 1228
rect 4371 1177 4527 1181
rect 4371 1159 4489 1177
rect 4507 1159 4527 1177
rect 4371 1138 4527 1159
rect 4371 1137 4471 1138
rect 4372 1101 4414 1137
rect 8401 1208 8462 1224
rect 8843 1193 8904 1209
rect 12891 1280 12933 1316
rect 13119 1309 13161 1345
rect 17148 1416 17209 1432
rect 17146 1370 17203 1389
rect 13119 1286 13270 1309
rect 12834 1279 12934 1280
rect 12778 1258 12934 1279
rect 13119 1271 13234 1286
rect 12778 1240 12798 1258
rect 12816 1240 12934 1258
rect 13213 1268 13234 1271
rect 13252 1268 13270 1286
rect 17146 1352 17164 1370
rect 17182 1367 17203 1370
rect 17182 1352 17297 1367
rect 17479 1363 17540 1379
rect 21527 1450 21569 1486
rect 25782 1540 25839 1559
rect 25782 1522 25800 1540
rect 25818 1537 25839 1540
rect 30162 1653 30182 1671
rect 30200 1653 30318 1671
rect 30162 1649 30318 1653
rect 30162 1633 30223 1649
rect 30495 1645 30537 1681
rect 30495 1622 30646 1645
rect 34530 1742 34681 1765
rect 34639 1706 34681 1742
rect 34582 1705 34682 1706
rect 34526 1684 34682 1705
rect 30495 1607 30610 1622
rect 30589 1604 30610 1607
rect 30628 1604 30646 1622
rect 30589 1585 30646 1604
rect 25818 1522 25933 1537
rect 25782 1499 25933 1522
rect 21470 1449 21570 1450
rect 21414 1428 21570 1449
rect 21414 1410 21434 1428
rect 21452 1410 21570 1428
rect 21414 1406 21570 1410
rect 17146 1329 17297 1352
rect 13213 1249 13270 1268
rect 12778 1236 12934 1240
rect 8748 1189 8904 1193
rect 8748 1171 8866 1189
rect 8884 1171 8904 1189
rect 8748 1150 8904 1171
rect 8748 1149 8848 1150
rect 8749 1113 8791 1149
rect 12778 1220 12839 1236
rect 13207 1206 13268 1222
rect 17255 1293 17297 1329
rect 17384 1359 17540 1363
rect 17384 1341 17502 1359
rect 17520 1341 17540 1359
rect 17384 1320 17540 1341
rect 17384 1319 17484 1320
rect 17198 1292 17298 1293
rect 17142 1271 17298 1292
rect 17142 1253 17162 1271
rect 17180 1253 17298 1271
rect 17142 1249 17298 1253
rect 17385 1283 17427 1319
rect 21414 1390 21475 1406
rect 21843 1376 21904 1392
rect 25891 1463 25933 1499
rect 30159 1552 30216 1571
rect 34526 1666 34546 1684
rect 34564 1666 34682 1684
rect 34526 1662 34682 1666
rect 34526 1646 34587 1662
rect 30159 1534 30177 1552
rect 30195 1549 30216 1552
rect 30195 1534 30310 1549
rect 30159 1511 30310 1534
rect 25834 1462 25934 1463
rect 25778 1441 25934 1462
rect 25778 1423 25798 1441
rect 25816 1423 25934 1441
rect 25778 1419 25934 1423
rect 21748 1372 21904 1376
rect 21412 1344 21469 1363
rect 17385 1260 17536 1283
rect 13112 1202 13268 1206
rect 13112 1184 13230 1202
rect 13248 1184 13268 1202
rect 13112 1163 13268 1184
rect 13112 1162 13212 1163
rect 13113 1126 13155 1162
rect 17142 1233 17203 1249
rect 17385 1245 17500 1260
rect 17479 1242 17500 1245
rect 17518 1242 17536 1260
rect 21412 1326 21430 1344
rect 21448 1341 21469 1344
rect 21748 1354 21866 1372
rect 21884 1354 21904 1372
rect 21448 1326 21563 1341
rect 21748 1333 21904 1354
rect 21748 1332 21848 1333
rect 21412 1303 21563 1326
rect 17479 1223 17536 1242
rect 17473 1180 17534 1196
rect 21521 1267 21563 1303
rect 21749 1296 21791 1332
rect 25778 1403 25839 1419
rect 26220 1388 26281 1404
rect 30268 1475 30310 1511
rect 34523 1565 34580 1584
rect 34523 1547 34541 1565
rect 34559 1562 34580 1565
rect 34559 1547 34674 1562
rect 34523 1524 34674 1547
rect 30211 1474 30311 1475
rect 30155 1453 30311 1474
rect 30155 1435 30175 1453
rect 30193 1435 30311 1453
rect 30155 1431 30311 1435
rect 26125 1384 26281 1388
rect 25776 1357 25833 1376
rect 21749 1273 21900 1296
rect 21464 1266 21564 1267
rect 21408 1245 21564 1266
rect 21749 1258 21864 1273
rect 21408 1227 21428 1245
rect 21446 1227 21564 1245
rect 21843 1255 21864 1258
rect 21882 1255 21900 1273
rect 25776 1339 25794 1357
rect 25812 1354 25833 1357
rect 26125 1366 26243 1384
rect 26261 1366 26281 1384
rect 25812 1339 25927 1354
rect 26125 1345 26281 1366
rect 26125 1344 26225 1345
rect 25776 1316 25927 1339
rect 21843 1236 21900 1255
rect 21408 1223 21564 1227
rect 17378 1176 17534 1180
rect 17378 1158 17496 1176
rect 17514 1158 17534 1176
rect 17378 1137 17534 1158
rect 17378 1136 17478 1137
rect 8 1065 159 1088
rect 8 1050 123 1065
rect 102 1047 123 1050
rect 141 1047 159 1065
rect 102 1028 159 1047
rect 4372 1078 4523 1101
rect 4372 1063 4487 1078
rect 4466 1060 4487 1063
rect 4505 1060 4523 1078
rect 95 950 156 966
rect 0 946 156 950
rect 0 928 118 946
rect 136 928 156 946
rect 4466 1041 4523 1060
rect 8749 1090 8900 1113
rect 8749 1075 8864 1090
rect 8843 1072 8864 1075
rect 8882 1072 8900 1090
rect 4036 1008 4093 1027
rect 4036 990 4054 1008
rect 4072 1005 4093 1008
rect 4072 990 4187 1005
rect 4036 967 4187 990
rect 0 907 156 928
rect 0 906 100 907
rect 1 870 43 906
rect 1 847 152 870
rect 4145 931 4187 967
rect 4459 963 4520 979
rect 4364 959 4520 963
rect 4364 941 4482 959
rect 4500 941 4520 959
rect 8843 1053 8900 1072
rect 13113 1103 13264 1126
rect 13113 1088 13228 1103
rect 13207 1085 13228 1088
rect 13246 1085 13264 1103
rect 8400 1021 8457 1040
rect 8400 1003 8418 1021
rect 8436 1018 8457 1021
rect 8436 1003 8551 1018
rect 8400 980 8551 1003
rect 4088 930 4188 931
rect 4032 909 4188 930
rect 4364 920 4520 941
rect 4364 919 4464 920
rect 4032 891 4052 909
rect 4070 891 4188 909
rect 4032 887 4188 891
rect 4032 871 4093 887
rect 4365 883 4407 919
rect 1 832 116 847
rect 95 829 116 832
rect 134 829 152 847
rect 95 810 152 829
rect 4365 860 4516 883
rect 8509 944 8551 980
rect 8836 975 8897 991
rect 8741 971 8897 975
rect 8741 953 8859 971
rect 8877 953 8897 971
rect 13207 1066 13264 1085
rect 17379 1100 17421 1136
rect 21408 1207 21469 1223
rect 21837 1193 21898 1209
rect 25885 1280 25927 1316
rect 26126 1308 26168 1344
rect 30155 1415 30216 1431
rect 30584 1401 30645 1417
rect 34632 1488 34674 1524
rect 34575 1487 34675 1488
rect 34519 1466 34675 1487
rect 34519 1448 34539 1466
rect 34557 1448 34675 1466
rect 34519 1444 34675 1448
rect 30489 1397 30645 1401
rect 30153 1369 30210 1388
rect 26126 1285 26277 1308
rect 25828 1279 25928 1280
rect 25772 1258 25928 1279
rect 26126 1270 26241 1285
rect 25772 1240 25792 1258
rect 25810 1240 25928 1258
rect 26220 1267 26241 1270
rect 26259 1267 26277 1285
rect 30153 1351 30171 1369
rect 30189 1366 30210 1369
rect 30489 1379 30607 1397
rect 30625 1379 30645 1397
rect 30189 1351 30304 1366
rect 30489 1358 30645 1379
rect 30489 1357 30589 1358
rect 30153 1328 30304 1351
rect 26220 1248 26277 1267
rect 25772 1236 25928 1240
rect 21742 1189 21898 1193
rect 21742 1171 21860 1189
rect 21878 1171 21898 1189
rect 21742 1150 21898 1171
rect 21742 1149 21842 1150
rect 21743 1113 21785 1149
rect 25772 1220 25833 1236
rect 26214 1205 26275 1221
rect 30262 1292 30304 1328
rect 30490 1321 30532 1357
rect 34519 1428 34580 1444
rect 34517 1382 34574 1401
rect 30490 1298 30641 1321
rect 30205 1291 30305 1292
rect 30149 1270 30305 1291
rect 30490 1283 30605 1298
rect 30149 1252 30169 1270
rect 30187 1252 30305 1270
rect 30584 1280 30605 1283
rect 30623 1280 30641 1298
rect 34517 1364 34535 1382
rect 34553 1379 34574 1382
rect 34553 1364 34668 1379
rect 34517 1341 34668 1364
rect 30584 1261 30641 1280
rect 30149 1248 30305 1252
rect 26119 1201 26275 1205
rect 26119 1183 26237 1201
rect 26255 1183 26275 1201
rect 26119 1162 26275 1183
rect 26119 1161 26219 1162
rect 26120 1125 26162 1161
rect 30149 1232 30210 1248
rect 30578 1218 30639 1234
rect 34626 1305 34668 1341
rect 34569 1304 34669 1305
rect 34513 1283 34669 1304
rect 34513 1265 34533 1283
rect 34551 1265 34669 1283
rect 34513 1261 34669 1265
rect 30483 1214 30639 1218
rect 30483 1196 30601 1214
rect 30619 1196 30639 1214
rect 30483 1175 30639 1196
rect 30483 1174 30583 1175
rect 30484 1138 30526 1174
rect 34513 1245 34574 1261
rect 12777 1033 12834 1052
rect 12777 1015 12795 1033
rect 12813 1030 12834 1033
rect 12813 1015 12928 1030
rect 12777 992 12928 1015
rect 8452 943 8552 944
rect 8396 922 8552 943
rect 8741 932 8897 953
rect 8741 931 8841 932
rect 8396 904 8416 922
rect 8434 904 8552 922
rect 8396 900 8552 904
rect 8396 884 8457 900
rect 8742 895 8784 931
rect 4365 845 4480 860
rect 4459 842 4480 845
rect 4498 842 4516 860
rect 4459 823 4516 842
rect 8742 872 8893 895
rect 12886 956 12928 992
rect 13200 988 13261 1004
rect 13105 984 13261 988
rect 13105 966 13223 984
rect 13241 966 13261 984
rect 17379 1077 17530 1100
rect 17141 1046 17198 1065
rect 17379 1062 17494 1077
rect 17141 1028 17159 1046
rect 17177 1043 17198 1046
rect 17473 1059 17494 1062
rect 17512 1059 17530 1077
rect 17177 1028 17292 1043
rect 17473 1040 17530 1059
rect 21743 1090 21894 1113
rect 21743 1075 21858 1090
rect 21837 1072 21858 1075
rect 21876 1072 21894 1090
rect 17141 1005 17292 1028
rect 12829 955 12929 956
rect 12773 934 12929 955
rect 13105 945 13261 966
rect 13105 944 13205 945
rect 12773 916 12793 934
rect 12811 916 12929 934
rect 12773 912 12929 916
rect 12773 896 12834 912
rect 13106 908 13148 944
rect 8742 857 8857 872
rect 8836 854 8857 857
rect 8875 854 8893 872
rect 8836 835 8893 854
rect 13106 885 13257 908
rect 17250 969 17292 1005
rect 17193 968 17293 969
rect 17137 947 17293 968
rect 17466 962 17527 978
rect 17137 929 17157 947
rect 17175 929 17293 947
rect 17137 925 17293 929
rect 17378 958 17527 962
rect 17378 940 17489 958
rect 17507 940 17527 958
rect 21837 1053 21894 1072
rect 26120 1102 26271 1125
rect 26120 1087 26235 1102
rect 26214 1084 26235 1087
rect 26253 1084 26271 1102
rect 21407 1020 21464 1039
rect 21407 1002 21425 1020
rect 21443 1017 21464 1020
rect 21443 1002 21558 1017
rect 21407 979 21558 1002
rect 17137 909 17198 925
rect 17378 919 17527 940
rect 17378 918 17471 919
rect 13106 870 13221 885
rect 13200 867 13221 870
rect 13239 867 13257 885
rect 13200 848 13257 867
rect 17378 882 17414 918
rect 17378 859 17523 882
rect 21516 943 21558 979
rect 21830 975 21891 991
rect 21735 971 21891 975
rect 21735 953 21853 971
rect 21871 953 21891 971
rect 26214 1065 26271 1084
rect 30484 1115 30635 1138
rect 30484 1100 30599 1115
rect 30578 1097 30599 1100
rect 30617 1097 30635 1115
rect 25771 1033 25828 1052
rect 25771 1015 25789 1033
rect 25807 1030 25828 1033
rect 25807 1015 25922 1030
rect 25771 992 25922 1015
rect 21459 942 21559 943
rect 21403 921 21559 942
rect 21735 932 21891 953
rect 21735 931 21835 932
rect 21403 903 21423 921
rect 21441 903 21559 921
rect 21403 899 21559 903
rect 21403 883 21464 899
rect 21736 895 21778 931
rect 17378 844 17487 859
rect 17466 841 17487 844
rect 17505 841 17523 859
rect 17466 822 17523 841
rect 21736 872 21887 895
rect 25880 956 25922 992
rect 26207 987 26268 1003
rect 26112 983 26268 987
rect 26112 965 26230 983
rect 26248 965 26268 983
rect 30578 1078 30635 1097
rect 30148 1045 30205 1064
rect 30148 1027 30166 1045
rect 30184 1042 30205 1045
rect 30184 1027 30299 1042
rect 30148 1004 30299 1027
rect 25823 955 25923 956
rect 25767 934 25923 955
rect 26112 944 26268 965
rect 26112 943 26212 944
rect 25767 916 25787 934
rect 25805 916 25923 934
rect 25767 912 25923 916
rect 25767 896 25828 912
rect 26113 907 26155 943
rect 21736 857 21851 872
rect 21830 854 21851 857
rect 21869 854 21887 872
rect 21830 835 21887 854
rect 26113 884 26264 907
rect 30257 968 30299 1004
rect 30571 1000 30632 1016
rect 30476 996 30632 1000
rect 30476 978 30594 996
rect 30612 978 30632 996
rect 34512 1058 34569 1077
rect 34512 1040 34530 1058
rect 34548 1055 34569 1058
rect 34548 1040 34663 1055
rect 34512 1017 34663 1040
rect 30200 967 30300 968
rect 30144 946 30300 967
rect 30476 957 30632 978
rect 30476 956 30576 957
rect 30144 928 30164 946
rect 30182 928 30300 946
rect 30144 924 30300 928
rect 30144 908 30205 924
rect 30477 920 30519 956
rect 26113 869 26228 884
rect 26207 866 26228 869
rect 26246 866 26264 884
rect 26207 847 26264 866
rect 30477 897 30628 920
rect 34621 981 34663 1017
rect 34564 980 34664 981
rect 34508 959 34664 980
rect 34508 941 34528 959
rect 34546 941 34664 959
rect 34508 937 34664 941
rect 34508 921 34569 937
rect 30477 882 30592 897
rect 30571 879 30592 882
rect 30610 879 30628 897
rect 30571 860 30628 879
<< locali >>
rect 25917 9041 25958 9044
rect 16890 9037 16929 9038
rect 8546 9029 8587 9032
rect 2875 8938 2915 8946
rect 2875 8916 2883 8938
rect 2907 8916 2915 8938
rect 3779 8941 4235 8976
rect 8146 8969 9041 9029
rect 16889 9004 17670 9037
rect 8146 8968 8593 8969
rect 7239 8951 7279 8959
rect 253 8797 300 8913
rect 253 8779 263 8797
rect 281 8779 300 8797
rect 253 8775 300 8779
rect 254 8770 291 8775
rect 242 8708 294 8710
rect 240 8704 673 8708
rect 240 8698 679 8704
rect 240 8680 261 8698
rect 279 8680 679 8698
rect 240 8662 679 8680
rect 242 8473 294 8662
rect 640 8637 679 8662
rect 2480 8687 2517 8693
rect 2480 8668 2488 8687
rect 2509 8668 2517 8687
rect 2480 8660 2517 8668
rect 424 8612 611 8636
rect 640 8617 1035 8637
rect 1055 8617 1058 8637
rect 640 8612 1058 8617
rect 424 8541 461 8612
rect 640 8611 983 8612
rect 640 8608 679 8611
rect 945 8610 982 8611
rect 576 8551 607 8552
rect 424 8521 433 8541
rect 453 8521 461 8541
rect 424 8511 461 8521
rect 520 8541 607 8551
rect 520 8521 529 8541
rect 549 8521 607 8541
rect 520 8512 607 8521
rect 520 8511 557 8512
rect 242 8455 258 8473
rect 276 8455 294 8473
rect 576 8461 607 8512
rect 642 8541 679 8608
rect 794 8551 830 8552
rect 642 8521 651 8541
rect 671 8521 679 8541
rect 642 8511 679 8521
rect 738 8541 886 8551
rect 986 8548 1082 8550
rect 738 8521 747 8541
rect 767 8521 857 8541
rect 877 8521 886 8541
rect 738 8512 886 8521
rect 944 8541 1082 8548
rect 944 8521 953 8541
rect 973 8521 1082 8541
rect 944 8512 1082 8521
rect 738 8511 775 8512
rect 468 8458 509 8459
rect 242 8437 294 8455
rect 360 8451 509 8458
rect 360 8431 419 8451
rect 439 8431 478 8451
rect 498 8431 509 8451
rect 360 8423 509 8431
rect 576 8454 733 8461
rect 576 8434 696 8454
rect 716 8434 733 8454
rect 576 8424 733 8434
rect 576 8423 611 8424
rect 576 8402 607 8423
rect 794 8402 830 8512
rect 849 8511 886 8512
rect 945 8511 982 8512
rect 905 8452 995 8458
rect 905 8432 914 8452
rect 934 8450 995 8452
rect 934 8432 959 8450
rect 905 8430 959 8432
rect 979 8430 995 8450
rect 905 8424 995 8430
rect 419 8401 456 8402
rect 418 8392 456 8401
rect 246 8374 286 8384
rect 246 8356 256 8374
rect 274 8356 286 8374
rect 418 8372 427 8392
rect 447 8372 456 8392
rect 418 8364 456 8372
rect 522 8396 607 8402
rect 637 8401 674 8402
rect 522 8376 530 8396
rect 550 8376 607 8396
rect 522 8368 607 8376
rect 636 8392 674 8401
rect 636 8372 645 8392
rect 665 8372 674 8392
rect 522 8367 558 8368
rect 636 8364 674 8372
rect 740 8396 884 8402
rect 740 8376 748 8396
rect 768 8376 801 8396
rect 821 8376 856 8396
rect 876 8376 884 8396
rect 740 8368 884 8376
rect 740 8367 776 8368
rect 848 8367 884 8368
rect 950 8401 987 8402
rect 950 8400 988 8401
rect 950 8392 1014 8400
rect 950 8372 959 8392
rect 979 8378 1014 8392
rect 1034 8378 1037 8398
rect 979 8373 1037 8378
rect 979 8372 1014 8373
rect 246 8300 286 8356
rect 419 8335 456 8364
rect 420 8333 456 8335
rect 420 8311 611 8333
rect 637 8332 674 8364
rect 950 8360 1014 8372
rect 1054 8334 1081 8512
rect 913 8332 1081 8334
rect 637 8322 1081 8332
rect 1222 8428 1409 8452
rect 1440 8433 1833 8453
rect 1853 8433 1856 8453
rect 1440 8428 1856 8433
rect 1222 8357 1259 8428
rect 1440 8427 1781 8428
rect 1374 8367 1405 8368
rect 1222 8337 1231 8357
rect 1251 8337 1259 8357
rect 1222 8327 1259 8337
rect 1318 8357 1405 8367
rect 1318 8337 1327 8357
rect 1347 8337 1405 8357
rect 1318 8328 1405 8337
rect 1318 8327 1355 8328
rect 243 8295 286 8300
rect 634 8306 1081 8322
rect 634 8300 662 8306
rect 913 8305 1081 8306
rect 243 8292 393 8295
rect 634 8292 661 8300
rect 243 8290 661 8292
rect 243 8272 252 8290
rect 270 8272 661 8290
rect 1374 8277 1405 8328
rect 1440 8357 1477 8427
rect 1743 8426 1780 8427
rect 1592 8367 1628 8368
rect 1440 8337 1449 8357
rect 1469 8337 1477 8357
rect 1440 8327 1477 8337
rect 1536 8357 1684 8367
rect 1784 8364 1880 8366
rect 1536 8337 1545 8357
rect 1565 8337 1655 8357
rect 1675 8337 1684 8357
rect 1536 8328 1684 8337
rect 1742 8357 1880 8364
rect 1742 8337 1751 8357
rect 1771 8337 1880 8357
rect 1742 8328 1880 8337
rect 1536 8327 1573 8328
rect 1266 8274 1307 8275
rect 243 8269 661 8272
rect 243 8263 286 8269
rect 246 8260 286 8263
rect 1158 8267 1307 8274
rect 643 8251 683 8252
rect 354 8234 683 8251
rect 1158 8247 1217 8267
rect 1237 8247 1276 8267
rect 1296 8247 1307 8267
rect 1158 8239 1307 8247
rect 1374 8270 1531 8277
rect 1374 8250 1494 8270
rect 1514 8250 1531 8270
rect 1374 8240 1531 8250
rect 1374 8239 1409 8240
rect 238 8191 281 8202
rect 238 8173 250 8191
rect 268 8173 281 8191
rect 238 8147 281 8173
rect 354 8147 381 8234
rect 643 8225 683 8234
rect 238 8126 381 8147
rect 425 8199 459 8215
rect 643 8205 1036 8225
rect 1056 8205 1059 8225
rect 1374 8218 1405 8239
rect 1592 8218 1628 8328
rect 1647 8327 1684 8328
rect 1743 8327 1780 8328
rect 1703 8268 1793 8274
rect 1703 8248 1712 8268
rect 1732 8266 1793 8268
rect 1732 8248 1757 8266
rect 1703 8246 1757 8248
rect 1777 8246 1793 8266
rect 1703 8240 1793 8246
rect 1217 8217 1254 8218
rect 643 8200 1059 8205
rect 1216 8208 1254 8217
rect 643 8199 984 8200
rect 425 8129 462 8199
rect 577 8139 608 8140
rect 238 8124 375 8126
rect 238 8082 281 8124
rect 425 8109 434 8129
rect 454 8109 462 8129
rect 425 8099 462 8109
rect 521 8129 608 8139
rect 521 8109 530 8129
rect 550 8109 608 8129
rect 521 8100 608 8109
rect 521 8099 558 8100
rect 236 8072 281 8082
rect 236 8054 245 8072
rect 263 8054 281 8072
rect 236 8048 281 8054
rect 577 8049 608 8100
rect 643 8129 680 8199
rect 946 8198 983 8199
rect 1216 8188 1225 8208
rect 1245 8188 1254 8208
rect 1216 8180 1254 8188
rect 1320 8212 1405 8218
rect 1435 8217 1472 8218
rect 1320 8192 1328 8212
rect 1348 8192 1405 8212
rect 1320 8184 1405 8192
rect 1434 8208 1472 8217
rect 1434 8188 1443 8208
rect 1463 8188 1472 8208
rect 1320 8183 1356 8184
rect 1434 8180 1472 8188
rect 1538 8212 1682 8218
rect 1538 8192 1546 8212
rect 1566 8193 1598 8212
rect 1619 8193 1654 8212
rect 1566 8192 1654 8193
rect 1674 8192 1682 8212
rect 1538 8184 1682 8192
rect 1538 8183 1574 8184
rect 1646 8183 1682 8184
rect 1748 8217 1785 8218
rect 1748 8216 1786 8217
rect 1748 8208 1812 8216
rect 1748 8188 1757 8208
rect 1777 8194 1812 8208
rect 1832 8194 1835 8214
rect 1777 8189 1835 8194
rect 1777 8188 1812 8189
rect 1217 8151 1254 8180
rect 1218 8149 1254 8151
rect 795 8139 831 8140
rect 643 8109 652 8129
rect 672 8109 680 8129
rect 643 8099 680 8109
rect 739 8129 887 8139
rect 987 8136 1083 8138
rect 739 8109 748 8129
rect 768 8109 858 8129
rect 878 8109 887 8129
rect 739 8100 887 8109
rect 945 8129 1083 8136
rect 945 8109 954 8129
rect 974 8109 1083 8129
rect 1218 8127 1409 8149
rect 1435 8148 1472 8180
rect 1748 8176 1812 8188
rect 1852 8150 1879 8328
rect 2484 8327 2517 8660
rect 2581 8692 2749 8693
rect 2875 8692 2915 8916
rect 3378 8920 3546 8921
rect 3779 8920 3824 8941
rect 3378 8894 3824 8920
rect 3378 8892 3546 8894
rect 3742 8893 3824 8894
rect 3959 8893 4040 8919
rect 4184 8906 4665 8941
rect 7239 8929 7247 8951
rect 7271 8929 7279 8951
rect 3378 8714 3405 8892
rect 3445 8854 3509 8866
rect 3785 8862 3822 8893
rect 4003 8862 4040 8893
rect 4187 8887 4226 8906
rect 4185 8868 4226 8887
rect 3445 8853 3480 8854
rect 3422 8848 3480 8853
rect 3422 8828 3425 8848
rect 3445 8834 3480 8848
rect 3500 8834 3509 8854
rect 3445 8826 3509 8834
rect 3471 8825 3509 8826
rect 3472 8824 3509 8825
rect 3575 8858 3611 8859
rect 3683 8858 3719 8859
rect 3575 8850 3719 8858
rect 3575 8830 3583 8850
rect 3603 8846 3691 8850
rect 3603 8830 3647 8846
rect 3575 8826 3647 8830
rect 3667 8830 3691 8846
rect 3711 8830 3719 8850
rect 3667 8826 3719 8830
rect 3575 8824 3719 8826
rect 3785 8854 3823 8862
rect 3901 8858 3937 8859
rect 3785 8834 3794 8854
rect 3814 8834 3823 8854
rect 3785 8825 3823 8834
rect 3852 8850 3937 8858
rect 3852 8830 3909 8850
rect 3929 8830 3937 8850
rect 3785 8824 3822 8825
rect 3852 8824 3937 8830
rect 4003 8854 4041 8862
rect 4003 8834 4012 8854
rect 4032 8834 4041 8854
rect 4003 8825 4041 8834
rect 4185 8859 4227 8868
rect 4185 8841 4199 8859
rect 4217 8841 4227 8859
rect 4185 8833 4227 8841
rect 4190 8831 4227 8833
rect 4003 8824 4040 8825
rect 3464 8796 3554 8802
rect 3464 8776 3480 8796
rect 3500 8794 3554 8796
rect 3500 8776 3525 8794
rect 3464 8774 3525 8776
rect 3545 8774 3554 8794
rect 3464 8768 3554 8774
rect 3477 8714 3514 8715
rect 3573 8714 3610 8715
rect 3629 8714 3665 8824
rect 3852 8803 3883 8824
rect 4617 8810 4664 8906
rect 3848 8802 3883 8803
rect 3726 8792 3883 8802
rect 3726 8772 3743 8792
rect 3763 8772 3883 8792
rect 3726 8765 3883 8772
rect 3950 8795 4099 8803
rect 3950 8775 3961 8795
rect 3981 8775 4020 8795
rect 4040 8775 4099 8795
rect 4617 8792 4627 8810
rect 4645 8792 4664 8810
rect 4617 8788 4664 8792
rect 4618 8783 4655 8788
rect 3950 8768 4099 8775
rect 3950 8767 3991 8768
rect 4187 8766 4224 8769
rect 3684 8714 3721 8715
rect 3377 8705 3515 8714
rect 2581 8666 3025 8692
rect 2581 8664 2749 8666
rect 2581 8486 2608 8664
rect 2648 8626 2712 8638
rect 2988 8634 3025 8666
rect 3051 8665 3242 8687
rect 3377 8685 3486 8705
rect 3506 8685 3515 8705
rect 3377 8678 3515 8685
rect 3573 8705 3721 8714
rect 3573 8685 3582 8705
rect 3602 8685 3692 8705
rect 3712 8685 3721 8705
rect 3377 8676 3473 8678
rect 3573 8675 3721 8685
rect 3780 8705 3817 8715
rect 3780 8685 3788 8705
rect 3808 8685 3817 8705
rect 3629 8674 3665 8675
rect 3206 8663 3242 8665
rect 3206 8634 3243 8663
rect 2648 8625 2683 8626
rect 2625 8620 2683 8625
rect 2625 8600 2628 8620
rect 2648 8606 2683 8620
rect 2703 8606 2712 8626
rect 2648 8600 2712 8606
rect 2625 8598 2712 8600
rect 2625 8594 2652 8598
rect 2674 8597 2712 8598
rect 2675 8596 2712 8597
rect 2778 8630 2814 8631
rect 2886 8630 2922 8631
rect 2778 8623 2922 8630
rect 2778 8622 2840 8623
rect 2778 8602 2786 8622
rect 2806 8605 2840 8622
rect 2859 8622 2922 8623
rect 2859 8605 2894 8622
rect 2806 8602 2894 8605
rect 2914 8602 2922 8622
rect 2778 8596 2922 8602
rect 2988 8626 3026 8634
rect 3104 8630 3140 8631
rect 2988 8606 2997 8626
rect 3017 8606 3026 8626
rect 2988 8597 3026 8606
rect 3055 8622 3140 8630
rect 3055 8602 3112 8622
rect 3132 8602 3140 8622
rect 2988 8596 3025 8597
rect 3055 8596 3140 8602
rect 3206 8626 3244 8634
rect 3206 8606 3215 8626
rect 3235 8606 3244 8626
rect 3477 8615 3514 8616
rect 3780 8615 3817 8685
rect 3852 8714 3883 8765
rect 4179 8760 4224 8766
rect 4179 8742 4197 8760
rect 4215 8742 4224 8760
rect 4179 8732 4224 8742
rect 3902 8714 3939 8715
rect 3852 8705 3939 8714
rect 3852 8685 3910 8705
rect 3930 8685 3939 8705
rect 3852 8675 3939 8685
rect 3998 8705 4035 8715
rect 3998 8685 4006 8705
rect 4026 8685 4035 8705
rect 4179 8690 4222 8732
rect 4606 8721 4658 8723
rect 4085 8688 4222 8690
rect 3852 8674 3883 8675
rect 3998 8615 4035 8685
rect 3476 8614 3817 8615
rect 3206 8597 3244 8606
rect 3401 8609 3817 8614
rect 3206 8596 3243 8597
rect 2667 8568 2757 8574
rect 2667 8548 2683 8568
rect 2703 8566 2757 8568
rect 2703 8548 2728 8566
rect 2667 8546 2728 8548
rect 2748 8546 2757 8566
rect 2667 8540 2757 8546
rect 2680 8486 2717 8487
rect 2776 8486 2813 8487
rect 2832 8486 2868 8596
rect 3055 8575 3086 8596
rect 3401 8589 3404 8609
rect 3424 8589 3817 8609
rect 4001 8599 4035 8615
rect 4079 8667 4222 8688
rect 4604 8717 5037 8721
rect 4604 8711 5043 8717
rect 4604 8693 4625 8711
rect 4643 8693 5043 8711
rect 4604 8675 5043 8693
rect 3777 8580 3817 8589
rect 4079 8580 4106 8667
rect 4179 8641 4222 8667
rect 4179 8623 4192 8641
rect 4210 8623 4222 8641
rect 4179 8612 4222 8623
rect 3051 8574 3086 8575
rect 2929 8564 3086 8574
rect 2929 8544 2946 8564
rect 2966 8544 3086 8564
rect 2929 8537 3086 8544
rect 3153 8567 3299 8575
rect 3153 8547 3164 8567
rect 3184 8547 3223 8567
rect 3243 8547 3299 8567
rect 3777 8563 4106 8580
rect 3777 8562 3817 8563
rect 3153 8540 3299 8547
rect 4174 8551 4214 8554
rect 4174 8545 4217 8551
rect 3799 8542 4217 8545
rect 3153 8539 3194 8540
rect 2887 8486 2924 8487
rect 2580 8477 2718 8486
rect 2580 8457 2689 8477
rect 2709 8457 2718 8477
rect 2580 8450 2718 8457
rect 2776 8477 2924 8486
rect 2776 8457 2785 8477
rect 2805 8457 2895 8477
rect 2915 8457 2924 8477
rect 2580 8448 2676 8450
rect 2776 8447 2924 8457
rect 2983 8477 3020 8487
rect 2983 8457 2991 8477
rect 3011 8457 3020 8477
rect 2832 8446 2868 8447
rect 2680 8387 2717 8388
rect 2983 8387 3020 8457
rect 3055 8486 3086 8537
rect 3799 8524 4190 8542
rect 4208 8524 4217 8542
rect 3799 8522 4217 8524
rect 3799 8514 3826 8522
rect 4067 8519 4217 8522
rect 3379 8508 3547 8509
rect 3798 8508 3826 8514
rect 3379 8492 3826 8508
rect 4174 8514 4217 8519
rect 3105 8486 3142 8487
rect 3055 8477 3142 8486
rect 3055 8457 3113 8477
rect 3133 8457 3142 8477
rect 3055 8447 3142 8457
rect 3201 8477 3238 8487
rect 3201 8457 3209 8477
rect 3229 8457 3238 8477
rect 3055 8446 3086 8447
rect 2679 8386 3020 8387
rect 3201 8386 3238 8457
rect 2604 8381 3020 8386
rect 2604 8361 2607 8381
rect 2627 8361 3020 8381
rect 3051 8362 3238 8386
rect 3379 8482 3823 8492
rect 3379 8480 3547 8482
rect 2479 8282 2521 8327
rect 3379 8302 3406 8480
rect 3446 8442 3510 8454
rect 3786 8450 3823 8482
rect 3849 8481 4040 8503
rect 4004 8479 4040 8481
rect 4004 8450 4041 8479
rect 4174 8458 4214 8514
rect 3446 8441 3481 8442
rect 3423 8436 3481 8441
rect 3423 8416 3426 8436
rect 3446 8422 3481 8436
rect 3501 8422 3510 8442
rect 3446 8414 3510 8422
rect 3472 8413 3510 8414
rect 3473 8412 3510 8413
rect 3576 8446 3612 8447
rect 3684 8446 3720 8447
rect 3576 8438 3720 8446
rect 3576 8418 3584 8438
rect 3604 8418 3639 8438
rect 3659 8418 3692 8438
rect 3712 8418 3720 8438
rect 3576 8412 3720 8418
rect 3786 8442 3824 8450
rect 3902 8446 3938 8447
rect 3786 8422 3795 8442
rect 3815 8422 3824 8442
rect 3786 8413 3824 8422
rect 3853 8438 3938 8446
rect 3853 8418 3910 8438
rect 3930 8418 3938 8438
rect 3786 8412 3823 8413
rect 3853 8412 3938 8418
rect 4004 8442 4042 8450
rect 4004 8422 4013 8442
rect 4033 8422 4042 8442
rect 4174 8440 4186 8458
rect 4204 8440 4214 8458
rect 4606 8486 4658 8675
rect 5004 8650 5043 8675
rect 6844 8700 6881 8706
rect 6844 8681 6852 8700
rect 6873 8681 6881 8700
rect 6844 8673 6881 8681
rect 4788 8625 4975 8649
rect 5004 8630 5399 8650
rect 5419 8630 5422 8650
rect 5004 8625 5422 8630
rect 4788 8554 4825 8625
rect 5004 8624 5347 8625
rect 5004 8621 5043 8624
rect 5309 8623 5346 8624
rect 4940 8564 4971 8565
rect 4788 8534 4797 8554
rect 4817 8534 4825 8554
rect 4788 8524 4825 8534
rect 4884 8554 4971 8564
rect 4884 8534 4893 8554
rect 4913 8534 4971 8554
rect 4884 8525 4971 8534
rect 4884 8524 4921 8525
rect 4606 8468 4622 8486
rect 4640 8468 4658 8486
rect 4940 8474 4971 8525
rect 5006 8554 5043 8621
rect 5158 8564 5194 8565
rect 5006 8534 5015 8554
rect 5035 8534 5043 8554
rect 5006 8524 5043 8534
rect 5102 8554 5250 8564
rect 5350 8561 5446 8563
rect 5102 8534 5111 8554
rect 5131 8534 5221 8554
rect 5241 8534 5250 8554
rect 5102 8525 5250 8534
rect 5308 8554 5446 8561
rect 5308 8534 5317 8554
rect 5337 8534 5446 8554
rect 5308 8525 5446 8534
rect 5102 8524 5139 8525
rect 4832 8471 4873 8472
rect 4606 8450 4658 8468
rect 4724 8464 4873 8471
rect 4174 8430 4214 8440
rect 4724 8444 4783 8464
rect 4803 8444 4842 8464
rect 4862 8444 4873 8464
rect 4724 8436 4873 8444
rect 4940 8467 5097 8474
rect 4940 8447 5060 8467
rect 5080 8447 5097 8467
rect 4940 8437 5097 8447
rect 4940 8436 4975 8437
rect 4004 8413 4042 8422
rect 4940 8415 4971 8436
rect 5158 8415 5194 8525
rect 5213 8524 5250 8525
rect 5309 8524 5346 8525
rect 5269 8465 5359 8471
rect 5269 8445 5278 8465
rect 5298 8463 5359 8465
rect 5298 8445 5323 8463
rect 5269 8443 5323 8445
rect 5343 8443 5359 8463
rect 5269 8437 5359 8443
rect 4783 8414 4820 8415
rect 4004 8412 4041 8413
rect 3465 8384 3555 8390
rect 3465 8364 3481 8384
rect 3501 8382 3555 8384
rect 3501 8364 3526 8382
rect 3465 8362 3526 8364
rect 3546 8362 3555 8382
rect 3465 8356 3555 8362
rect 3478 8302 3515 8303
rect 3574 8302 3611 8303
rect 3630 8302 3666 8412
rect 3853 8391 3884 8412
rect 4782 8405 4820 8414
rect 3849 8390 3884 8391
rect 3727 8380 3884 8390
rect 3727 8360 3744 8380
rect 3764 8360 3884 8380
rect 3727 8353 3884 8360
rect 3951 8383 4100 8391
rect 3951 8363 3962 8383
rect 3982 8363 4021 8383
rect 4041 8363 4100 8383
rect 4610 8387 4650 8397
rect 3951 8356 4100 8363
rect 4166 8359 4218 8377
rect 3951 8355 3992 8356
rect 3685 8302 3722 8303
rect 3378 8293 3516 8302
rect 2850 8282 2883 8284
rect 2479 8270 2926 8282
rect 1711 8148 1879 8150
rect 1435 8122 1879 8148
rect 945 8100 1083 8109
rect 739 8099 776 8100
rect 236 8045 273 8048
rect 469 8046 510 8047
rect 361 8039 510 8046
rect 361 8019 420 8039
rect 440 8019 479 8039
rect 499 8019 510 8039
rect 361 8011 510 8019
rect 577 8042 734 8049
rect 577 8022 697 8042
rect 717 8022 734 8042
rect 577 8012 734 8022
rect 577 8011 612 8012
rect 577 7990 608 8011
rect 795 7990 831 8100
rect 850 8099 887 8100
rect 946 8099 983 8100
rect 906 8040 996 8046
rect 906 8020 915 8040
rect 935 8038 996 8040
rect 935 8020 960 8038
rect 906 8018 960 8020
rect 980 8018 996 8038
rect 906 8012 996 8018
rect 420 7989 457 7990
rect 233 7981 270 7983
rect 233 7973 275 7981
rect 233 7955 243 7973
rect 261 7955 275 7973
rect 233 7946 275 7955
rect 419 7980 457 7989
rect 419 7960 428 7980
rect 448 7960 457 7980
rect 419 7952 457 7960
rect 523 7984 608 7990
rect 638 7989 675 7990
rect 523 7964 531 7984
rect 551 7964 608 7984
rect 523 7956 608 7964
rect 637 7980 675 7989
rect 637 7960 646 7980
rect 666 7960 675 7980
rect 523 7955 559 7956
rect 637 7952 675 7960
rect 741 7988 885 7990
rect 741 7984 793 7988
rect 741 7964 749 7984
rect 769 7968 793 7984
rect 813 7984 885 7988
rect 813 7968 857 7984
rect 769 7964 857 7968
rect 877 7964 885 7984
rect 741 7956 885 7964
rect 741 7955 777 7956
rect 849 7955 885 7956
rect 951 7989 988 7990
rect 951 7988 989 7989
rect 951 7980 1015 7988
rect 951 7960 960 7980
rect 980 7966 1015 7980
rect 1035 7966 1038 7986
rect 980 7961 1038 7966
rect 980 7960 1015 7961
rect 234 7921 275 7946
rect 420 7921 457 7952
rect 638 7921 675 7952
rect 951 7948 1015 7960
rect 1055 7922 1082 8100
rect 234 7894 283 7921
rect 419 7895 468 7921
rect 637 7920 718 7921
rect 914 7920 1082 7922
rect 637 7895 1082 7920
rect 638 7894 1082 7895
rect 236 7861 283 7894
rect 639 7861 679 7894
rect 914 7893 1082 7894
rect 1545 7898 1585 8122
rect 1711 8121 1879 8122
rect 2482 8256 2926 8270
rect 2482 8254 2650 8256
rect 2482 8076 2509 8254
rect 2549 8216 2613 8228
rect 2889 8224 2926 8256
rect 2952 8255 3143 8277
rect 3378 8273 3487 8293
rect 3507 8273 3516 8293
rect 3378 8266 3516 8273
rect 3574 8293 3722 8302
rect 3574 8273 3583 8293
rect 3603 8273 3693 8293
rect 3713 8273 3722 8293
rect 3378 8264 3474 8266
rect 3574 8263 3722 8273
rect 3781 8293 3818 8303
rect 3781 8273 3789 8293
rect 3809 8273 3818 8293
rect 3630 8262 3666 8263
rect 3107 8253 3143 8255
rect 3107 8224 3144 8253
rect 2549 8215 2584 8216
rect 2526 8210 2584 8215
rect 2526 8190 2529 8210
rect 2549 8196 2584 8210
rect 2604 8196 2613 8216
rect 2549 8188 2613 8196
rect 2575 8187 2613 8188
rect 2576 8186 2613 8187
rect 2679 8220 2715 8221
rect 2787 8220 2823 8221
rect 2679 8214 2823 8220
rect 2679 8212 2740 8214
rect 2679 8192 2687 8212
rect 2707 8197 2740 8212
rect 2759 8212 2823 8214
rect 2759 8197 2795 8212
rect 2707 8192 2795 8197
rect 2815 8192 2823 8212
rect 2679 8186 2823 8192
rect 2889 8216 2927 8224
rect 3005 8220 3041 8221
rect 2889 8196 2898 8216
rect 2918 8196 2927 8216
rect 2889 8187 2927 8196
rect 2956 8212 3041 8220
rect 2956 8192 3013 8212
rect 3033 8192 3041 8212
rect 2889 8186 2926 8187
rect 2956 8186 3041 8192
rect 3107 8216 3145 8224
rect 3107 8196 3116 8216
rect 3136 8196 3145 8216
rect 3781 8206 3818 8273
rect 3853 8302 3884 8353
rect 4166 8341 4184 8359
rect 4202 8341 4218 8359
rect 3903 8302 3940 8303
rect 3853 8293 3940 8302
rect 3853 8273 3911 8293
rect 3931 8273 3940 8293
rect 3853 8263 3940 8273
rect 3999 8293 4036 8303
rect 3999 8273 4007 8293
rect 4027 8273 4036 8293
rect 3853 8262 3884 8263
rect 3478 8203 3515 8204
rect 3781 8203 3820 8206
rect 3477 8202 3820 8203
rect 3999 8202 4036 8273
rect 3107 8187 3145 8196
rect 3402 8197 3820 8202
rect 3107 8186 3144 8187
rect 2568 8158 2658 8164
rect 2568 8138 2584 8158
rect 2604 8156 2658 8158
rect 2604 8138 2629 8156
rect 2568 8136 2629 8138
rect 2649 8136 2658 8156
rect 2568 8130 2658 8136
rect 2581 8076 2618 8077
rect 2677 8076 2714 8077
rect 2733 8076 2769 8186
rect 2956 8165 2987 8186
rect 3402 8177 3405 8197
rect 3425 8177 3820 8197
rect 3849 8178 4036 8202
rect 2952 8164 2987 8165
rect 2830 8154 2987 8164
rect 2830 8134 2847 8154
rect 2867 8134 2987 8154
rect 2830 8127 2987 8134
rect 3054 8157 3203 8165
rect 3054 8137 3065 8157
rect 3085 8137 3124 8157
rect 3144 8137 3203 8157
rect 3054 8130 3203 8137
rect 3781 8152 3820 8177
rect 4166 8152 4218 8341
rect 4610 8369 4620 8387
rect 4638 8369 4650 8387
rect 4782 8385 4791 8405
rect 4811 8385 4820 8405
rect 4782 8377 4820 8385
rect 4886 8409 4971 8415
rect 5001 8414 5038 8415
rect 4886 8389 4894 8409
rect 4914 8389 4971 8409
rect 4886 8381 4971 8389
rect 5000 8405 5038 8414
rect 5000 8385 5009 8405
rect 5029 8385 5038 8405
rect 4886 8380 4922 8381
rect 5000 8377 5038 8385
rect 5104 8409 5248 8415
rect 5104 8389 5112 8409
rect 5132 8389 5165 8409
rect 5185 8389 5220 8409
rect 5240 8389 5248 8409
rect 5104 8381 5248 8389
rect 5104 8380 5140 8381
rect 5212 8380 5248 8381
rect 5314 8414 5351 8415
rect 5314 8413 5352 8414
rect 5314 8405 5378 8413
rect 5314 8385 5323 8405
rect 5343 8391 5378 8405
rect 5398 8391 5401 8411
rect 5343 8386 5401 8391
rect 5343 8385 5378 8386
rect 4610 8313 4650 8369
rect 4783 8348 4820 8377
rect 4784 8346 4820 8348
rect 4784 8324 4975 8346
rect 5001 8345 5038 8377
rect 5314 8373 5378 8385
rect 5418 8347 5445 8525
rect 5277 8345 5445 8347
rect 5001 8335 5445 8345
rect 5586 8441 5773 8465
rect 5804 8446 6197 8466
rect 6217 8446 6220 8466
rect 5804 8441 6220 8446
rect 5586 8370 5623 8441
rect 5804 8440 6145 8441
rect 5738 8380 5769 8381
rect 5586 8350 5595 8370
rect 5615 8350 5623 8370
rect 5586 8340 5623 8350
rect 5682 8370 5769 8380
rect 5682 8350 5691 8370
rect 5711 8350 5769 8370
rect 5682 8341 5769 8350
rect 5682 8340 5719 8341
rect 4607 8308 4650 8313
rect 4998 8319 5445 8335
rect 4998 8313 5026 8319
rect 5277 8318 5445 8319
rect 4607 8305 4757 8308
rect 4998 8305 5025 8313
rect 4607 8303 5025 8305
rect 4607 8285 4616 8303
rect 4634 8285 5025 8303
rect 5738 8290 5769 8341
rect 5804 8370 5841 8440
rect 6107 8439 6144 8440
rect 5956 8380 5992 8381
rect 5804 8350 5813 8370
rect 5833 8350 5841 8370
rect 5804 8340 5841 8350
rect 5900 8370 6048 8380
rect 6148 8377 6244 8379
rect 5900 8350 5909 8370
rect 5929 8350 6019 8370
rect 6039 8350 6048 8370
rect 5900 8341 6048 8350
rect 6106 8370 6244 8377
rect 6106 8350 6115 8370
rect 6135 8350 6244 8370
rect 6106 8341 6244 8350
rect 5900 8340 5937 8341
rect 5630 8287 5671 8288
rect 4607 8282 5025 8285
rect 4607 8276 4650 8282
rect 4610 8273 4650 8276
rect 5522 8280 5671 8287
rect 5007 8264 5047 8265
rect 4718 8247 5047 8264
rect 5522 8260 5581 8280
rect 5601 8260 5640 8280
rect 5660 8260 5671 8280
rect 5522 8252 5671 8260
rect 5738 8283 5895 8290
rect 5738 8263 5858 8283
rect 5878 8263 5895 8283
rect 5738 8253 5895 8263
rect 5738 8252 5773 8253
rect 4602 8204 4645 8215
rect 4602 8186 4614 8204
rect 4632 8186 4645 8204
rect 4602 8160 4645 8186
rect 4718 8160 4745 8247
rect 5007 8238 5047 8247
rect 3781 8134 4220 8152
rect 3054 8129 3095 8130
rect 2788 8076 2825 8077
rect 2481 8067 2619 8076
rect 2481 8047 2590 8067
rect 2610 8047 2619 8067
rect 2481 8040 2619 8047
rect 2677 8067 2825 8076
rect 2677 8047 2686 8067
rect 2706 8047 2796 8067
rect 2816 8047 2825 8067
rect 2481 8038 2577 8040
rect 2677 8037 2825 8047
rect 2884 8067 2921 8077
rect 2884 8047 2892 8067
rect 2912 8047 2921 8067
rect 2733 8036 2769 8037
rect 2581 7977 2618 7978
rect 2884 7977 2921 8047
rect 2956 8076 2987 8127
rect 3781 8116 4181 8134
rect 4199 8116 4220 8134
rect 3781 8110 4220 8116
rect 3787 8106 4220 8110
rect 4602 8139 4745 8160
rect 4789 8212 4823 8228
rect 5007 8218 5400 8238
rect 5420 8218 5423 8238
rect 5738 8231 5769 8252
rect 5956 8231 5992 8341
rect 6011 8340 6048 8341
rect 6107 8340 6144 8341
rect 6067 8281 6157 8287
rect 6067 8261 6076 8281
rect 6096 8279 6157 8281
rect 6096 8261 6121 8279
rect 6067 8259 6121 8261
rect 6141 8259 6157 8279
rect 6067 8253 6157 8259
rect 5581 8230 5618 8231
rect 5007 8213 5423 8218
rect 5580 8221 5618 8230
rect 5007 8212 5348 8213
rect 4789 8142 4826 8212
rect 4941 8152 4972 8153
rect 4602 8137 4739 8139
rect 4166 8104 4218 8106
rect 4602 8095 4645 8137
rect 4789 8122 4798 8142
rect 4818 8122 4826 8142
rect 4789 8112 4826 8122
rect 4885 8142 4972 8152
rect 4885 8122 4894 8142
rect 4914 8122 4972 8142
rect 4885 8113 4972 8122
rect 4885 8112 4922 8113
rect 4600 8085 4645 8095
rect 3006 8076 3043 8077
rect 2956 8067 3043 8076
rect 2956 8047 3014 8067
rect 3034 8047 3043 8067
rect 2956 8037 3043 8047
rect 3102 8067 3139 8077
rect 3102 8047 3110 8067
rect 3130 8047 3139 8067
rect 4600 8067 4609 8085
rect 4627 8067 4645 8085
rect 4600 8061 4645 8067
rect 4941 8062 4972 8113
rect 5007 8142 5044 8212
rect 5310 8211 5347 8212
rect 5580 8201 5589 8221
rect 5609 8201 5618 8221
rect 5580 8193 5618 8201
rect 5684 8225 5769 8231
rect 5799 8230 5836 8231
rect 5684 8205 5692 8225
rect 5712 8205 5769 8225
rect 5684 8197 5769 8205
rect 5798 8221 5836 8230
rect 5798 8201 5807 8221
rect 5827 8201 5836 8221
rect 5684 8196 5720 8197
rect 5798 8193 5836 8201
rect 5902 8225 6046 8231
rect 5902 8205 5910 8225
rect 5930 8206 5962 8225
rect 5983 8206 6018 8225
rect 5930 8205 6018 8206
rect 6038 8205 6046 8225
rect 5902 8197 6046 8205
rect 5902 8196 5938 8197
rect 6010 8196 6046 8197
rect 6112 8230 6149 8231
rect 6112 8229 6150 8230
rect 6112 8221 6176 8229
rect 6112 8201 6121 8221
rect 6141 8207 6176 8221
rect 6196 8207 6199 8227
rect 6141 8202 6199 8207
rect 6141 8201 6176 8202
rect 5581 8164 5618 8193
rect 5582 8162 5618 8164
rect 5159 8152 5195 8153
rect 5007 8122 5016 8142
rect 5036 8122 5044 8142
rect 5007 8112 5044 8122
rect 5103 8142 5251 8152
rect 5351 8149 5447 8151
rect 5103 8122 5112 8142
rect 5132 8122 5222 8142
rect 5242 8122 5251 8142
rect 5103 8113 5251 8122
rect 5309 8142 5447 8149
rect 5309 8122 5318 8142
rect 5338 8122 5447 8142
rect 5582 8140 5773 8162
rect 5799 8161 5836 8193
rect 6112 8189 6176 8201
rect 6216 8163 6243 8341
rect 6848 8340 6881 8673
rect 6945 8705 7113 8706
rect 7239 8705 7279 8929
rect 7742 8933 7910 8934
rect 8146 8933 8195 8968
rect 7742 8907 8195 8933
rect 7742 8905 7910 8907
rect 8106 8906 8188 8907
rect 8328 8906 8406 8932
rect 8546 8910 8593 8968
rect 8994 8964 9041 8969
rect 7742 8727 7769 8905
rect 7809 8867 7873 8879
rect 8149 8875 8186 8906
rect 8367 8875 8404 8906
rect 8546 8897 8594 8910
rect 7809 8866 7844 8867
rect 7786 8861 7844 8866
rect 7786 8841 7789 8861
rect 7809 8847 7844 8861
rect 7864 8847 7873 8867
rect 7809 8839 7873 8847
rect 7835 8838 7873 8839
rect 7836 8837 7873 8838
rect 7939 8871 7975 8872
rect 8047 8871 8083 8872
rect 7939 8863 8083 8871
rect 7939 8843 7947 8863
rect 7967 8859 8055 8863
rect 7967 8843 8011 8859
rect 7939 8839 8011 8843
rect 8031 8843 8055 8859
rect 8075 8843 8083 8863
rect 8031 8839 8083 8843
rect 7939 8837 8083 8839
rect 8149 8867 8187 8875
rect 8265 8871 8301 8872
rect 8149 8847 8158 8867
rect 8178 8847 8187 8867
rect 8149 8838 8187 8847
rect 8216 8863 8301 8871
rect 8216 8843 8273 8863
rect 8293 8843 8301 8863
rect 8149 8837 8186 8838
rect 8216 8837 8301 8843
rect 8367 8867 8405 8875
rect 8367 8847 8376 8867
rect 8396 8847 8405 8867
rect 8367 8838 8405 8847
rect 8549 8872 8594 8897
rect 8549 8854 8563 8872
rect 8581 8854 8594 8872
rect 8549 8846 8594 8854
rect 8554 8844 8594 8846
rect 8994 8902 9042 8964
rect 11616 8963 11656 8971
rect 11616 8941 11624 8963
rect 11648 8941 11656 8963
rect 12520 8966 12976 9001
rect 15980 8976 16020 8984
rect 8367 8837 8404 8838
rect 7828 8809 7918 8815
rect 7828 8789 7844 8809
rect 7864 8807 7918 8809
rect 7864 8789 7889 8807
rect 7828 8787 7889 8789
rect 7909 8787 7918 8807
rect 7828 8781 7918 8787
rect 7841 8727 7878 8728
rect 7937 8727 7974 8728
rect 7993 8727 8029 8837
rect 8216 8816 8247 8837
rect 8994 8822 9041 8902
rect 8212 8815 8247 8816
rect 8090 8805 8247 8815
rect 8090 8785 8107 8805
rect 8127 8785 8247 8805
rect 8090 8778 8247 8785
rect 8314 8808 8463 8816
rect 8314 8788 8325 8808
rect 8345 8788 8384 8808
rect 8404 8788 8463 8808
rect 8994 8804 9004 8822
rect 9022 8804 9041 8822
rect 8994 8800 9041 8804
rect 8995 8795 9032 8800
rect 8314 8781 8463 8788
rect 8314 8780 8355 8781
rect 8551 8779 8588 8782
rect 8048 8727 8085 8728
rect 7741 8718 7879 8727
rect 6945 8679 7389 8705
rect 6945 8677 7113 8679
rect 6945 8499 6972 8677
rect 7012 8639 7076 8651
rect 7352 8647 7389 8679
rect 7415 8678 7606 8700
rect 7741 8698 7850 8718
rect 7870 8698 7879 8718
rect 7741 8691 7879 8698
rect 7937 8718 8085 8727
rect 7937 8698 7946 8718
rect 7966 8698 8056 8718
rect 8076 8698 8085 8718
rect 7741 8689 7837 8691
rect 7937 8688 8085 8698
rect 8144 8718 8181 8728
rect 8144 8698 8152 8718
rect 8172 8698 8181 8718
rect 7993 8687 8029 8688
rect 7570 8676 7606 8678
rect 7570 8647 7607 8676
rect 7012 8638 7047 8639
rect 6989 8633 7047 8638
rect 6989 8613 6992 8633
rect 7012 8619 7047 8633
rect 7067 8619 7076 8639
rect 7012 8613 7076 8619
rect 6989 8611 7076 8613
rect 6989 8607 7016 8611
rect 7038 8610 7076 8611
rect 7039 8609 7076 8610
rect 7142 8643 7178 8644
rect 7250 8643 7286 8644
rect 7142 8636 7286 8643
rect 7142 8635 7204 8636
rect 7142 8615 7150 8635
rect 7170 8618 7204 8635
rect 7223 8635 7286 8636
rect 7223 8618 7258 8635
rect 7170 8615 7258 8618
rect 7278 8615 7286 8635
rect 7142 8609 7286 8615
rect 7352 8639 7390 8647
rect 7468 8643 7504 8644
rect 7352 8619 7361 8639
rect 7381 8619 7390 8639
rect 7352 8610 7390 8619
rect 7419 8635 7504 8643
rect 7419 8615 7476 8635
rect 7496 8615 7504 8635
rect 7352 8609 7389 8610
rect 7419 8609 7504 8615
rect 7570 8639 7608 8647
rect 7570 8619 7579 8639
rect 7599 8619 7608 8639
rect 7841 8628 7878 8629
rect 8144 8628 8181 8698
rect 8216 8727 8247 8778
rect 8543 8773 8588 8779
rect 8543 8755 8561 8773
rect 8579 8755 8588 8773
rect 8543 8745 8588 8755
rect 8266 8727 8303 8728
rect 8216 8718 8303 8727
rect 8216 8698 8274 8718
rect 8294 8698 8303 8718
rect 8216 8688 8303 8698
rect 8362 8718 8399 8728
rect 8362 8698 8370 8718
rect 8390 8698 8399 8718
rect 8543 8703 8586 8745
rect 8983 8733 9035 8735
rect 8449 8701 8586 8703
rect 8216 8687 8247 8688
rect 8362 8628 8399 8698
rect 7840 8627 8181 8628
rect 7570 8610 7608 8619
rect 7765 8622 8181 8627
rect 7570 8609 7607 8610
rect 7031 8581 7121 8587
rect 7031 8561 7047 8581
rect 7067 8579 7121 8581
rect 7067 8561 7092 8579
rect 7031 8559 7092 8561
rect 7112 8559 7121 8579
rect 7031 8553 7121 8559
rect 7044 8499 7081 8500
rect 7140 8499 7177 8500
rect 7196 8499 7232 8609
rect 7419 8588 7450 8609
rect 7765 8602 7768 8622
rect 7788 8602 8181 8622
rect 8365 8612 8399 8628
rect 8443 8680 8586 8701
rect 8981 8729 9414 8733
rect 8981 8723 9420 8729
rect 8981 8705 9002 8723
rect 9020 8705 9420 8723
rect 8981 8687 9420 8705
rect 8141 8593 8181 8602
rect 8443 8593 8470 8680
rect 8543 8654 8586 8680
rect 8543 8636 8556 8654
rect 8574 8636 8586 8654
rect 8543 8625 8586 8636
rect 7415 8587 7450 8588
rect 7293 8577 7450 8587
rect 7293 8557 7310 8577
rect 7330 8557 7450 8577
rect 7293 8550 7450 8557
rect 7517 8580 7663 8588
rect 7517 8560 7528 8580
rect 7548 8560 7587 8580
rect 7607 8560 7663 8580
rect 8141 8576 8470 8593
rect 8141 8575 8181 8576
rect 7517 8553 7663 8560
rect 8538 8564 8578 8567
rect 8538 8558 8581 8564
rect 8163 8555 8581 8558
rect 7517 8552 7558 8553
rect 7251 8499 7288 8500
rect 6944 8490 7082 8499
rect 6944 8470 7053 8490
rect 7073 8470 7082 8490
rect 6944 8463 7082 8470
rect 7140 8490 7288 8499
rect 7140 8470 7149 8490
rect 7169 8470 7259 8490
rect 7279 8470 7288 8490
rect 6944 8461 7040 8463
rect 7140 8460 7288 8470
rect 7347 8490 7384 8500
rect 7347 8470 7355 8490
rect 7375 8470 7384 8490
rect 7196 8459 7232 8460
rect 7044 8400 7081 8401
rect 7347 8400 7384 8470
rect 7419 8499 7450 8550
rect 8163 8537 8554 8555
rect 8572 8537 8581 8555
rect 8163 8535 8581 8537
rect 8163 8527 8190 8535
rect 8431 8532 8581 8535
rect 7743 8521 7911 8522
rect 8162 8521 8190 8527
rect 7743 8505 8190 8521
rect 8538 8527 8581 8532
rect 7469 8499 7506 8500
rect 7419 8490 7506 8499
rect 7419 8470 7477 8490
rect 7497 8470 7506 8490
rect 7419 8460 7506 8470
rect 7565 8490 7602 8500
rect 7565 8470 7573 8490
rect 7593 8470 7602 8490
rect 7419 8459 7450 8460
rect 7043 8399 7384 8400
rect 7565 8399 7602 8470
rect 6968 8394 7384 8399
rect 6968 8374 6971 8394
rect 6991 8374 7384 8394
rect 7415 8375 7602 8399
rect 7743 8495 8187 8505
rect 7743 8493 7911 8495
rect 6843 8295 6885 8340
rect 7743 8315 7770 8493
rect 7810 8455 7874 8467
rect 8150 8463 8187 8495
rect 8213 8494 8404 8516
rect 8368 8492 8404 8494
rect 8368 8463 8405 8492
rect 8538 8471 8578 8527
rect 7810 8454 7845 8455
rect 7787 8449 7845 8454
rect 7787 8429 7790 8449
rect 7810 8435 7845 8449
rect 7865 8435 7874 8455
rect 7810 8427 7874 8435
rect 7836 8426 7874 8427
rect 7837 8425 7874 8426
rect 7940 8459 7976 8460
rect 8048 8459 8084 8460
rect 7940 8451 8084 8459
rect 7940 8431 7948 8451
rect 7968 8431 8003 8451
rect 8023 8431 8056 8451
rect 8076 8431 8084 8451
rect 7940 8425 8084 8431
rect 8150 8455 8188 8463
rect 8266 8459 8302 8460
rect 8150 8435 8159 8455
rect 8179 8435 8188 8455
rect 8150 8426 8188 8435
rect 8217 8451 8302 8459
rect 8217 8431 8274 8451
rect 8294 8431 8302 8451
rect 8150 8425 8187 8426
rect 8217 8425 8302 8431
rect 8368 8455 8406 8463
rect 8368 8435 8377 8455
rect 8397 8435 8406 8455
rect 8538 8453 8550 8471
rect 8568 8453 8578 8471
rect 8983 8498 9035 8687
rect 9381 8662 9420 8687
rect 11221 8712 11258 8718
rect 11221 8693 11229 8712
rect 11250 8693 11258 8712
rect 11221 8685 11258 8693
rect 9165 8637 9352 8661
rect 9381 8642 9776 8662
rect 9796 8642 9799 8662
rect 9381 8637 9799 8642
rect 9165 8566 9202 8637
rect 9381 8636 9724 8637
rect 9381 8633 9420 8636
rect 9686 8635 9723 8636
rect 9317 8576 9348 8577
rect 9165 8546 9174 8566
rect 9194 8546 9202 8566
rect 9165 8536 9202 8546
rect 9261 8566 9348 8576
rect 9261 8546 9270 8566
rect 9290 8546 9348 8566
rect 9261 8537 9348 8546
rect 9261 8536 9298 8537
rect 8983 8480 8999 8498
rect 9017 8480 9035 8498
rect 9317 8486 9348 8537
rect 9383 8566 9420 8633
rect 9535 8576 9571 8577
rect 9383 8546 9392 8566
rect 9412 8546 9420 8566
rect 9383 8536 9420 8546
rect 9479 8566 9627 8576
rect 9727 8573 9823 8575
rect 9479 8546 9488 8566
rect 9508 8546 9598 8566
rect 9618 8546 9627 8566
rect 9479 8537 9627 8546
rect 9685 8566 9823 8573
rect 9685 8546 9694 8566
rect 9714 8546 9823 8566
rect 9685 8537 9823 8546
rect 9479 8536 9516 8537
rect 9209 8483 9250 8484
rect 8983 8462 9035 8480
rect 9101 8476 9250 8483
rect 8538 8443 8578 8453
rect 9101 8456 9160 8476
rect 9180 8456 9219 8476
rect 9239 8456 9250 8476
rect 9101 8448 9250 8456
rect 9317 8479 9474 8486
rect 9317 8459 9437 8479
rect 9457 8459 9474 8479
rect 9317 8449 9474 8459
rect 9317 8448 9352 8449
rect 8368 8426 8406 8435
rect 9317 8427 9348 8448
rect 9535 8427 9571 8537
rect 9590 8536 9627 8537
rect 9686 8536 9723 8537
rect 9646 8477 9736 8483
rect 9646 8457 9655 8477
rect 9675 8475 9736 8477
rect 9675 8457 9700 8475
rect 9646 8455 9700 8457
rect 9720 8455 9736 8475
rect 9646 8449 9736 8455
rect 9160 8426 9197 8427
rect 8368 8425 8405 8426
rect 7829 8397 7919 8403
rect 7829 8377 7845 8397
rect 7865 8395 7919 8397
rect 7865 8377 7890 8395
rect 7829 8375 7890 8377
rect 7910 8375 7919 8395
rect 7829 8369 7919 8375
rect 7842 8315 7879 8316
rect 7938 8315 7975 8316
rect 7994 8315 8030 8425
rect 8217 8404 8248 8425
rect 9159 8417 9197 8426
rect 8213 8403 8248 8404
rect 8091 8393 8248 8403
rect 8091 8373 8108 8393
rect 8128 8373 8248 8393
rect 8091 8366 8248 8373
rect 8315 8396 8464 8404
rect 8315 8376 8326 8396
rect 8346 8376 8385 8396
rect 8405 8376 8464 8396
rect 8987 8399 9027 8409
rect 8315 8369 8464 8376
rect 8530 8372 8582 8390
rect 8315 8368 8356 8369
rect 8049 8315 8086 8316
rect 7742 8306 7880 8315
rect 7214 8295 7247 8297
rect 6843 8283 7290 8295
rect 6075 8161 6243 8163
rect 5799 8135 6243 8161
rect 5309 8113 5447 8122
rect 5103 8112 5140 8113
rect 4600 8058 4637 8061
rect 4833 8059 4874 8060
rect 2956 8036 2987 8037
rect 2580 7976 2921 7977
rect 3102 7976 3139 8047
rect 4725 8052 4874 8059
rect 4169 8039 4206 8044
rect 4160 8035 4207 8039
rect 4160 8017 4179 8035
rect 4197 8017 4207 8035
rect 4725 8032 4784 8052
rect 4804 8032 4843 8052
rect 4863 8032 4874 8052
rect 4725 8024 4874 8032
rect 4941 8055 5098 8062
rect 4941 8035 5061 8055
rect 5081 8035 5098 8055
rect 4941 8025 5098 8035
rect 4941 8024 4976 8025
rect 2505 7971 2921 7976
rect 2505 7951 2508 7971
rect 2528 7951 2921 7971
rect 2952 7952 3139 7976
rect 3764 7974 3804 7979
rect 4160 7974 4207 8017
rect 4941 8003 4972 8024
rect 5159 8003 5195 8113
rect 5214 8112 5251 8113
rect 5310 8112 5347 8113
rect 5270 8053 5360 8059
rect 5270 8033 5279 8053
rect 5299 8051 5360 8053
rect 5299 8033 5324 8051
rect 5270 8031 5324 8033
rect 5344 8031 5360 8051
rect 5270 8025 5360 8031
rect 4784 8002 4821 8003
rect 3764 7935 4207 7974
rect 4597 7994 4634 7996
rect 4597 7986 4639 7994
rect 4597 7968 4607 7986
rect 4625 7968 4639 7986
rect 4597 7959 4639 7968
rect 4783 7993 4821 8002
rect 4783 7973 4792 7993
rect 4812 7973 4821 7993
rect 4783 7965 4821 7973
rect 4887 7997 4972 8003
rect 5002 8002 5039 8003
rect 4887 7977 4895 7997
rect 4915 7977 4972 7997
rect 4887 7969 4972 7977
rect 5001 7993 5039 8002
rect 5001 7973 5010 7993
rect 5030 7973 5039 7993
rect 4887 7968 4923 7969
rect 5001 7965 5039 7973
rect 5105 8001 5249 8003
rect 5105 7997 5157 8001
rect 5105 7977 5113 7997
rect 5133 7981 5157 7997
rect 5177 7997 5249 8001
rect 5177 7981 5221 7997
rect 5133 7977 5221 7981
rect 5241 7977 5249 7997
rect 5105 7969 5249 7977
rect 5105 7968 5141 7969
rect 5213 7968 5249 7969
rect 5315 8002 5352 8003
rect 5315 8001 5353 8002
rect 5315 7993 5379 8001
rect 5315 7973 5324 7993
rect 5344 7979 5379 7993
rect 5399 7979 5402 7999
rect 5344 7974 5402 7979
rect 5344 7973 5379 7974
rect 1545 7876 1553 7898
rect 1577 7876 1585 7898
rect 1545 7868 1585 7876
rect 2858 7920 2898 7928
rect 2858 7898 2866 7920
rect 2890 7898 2898 7920
rect 236 7822 679 7861
rect 236 7779 283 7822
rect 639 7817 679 7822
rect 1304 7820 1491 7844
rect 1522 7825 1915 7845
rect 1935 7825 1938 7845
rect 1522 7820 1938 7825
rect 236 7761 246 7779
rect 264 7761 283 7779
rect 236 7757 283 7761
rect 237 7752 274 7757
rect 1304 7749 1341 7820
rect 1522 7819 1863 7820
rect 1456 7759 1487 7760
rect 1304 7729 1313 7749
rect 1333 7729 1341 7749
rect 1304 7719 1341 7729
rect 1400 7749 1487 7759
rect 1400 7729 1409 7749
rect 1429 7729 1487 7749
rect 1400 7720 1487 7729
rect 1400 7719 1437 7720
rect 225 7690 277 7692
rect 223 7686 656 7690
rect 223 7680 662 7686
rect 223 7662 244 7680
rect 262 7662 662 7680
rect 1456 7669 1487 7720
rect 1522 7749 1559 7819
rect 1825 7818 1862 7819
rect 1674 7759 1710 7760
rect 1522 7729 1531 7749
rect 1551 7729 1559 7749
rect 1522 7719 1559 7729
rect 1618 7749 1766 7759
rect 1866 7756 1962 7758
rect 1618 7729 1627 7749
rect 1647 7729 1737 7749
rect 1757 7729 1766 7749
rect 1618 7720 1766 7729
rect 1824 7749 1962 7756
rect 1824 7729 1833 7749
rect 1853 7729 1962 7749
rect 1824 7720 1962 7729
rect 1618 7719 1655 7720
rect 1348 7666 1389 7667
rect 223 7644 662 7662
rect 225 7455 277 7644
rect 623 7619 662 7644
rect 1240 7659 1389 7666
rect 1240 7639 1299 7659
rect 1319 7639 1358 7659
rect 1378 7639 1389 7659
rect 1240 7631 1389 7639
rect 1456 7662 1613 7669
rect 1456 7642 1576 7662
rect 1596 7642 1613 7662
rect 1456 7632 1613 7642
rect 1456 7631 1491 7632
rect 407 7594 594 7618
rect 623 7599 1018 7619
rect 1038 7599 1041 7619
rect 1456 7610 1487 7631
rect 1674 7610 1710 7720
rect 1729 7719 1766 7720
rect 1825 7719 1862 7720
rect 1785 7660 1875 7666
rect 1785 7640 1794 7660
rect 1814 7658 1875 7660
rect 1814 7640 1839 7658
rect 1785 7638 1839 7640
rect 1859 7638 1875 7658
rect 1785 7632 1875 7638
rect 1299 7609 1336 7610
rect 623 7594 1041 7599
rect 1298 7600 1336 7609
rect 407 7523 444 7594
rect 623 7593 966 7594
rect 623 7590 662 7593
rect 928 7592 965 7593
rect 559 7533 590 7534
rect 407 7503 416 7523
rect 436 7503 444 7523
rect 407 7493 444 7503
rect 503 7523 590 7533
rect 503 7503 512 7523
rect 532 7503 590 7523
rect 503 7494 590 7503
rect 503 7493 540 7494
rect 225 7437 241 7455
rect 259 7437 277 7455
rect 559 7443 590 7494
rect 625 7523 662 7590
rect 1298 7580 1307 7600
rect 1327 7580 1336 7600
rect 1298 7572 1336 7580
rect 1402 7604 1487 7610
rect 1517 7609 1554 7610
rect 1402 7584 1410 7604
rect 1430 7584 1487 7604
rect 1402 7576 1487 7584
rect 1516 7600 1554 7609
rect 1516 7580 1525 7600
rect 1545 7580 1554 7600
rect 1402 7575 1438 7576
rect 1516 7572 1554 7580
rect 1620 7605 1764 7610
rect 1620 7604 1682 7605
rect 1620 7584 1628 7604
rect 1648 7586 1682 7604
rect 1703 7604 1764 7605
rect 1703 7586 1736 7604
rect 1648 7584 1736 7586
rect 1756 7584 1764 7604
rect 1620 7576 1764 7584
rect 1620 7575 1656 7576
rect 1728 7575 1764 7576
rect 1830 7609 1867 7610
rect 1830 7608 1868 7609
rect 1830 7600 1894 7608
rect 1830 7580 1839 7600
rect 1859 7586 1894 7600
rect 1914 7586 1917 7606
rect 1859 7581 1917 7586
rect 1859 7580 1894 7581
rect 1299 7543 1336 7572
rect 1300 7541 1336 7543
rect 777 7533 813 7534
rect 625 7503 634 7523
rect 654 7503 662 7523
rect 625 7493 662 7503
rect 721 7523 869 7533
rect 969 7530 1065 7532
rect 721 7503 730 7523
rect 750 7503 840 7523
rect 860 7503 869 7523
rect 721 7494 869 7503
rect 927 7523 1065 7530
rect 927 7503 936 7523
rect 956 7503 1065 7523
rect 1300 7519 1491 7541
rect 1517 7540 1554 7572
rect 1830 7568 1894 7580
rect 1934 7542 1961 7720
rect 1793 7540 1961 7542
rect 1517 7526 1961 7540
rect 2564 7674 2732 7675
rect 2858 7674 2898 7898
rect 3361 7902 3529 7903
rect 3764 7902 3804 7935
rect 4160 7902 4207 7935
rect 4598 7934 4639 7959
rect 4784 7934 4821 7965
rect 5002 7934 5039 7965
rect 5315 7961 5379 7973
rect 5419 7935 5446 8113
rect 4598 7907 4647 7934
rect 4783 7908 4832 7934
rect 5001 7933 5082 7934
rect 5278 7933 5446 7935
rect 5001 7908 5446 7933
rect 5002 7907 5446 7908
rect 3361 7901 3805 7902
rect 3361 7876 3806 7901
rect 3361 7874 3529 7876
rect 3725 7875 3806 7876
rect 3975 7875 4024 7901
rect 4160 7875 4209 7902
rect 3361 7696 3388 7874
rect 3428 7836 3492 7848
rect 3768 7844 3805 7875
rect 3986 7844 4023 7875
rect 4168 7850 4209 7875
rect 4600 7874 4647 7907
rect 5003 7874 5043 7907
rect 5278 7906 5446 7907
rect 5909 7911 5949 8135
rect 6075 8134 6243 8135
rect 6846 8269 7290 8283
rect 6846 8267 7014 8269
rect 6846 8089 6873 8267
rect 6913 8229 6977 8241
rect 7253 8237 7290 8269
rect 7316 8268 7507 8290
rect 7742 8286 7851 8306
rect 7871 8286 7880 8306
rect 7742 8279 7880 8286
rect 7938 8306 8086 8315
rect 7938 8286 7947 8306
rect 7967 8286 8057 8306
rect 8077 8286 8086 8306
rect 7742 8277 7838 8279
rect 7938 8276 8086 8286
rect 8145 8306 8182 8316
rect 8145 8286 8153 8306
rect 8173 8286 8182 8306
rect 7994 8275 8030 8276
rect 7471 8266 7507 8268
rect 7471 8237 7508 8266
rect 6913 8228 6948 8229
rect 6890 8223 6948 8228
rect 6890 8203 6893 8223
rect 6913 8209 6948 8223
rect 6968 8209 6977 8229
rect 6913 8201 6977 8209
rect 6939 8200 6977 8201
rect 6940 8199 6977 8200
rect 7043 8233 7079 8234
rect 7151 8233 7187 8234
rect 7043 8227 7187 8233
rect 7043 8225 7104 8227
rect 7043 8205 7051 8225
rect 7071 8210 7104 8225
rect 7123 8225 7187 8227
rect 7123 8210 7159 8225
rect 7071 8205 7159 8210
rect 7179 8205 7187 8225
rect 7043 8199 7187 8205
rect 7253 8229 7291 8237
rect 7369 8233 7405 8234
rect 7253 8209 7262 8229
rect 7282 8209 7291 8229
rect 7253 8200 7291 8209
rect 7320 8225 7405 8233
rect 7320 8205 7377 8225
rect 7397 8205 7405 8225
rect 7253 8199 7290 8200
rect 7320 8199 7405 8205
rect 7471 8229 7509 8237
rect 7471 8209 7480 8229
rect 7500 8209 7509 8229
rect 8145 8219 8182 8286
rect 8217 8315 8248 8366
rect 8530 8354 8548 8372
rect 8566 8354 8582 8372
rect 8267 8315 8304 8316
rect 8217 8306 8304 8315
rect 8217 8286 8275 8306
rect 8295 8286 8304 8306
rect 8217 8276 8304 8286
rect 8363 8306 8400 8316
rect 8363 8286 8371 8306
rect 8391 8286 8400 8306
rect 8217 8275 8248 8276
rect 7842 8216 7879 8217
rect 8145 8216 8184 8219
rect 7841 8215 8184 8216
rect 8363 8215 8400 8286
rect 7471 8200 7509 8209
rect 7766 8210 8184 8215
rect 7471 8199 7508 8200
rect 6932 8171 7022 8177
rect 6932 8151 6948 8171
rect 6968 8169 7022 8171
rect 6968 8151 6993 8169
rect 6932 8149 6993 8151
rect 7013 8149 7022 8169
rect 6932 8143 7022 8149
rect 6945 8089 6982 8090
rect 7041 8089 7078 8090
rect 7097 8089 7133 8199
rect 7320 8178 7351 8199
rect 7766 8190 7769 8210
rect 7789 8190 8184 8210
rect 8213 8191 8400 8215
rect 7316 8177 7351 8178
rect 7194 8167 7351 8177
rect 7194 8147 7211 8167
rect 7231 8147 7351 8167
rect 7194 8140 7351 8147
rect 7418 8170 7567 8178
rect 7418 8150 7429 8170
rect 7449 8150 7488 8170
rect 7508 8150 7567 8170
rect 7418 8143 7567 8150
rect 8145 8165 8184 8190
rect 8530 8165 8582 8354
rect 8987 8381 8997 8399
rect 9015 8381 9027 8399
rect 9159 8397 9168 8417
rect 9188 8397 9197 8417
rect 9159 8389 9197 8397
rect 9263 8421 9348 8427
rect 9378 8426 9415 8427
rect 9263 8401 9271 8421
rect 9291 8401 9348 8421
rect 9263 8393 9348 8401
rect 9377 8417 9415 8426
rect 9377 8397 9386 8417
rect 9406 8397 9415 8417
rect 9263 8392 9299 8393
rect 9377 8389 9415 8397
rect 9481 8421 9625 8427
rect 9481 8401 9489 8421
rect 9509 8401 9542 8421
rect 9562 8401 9597 8421
rect 9617 8401 9625 8421
rect 9481 8393 9625 8401
rect 9481 8392 9517 8393
rect 9589 8392 9625 8393
rect 9691 8426 9728 8427
rect 9691 8425 9729 8426
rect 9691 8417 9755 8425
rect 9691 8397 9700 8417
rect 9720 8403 9755 8417
rect 9775 8403 9778 8423
rect 9720 8398 9778 8403
rect 9720 8397 9755 8398
rect 8987 8325 9027 8381
rect 9160 8360 9197 8389
rect 9161 8358 9197 8360
rect 9161 8336 9352 8358
rect 9378 8357 9415 8389
rect 9691 8385 9755 8397
rect 9795 8359 9822 8537
rect 9654 8357 9822 8359
rect 9378 8347 9822 8357
rect 9963 8453 10150 8477
rect 10181 8458 10574 8478
rect 10594 8458 10597 8478
rect 10181 8453 10597 8458
rect 9963 8382 10000 8453
rect 10181 8452 10522 8453
rect 10115 8392 10146 8393
rect 9963 8362 9972 8382
rect 9992 8362 10000 8382
rect 9963 8352 10000 8362
rect 10059 8382 10146 8392
rect 10059 8362 10068 8382
rect 10088 8362 10146 8382
rect 10059 8353 10146 8362
rect 10059 8352 10096 8353
rect 8984 8320 9027 8325
rect 9375 8331 9822 8347
rect 9375 8325 9403 8331
rect 9654 8330 9822 8331
rect 8984 8317 9134 8320
rect 9375 8317 9402 8325
rect 8984 8315 9402 8317
rect 8984 8297 8993 8315
rect 9011 8297 9402 8315
rect 10115 8302 10146 8353
rect 10181 8382 10218 8452
rect 10484 8451 10521 8452
rect 10333 8392 10369 8393
rect 10181 8362 10190 8382
rect 10210 8362 10218 8382
rect 10181 8352 10218 8362
rect 10277 8382 10425 8392
rect 10525 8389 10621 8391
rect 10277 8362 10286 8382
rect 10306 8362 10396 8382
rect 10416 8362 10425 8382
rect 10277 8353 10425 8362
rect 10483 8382 10621 8389
rect 10483 8362 10492 8382
rect 10512 8362 10621 8382
rect 10483 8353 10621 8362
rect 10277 8352 10314 8353
rect 10007 8299 10048 8300
rect 8984 8294 9402 8297
rect 8984 8288 9027 8294
rect 8987 8285 9027 8288
rect 9899 8292 10048 8299
rect 9384 8276 9424 8277
rect 9095 8259 9424 8276
rect 9899 8272 9958 8292
rect 9978 8272 10017 8292
rect 10037 8272 10048 8292
rect 9899 8264 10048 8272
rect 10115 8295 10272 8302
rect 10115 8275 10235 8295
rect 10255 8275 10272 8295
rect 10115 8265 10272 8275
rect 10115 8264 10150 8265
rect 8979 8216 9022 8227
rect 8979 8198 8991 8216
rect 9009 8198 9022 8216
rect 8979 8172 9022 8198
rect 9095 8172 9122 8259
rect 9384 8250 9424 8259
rect 8145 8147 8584 8165
rect 7418 8142 7459 8143
rect 7152 8089 7189 8090
rect 6845 8080 6983 8089
rect 6845 8060 6954 8080
rect 6974 8060 6983 8080
rect 6845 8053 6983 8060
rect 7041 8080 7189 8089
rect 7041 8060 7050 8080
rect 7070 8060 7160 8080
rect 7180 8060 7189 8080
rect 6845 8051 6941 8053
rect 7041 8050 7189 8060
rect 7248 8080 7285 8090
rect 7248 8060 7256 8080
rect 7276 8060 7285 8080
rect 7097 8049 7133 8050
rect 6945 7990 6982 7991
rect 7248 7990 7285 8060
rect 7320 8089 7351 8140
rect 8145 8129 8545 8147
rect 8563 8129 8584 8147
rect 8145 8123 8584 8129
rect 8151 8119 8584 8123
rect 8979 8151 9122 8172
rect 9166 8224 9200 8240
rect 9384 8230 9777 8250
rect 9797 8230 9800 8250
rect 10115 8243 10146 8264
rect 10333 8243 10369 8353
rect 10388 8352 10425 8353
rect 10484 8352 10521 8353
rect 10444 8293 10534 8299
rect 10444 8273 10453 8293
rect 10473 8291 10534 8293
rect 10473 8273 10498 8291
rect 10444 8271 10498 8273
rect 10518 8271 10534 8291
rect 10444 8265 10534 8271
rect 9958 8242 9995 8243
rect 9384 8225 9800 8230
rect 9957 8233 9995 8242
rect 9384 8224 9725 8225
rect 9166 8154 9203 8224
rect 9318 8164 9349 8165
rect 8979 8149 9116 8151
rect 8530 8117 8582 8119
rect 8979 8107 9022 8149
rect 9166 8134 9175 8154
rect 9195 8134 9203 8154
rect 9166 8124 9203 8134
rect 9262 8154 9349 8164
rect 9262 8134 9271 8154
rect 9291 8134 9349 8154
rect 9262 8125 9349 8134
rect 9262 8124 9299 8125
rect 8977 8097 9022 8107
rect 7370 8089 7407 8090
rect 7320 8080 7407 8089
rect 7320 8060 7378 8080
rect 7398 8060 7407 8080
rect 7320 8050 7407 8060
rect 7466 8080 7503 8090
rect 7466 8060 7474 8080
rect 7494 8060 7503 8080
rect 8977 8079 8986 8097
rect 9004 8079 9022 8097
rect 8977 8073 9022 8079
rect 9318 8074 9349 8125
rect 9384 8154 9421 8224
rect 9687 8223 9724 8224
rect 9957 8213 9966 8233
rect 9986 8213 9995 8233
rect 9957 8205 9995 8213
rect 10061 8237 10146 8243
rect 10176 8242 10213 8243
rect 10061 8217 10069 8237
rect 10089 8217 10146 8237
rect 10061 8209 10146 8217
rect 10175 8233 10213 8242
rect 10175 8213 10184 8233
rect 10204 8213 10213 8233
rect 10061 8208 10097 8209
rect 10175 8205 10213 8213
rect 10279 8237 10423 8243
rect 10279 8217 10287 8237
rect 10307 8218 10339 8237
rect 10360 8218 10395 8237
rect 10307 8217 10395 8218
rect 10415 8217 10423 8237
rect 10279 8209 10423 8217
rect 10279 8208 10315 8209
rect 10387 8208 10423 8209
rect 10489 8242 10526 8243
rect 10489 8241 10527 8242
rect 10489 8233 10553 8241
rect 10489 8213 10498 8233
rect 10518 8219 10553 8233
rect 10573 8219 10576 8239
rect 10518 8214 10576 8219
rect 10518 8213 10553 8214
rect 9958 8176 9995 8205
rect 9959 8174 9995 8176
rect 9536 8164 9572 8165
rect 9384 8134 9393 8154
rect 9413 8134 9421 8154
rect 9384 8124 9421 8134
rect 9480 8154 9628 8164
rect 9728 8161 9824 8163
rect 9480 8134 9489 8154
rect 9509 8134 9599 8154
rect 9619 8134 9628 8154
rect 9480 8125 9628 8134
rect 9686 8154 9824 8161
rect 9686 8134 9695 8154
rect 9715 8134 9824 8154
rect 9959 8152 10150 8174
rect 10176 8173 10213 8205
rect 10489 8201 10553 8213
rect 10593 8175 10620 8353
rect 11225 8352 11258 8685
rect 11322 8717 11490 8718
rect 11616 8717 11656 8941
rect 12119 8945 12287 8946
rect 12520 8945 12565 8966
rect 12119 8919 12565 8945
rect 12119 8917 12287 8919
rect 12483 8918 12565 8919
rect 12700 8918 12781 8944
rect 12925 8931 13406 8966
rect 15980 8954 15988 8976
rect 16012 8954 16020 8976
rect 12119 8739 12146 8917
rect 12186 8879 12250 8891
rect 12526 8887 12563 8918
rect 12744 8887 12781 8918
rect 12928 8912 12967 8931
rect 12926 8893 12967 8912
rect 12186 8878 12221 8879
rect 12163 8873 12221 8878
rect 12163 8853 12166 8873
rect 12186 8859 12221 8873
rect 12241 8859 12250 8879
rect 12186 8851 12250 8859
rect 12212 8850 12250 8851
rect 12213 8849 12250 8850
rect 12316 8883 12352 8884
rect 12424 8883 12460 8884
rect 12316 8875 12460 8883
rect 12316 8855 12324 8875
rect 12344 8871 12432 8875
rect 12344 8855 12388 8871
rect 12316 8851 12388 8855
rect 12408 8855 12432 8871
rect 12452 8855 12460 8875
rect 12408 8851 12460 8855
rect 12316 8849 12460 8851
rect 12526 8879 12564 8887
rect 12642 8883 12678 8884
rect 12526 8859 12535 8879
rect 12555 8859 12564 8879
rect 12526 8850 12564 8859
rect 12593 8875 12678 8883
rect 12593 8855 12650 8875
rect 12670 8855 12678 8875
rect 12526 8849 12563 8850
rect 12593 8849 12678 8855
rect 12744 8879 12782 8887
rect 12744 8859 12753 8879
rect 12773 8859 12782 8879
rect 12744 8850 12782 8859
rect 12926 8884 12968 8893
rect 12926 8866 12940 8884
rect 12958 8866 12968 8884
rect 12926 8858 12968 8866
rect 12931 8856 12968 8858
rect 12744 8849 12781 8850
rect 12205 8821 12295 8827
rect 12205 8801 12221 8821
rect 12241 8819 12295 8821
rect 12241 8801 12266 8819
rect 12205 8799 12266 8801
rect 12286 8799 12295 8819
rect 12205 8793 12295 8799
rect 12218 8739 12255 8740
rect 12314 8739 12351 8740
rect 12370 8739 12406 8849
rect 12593 8828 12624 8849
rect 13358 8835 13405 8931
rect 12589 8827 12624 8828
rect 12467 8817 12624 8827
rect 12467 8797 12484 8817
rect 12504 8797 12624 8817
rect 12467 8790 12624 8797
rect 12691 8820 12840 8828
rect 12691 8800 12702 8820
rect 12722 8800 12761 8820
rect 12781 8800 12840 8820
rect 13358 8817 13368 8835
rect 13386 8817 13405 8835
rect 13358 8813 13405 8817
rect 13359 8808 13396 8813
rect 12691 8793 12840 8800
rect 12691 8792 12732 8793
rect 12928 8791 12965 8794
rect 12425 8739 12462 8740
rect 12118 8730 12256 8739
rect 11322 8691 11766 8717
rect 11322 8689 11490 8691
rect 11322 8511 11349 8689
rect 11389 8651 11453 8663
rect 11729 8659 11766 8691
rect 11792 8690 11983 8712
rect 12118 8710 12227 8730
rect 12247 8710 12256 8730
rect 12118 8703 12256 8710
rect 12314 8730 12462 8739
rect 12314 8710 12323 8730
rect 12343 8710 12433 8730
rect 12453 8710 12462 8730
rect 12118 8701 12214 8703
rect 12314 8700 12462 8710
rect 12521 8730 12558 8740
rect 12521 8710 12529 8730
rect 12549 8710 12558 8730
rect 12370 8699 12406 8700
rect 11947 8688 11983 8690
rect 11947 8659 11984 8688
rect 11389 8650 11424 8651
rect 11366 8645 11424 8650
rect 11366 8625 11369 8645
rect 11389 8631 11424 8645
rect 11444 8631 11453 8651
rect 11389 8625 11453 8631
rect 11366 8623 11453 8625
rect 11366 8619 11393 8623
rect 11415 8622 11453 8623
rect 11416 8621 11453 8622
rect 11519 8655 11555 8656
rect 11627 8655 11663 8656
rect 11519 8648 11663 8655
rect 11519 8647 11581 8648
rect 11519 8627 11527 8647
rect 11547 8630 11581 8647
rect 11600 8647 11663 8648
rect 11600 8630 11635 8647
rect 11547 8627 11635 8630
rect 11655 8627 11663 8647
rect 11519 8621 11663 8627
rect 11729 8651 11767 8659
rect 11845 8655 11881 8656
rect 11729 8631 11738 8651
rect 11758 8631 11767 8651
rect 11729 8622 11767 8631
rect 11796 8647 11881 8655
rect 11796 8627 11853 8647
rect 11873 8627 11881 8647
rect 11729 8621 11766 8622
rect 11796 8621 11881 8627
rect 11947 8651 11985 8659
rect 11947 8631 11956 8651
rect 11976 8631 11985 8651
rect 12218 8640 12255 8641
rect 12521 8640 12558 8710
rect 12593 8739 12624 8790
rect 12920 8785 12965 8791
rect 12920 8767 12938 8785
rect 12956 8767 12965 8785
rect 12920 8757 12965 8767
rect 12643 8739 12680 8740
rect 12593 8730 12680 8739
rect 12593 8710 12651 8730
rect 12671 8710 12680 8730
rect 12593 8700 12680 8710
rect 12739 8730 12776 8740
rect 12739 8710 12747 8730
rect 12767 8710 12776 8730
rect 12920 8715 12963 8757
rect 13347 8746 13399 8748
rect 12826 8713 12963 8715
rect 12593 8699 12624 8700
rect 12739 8640 12776 8710
rect 12217 8639 12558 8640
rect 11947 8622 11985 8631
rect 12142 8634 12558 8639
rect 11947 8621 11984 8622
rect 11408 8593 11498 8599
rect 11408 8573 11424 8593
rect 11444 8591 11498 8593
rect 11444 8573 11469 8591
rect 11408 8571 11469 8573
rect 11489 8571 11498 8591
rect 11408 8565 11498 8571
rect 11421 8511 11458 8512
rect 11517 8511 11554 8512
rect 11573 8511 11609 8621
rect 11796 8600 11827 8621
rect 12142 8614 12145 8634
rect 12165 8614 12558 8634
rect 12742 8624 12776 8640
rect 12820 8692 12963 8713
rect 13345 8742 13778 8746
rect 13345 8736 13784 8742
rect 13345 8718 13366 8736
rect 13384 8718 13784 8736
rect 13345 8700 13784 8718
rect 12518 8605 12558 8614
rect 12820 8605 12847 8692
rect 12920 8666 12963 8692
rect 12920 8648 12933 8666
rect 12951 8648 12963 8666
rect 12920 8637 12963 8648
rect 11792 8599 11827 8600
rect 11670 8589 11827 8599
rect 11670 8569 11687 8589
rect 11707 8569 11827 8589
rect 11670 8562 11827 8569
rect 11894 8592 12040 8600
rect 11894 8572 11905 8592
rect 11925 8572 11964 8592
rect 11984 8572 12040 8592
rect 12518 8588 12847 8605
rect 12518 8587 12558 8588
rect 11894 8565 12040 8572
rect 12915 8576 12955 8579
rect 12915 8570 12958 8576
rect 12540 8567 12958 8570
rect 11894 8564 11935 8565
rect 11628 8511 11665 8512
rect 11321 8502 11459 8511
rect 11321 8482 11430 8502
rect 11450 8482 11459 8502
rect 11321 8475 11459 8482
rect 11517 8502 11665 8511
rect 11517 8482 11526 8502
rect 11546 8482 11636 8502
rect 11656 8482 11665 8502
rect 11321 8473 11417 8475
rect 11517 8472 11665 8482
rect 11724 8502 11761 8512
rect 11724 8482 11732 8502
rect 11752 8482 11761 8502
rect 11573 8471 11609 8472
rect 11421 8412 11458 8413
rect 11724 8412 11761 8482
rect 11796 8511 11827 8562
rect 12540 8549 12931 8567
rect 12949 8549 12958 8567
rect 12540 8547 12958 8549
rect 12540 8539 12567 8547
rect 12808 8544 12958 8547
rect 12120 8533 12288 8534
rect 12539 8533 12567 8539
rect 12120 8517 12567 8533
rect 12915 8539 12958 8544
rect 11846 8511 11883 8512
rect 11796 8502 11883 8511
rect 11796 8482 11854 8502
rect 11874 8482 11883 8502
rect 11796 8472 11883 8482
rect 11942 8502 11979 8512
rect 11942 8482 11950 8502
rect 11970 8482 11979 8502
rect 11796 8471 11827 8472
rect 11420 8411 11761 8412
rect 11942 8411 11979 8482
rect 11345 8406 11761 8411
rect 11345 8386 11348 8406
rect 11368 8386 11761 8406
rect 11792 8387 11979 8411
rect 12120 8507 12564 8517
rect 12120 8505 12288 8507
rect 11220 8307 11262 8352
rect 12120 8327 12147 8505
rect 12187 8467 12251 8479
rect 12527 8475 12564 8507
rect 12590 8506 12781 8528
rect 12745 8504 12781 8506
rect 12745 8475 12782 8504
rect 12915 8483 12955 8539
rect 12187 8466 12222 8467
rect 12164 8461 12222 8466
rect 12164 8441 12167 8461
rect 12187 8447 12222 8461
rect 12242 8447 12251 8467
rect 12187 8439 12251 8447
rect 12213 8438 12251 8439
rect 12214 8437 12251 8438
rect 12317 8471 12353 8472
rect 12425 8471 12461 8472
rect 12317 8463 12461 8471
rect 12317 8443 12325 8463
rect 12345 8443 12380 8463
rect 12400 8443 12433 8463
rect 12453 8443 12461 8463
rect 12317 8437 12461 8443
rect 12527 8467 12565 8475
rect 12643 8471 12679 8472
rect 12527 8447 12536 8467
rect 12556 8447 12565 8467
rect 12527 8438 12565 8447
rect 12594 8463 12679 8471
rect 12594 8443 12651 8463
rect 12671 8443 12679 8463
rect 12527 8437 12564 8438
rect 12594 8437 12679 8443
rect 12745 8467 12783 8475
rect 12745 8447 12754 8467
rect 12774 8447 12783 8467
rect 12915 8465 12927 8483
rect 12945 8465 12955 8483
rect 13347 8511 13399 8700
rect 13745 8675 13784 8700
rect 15585 8725 15622 8731
rect 15585 8706 15593 8725
rect 15614 8706 15622 8725
rect 15585 8698 15622 8706
rect 13529 8650 13716 8674
rect 13745 8655 14140 8675
rect 14160 8655 14163 8675
rect 13745 8650 14163 8655
rect 13529 8579 13566 8650
rect 13745 8649 14088 8650
rect 13745 8646 13784 8649
rect 14050 8648 14087 8649
rect 13681 8589 13712 8590
rect 13529 8559 13538 8579
rect 13558 8559 13566 8579
rect 13529 8549 13566 8559
rect 13625 8579 13712 8589
rect 13625 8559 13634 8579
rect 13654 8559 13712 8579
rect 13625 8550 13712 8559
rect 13625 8549 13662 8550
rect 13347 8493 13363 8511
rect 13381 8493 13399 8511
rect 13681 8499 13712 8550
rect 13747 8579 13784 8646
rect 13899 8589 13935 8590
rect 13747 8559 13756 8579
rect 13776 8559 13784 8579
rect 13747 8549 13784 8559
rect 13843 8579 13991 8589
rect 14091 8586 14187 8588
rect 13843 8559 13852 8579
rect 13872 8559 13962 8579
rect 13982 8559 13991 8579
rect 13843 8550 13991 8559
rect 14049 8579 14187 8586
rect 14049 8559 14058 8579
rect 14078 8559 14187 8579
rect 14049 8550 14187 8559
rect 13843 8549 13880 8550
rect 13573 8496 13614 8497
rect 13347 8475 13399 8493
rect 13465 8489 13614 8496
rect 12915 8455 12955 8465
rect 13465 8469 13524 8489
rect 13544 8469 13583 8489
rect 13603 8469 13614 8489
rect 13465 8461 13614 8469
rect 13681 8492 13838 8499
rect 13681 8472 13801 8492
rect 13821 8472 13838 8492
rect 13681 8462 13838 8472
rect 13681 8461 13716 8462
rect 12745 8438 12783 8447
rect 13681 8440 13712 8461
rect 13899 8440 13935 8550
rect 13954 8549 13991 8550
rect 14050 8549 14087 8550
rect 14010 8490 14100 8496
rect 14010 8470 14019 8490
rect 14039 8488 14100 8490
rect 14039 8470 14064 8488
rect 14010 8468 14064 8470
rect 14084 8468 14100 8488
rect 14010 8462 14100 8468
rect 13524 8439 13561 8440
rect 12745 8437 12782 8438
rect 12206 8409 12296 8415
rect 12206 8389 12222 8409
rect 12242 8407 12296 8409
rect 12242 8389 12267 8407
rect 12206 8387 12267 8389
rect 12287 8387 12296 8407
rect 12206 8381 12296 8387
rect 12219 8327 12256 8328
rect 12315 8327 12352 8328
rect 12371 8327 12407 8437
rect 12594 8416 12625 8437
rect 13523 8430 13561 8439
rect 12590 8415 12625 8416
rect 12468 8405 12625 8415
rect 12468 8385 12485 8405
rect 12505 8385 12625 8405
rect 12468 8378 12625 8385
rect 12692 8408 12841 8416
rect 12692 8388 12703 8408
rect 12723 8388 12762 8408
rect 12782 8388 12841 8408
rect 13351 8412 13391 8422
rect 12692 8381 12841 8388
rect 12907 8384 12959 8402
rect 12692 8380 12733 8381
rect 12426 8327 12463 8328
rect 12119 8318 12257 8327
rect 11591 8307 11624 8309
rect 11220 8295 11667 8307
rect 10452 8173 10620 8175
rect 10176 8147 10620 8173
rect 9686 8125 9824 8134
rect 9480 8124 9517 8125
rect 8977 8070 9014 8073
rect 9210 8071 9251 8072
rect 7320 8049 7351 8050
rect 6944 7989 7285 7990
rect 7466 7989 7503 8060
rect 9102 8064 9251 8071
rect 8533 8052 8570 8057
rect 8524 8048 8571 8052
rect 8524 8030 8543 8048
rect 8561 8030 8571 8048
rect 9102 8044 9161 8064
rect 9181 8044 9220 8064
rect 9240 8044 9251 8064
rect 9102 8036 9251 8044
rect 9318 8067 9475 8074
rect 9318 8047 9438 8067
rect 9458 8047 9475 8067
rect 9318 8037 9475 8047
rect 9318 8036 9353 8037
rect 6869 7984 7285 7989
rect 6869 7964 6872 7984
rect 6892 7964 7285 7984
rect 7316 7965 7503 7989
rect 8128 7987 8168 7992
rect 8524 7987 8571 8030
rect 9318 8015 9349 8036
rect 9536 8015 9572 8125
rect 9591 8124 9628 8125
rect 9687 8124 9724 8125
rect 9647 8065 9737 8071
rect 9647 8045 9656 8065
rect 9676 8063 9737 8065
rect 9676 8045 9701 8063
rect 9647 8043 9701 8045
rect 9721 8043 9737 8063
rect 9647 8037 9737 8043
rect 9161 8014 9198 8015
rect 8128 7948 8571 7987
rect 8974 8006 9011 8008
rect 8974 7998 9016 8006
rect 8974 7980 8984 7998
rect 9002 7980 9016 7998
rect 8974 7971 9016 7980
rect 9160 8005 9198 8014
rect 9160 7985 9169 8005
rect 9189 7985 9198 8005
rect 9160 7977 9198 7985
rect 9264 8009 9349 8015
rect 9379 8014 9416 8015
rect 9264 7989 9272 8009
rect 9292 7989 9349 8009
rect 9264 7981 9349 7989
rect 9378 8005 9416 8014
rect 9378 7985 9387 8005
rect 9407 7985 9416 8005
rect 9264 7980 9300 7981
rect 9378 7977 9416 7985
rect 9482 8013 9626 8015
rect 9482 8009 9534 8013
rect 9482 7989 9490 8009
rect 9510 7993 9534 8009
rect 9554 8009 9626 8013
rect 9554 7993 9598 8009
rect 9510 7989 9598 7993
rect 9618 7989 9626 8009
rect 9482 7981 9626 7989
rect 9482 7980 9518 7981
rect 9590 7980 9626 7981
rect 9692 8014 9729 8015
rect 9692 8013 9730 8014
rect 9692 8005 9756 8013
rect 9692 7985 9701 8005
rect 9721 7991 9756 8005
rect 9776 7991 9779 8011
rect 9721 7986 9779 7991
rect 9721 7985 9756 7986
rect 5909 7889 5917 7911
rect 5941 7889 5949 7911
rect 5909 7881 5949 7889
rect 7222 7933 7262 7941
rect 7222 7911 7230 7933
rect 7254 7911 7262 7933
rect 3428 7835 3463 7836
rect 3405 7830 3463 7835
rect 3405 7810 3408 7830
rect 3428 7816 3463 7830
rect 3483 7816 3492 7836
rect 3428 7808 3492 7816
rect 3454 7807 3492 7808
rect 3455 7806 3492 7807
rect 3558 7840 3594 7841
rect 3666 7840 3702 7841
rect 3558 7832 3702 7840
rect 3558 7812 3566 7832
rect 3586 7828 3674 7832
rect 3586 7812 3630 7828
rect 3558 7808 3630 7812
rect 3650 7812 3674 7828
rect 3694 7812 3702 7832
rect 3650 7808 3702 7812
rect 3558 7806 3702 7808
rect 3768 7836 3806 7844
rect 3884 7840 3920 7841
rect 3768 7816 3777 7836
rect 3797 7816 3806 7836
rect 3768 7807 3806 7816
rect 3835 7832 3920 7840
rect 3835 7812 3892 7832
rect 3912 7812 3920 7832
rect 3768 7806 3805 7807
rect 3835 7806 3920 7812
rect 3986 7836 4024 7844
rect 3986 7816 3995 7836
rect 4015 7816 4024 7836
rect 3986 7807 4024 7816
rect 4168 7841 4210 7850
rect 4168 7823 4182 7841
rect 4200 7823 4210 7841
rect 4168 7815 4210 7823
rect 4173 7813 4210 7815
rect 4600 7835 5043 7874
rect 3986 7806 4023 7807
rect 3447 7778 3537 7784
rect 3447 7758 3463 7778
rect 3483 7776 3537 7778
rect 3483 7758 3508 7776
rect 3447 7756 3508 7758
rect 3528 7756 3537 7776
rect 3447 7750 3537 7756
rect 3460 7696 3497 7697
rect 3556 7696 3593 7697
rect 3612 7696 3648 7806
rect 3835 7785 3866 7806
rect 4600 7792 4647 7835
rect 5003 7830 5043 7835
rect 5668 7833 5855 7857
rect 5886 7838 6279 7858
rect 6299 7838 6302 7858
rect 5886 7833 6302 7838
rect 3831 7784 3866 7785
rect 3709 7774 3866 7784
rect 3709 7754 3726 7774
rect 3746 7754 3866 7774
rect 3709 7747 3866 7754
rect 3933 7777 4082 7785
rect 3933 7757 3944 7777
rect 3964 7757 4003 7777
rect 4023 7757 4082 7777
rect 4600 7774 4610 7792
rect 4628 7774 4647 7792
rect 4600 7770 4647 7774
rect 4601 7765 4638 7770
rect 3933 7750 4082 7757
rect 5668 7762 5705 7833
rect 5886 7832 6227 7833
rect 5820 7772 5851 7773
rect 3933 7749 3974 7750
rect 4170 7748 4207 7751
rect 3667 7696 3704 7697
rect 3360 7687 3498 7696
rect 2564 7648 3008 7674
rect 2564 7646 2732 7648
rect 1517 7514 1964 7526
rect 1560 7512 1593 7514
rect 927 7494 1065 7503
rect 721 7493 758 7494
rect 451 7440 492 7441
rect 225 7419 277 7437
rect 343 7433 492 7440
rect 343 7413 402 7433
rect 422 7413 461 7433
rect 481 7413 492 7433
rect 343 7405 492 7413
rect 559 7436 716 7443
rect 559 7416 679 7436
rect 699 7416 716 7436
rect 559 7406 716 7416
rect 559 7405 594 7406
rect 559 7384 590 7405
rect 777 7384 813 7494
rect 832 7493 869 7494
rect 928 7493 965 7494
rect 888 7434 978 7440
rect 888 7414 897 7434
rect 917 7432 978 7434
rect 917 7414 942 7432
rect 888 7412 942 7414
rect 962 7412 978 7432
rect 888 7406 978 7412
rect 402 7383 439 7384
rect 401 7374 439 7383
rect 229 7356 269 7366
rect 229 7338 239 7356
rect 257 7338 269 7356
rect 401 7354 410 7374
rect 430 7354 439 7374
rect 401 7346 439 7354
rect 505 7378 590 7384
rect 620 7383 657 7384
rect 505 7358 513 7378
rect 533 7358 590 7378
rect 505 7350 590 7358
rect 619 7374 657 7383
rect 619 7354 628 7374
rect 648 7354 657 7374
rect 505 7349 541 7350
rect 619 7346 657 7354
rect 723 7378 867 7384
rect 723 7358 731 7378
rect 751 7358 784 7378
rect 804 7358 839 7378
rect 859 7358 867 7378
rect 723 7350 867 7358
rect 723 7349 759 7350
rect 831 7349 867 7350
rect 933 7383 970 7384
rect 933 7382 971 7383
rect 933 7374 997 7382
rect 933 7354 942 7374
rect 962 7360 997 7374
rect 1017 7360 1020 7380
rect 962 7355 1020 7360
rect 962 7354 997 7355
rect 229 7282 269 7338
rect 402 7317 439 7346
rect 403 7315 439 7317
rect 403 7293 594 7315
rect 620 7314 657 7346
rect 933 7342 997 7354
rect 1037 7316 1064 7494
rect 1922 7469 1964 7514
rect 896 7314 1064 7316
rect 620 7304 1064 7314
rect 1205 7410 1392 7434
rect 1423 7415 1816 7435
rect 1836 7415 1839 7435
rect 1423 7410 1839 7415
rect 1205 7339 1242 7410
rect 1423 7409 1764 7410
rect 1357 7349 1388 7350
rect 1205 7319 1214 7339
rect 1234 7319 1242 7339
rect 1205 7309 1242 7319
rect 1301 7339 1388 7349
rect 1301 7319 1310 7339
rect 1330 7319 1388 7339
rect 1301 7310 1388 7319
rect 1301 7309 1338 7310
rect 226 7277 269 7282
rect 617 7288 1064 7304
rect 617 7282 645 7288
rect 896 7287 1064 7288
rect 226 7274 376 7277
rect 617 7274 644 7282
rect 226 7272 644 7274
rect 226 7254 235 7272
rect 253 7254 644 7272
rect 1357 7259 1388 7310
rect 1423 7339 1460 7409
rect 1726 7408 1763 7409
rect 1575 7349 1611 7350
rect 1423 7319 1432 7339
rect 1452 7319 1460 7339
rect 1423 7309 1460 7319
rect 1519 7339 1667 7349
rect 1767 7346 1863 7348
rect 1519 7319 1528 7339
rect 1548 7319 1638 7339
rect 1658 7319 1667 7339
rect 1519 7310 1667 7319
rect 1725 7339 1863 7346
rect 1725 7319 1734 7339
rect 1754 7319 1863 7339
rect 1725 7310 1863 7319
rect 1519 7309 1556 7310
rect 1249 7256 1290 7257
rect 226 7251 644 7254
rect 226 7245 269 7251
rect 229 7242 269 7245
rect 1144 7249 1290 7256
rect 626 7233 666 7234
rect 337 7216 666 7233
rect 1144 7229 1200 7249
rect 1220 7229 1259 7249
rect 1279 7229 1290 7249
rect 1144 7221 1290 7229
rect 1357 7252 1514 7259
rect 1357 7232 1477 7252
rect 1497 7232 1514 7252
rect 1357 7222 1514 7232
rect 1357 7221 1392 7222
rect 221 7173 264 7184
rect 221 7155 233 7173
rect 251 7155 264 7173
rect 221 7129 264 7155
rect 337 7129 364 7216
rect 626 7207 666 7216
rect 221 7108 364 7129
rect 408 7181 442 7197
rect 626 7187 1019 7207
rect 1039 7187 1042 7207
rect 1357 7200 1388 7221
rect 1575 7200 1611 7310
rect 1630 7309 1667 7310
rect 1726 7309 1763 7310
rect 1686 7250 1776 7256
rect 1686 7230 1695 7250
rect 1715 7248 1776 7250
rect 1715 7230 1740 7248
rect 1686 7228 1740 7230
rect 1760 7228 1776 7248
rect 1686 7222 1776 7228
rect 1200 7199 1237 7200
rect 626 7182 1042 7187
rect 1199 7190 1237 7199
rect 626 7181 967 7182
rect 408 7111 445 7181
rect 560 7121 591 7122
rect 221 7106 358 7108
rect 221 7064 264 7106
rect 408 7091 417 7111
rect 437 7091 445 7111
rect 408 7081 445 7091
rect 504 7111 591 7121
rect 504 7091 513 7111
rect 533 7091 591 7111
rect 504 7082 591 7091
rect 504 7081 541 7082
rect 219 7054 264 7064
rect 219 7036 228 7054
rect 246 7036 264 7054
rect 219 7030 264 7036
rect 560 7031 591 7082
rect 626 7111 663 7181
rect 929 7180 966 7181
rect 1199 7170 1208 7190
rect 1228 7170 1237 7190
rect 1199 7162 1237 7170
rect 1303 7194 1388 7200
rect 1418 7199 1455 7200
rect 1303 7174 1311 7194
rect 1331 7174 1388 7194
rect 1303 7166 1388 7174
rect 1417 7190 1455 7199
rect 1417 7170 1426 7190
rect 1446 7170 1455 7190
rect 1303 7165 1339 7166
rect 1417 7162 1455 7170
rect 1521 7194 1665 7200
rect 1521 7174 1529 7194
rect 1549 7191 1637 7194
rect 1549 7174 1584 7191
rect 1521 7173 1584 7174
rect 1603 7174 1637 7191
rect 1657 7174 1665 7194
rect 1603 7173 1665 7174
rect 1521 7166 1665 7173
rect 1521 7165 1557 7166
rect 1629 7165 1665 7166
rect 1731 7199 1768 7200
rect 1731 7198 1769 7199
rect 1791 7198 1818 7202
rect 1731 7196 1818 7198
rect 1731 7190 1795 7196
rect 1731 7170 1740 7190
rect 1760 7176 1795 7190
rect 1815 7176 1818 7196
rect 1760 7171 1818 7176
rect 1760 7170 1795 7171
rect 1200 7133 1237 7162
rect 1201 7131 1237 7133
rect 778 7121 814 7122
rect 626 7091 635 7111
rect 655 7091 663 7111
rect 626 7081 663 7091
rect 722 7111 870 7121
rect 970 7118 1066 7120
rect 722 7091 731 7111
rect 751 7091 841 7111
rect 861 7091 870 7111
rect 722 7082 870 7091
rect 928 7111 1066 7118
rect 928 7091 937 7111
rect 957 7091 1066 7111
rect 1201 7109 1392 7131
rect 1418 7130 1455 7162
rect 1731 7158 1795 7170
rect 1835 7132 1862 7310
rect 1694 7130 1862 7132
rect 1418 7104 1862 7130
rect 928 7082 1066 7091
rect 722 7081 759 7082
rect 219 7027 256 7030
rect 452 7028 493 7029
rect 344 7021 493 7028
rect 344 7001 403 7021
rect 423 7001 462 7021
rect 482 7001 493 7021
rect 344 6993 493 7001
rect 560 7024 717 7031
rect 560 7004 680 7024
rect 700 7004 717 7024
rect 560 6994 717 7004
rect 560 6993 595 6994
rect 560 6972 591 6993
rect 778 6972 814 7082
rect 833 7081 870 7082
rect 929 7081 966 7082
rect 889 7022 979 7028
rect 889 7002 898 7022
rect 918 7020 979 7022
rect 918 7002 943 7020
rect 889 7000 943 7002
rect 963 7000 979 7020
rect 889 6994 979 7000
rect 403 6971 440 6972
rect 215 6963 253 6965
rect 215 6955 258 6963
rect 215 6937 226 6955
rect 244 6937 258 6955
rect 215 6910 258 6937
rect 402 6962 440 6971
rect 402 6942 411 6962
rect 431 6942 440 6962
rect 402 6934 440 6942
rect 506 6966 591 6972
rect 621 6971 658 6972
rect 506 6946 514 6966
rect 534 6946 591 6966
rect 506 6938 591 6946
rect 620 6962 658 6971
rect 620 6942 629 6962
rect 649 6942 658 6962
rect 506 6937 542 6938
rect 620 6934 658 6942
rect 724 6970 868 6972
rect 724 6966 776 6970
rect 724 6946 732 6966
rect 752 6950 776 6966
rect 796 6966 868 6970
rect 796 6950 840 6966
rect 752 6946 840 6950
rect 860 6946 868 6966
rect 724 6938 868 6946
rect 724 6937 760 6938
rect 832 6937 868 6938
rect 934 6971 971 6972
rect 934 6970 972 6971
rect 934 6962 998 6970
rect 934 6942 943 6962
rect 963 6948 998 6962
rect 1018 6948 1021 6968
rect 963 6943 1021 6948
rect 963 6942 998 6943
rect 216 6903 258 6910
rect 403 6903 440 6934
rect 621 6903 658 6934
rect 934 6930 998 6942
rect 1038 6904 1065 7082
rect 216 6863 261 6903
rect 403 6878 548 6903
rect 621 6902 701 6903
rect 897 6902 1065 6904
rect 621 6886 1065 6902
rect 405 6877 548 6878
rect 620 6876 1065 6886
rect 216 6842 263 6863
rect 620 6842 661 6876
rect 897 6875 1065 6876
rect 1528 6880 1568 7104
rect 1694 7103 1862 7104
rect 1926 7136 1959 7469
rect 2564 7468 2591 7646
rect 2631 7608 2695 7620
rect 2971 7616 3008 7648
rect 3034 7647 3225 7669
rect 3360 7667 3469 7687
rect 3489 7667 3498 7687
rect 3360 7660 3498 7667
rect 3556 7687 3704 7696
rect 3556 7667 3565 7687
rect 3585 7667 3675 7687
rect 3695 7667 3704 7687
rect 3360 7658 3456 7660
rect 3556 7657 3704 7667
rect 3763 7687 3800 7697
rect 3763 7667 3771 7687
rect 3791 7667 3800 7687
rect 3612 7656 3648 7657
rect 3189 7645 3225 7647
rect 3189 7616 3226 7645
rect 2631 7607 2666 7608
rect 2608 7602 2666 7607
rect 2608 7582 2611 7602
rect 2631 7588 2666 7602
rect 2686 7588 2695 7608
rect 2631 7580 2695 7588
rect 2657 7579 2695 7580
rect 2658 7578 2695 7579
rect 2761 7612 2797 7613
rect 2869 7612 2905 7613
rect 2761 7604 2905 7612
rect 2761 7584 2769 7604
rect 2789 7603 2877 7604
rect 2789 7584 2824 7603
rect 2845 7584 2877 7603
rect 2897 7584 2905 7604
rect 2761 7578 2905 7584
rect 2971 7608 3009 7616
rect 3087 7612 3123 7613
rect 2971 7588 2980 7608
rect 3000 7588 3009 7608
rect 2971 7579 3009 7588
rect 3038 7604 3123 7612
rect 3038 7584 3095 7604
rect 3115 7584 3123 7604
rect 2971 7578 3008 7579
rect 3038 7578 3123 7584
rect 3189 7608 3227 7616
rect 3189 7588 3198 7608
rect 3218 7588 3227 7608
rect 3460 7597 3497 7598
rect 3763 7597 3800 7667
rect 3835 7696 3866 7747
rect 4162 7742 4207 7748
rect 4162 7724 4180 7742
rect 4198 7724 4207 7742
rect 5668 7742 5677 7762
rect 5697 7742 5705 7762
rect 5668 7732 5705 7742
rect 5764 7762 5851 7772
rect 5764 7742 5773 7762
rect 5793 7742 5851 7762
rect 5764 7733 5851 7742
rect 5764 7732 5801 7733
rect 4162 7714 4207 7724
rect 3885 7696 3922 7697
rect 3835 7687 3922 7696
rect 3835 7667 3893 7687
rect 3913 7667 3922 7687
rect 3835 7657 3922 7667
rect 3981 7687 4018 7697
rect 3981 7667 3989 7687
rect 4009 7667 4018 7687
rect 4162 7672 4205 7714
rect 4589 7703 4641 7705
rect 4068 7670 4205 7672
rect 3835 7656 3866 7657
rect 3981 7597 4018 7667
rect 3459 7596 3800 7597
rect 3189 7579 3227 7588
rect 3384 7591 3800 7596
rect 3189 7578 3226 7579
rect 2650 7550 2740 7556
rect 2650 7530 2666 7550
rect 2686 7548 2740 7550
rect 2686 7530 2711 7548
rect 2650 7528 2711 7530
rect 2731 7528 2740 7548
rect 2650 7522 2740 7528
rect 2663 7468 2700 7469
rect 2759 7468 2796 7469
rect 2815 7468 2851 7578
rect 3038 7557 3069 7578
rect 3384 7571 3387 7591
rect 3407 7571 3800 7591
rect 3984 7581 4018 7597
rect 4062 7649 4205 7670
rect 4587 7699 5020 7703
rect 4587 7693 5026 7699
rect 4587 7675 4608 7693
rect 4626 7675 5026 7693
rect 5820 7682 5851 7733
rect 5886 7762 5923 7832
rect 6189 7831 6226 7832
rect 6038 7772 6074 7773
rect 5886 7742 5895 7762
rect 5915 7742 5923 7762
rect 5886 7732 5923 7742
rect 5982 7762 6130 7772
rect 6230 7769 6326 7771
rect 5982 7742 5991 7762
rect 6011 7742 6101 7762
rect 6121 7742 6130 7762
rect 5982 7733 6130 7742
rect 6188 7762 6326 7769
rect 6188 7742 6197 7762
rect 6217 7742 6326 7762
rect 6188 7733 6326 7742
rect 5982 7732 6019 7733
rect 5712 7679 5753 7680
rect 4587 7657 5026 7675
rect 3760 7562 3800 7571
rect 4062 7562 4089 7649
rect 4162 7623 4205 7649
rect 4162 7605 4175 7623
rect 4193 7605 4205 7623
rect 4162 7594 4205 7605
rect 3034 7556 3069 7557
rect 2912 7546 3069 7556
rect 2912 7526 2929 7546
rect 2949 7526 3069 7546
rect 2912 7519 3069 7526
rect 3136 7549 3285 7557
rect 3136 7529 3147 7549
rect 3167 7529 3206 7549
rect 3226 7529 3285 7549
rect 3760 7545 4089 7562
rect 3760 7544 3800 7545
rect 3136 7522 3285 7529
rect 4157 7533 4197 7536
rect 4157 7527 4200 7533
rect 3782 7524 4200 7527
rect 3136 7521 3177 7522
rect 2870 7468 2907 7469
rect 2563 7459 2701 7468
rect 2426 7449 2462 7455
rect 2426 7431 2431 7449
rect 2453 7431 2462 7449
rect 2426 7427 2462 7431
rect 2563 7439 2672 7459
rect 2692 7439 2701 7459
rect 2563 7432 2701 7439
rect 2759 7459 2907 7468
rect 2759 7439 2768 7459
rect 2788 7439 2878 7459
rect 2898 7439 2907 7459
rect 2563 7430 2659 7432
rect 2759 7429 2907 7439
rect 2966 7459 3003 7469
rect 2966 7439 2974 7459
rect 2994 7439 3003 7459
rect 2815 7428 2851 7429
rect 2429 7268 2462 7427
rect 2663 7369 2700 7370
rect 2966 7369 3003 7439
rect 3038 7468 3069 7519
rect 3782 7506 4173 7524
rect 4191 7506 4200 7524
rect 3782 7504 4200 7506
rect 3782 7496 3809 7504
rect 4050 7501 4200 7504
rect 3362 7490 3530 7491
rect 3781 7490 3809 7496
rect 3362 7474 3809 7490
rect 4157 7496 4200 7501
rect 3088 7468 3125 7469
rect 3038 7459 3125 7468
rect 3038 7439 3096 7459
rect 3116 7439 3125 7459
rect 3038 7429 3125 7439
rect 3184 7459 3221 7469
rect 3184 7439 3192 7459
rect 3212 7439 3221 7459
rect 3038 7428 3069 7429
rect 2662 7368 3003 7369
rect 3184 7368 3221 7439
rect 2587 7363 3003 7368
rect 2587 7343 2590 7363
rect 2610 7343 3003 7363
rect 3034 7344 3221 7368
rect 3362 7464 3806 7474
rect 3362 7462 3530 7464
rect 3362 7284 3389 7462
rect 3429 7424 3493 7436
rect 3769 7432 3806 7464
rect 3832 7463 4023 7485
rect 3987 7461 4023 7463
rect 3987 7432 4024 7461
rect 4157 7440 4197 7496
rect 3429 7423 3464 7424
rect 3406 7418 3464 7423
rect 3406 7398 3409 7418
rect 3429 7404 3464 7418
rect 3484 7404 3493 7424
rect 3429 7396 3493 7404
rect 3455 7395 3493 7396
rect 3456 7394 3493 7395
rect 3559 7428 3595 7429
rect 3667 7428 3703 7429
rect 3559 7420 3703 7428
rect 3559 7400 3567 7420
rect 3587 7400 3622 7420
rect 3642 7400 3675 7420
rect 3695 7400 3703 7420
rect 3559 7394 3703 7400
rect 3769 7424 3807 7432
rect 3885 7428 3921 7429
rect 3769 7404 3778 7424
rect 3798 7404 3807 7424
rect 3769 7395 3807 7404
rect 3836 7420 3921 7428
rect 3836 7400 3893 7420
rect 3913 7400 3921 7420
rect 3769 7394 3806 7395
rect 3836 7394 3921 7400
rect 3987 7424 4025 7432
rect 3987 7404 3996 7424
rect 4016 7404 4025 7424
rect 4157 7422 4169 7440
rect 4187 7422 4197 7440
rect 4589 7468 4641 7657
rect 4987 7632 5026 7657
rect 5604 7672 5753 7679
rect 5604 7652 5663 7672
rect 5683 7652 5722 7672
rect 5742 7652 5753 7672
rect 5604 7644 5753 7652
rect 5820 7675 5977 7682
rect 5820 7655 5940 7675
rect 5960 7655 5977 7675
rect 5820 7645 5977 7655
rect 5820 7644 5855 7645
rect 4771 7607 4958 7631
rect 4987 7612 5382 7632
rect 5402 7612 5405 7632
rect 5820 7623 5851 7644
rect 6038 7623 6074 7733
rect 6093 7732 6130 7733
rect 6189 7732 6226 7733
rect 6149 7673 6239 7679
rect 6149 7653 6158 7673
rect 6178 7671 6239 7673
rect 6178 7653 6203 7671
rect 6149 7651 6203 7653
rect 6223 7651 6239 7671
rect 6149 7645 6239 7651
rect 5663 7622 5700 7623
rect 4987 7607 5405 7612
rect 5662 7613 5700 7622
rect 4771 7536 4808 7607
rect 4987 7606 5330 7607
rect 4987 7603 5026 7606
rect 5292 7605 5329 7606
rect 4923 7546 4954 7547
rect 4771 7516 4780 7536
rect 4800 7516 4808 7536
rect 4771 7506 4808 7516
rect 4867 7536 4954 7546
rect 4867 7516 4876 7536
rect 4896 7516 4954 7536
rect 4867 7507 4954 7516
rect 4867 7506 4904 7507
rect 4589 7450 4605 7468
rect 4623 7450 4641 7468
rect 4923 7456 4954 7507
rect 4989 7536 5026 7603
rect 5662 7593 5671 7613
rect 5691 7593 5700 7613
rect 5662 7585 5700 7593
rect 5766 7617 5851 7623
rect 5881 7622 5918 7623
rect 5766 7597 5774 7617
rect 5794 7597 5851 7617
rect 5766 7589 5851 7597
rect 5880 7613 5918 7622
rect 5880 7593 5889 7613
rect 5909 7593 5918 7613
rect 5766 7588 5802 7589
rect 5880 7585 5918 7593
rect 5984 7618 6128 7623
rect 5984 7617 6046 7618
rect 5984 7597 5992 7617
rect 6012 7599 6046 7617
rect 6067 7617 6128 7618
rect 6067 7599 6100 7617
rect 6012 7597 6100 7599
rect 6120 7597 6128 7617
rect 5984 7589 6128 7597
rect 5984 7588 6020 7589
rect 6092 7588 6128 7589
rect 6194 7622 6231 7623
rect 6194 7621 6232 7622
rect 6194 7613 6258 7621
rect 6194 7593 6203 7613
rect 6223 7599 6258 7613
rect 6278 7599 6281 7619
rect 6223 7594 6281 7599
rect 6223 7593 6258 7594
rect 5663 7556 5700 7585
rect 5664 7554 5700 7556
rect 5141 7546 5177 7547
rect 4989 7516 4998 7536
rect 5018 7516 5026 7536
rect 4989 7506 5026 7516
rect 5085 7536 5233 7546
rect 5333 7543 5429 7545
rect 5085 7516 5094 7536
rect 5114 7516 5204 7536
rect 5224 7516 5233 7536
rect 5085 7507 5233 7516
rect 5291 7536 5429 7543
rect 5291 7516 5300 7536
rect 5320 7516 5429 7536
rect 5664 7532 5855 7554
rect 5881 7553 5918 7585
rect 6194 7581 6258 7593
rect 6298 7555 6325 7733
rect 6157 7553 6325 7555
rect 5881 7539 6325 7553
rect 6928 7687 7096 7688
rect 7222 7687 7262 7911
rect 7725 7915 7893 7916
rect 8128 7915 8168 7948
rect 8524 7915 8571 7948
rect 8975 7946 9016 7971
rect 9161 7946 9198 7977
rect 9379 7946 9416 7977
rect 9692 7973 9756 7985
rect 9796 7947 9823 8125
rect 8975 7919 9024 7946
rect 9160 7920 9209 7946
rect 9378 7945 9459 7946
rect 9655 7945 9823 7947
rect 9378 7920 9823 7945
rect 9379 7919 9823 7920
rect 7725 7914 8169 7915
rect 7725 7889 8170 7914
rect 7725 7887 7893 7889
rect 8089 7888 8170 7889
rect 8339 7888 8388 7914
rect 8524 7888 8573 7915
rect 7725 7709 7752 7887
rect 7792 7849 7856 7861
rect 8132 7857 8169 7888
rect 8350 7857 8387 7888
rect 8532 7863 8573 7888
rect 8977 7886 9024 7919
rect 9380 7886 9420 7919
rect 9655 7918 9823 7919
rect 10286 7923 10326 8147
rect 10452 8146 10620 8147
rect 11223 8281 11667 8295
rect 11223 8279 11391 8281
rect 11223 8101 11250 8279
rect 11290 8241 11354 8253
rect 11630 8249 11667 8281
rect 11693 8280 11884 8302
rect 12119 8298 12228 8318
rect 12248 8298 12257 8318
rect 12119 8291 12257 8298
rect 12315 8318 12463 8327
rect 12315 8298 12324 8318
rect 12344 8298 12434 8318
rect 12454 8298 12463 8318
rect 12119 8289 12215 8291
rect 12315 8288 12463 8298
rect 12522 8318 12559 8328
rect 12522 8298 12530 8318
rect 12550 8298 12559 8318
rect 12371 8287 12407 8288
rect 11848 8278 11884 8280
rect 11848 8249 11885 8278
rect 11290 8240 11325 8241
rect 11267 8235 11325 8240
rect 11267 8215 11270 8235
rect 11290 8221 11325 8235
rect 11345 8221 11354 8241
rect 11290 8213 11354 8221
rect 11316 8212 11354 8213
rect 11317 8211 11354 8212
rect 11420 8245 11456 8246
rect 11528 8245 11564 8246
rect 11420 8239 11564 8245
rect 11420 8237 11481 8239
rect 11420 8217 11428 8237
rect 11448 8222 11481 8237
rect 11500 8237 11564 8239
rect 11500 8222 11536 8237
rect 11448 8217 11536 8222
rect 11556 8217 11564 8237
rect 11420 8211 11564 8217
rect 11630 8241 11668 8249
rect 11746 8245 11782 8246
rect 11630 8221 11639 8241
rect 11659 8221 11668 8241
rect 11630 8212 11668 8221
rect 11697 8237 11782 8245
rect 11697 8217 11754 8237
rect 11774 8217 11782 8237
rect 11630 8211 11667 8212
rect 11697 8211 11782 8217
rect 11848 8241 11886 8249
rect 11848 8221 11857 8241
rect 11877 8221 11886 8241
rect 12522 8231 12559 8298
rect 12594 8327 12625 8378
rect 12907 8366 12925 8384
rect 12943 8366 12959 8384
rect 12644 8327 12681 8328
rect 12594 8318 12681 8327
rect 12594 8298 12652 8318
rect 12672 8298 12681 8318
rect 12594 8288 12681 8298
rect 12740 8318 12777 8328
rect 12740 8298 12748 8318
rect 12768 8298 12777 8318
rect 12594 8287 12625 8288
rect 12219 8228 12256 8229
rect 12522 8228 12561 8231
rect 12218 8227 12561 8228
rect 12740 8227 12777 8298
rect 11848 8212 11886 8221
rect 12143 8222 12561 8227
rect 11848 8211 11885 8212
rect 11309 8183 11399 8189
rect 11309 8163 11325 8183
rect 11345 8181 11399 8183
rect 11345 8163 11370 8181
rect 11309 8161 11370 8163
rect 11390 8161 11399 8181
rect 11309 8155 11399 8161
rect 11322 8101 11359 8102
rect 11418 8101 11455 8102
rect 11474 8101 11510 8211
rect 11697 8190 11728 8211
rect 12143 8202 12146 8222
rect 12166 8202 12561 8222
rect 12590 8203 12777 8227
rect 11693 8189 11728 8190
rect 11571 8179 11728 8189
rect 11571 8159 11588 8179
rect 11608 8159 11728 8179
rect 11571 8152 11728 8159
rect 11795 8182 11944 8190
rect 11795 8162 11806 8182
rect 11826 8162 11865 8182
rect 11885 8162 11944 8182
rect 11795 8155 11944 8162
rect 12522 8177 12561 8202
rect 12907 8177 12959 8366
rect 13351 8394 13361 8412
rect 13379 8394 13391 8412
rect 13523 8410 13532 8430
rect 13552 8410 13561 8430
rect 13523 8402 13561 8410
rect 13627 8434 13712 8440
rect 13742 8439 13779 8440
rect 13627 8414 13635 8434
rect 13655 8414 13712 8434
rect 13627 8406 13712 8414
rect 13741 8430 13779 8439
rect 13741 8410 13750 8430
rect 13770 8410 13779 8430
rect 13627 8405 13663 8406
rect 13741 8402 13779 8410
rect 13845 8434 13989 8440
rect 13845 8414 13853 8434
rect 13873 8414 13906 8434
rect 13926 8414 13961 8434
rect 13981 8414 13989 8434
rect 13845 8406 13989 8414
rect 13845 8405 13881 8406
rect 13953 8405 13989 8406
rect 14055 8439 14092 8440
rect 14055 8438 14093 8439
rect 14055 8430 14119 8438
rect 14055 8410 14064 8430
rect 14084 8416 14119 8430
rect 14139 8416 14142 8436
rect 14084 8411 14142 8416
rect 14084 8410 14119 8411
rect 13351 8338 13391 8394
rect 13524 8373 13561 8402
rect 13525 8371 13561 8373
rect 13525 8349 13716 8371
rect 13742 8370 13779 8402
rect 14055 8398 14119 8410
rect 14159 8372 14186 8550
rect 14018 8370 14186 8372
rect 13742 8360 14186 8370
rect 14327 8466 14514 8490
rect 14545 8471 14938 8491
rect 14958 8471 14961 8491
rect 14545 8466 14961 8471
rect 14327 8395 14364 8466
rect 14545 8465 14886 8466
rect 14479 8405 14510 8406
rect 14327 8375 14336 8395
rect 14356 8375 14364 8395
rect 14327 8365 14364 8375
rect 14423 8395 14510 8405
rect 14423 8375 14432 8395
rect 14452 8375 14510 8395
rect 14423 8366 14510 8375
rect 14423 8365 14460 8366
rect 13348 8333 13391 8338
rect 13739 8344 14186 8360
rect 13739 8338 13767 8344
rect 14018 8343 14186 8344
rect 13348 8330 13498 8333
rect 13739 8330 13766 8338
rect 13348 8328 13766 8330
rect 13348 8310 13357 8328
rect 13375 8310 13766 8328
rect 14479 8315 14510 8366
rect 14545 8395 14582 8465
rect 14848 8464 14885 8465
rect 14697 8405 14733 8406
rect 14545 8375 14554 8395
rect 14574 8375 14582 8395
rect 14545 8365 14582 8375
rect 14641 8395 14789 8405
rect 14889 8402 14985 8404
rect 14641 8375 14650 8395
rect 14670 8375 14760 8395
rect 14780 8375 14789 8395
rect 14641 8366 14789 8375
rect 14847 8395 14985 8402
rect 14847 8375 14856 8395
rect 14876 8375 14985 8395
rect 14847 8366 14985 8375
rect 14641 8365 14678 8366
rect 14371 8312 14412 8313
rect 13348 8307 13766 8310
rect 13348 8301 13391 8307
rect 13351 8298 13391 8301
rect 14263 8305 14412 8312
rect 13748 8289 13788 8290
rect 13459 8272 13788 8289
rect 14263 8285 14322 8305
rect 14342 8285 14381 8305
rect 14401 8285 14412 8305
rect 14263 8277 14412 8285
rect 14479 8308 14636 8315
rect 14479 8288 14599 8308
rect 14619 8288 14636 8308
rect 14479 8278 14636 8288
rect 14479 8277 14514 8278
rect 13343 8229 13386 8240
rect 13343 8211 13355 8229
rect 13373 8211 13386 8229
rect 13343 8185 13386 8211
rect 13459 8185 13486 8272
rect 13748 8263 13788 8272
rect 12522 8159 12961 8177
rect 11795 8154 11836 8155
rect 11529 8101 11566 8102
rect 11222 8092 11360 8101
rect 11222 8072 11331 8092
rect 11351 8072 11360 8092
rect 11222 8065 11360 8072
rect 11418 8092 11566 8101
rect 11418 8072 11427 8092
rect 11447 8072 11537 8092
rect 11557 8072 11566 8092
rect 11222 8063 11318 8065
rect 11418 8062 11566 8072
rect 11625 8092 11662 8102
rect 11625 8072 11633 8092
rect 11653 8072 11662 8092
rect 11474 8061 11510 8062
rect 11322 8002 11359 8003
rect 11625 8002 11662 8072
rect 11697 8101 11728 8152
rect 12522 8141 12922 8159
rect 12940 8141 12961 8159
rect 12522 8135 12961 8141
rect 12528 8131 12961 8135
rect 13343 8164 13486 8185
rect 13530 8237 13564 8253
rect 13748 8243 14141 8263
rect 14161 8243 14164 8263
rect 14479 8256 14510 8277
rect 14697 8256 14733 8366
rect 14752 8365 14789 8366
rect 14848 8365 14885 8366
rect 14808 8306 14898 8312
rect 14808 8286 14817 8306
rect 14837 8304 14898 8306
rect 14837 8286 14862 8304
rect 14808 8284 14862 8286
rect 14882 8284 14898 8304
rect 14808 8278 14898 8284
rect 14322 8255 14359 8256
rect 13748 8238 14164 8243
rect 14321 8246 14359 8255
rect 13748 8237 14089 8238
rect 13530 8167 13567 8237
rect 13682 8177 13713 8178
rect 13343 8162 13480 8164
rect 12907 8129 12959 8131
rect 13343 8120 13386 8162
rect 13530 8147 13539 8167
rect 13559 8147 13567 8167
rect 13530 8137 13567 8147
rect 13626 8167 13713 8177
rect 13626 8147 13635 8167
rect 13655 8147 13713 8167
rect 13626 8138 13713 8147
rect 13626 8137 13663 8138
rect 13341 8110 13386 8120
rect 11747 8101 11784 8102
rect 11697 8092 11784 8101
rect 11697 8072 11755 8092
rect 11775 8072 11784 8092
rect 11697 8062 11784 8072
rect 11843 8092 11880 8102
rect 11843 8072 11851 8092
rect 11871 8072 11880 8092
rect 13341 8092 13350 8110
rect 13368 8092 13386 8110
rect 13341 8086 13386 8092
rect 13682 8087 13713 8138
rect 13748 8167 13785 8237
rect 14051 8236 14088 8237
rect 14321 8226 14330 8246
rect 14350 8226 14359 8246
rect 14321 8218 14359 8226
rect 14425 8250 14510 8256
rect 14540 8255 14577 8256
rect 14425 8230 14433 8250
rect 14453 8230 14510 8250
rect 14425 8222 14510 8230
rect 14539 8246 14577 8255
rect 14539 8226 14548 8246
rect 14568 8226 14577 8246
rect 14425 8221 14461 8222
rect 14539 8218 14577 8226
rect 14643 8250 14787 8256
rect 14643 8230 14651 8250
rect 14671 8231 14703 8250
rect 14724 8231 14759 8250
rect 14671 8230 14759 8231
rect 14779 8230 14787 8250
rect 14643 8222 14787 8230
rect 14643 8221 14679 8222
rect 14751 8221 14787 8222
rect 14853 8255 14890 8256
rect 14853 8254 14891 8255
rect 14853 8246 14917 8254
rect 14853 8226 14862 8246
rect 14882 8232 14917 8246
rect 14937 8232 14940 8252
rect 14882 8227 14940 8232
rect 14882 8226 14917 8227
rect 14322 8189 14359 8218
rect 14323 8187 14359 8189
rect 13900 8177 13936 8178
rect 13748 8147 13757 8167
rect 13777 8147 13785 8167
rect 13748 8137 13785 8147
rect 13844 8167 13992 8177
rect 14092 8174 14188 8176
rect 13844 8147 13853 8167
rect 13873 8147 13963 8167
rect 13983 8147 13992 8167
rect 13844 8138 13992 8147
rect 14050 8167 14188 8174
rect 14050 8147 14059 8167
rect 14079 8147 14188 8167
rect 14323 8165 14514 8187
rect 14540 8186 14577 8218
rect 14853 8214 14917 8226
rect 14957 8188 14984 8366
rect 15589 8365 15622 8698
rect 15686 8730 15854 8731
rect 15980 8730 16020 8954
rect 16483 8958 16651 8959
rect 16890 8958 16929 9004
rect 16483 8932 16929 8958
rect 16483 8930 16651 8932
rect 16847 8931 16929 8932
rect 17068 8931 17147 8957
rect 17289 8938 17332 9004
rect 16483 8752 16510 8930
rect 16550 8892 16614 8904
rect 16890 8900 16927 8931
rect 17108 8900 17145 8931
rect 17289 8921 17331 8938
rect 17626 8925 17669 9004
rect 20246 8950 20286 8958
rect 20246 8928 20254 8950
rect 20278 8928 20286 8950
rect 21150 8953 21606 8988
rect 25517 8981 26412 9041
rect 25517 8980 25964 8981
rect 24610 8963 24650 8971
rect 17290 8906 17331 8921
rect 16550 8891 16585 8892
rect 16527 8886 16585 8891
rect 16527 8866 16530 8886
rect 16550 8872 16585 8886
rect 16605 8872 16614 8892
rect 16550 8864 16614 8872
rect 16576 8863 16614 8864
rect 16577 8862 16614 8863
rect 16680 8896 16716 8897
rect 16788 8896 16824 8897
rect 16680 8888 16824 8896
rect 16680 8868 16688 8888
rect 16708 8884 16796 8888
rect 16708 8868 16752 8884
rect 16680 8864 16752 8868
rect 16772 8868 16796 8884
rect 16816 8868 16824 8888
rect 16772 8864 16824 8868
rect 16680 8862 16824 8864
rect 16890 8892 16928 8900
rect 17006 8896 17042 8897
rect 16890 8872 16899 8892
rect 16919 8872 16928 8892
rect 16890 8863 16928 8872
rect 16957 8888 17042 8896
rect 16957 8868 17014 8888
rect 17034 8868 17042 8888
rect 16890 8862 16927 8863
rect 16957 8862 17042 8868
rect 17108 8892 17146 8900
rect 17108 8872 17117 8892
rect 17137 8872 17146 8892
rect 17108 8863 17146 8872
rect 17290 8897 17332 8906
rect 17290 8879 17304 8897
rect 17322 8879 17332 8897
rect 17290 8871 17332 8879
rect 17295 8869 17332 8871
rect 17108 8862 17145 8863
rect 16569 8834 16659 8840
rect 16569 8814 16585 8834
rect 16605 8832 16659 8834
rect 16605 8814 16630 8832
rect 16569 8812 16630 8814
rect 16650 8812 16659 8832
rect 16569 8806 16659 8812
rect 16582 8752 16619 8753
rect 16678 8752 16715 8753
rect 16734 8752 16770 8862
rect 16957 8841 16988 8862
rect 16953 8840 16988 8841
rect 16831 8830 16988 8840
rect 16831 8810 16848 8830
rect 16868 8810 16988 8830
rect 16831 8803 16988 8810
rect 17055 8833 17204 8841
rect 17055 8813 17066 8833
rect 17086 8813 17125 8833
rect 17145 8813 17204 8833
rect 17055 8806 17204 8813
rect 17624 8809 17671 8925
rect 17055 8805 17096 8806
rect 17292 8804 17329 8807
rect 16789 8752 16826 8753
rect 16482 8743 16620 8752
rect 15686 8704 16130 8730
rect 15686 8702 15854 8704
rect 15686 8524 15713 8702
rect 15753 8664 15817 8676
rect 16093 8672 16130 8704
rect 16156 8703 16347 8725
rect 16482 8723 16591 8743
rect 16611 8723 16620 8743
rect 16482 8716 16620 8723
rect 16678 8743 16826 8752
rect 16678 8723 16687 8743
rect 16707 8723 16797 8743
rect 16817 8723 16826 8743
rect 16482 8714 16578 8716
rect 16678 8713 16826 8723
rect 16885 8743 16922 8753
rect 16885 8723 16893 8743
rect 16913 8723 16922 8743
rect 16734 8712 16770 8713
rect 16311 8701 16347 8703
rect 16311 8672 16348 8701
rect 15753 8663 15788 8664
rect 15730 8658 15788 8663
rect 15730 8638 15733 8658
rect 15753 8644 15788 8658
rect 15808 8644 15817 8664
rect 15753 8638 15817 8644
rect 15730 8636 15817 8638
rect 15730 8632 15757 8636
rect 15779 8635 15817 8636
rect 15780 8634 15817 8635
rect 15883 8668 15919 8669
rect 15991 8668 16027 8669
rect 15883 8661 16027 8668
rect 15883 8660 15945 8661
rect 15883 8640 15891 8660
rect 15911 8643 15945 8660
rect 15964 8660 16027 8661
rect 15964 8643 15999 8660
rect 15911 8640 15999 8643
rect 16019 8640 16027 8660
rect 15883 8634 16027 8640
rect 16093 8664 16131 8672
rect 16209 8668 16245 8669
rect 16093 8644 16102 8664
rect 16122 8644 16131 8664
rect 16093 8635 16131 8644
rect 16160 8660 16245 8668
rect 16160 8640 16217 8660
rect 16237 8640 16245 8660
rect 16093 8634 16130 8635
rect 16160 8634 16245 8640
rect 16311 8664 16349 8672
rect 16311 8644 16320 8664
rect 16340 8644 16349 8664
rect 16582 8653 16619 8654
rect 16885 8653 16922 8723
rect 16957 8752 16988 8803
rect 17284 8798 17329 8804
rect 17284 8780 17302 8798
rect 17320 8780 17329 8798
rect 17624 8791 17634 8809
rect 17652 8791 17671 8809
rect 17624 8787 17671 8791
rect 17625 8782 17662 8787
rect 17284 8770 17329 8780
rect 17007 8752 17044 8753
rect 16957 8743 17044 8752
rect 16957 8723 17015 8743
rect 17035 8723 17044 8743
rect 16957 8713 17044 8723
rect 17103 8743 17140 8753
rect 17103 8723 17111 8743
rect 17131 8723 17140 8743
rect 17284 8728 17327 8770
rect 17190 8726 17327 8728
rect 16957 8712 16988 8713
rect 17103 8653 17140 8723
rect 16581 8652 16922 8653
rect 16311 8635 16349 8644
rect 16506 8647 16922 8652
rect 16311 8634 16348 8635
rect 15772 8606 15862 8612
rect 15772 8586 15788 8606
rect 15808 8604 15862 8606
rect 15808 8586 15833 8604
rect 15772 8584 15833 8586
rect 15853 8584 15862 8604
rect 15772 8578 15862 8584
rect 15785 8524 15822 8525
rect 15881 8524 15918 8525
rect 15937 8524 15973 8634
rect 16160 8613 16191 8634
rect 16506 8627 16509 8647
rect 16529 8627 16922 8647
rect 17106 8637 17140 8653
rect 17184 8705 17327 8726
rect 17613 8720 17665 8722
rect 16882 8618 16922 8627
rect 17184 8618 17211 8705
rect 17284 8679 17327 8705
rect 17284 8661 17297 8679
rect 17315 8661 17327 8679
rect 17611 8716 18044 8720
rect 17611 8710 18050 8716
rect 17611 8692 17632 8710
rect 17650 8692 18050 8710
rect 17611 8674 18050 8692
rect 17284 8650 17327 8661
rect 16156 8612 16191 8613
rect 16034 8602 16191 8612
rect 16034 8582 16051 8602
rect 16071 8582 16191 8602
rect 16034 8575 16191 8582
rect 16258 8605 16404 8613
rect 16258 8585 16269 8605
rect 16289 8585 16328 8605
rect 16348 8585 16404 8605
rect 16882 8601 17211 8618
rect 16882 8600 16922 8601
rect 16258 8578 16404 8585
rect 17279 8589 17319 8592
rect 17279 8583 17322 8589
rect 16904 8580 17322 8583
rect 16258 8577 16299 8578
rect 15992 8524 16029 8525
rect 15685 8515 15823 8524
rect 15685 8495 15794 8515
rect 15814 8495 15823 8515
rect 15685 8488 15823 8495
rect 15881 8515 16029 8524
rect 15881 8495 15890 8515
rect 15910 8495 16000 8515
rect 16020 8495 16029 8515
rect 15685 8486 15781 8488
rect 15881 8485 16029 8495
rect 16088 8515 16125 8525
rect 16088 8495 16096 8515
rect 16116 8495 16125 8515
rect 15937 8484 15973 8485
rect 15785 8425 15822 8426
rect 16088 8425 16125 8495
rect 16160 8524 16191 8575
rect 16904 8562 17295 8580
rect 17313 8562 17322 8580
rect 16904 8560 17322 8562
rect 16904 8552 16931 8560
rect 17172 8557 17322 8560
rect 16484 8546 16652 8547
rect 16903 8546 16931 8552
rect 16484 8530 16931 8546
rect 17279 8552 17322 8557
rect 16210 8524 16247 8525
rect 16160 8515 16247 8524
rect 16160 8495 16218 8515
rect 16238 8495 16247 8515
rect 16160 8485 16247 8495
rect 16306 8515 16343 8525
rect 16306 8495 16314 8515
rect 16334 8495 16343 8515
rect 16160 8484 16191 8485
rect 15784 8424 16125 8425
rect 16306 8424 16343 8495
rect 15709 8419 16125 8424
rect 15709 8399 15712 8419
rect 15732 8399 16125 8419
rect 16156 8400 16343 8424
rect 16484 8520 16928 8530
rect 16484 8518 16652 8520
rect 15584 8320 15626 8365
rect 16484 8340 16511 8518
rect 16551 8480 16615 8492
rect 16891 8488 16928 8520
rect 16954 8519 17145 8541
rect 17109 8517 17145 8519
rect 17109 8488 17146 8517
rect 17279 8496 17319 8552
rect 16551 8479 16586 8480
rect 16528 8474 16586 8479
rect 16528 8454 16531 8474
rect 16551 8460 16586 8474
rect 16606 8460 16615 8480
rect 16551 8452 16615 8460
rect 16577 8451 16615 8452
rect 16578 8450 16615 8451
rect 16681 8484 16717 8485
rect 16789 8484 16825 8485
rect 16681 8476 16825 8484
rect 16681 8456 16689 8476
rect 16709 8456 16744 8476
rect 16764 8456 16797 8476
rect 16817 8456 16825 8476
rect 16681 8450 16825 8456
rect 16891 8480 16929 8488
rect 17007 8484 17043 8485
rect 16891 8460 16900 8480
rect 16920 8460 16929 8480
rect 16891 8451 16929 8460
rect 16958 8476 17043 8484
rect 16958 8456 17015 8476
rect 17035 8456 17043 8476
rect 16891 8450 16928 8451
rect 16958 8450 17043 8456
rect 17109 8480 17147 8488
rect 17109 8460 17118 8480
rect 17138 8460 17147 8480
rect 17279 8478 17291 8496
rect 17309 8478 17319 8496
rect 17279 8468 17319 8478
rect 17613 8485 17665 8674
rect 18011 8649 18050 8674
rect 19851 8699 19888 8705
rect 19851 8680 19859 8699
rect 19880 8680 19888 8699
rect 19851 8672 19888 8680
rect 17795 8624 17982 8648
rect 18011 8629 18406 8649
rect 18426 8629 18429 8649
rect 18011 8624 18429 8629
rect 17795 8553 17832 8624
rect 18011 8623 18354 8624
rect 18011 8620 18050 8623
rect 18316 8622 18353 8623
rect 17947 8563 17978 8564
rect 17795 8533 17804 8553
rect 17824 8533 17832 8553
rect 17795 8523 17832 8533
rect 17891 8553 17978 8563
rect 17891 8533 17900 8553
rect 17920 8533 17978 8553
rect 17891 8524 17978 8533
rect 17891 8523 17928 8524
rect 17109 8451 17147 8460
rect 17613 8467 17629 8485
rect 17647 8467 17665 8485
rect 17947 8473 17978 8524
rect 18013 8553 18050 8620
rect 18165 8563 18201 8564
rect 18013 8533 18022 8553
rect 18042 8533 18050 8553
rect 18013 8523 18050 8533
rect 18109 8553 18257 8563
rect 18357 8560 18453 8562
rect 18109 8533 18118 8553
rect 18138 8533 18228 8553
rect 18248 8533 18257 8553
rect 18109 8524 18257 8533
rect 18315 8553 18453 8560
rect 18315 8533 18324 8553
rect 18344 8533 18453 8553
rect 18315 8524 18453 8533
rect 18109 8523 18146 8524
rect 17839 8470 17880 8471
rect 17109 8450 17146 8451
rect 16570 8422 16660 8428
rect 16570 8402 16586 8422
rect 16606 8420 16660 8422
rect 16606 8402 16631 8420
rect 16570 8400 16631 8402
rect 16651 8400 16660 8420
rect 16570 8394 16660 8400
rect 16583 8340 16620 8341
rect 16679 8340 16716 8341
rect 16735 8340 16771 8450
rect 16958 8429 16989 8450
rect 17613 8449 17665 8467
rect 17731 8463 17880 8470
rect 17731 8443 17790 8463
rect 17810 8443 17849 8463
rect 17869 8443 17880 8463
rect 17731 8435 17880 8443
rect 17947 8466 18104 8473
rect 17947 8446 18067 8466
rect 18087 8446 18104 8466
rect 17947 8436 18104 8446
rect 17947 8435 17982 8436
rect 16954 8428 16989 8429
rect 16832 8418 16989 8428
rect 16832 8398 16849 8418
rect 16869 8398 16989 8418
rect 16832 8391 16989 8398
rect 17056 8421 17205 8429
rect 17056 8401 17067 8421
rect 17087 8401 17126 8421
rect 17146 8401 17205 8421
rect 17056 8394 17205 8401
rect 17271 8397 17323 8415
rect 17947 8414 17978 8435
rect 18165 8414 18201 8524
rect 18220 8523 18257 8524
rect 18316 8523 18353 8524
rect 18276 8464 18366 8470
rect 18276 8444 18285 8464
rect 18305 8462 18366 8464
rect 18305 8444 18330 8462
rect 18276 8442 18330 8444
rect 18350 8442 18366 8462
rect 18276 8436 18366 8442
rect 17790 8413 17827 8414
rect 17056 8393 17097 8394
rect 16790 8340 16827 8341
rect 16483 8331 16621 8340
rect 15955 8320 15988 8322
rect 15584 8308 16031 8320
rect 14816 8186 14984 8188
rect 14540 8160 14984 8186
rect 14050 8138 14188 8147
rect 13844 8137 13881 8138
rect 13341 8083 13378 8086
rect 13574 8084 13615 8085
rect 11697 8061 11728 8062
rect 11321 8001 11662 8002
rect 11843 8001 11880 8072
rect 13466 8077 13615 8084
rect 12910 8064 12947 8069
rect 12901 8060 12948 8064
rect 12901 8042 12920 8060
rect 12938 8042 12948 8060
rect 13466 8057 13525 8077
rect 13545 8057 13584 8077
rect 13604 8057 13615 8077
rect 13466 8049 13615 8057
rect 13682 8080 13839 8087
rect 13682 8060 13802 8080
rect 13822 8060 13839 8080
rect 13682 8050 13839 8060
rect 13682 8049 13717 8050
rect 11246 7996 11662 8001
rect 11246 7976 11249 7996
rect 11269 7976 11662 7996
rect 11693 7977 11880 8001
rect 12505 7999 12545 8004
rect 12901 7999 12948 8042
rect 13682 8028 13713 8049
rect 13900 8028 13936 8138
rect 13955 8137 13992 8138
rect 14051 8137 14088 8138
rect 14011 8078 14101 8084
rect 14011 8058 14020 8078
rect 14040 8076 14101 8078
rect 14040 8058 14065 8076
rect 14011 8056 14065 8058
rect 14085 8056 14101 8076
rect 14011 8050 14101 8056
rect 13525 8027 13562 8028
rect 12505 7960 12948 7999
rect 13338 8019 13375 8021
rect 13338 8011 13380 8019
rect 13338 7993 13348 8011
rect 13366 7993 13380 8011
rect 13338 7984 13380 7993
rect 13524 8018 13562 8027
rect 13524 7998 13533 8018
rect 13553 7998 13562 8018
rect 13524 7990 13562 7998
rect 13628 8022 13713 8028
rect 13743 8027 13780 8028
rect 13628 8002 13636 8022
rect 13656 8002 13713 8022
rect 13628 7994 13713 8002
rect 13742 8018 13780 8027
rect 13742 7998 13751 8018
rect 13771 7998 13780 8018
rect 13628 7993 13664 7994
rect 13742 7990 13780 7998
rect 13846 8026 13990 8028
rect 13846 8022 13898 8026
rect 13846 8002 13854 8022
rect 13874 8006 13898 8022
rect 13918 8022 13990 8026
rect 13918 8006 13962 8022
rect 13874 8002 13962 8006
rect 13982 8002 13990 8022
rect 13846 7994 13990 8002
rect 13846 7993 13882 7994
rect 13954 7993 13990 7994
rect 14056 8027 14093 8028
rect 14056 8026 14094 8027
rect 14056 8018 14120 8026
rect 14056 7998 14065 8018
rect 14085 8004 14120 8018
rect 14140 8004 14143 8024
rect 14085 7999 14143 8004
rect 14085 7998 14120 7999
rect 10286 7901 10294 7923
rect 10318 7901 10326 7923
rect 10286 7893 10326 7901
rect 11599 7945 11639 7953
rect 11599 7923 11607 7945
rect 11631 7923 11639 7945
rect 7792 7848 7827 7849
rect 7769 7843 7827 7848
rect 7769 7823 7772 7843
rect 7792 7829 7827 7843
rect 7847 7829 7856 7849
rect 7792 7821 7856 7829
rect 7818 7820 7856 7821
rect 7819 7819 7856 7820
rect 7922 7853 7958 7854
rect 8030 7853 8066 7854
rect 7922 7845 8066 7853
rect 7922 7825 7930 7845
rect 7950 7841 8038 7845
rect 7950 7825 7994 7841
rect 7922 7821 7994 7825
rect 8014 7825 8038 7841
rect 8058 7825 8066 7845
rect 8014 7821 8066 7825
rect 7922 7819 8066 7821
rect 8132 7849 8170 7857
rect 8248 7853 8284 7854
rect 8132 7829 8141 7849
rect 8161 7829 8170 7849
rect 8132 7820 8170 7829
rect 8199 7845 8284 7853
rect 8199 7825 8256 7845
rect 8276 7825 8284 7845
rect 8132 7819 8169 7820
rect 8199 7819 8284 7825
rect 8350 7849 8388 7857
rect 8350 7829 8359 7849
rect 8379 7829 8388 7849
rect 8350 7820 8388 7829
rect 8532 7854 8574 7863
rect 8532 7836 8546 7854
rect 8564 7836 8574 7854
rect 8532 7828 8574 7836
rect 8537 7826 8574 7828
rect 8977 7847 9420 7886
rect 8350 7819 8387 7820
rect 7811 7791 7901 7797
rect 7811 7771 7827 7791
rect 7847 7789 7901 7791
rect 7847 7771 7872 7789
rect 7811 7769 7872 7771
rect 7892 7769 7901 7789
rect 7811 7763 7901 7769
rect 7824 7709 7861 7710
rect 7920 7709 7957 7710
rect 7976 7709 8012 7819
rect 8199 7798 8230 7819
rect 8977 7804 9024 7847
rect 9380 7842 9420 7847
rect 10045 7845 10232 7869
rect 10263 7850 10656 7870
rect 10676 7850 10679 7870
rect 10263 7845 10679 7850
rect 8195 7797 8230 7798
rect 8073 7787 8230 7797
rect 8073 7767 8090 7787
rect 8110 7767 8230 7787
rect 8073 7760 8230 7767
rect 8297 7790 8446 7798
rect 8297 7770 8308 7790
rect 8328 7770 8367 7790
rect 8387 7770 8446 7790
rect 8977 7786 8987 7804
rect 9005 7786 9024 7804
rect 8977 7782 9024 7786
rect 8978 7777 9015 7782
rect 8297 7763 8446 7770
rect 10045 7774 10082 7845
rect 10263 7844 10604 7845
rect 10197 7784 10228 7785
rect 8297 7762 8338 7763
rect 8534 7761 8571 7764
rect 8031 7709 8068 7710
rect 7724 7700 7862 7709
rect 6928 7661 7372 7687
rect 6928 7659 7096 7661
rect 5881 7527 6328 7539
rect 5924 7525 5957 7527
rect 5291 7507 5429 7516
rect 5085 7506 5122 7507
rect 4815 7453 4856 7454
rect 4589 7432 4641 7450
rect 4707 7446 4856 7453
rect 4157 7412 4197 7422
rect 4707 7426 4766 7446
rect 4786 7426 4825 7446
rect 4845 7426 4856 7446
rect 4707 7418 4856 7426
rect 4923 7449 5080 7456
rect 4923 7429 5043 7449
rect 5063 7429 5080 7449
rect 4923 7419 5080 7429
rect 4923 7418 4958 7419
rect 3987 7395 4025 7404
rect 4923 7397 4954 7418
rect 5141 7397 5177 7507
rect 5196 7506 5233 7507
rect 5292 7506 5329 7507
rect 5252 7447 5342 7453
rect 5252 7427 5261 7447
rect 5281 7445 5342 7447
rect 5281 7427 5306 7445
rect 5252 7425 5306 7427
rect 5326 7425 5342 7445
rect 5252 7419 5342 7425
rect 4766 7396 4803 7397
rect 3987 7394 4024 7395
rect 3448 7366 3538 7372
rect 3448 7346 3464 7366
rect 3484 7364 3538 7366
rect 3484 7346 3509 7364
rect 3448 7344 3509 7346
rect 3529 7344 3538 7364
rect 3448 7338 3538 7344
rect 3461 7284 3498 7285
rect 3557 7284 3594 7285
rect 3613 7284 3649 7394
rect 3836 7373 3867 7394
rect 4765 7387 4803 7396
rect 3832 7372 3867 7373
rect 3710 7362 3867 7372
rect 3710 7342 3727 7362
rect 3747 7342 3867 7362
rect 3710 7335 3867 7342
rect 3934 7365 4083 7373
rect 3934 7345 3945 7365
rect 3965 7345 4004 7365
rect 4024 7345 4083 7365
rect 4593 7369 4633 7379
rect 3934 7338 4083 7345
rect 4149 7341 4201 7359
rect 3934 7337 3975 7338
rect 3668 7284 3705 7285
rect 3361 7275 3499 7284
rect 2428 7267 2465 7268
rect 2399 7266 2567 7267
rect 2693 7266 2733 7268
rect 2224 7257 2263 7263
rect 2224 7235 2232 7257
rect 2256 7235 2263 7257
rect 1926 7128 1963 7136
rect 1926 7109 1934 7128
rect 1955 7109 1963 7128
rect 1926 7103 1963 7109
rect 1528 6858 1536 6880
rect 1560 6858 1568 6880
rect 1528 6850 1568 6858
rect 216 6812 661 6842
rect 1699 6825 1764 6826
rect 216 6809 639 6812
rect 216 6761 263 6809
rect 216 6743 226 6761
rect 244 6743 263 6761
rect 216 6739 263 6743
rect 1350 6800 1537 6824
rect 1568 6805 1961 6825
rect 1981 6805 1984 6825
rect 1568 6800 1984 6805
rect 217 6734 254 6739
rect 1350 6729 1387 6800
rect 1568 6799 1909 6800
rect 1502 6739 1533 6740
rect 1350 6709 1359 6729
rect 1379 6709 1387 6729
rect 1350 6699 1387 6709
rect 1446 6729 1533 6739
rect 1446 6709 1455 6729
rect 1475 6709 1533 6729
rect 1446 6700 1533 6709
rect 1446 6699 1483 6700
rect 205 6672 257 6674
rect 203 6668 636 6672
rect 203 6662 642 6668
rect 203 6644 224 6662
rect 242 6644 642 6662
rect 1502 6649 1533 6700
rect 1568 6729 1605 6799
rect 1871 6798 1908 6799
rect 1720 6739 1756 6740
rect 1568 6709 1577 6729
rect 1597 6709 1605 6729
rect 1568 6699 1605 6709
rect 1664 6729 1812 6739
rect 1912 6736 2008 6738
rect 1664 6709 1673 6729
rect 1693 6709 1783 6729
rect 1803 6709 1812 6729
rect 1664 6700 1812 6709
rect 1870 6729 2008 6736
rect 1870 6709 1879 6729
rect 1899 6709 2008 6729
rect 1870 6700 2008 6709
rect 1664 6699 1701 6700
rect 1394 6646 1435 6647
rect 203 6626 642 6644
rect 205 6437 257 6626
rect 603 6601 642 6626
rect 1286 6639 1435 6646
rect 1286 6619 1345 6639
rect 1365 6619 1404 6639
rect 1424 6619 1435 6639
rect 1286 6611 1435 6619
rect 1502 6642 1659 6649
rect 1502 6622 1622 6642
rect 1642 6622 1659 6642
rect 1502 6612 1659 6622
rect 1502 6611 1537 6612
rect 387 6576 574 6600
rect 603 6581 998 6601
rect 1018 6581 1021 6601
rect 1502 6590 1533 6611
rect 1720 6590 1756 6700
rect 1775 6699 1812 6700
rect 1871 6699 1908 6700
rect 1831 6640 1921 6646
rect 1831 6620 1840 6640
rect 1860 6638 1921 6640
rect 1860 6620 1885 6638
rect 1831 6618 1885 6620
rect 1905 6618 1921 6638
rect 1831 6612 1921 6618
rect 1345 6589 1382 6590
rect 603 6576 1021 6581
rect 1344 6580 1382 6589
rect 387 6505 424 6576
rect 603 6575 946 6576
rect 603 6572 642 6575
rect 908 6574 945 6575
rect 539 6515 570 6516
rect 387 6485 396 6505
rect 416 6485 424 6505
rect 387 6475 424 6485
rect 483 6505 570 6515
rect 483 6485 492 6505
rect 512 6485 570 6505
rect 483 6476 570 6485
rect 483 6475 520 6476
rect 205 6419 221 6437
rect 239 6419 257 6437
rect 539 6425 570 6476
rect 605 6505 642 6572
rect 1344 6560 1353 6580
rect 1373 6560 1382 6580
rect 1344 6552 1382 6560
rect 1448 6584 1533 6590
rect 1563 6589 1600 6590
rect 1448 6564 1456 6584
rect 1476 6564 1533 6584
rect 1448 6556 1533 6564
rect 1562 6580 1600 6589
rect 1562 6560 1571 6580
rect 1591 6560 1600 6580
rect 1448 6555 1484 6556
rect 1562 6552 1600 6560
rect 1666 6584 1810 6590
rect 1666 6564 1674 6584
rect 1694 6583 1782 6584
rect 1694 6565 1729 6583
rect 1747 6565 1782 6583
rect 1694 6564 1782 6565
rect 1802 6564 1810 6584
rect 1666 6556 1810 6564
rect 1666 6555 1702 6556
rect 1774 6555 1810 6556
rect 1876 6589 1913 6590
rect 1876 6588 1914 6589
rect 1876 6580 1940 6588
rect 1876 6560 1885 6580
rect 1905 6566 1940 6580
rect 1960 6566 1963 6586
rect 1905 6561 1963 6566
rect 1905 6560 1940 6561
rect 1345 6523 1382 6552
rect 1346 6521 1382 6523
rect 757 6515 793 6516
rect 605 6485 614 6505
rect 634 6485 642 6505
rect 605 6475 642 6485
rect 701 6505 849 6515
rect 949 6512 1045 6514
rect 701 6485 710 6505
rect 730 6485 820 6505
rect 840 6485 849 6505
rect 701 6476 849 6485
rect 907 6505 1045 6512
rect 907 6485 916 6505
rect 936 6485 1045 6505
rect 1346 6499 1537 6521
rect 1563 6520 1600 6552
rect 1876 6548 1940 6560
rect 1980 6524 2007 6700
rect 1926 6522 2007 6524
rect 1839 6520 2007 6522
rect 1563 6494 2007 6520
rect 1673 6492 1713 6494
rect 1839 6493 2007 6494
rect 907 6476 1045 6485
rect 1948 6491 2007 6493
rect 701 6475 738 6476
rect 431 6422 472 6423
rect 205 6401 257 6419
rect 323 6415 472 6422
rect 323 6395 382 6415
rect 402 6395 441 6415
rect 461 6395 472 6415
rect 323 6387 472 6395
rect 539 6418 696 6425
rect 539 6398 659 6418
rect 679 6398 696 6418
rect 539 6388 696 6398
rect 539 6387 574 6388
rect 539 6366 570 6387
rect 757 6366 793 6476
rect 812 6475 849 6476
rect 908 6475 945 6476
rect 868 6416 958 6422
rect 868 6396 877 6416
rect 897 6414 958 6416
rect 897 6396 922 6414
rect 868 6394 922 6396
rect 942 6394 958 6414
rect 868 6388 958 6394
rect 382 6365 419 6366
rect 381 6356 419 6365
rect 209 6338 249 6348
rect 209 6320 219 6338
rect 237 6320 249 6338
rect 381 6336 390 6356
rect 410 6336 419 6356
rect 381 6328 419 6336
rect 485 6360 570 6366
rect 600 6365 637 6366
rect 485 6340 493 6360
rect 513 6340 570 6360
rect 485 6332 570 6340
rect 599 6356 637 6365
rect 599 6336 608 6356
rect 628 6336 637 6356
rect 485 6331 521 6332
rect 599 6328 637 6336
rect 703 6360 847 6366
rect 703 6340 711 6360
rect 731 6340 764 6360
rect 784 6340 819 6360
rect 839 6340 847 6360
rect 703 6332 847 6340
rect 703 6331 739 6332
rect 811 6331 847 6332
rect 913 6365 950 6366
rect 913 6364 951 6365
rect 913 6356 977 6364
rect 913 6336 922 6356
rect 942 6342 977 6356
rect 997 6342 1000 6362
rect 942 6337 1000 6342
rect 942 6336 977 6337
rect 209 6264 249 6320
rect 382 6299 419 6328
rect 383 6297 419 6299
rect 383 6275 574 6297
rect 600 6296 637 6328
rect 913 6324 977 6336
rect 1017 6298 1044 6476
rect 1948 6473 1977 6491
rect 876 6296 1044 6298
rect 600 6286 1044 6296
rect 1185 6392 1372 6416
rect 1403 6397 1796 6417
rect 1816 6397 1819 6417
rect 1403 6392 1819 6397
rect 1185 6321 1222 6392
rect 1403 6391 1744 6392
rect 1337 6331 1368 6332
rect 1185 6301 1194 6321
rect 1214 6301 1222 6321
rect 1185 6291 1222 6301
rect 1281 6321 1368 6331
rect 1281 6301 1290 6321
rect 1310 6301 1368 6321
rect 1281 6292 1368 6301
rect 1281 6291 1318 6292
rect 206 6259 249 6264
rect 597 6270 1044 6286
rect 597 6264 625 6270
rect 876 6269 1044 6270
rect 206 6256 356 6259
rect 597 6256 624 6264
rect 206 6254 624 6256
rect 206 6236 215 6254
rect 233 6236 624 6254
rect 1337 6241 1368 6292
rect 1403 6321 1440 6391
rect 1706 6390 1743 6391
rect 1555 6331 1591 6332
rect 1403 6301 1412 6321
rect 1432 6301 1440 6321
rect 1403 6291 1440 6301
rect 1499 6321 1647 6331
rect 1747 6328 1843 6330
rect 1499 6301 1508 6321
rect 1528 6301 1618 6321
rect 1638 6301 1647 6321
rect 1499 6292 1647 6301
rect 1705 6321 1843 6328
rect 1705 6301 1714 6321
rect 1734 6301 1843 6321
rect 1705 6292 1843 6301
rect 1499 6291 1536 6292
rect 1229 6238 1270 6239
rect 206 6233 624 6236
rect 206 6227 249 6233
rect 209 6224 249 6227
rect 1121 6231 1270 6238
rect 606 6215 646 6216
rect 317 6198 646 6215
rect 1121 6211 1180 6231
rect 1200 6211 1239 6231
rect 1259 6211 1270 6231
rect 1121 6203 1270 6211
rect 1337 6234 1494 6241
rect 1337 6214 1457 6234
rect 1477 6214 1494 6234
rect 1337 6204 1494 6214
rect 1337 6203 1372 6204
rect 201 6155 244 6166
rect 201 6137 213 6155
rect 231 6137 244 6155
rect 201 6111 244 6137
rect 317 6111 344 6198
rect 606 6189 646 6198
rect 201 6090 344 6111
rect 388 6163 422 6179
rect 606 6169 999 6189
rect 1019 6169 1022 6189
rect 1337 6182 1368 6203
rect 1555 6182 1591 6292
rect 1610 6291 1647 6292
rect 1706 6291 1743 6292
rect 1666 6232 1756 6238
rect 1666 6212 1675 6232
rect 1695 6230 1756 6232
rect 1695 6212 1720 6230
rect 1666 6210 1720 6212
rect 1740 6210 1756 6230
rect 1666 6204 1756 6210
rect 1180 6181 1217 6182
rect 606 6164 1022 6169
rect 1179 6172 1217 6181
rect 606 6163 947 6164
rect 388 6093 425 6163
rect 540 6103 571 6104
rect 201 6088 338 6090
rect 201 6046 244 6088
rect 388 6073 397 6093
rect 417 6073 425 6093
rect 388 6063 425 6073
rect 484 6093 571 6103
rect 484 6073 493 6093
rect 513 6073 571 6093
rect 484 6064 571 6073
rect 484 6063 521 6064
rect 199 6036 244 6046
rect 199 6018 208 6036
rect 226 6018 244 6036
rect 199 6012 244 6018
rect 540 6013 571 6064
rect 606 6093 643 6163
rect 909 6162 946 6163
rect 1179 6152 1188 6172
rect 1208 6152 1217 6172
rect 1179 6144 1217 6152
rect 1283 6176 1368 6182
rect 1398 6181 1435 6182
rect 1283 6156 1291 6176
rect 1311 6156 1368 6176
rect 1283 6148 1368 6156
rect 1397 6172 1435 6181
rect 1397 6152 1406 6172
rect 1426 6152 1435 6172
rect 1283 6147 1319 6148
rect 1397 6144 1435 6152
rect 1501 6176 1645 6182
rect 1501 6156 1509 6176
rect 1529 6157 1561 6176
rect 1582 6157 1617 6176
rect 1529 6156 1617 6157
rect 1637 6156 1645 6176
rect 1501 6148 1645 6156
rect 1501 6147 1537 6148
rect 1609 6147 1645 6148
rect 1711 6181 1748 6182
rect 1711 6180 1749 6181
rect 1711 6172 1775 6180
rect 1711 6152 1720 6172
rect 1740 6158 1775 6172
rect 1795 6158 1798 6178
rect 1740 6153 1798 6158
rect 1740 6152 1775 6153
rect 1180 6115 1217 6144
rect 1181 6113 1217 6115
rect 758 6103 794 6104
rect 606 6073 615 6093
rect 635 6073 643 6093
rect 606 6063 643 6073
rect 702 6093 850 6103
rect 950 6100 1046 6102
rect 702 6073 711 6093
rect 731 6073 821 6093
rect 841 6073 850 6093
rect 702 6064 850 6073
rect 908 6093 1046 6100
rect 908 6073 917 6093
rect 937 6073 1046 6093
rect 1181 6091 1372 6113
rect 1398 6112 1435 6144
rect 1711 6140 1775 6152
rect 1815 6114 1842 6292
rect 1674 6112 1842 6114
rect 1398 6086 1842 6112
rect 908 6064 1046 6073
rect 702 6063 739 6064
rect 199 6009 236 6012
rect 432 6010 473 6011
rect 324 6003 473 6010
rect 324 5983 383 6003
rect 403 5983 442 6003
rect 462 5983 473 6003
rect 324 5975 473 5983
rect 540 6006 697 6013
rect 540 5986 660 6006
rect 680 5986 697 6006
rect 540 5976 697 5986
rect 540 5975 575 5976
rect 540 5954 571 5975
rect 758 5954 794 6064
rect 813 6063 850 6064
rect 909 6063 946 6064
rect 869 6004 959 6010
rect 869 5984 878 6004
rect 898 6002 959 6004
rect 898 5984 923 6002
rect 869 5982 923 5984
rect 943 5982 959 6002
rect 869 5976 959 5982
rect 383 5953 420 5954
rect 196 5945 233 5947
rect 196 5937 238 5945
rect 196 5919 206 5937
rect 224 5919 238 5937
rect 196 5910 238 5919
rect 382 5944 420 5953
rect 382 5924 391 5944
rect 411 5924 420 5944
rect 382 5916 420 5924
rect 486 5948 571 5954
rect 601 5953 638 5954
rect 486 5928 494 5948
rect 514 5928 571 5948
rect 486 5920 571 5928
rect 600 5944 638 5953
rect 600 5924 609 5944
rect 629 5924 638 5944
rect 486 5919 522 5920
rect 600 5916 638 5924
rect 704 5952 848 5954
rect 704 5948 756 5952
rect 704 5928 712 5948
rect 732 5932 756 5948
rect 776 5948 848 5952
rect 776 5932 820 5948
rect 732 5928 820 5932
rect 840 5928 848 5948
rect 704 5920 848 5928
rect 704 5919 740 5920
rect 812 5919 848 5920
rect 914 5953 951 5954
rect 914 5952 952 5953
rect 914 5944 978 5952
rect 914 5924 923 5944
rect 943 5930 978 5944
rect 998 5930 1001 5950
rect 943 5925 1001 5930
rect 943 5924 978 5925
rect 197 5885 238 5910
rect 383 5885 420 5916
rect 601 5885 638 5916
rect 914 5912 978 5924
rect 1018 5886 1045 6064
rect 197 5858 246 5885
rect 382 5859 431 5885
rect 600 5884 681 5885
rect 877 5884 1045 5886
rect 600 5859 1045 5884
rect 601 5858 1045 5859
rect 199 5825 246 5858
rect 602 5825 642 5858
rect 877 5857 1045 5858
rect 1508 5862 1548 6086
rect 1674 6085 1842 6086
rect 1508 5840 1516 5862
rect 1540 5840 1548 5862
rect 1508 5832 1548 5840
rect 199 5786 642 5825
rect 199 5743 246 5786
rect 602 5781 642 5786
rect 1267 5784 1454 5808
rect 1485 5789 1878 5809
rect 1898 5789 1901 5809
rect 1485 5784 1901 5789
rect 199 5725 209 5743
rect 227 5725 246 5743
rect 199 5721 246 5725
rect 200 5716 237 5721
rect 1267 5713 1304 5784
rect 1485 5783 1826 5784
rect 1419 5723 1450 5724
rect 1267 5693 1276 5713
rect 1296 5693 1304 5713
rect 1267 5683 1304 5693
rect 1363 5713 1450 5723
rect 1363 5693 1372 5713
rect 1392 5693 1450 5713
rect 1363 5684 1450 5693
rect 1363 5683 1400 5684
rect 188 5654 240 5656
rect 186 5650 619 5654
rect 186 5644 625 5650
rect 186 5626 207 5644
rect 225 5626 625 5644
rect 1419 5633 1450 5684
rect 1485 5713 1522 5783
rect 1788 5782 1825 5783
rect 1637 5723 1673 5724
rect 1485 5693 1494 5713
rect 1514 5693 1522 5713
rect 1485 5683 1522 5693
rect 1581 5713 1729 5723
rect 1829 5720 1925 5722
rect 1581 5693 1590 5713
rect 1610 5693 1700 5713
rect 1720 5693 1729 5713
rect 1581 5684 1729 5693
rect 1787 5713 1925 5720
rect 1787 5693 1796 5713
rect 1816 5693 1925 5713
rect 1787 5684 1925 5693
rect 1581 5683 1618 5684
rect 1311 5630 1352 5631
rect 186 5608 625 5626
rect 188 5419 240 5608
rect 586 5583 625 5608
rect 1203 5623 1352 5630
rect 1203 5603 1262 5623
rect 1282 5603 1321 5623
rect 1341 5603 1352 5623
rect 1203 5595 1352 5603
rect 1419 5626 1576 5633
rect 1419 5606 1539 5626
rect 1559 5606 1576 5626
rect 1419 5596 1576 5606
rect 1419 5595 1454 5596
rect 370 5558 557 5582
rect 586 5563 981 5583
rect 1001 5563 1004 5583
rect 1419 5574 1450 5595
rect 1637 5574 1673 5684
rect 1692 5683 1729 5684
rect 1788 5683 1825 5684
rect 1748 5624 1838 5630
rect 1748 5604 1757 5624
rect 1777 5622 1838 5624
rect 1777 5604 1802 5622
rect 1748 5602 1802 5604
rect 1822 5602 1838 5622
rect 1748 5596 1838 5602
rect 1262 5573 1299 5574
rect 586 5558 1004 5563
rect 1261 5564 1299 5573
rect 370 5487 407 5558
rect 586 5557 929 5558
rect 586 5554 625 5557
rect 891 5556 928 5557
rect 522 5497 553 5498
rect 370 5467 379 5487
rect 399 5467 407 5487
rect 370 5457 407 5467
rect 466 5487 553 5497
rect 466 5467 475 5487
rect 495 5467 553 5487
rect 466 5458 553 5467
rect 466 5457 503 5458
rect 188 5401 204 5419
rect 222 5401 240 5419
rect 522 5407 553 5458
rect 588 5487 625 5554
rect 1261 5544 1270 5564
rect 1290 5544 1299 5564
rect 1261 5536 1299 5544
rect 1365 5568 1450 5574
rect 1480 5573 1517 5574
rect 1365 5548 1373 5568
rect 1393 5548 1450 5568
rect 1365 5540 1450 5548
rect 1479 5564 1517 5573
rect 1479 5544 1488 5564
rect 1508 5544 1517 5564
rect 1365 5539 1401 5540
rect 1479 5536 1517 5544
rect 1583 5568 1727 5574
rect 1583 5548 1591 5568
rect 1611 5563 1699 5568
rect 1611 5548 1647 5563
rect 1583 5546 1647 5548
rect 1666 5548 1699 5563
rect 1719 5548 1727 5568
rect 1666 5546 1727 5548
rect 1583 5540 1727 5546
rect 1583 5539 1619 5540
rect 1691 5539 1727 5540
rect 1793 5573 1830 5574
rect 1793 5572 1831 5573
rect 1793 5564 1857 5572
rect 1793 5544 1802 5564
rect 1822 5550 1857 5564
rect 1877 5550 1880 5570
rect 1822 5545 1880 5550
rect 1822 5544 1857 5545
rect 1262 5507 1299 5536
rect 1263 5505 1299 5507
rect 740 5497 776 5498
rect 588 5467 597 5487
rect 617 5467 625 5487
rect 588 5457 625 5467
rect 684 5487 832 5497
rect 932 5494 1028 5496
rect 684 5467 693 5487
rect 713 5467 803 5487
rect 823 5467 832 5487
rect 684 5458 832 5467
rect 890 5487 1028 5494
rect 890 5467 899 5487
rect 919 5467 1028 5487
rect 1263 5483 1454 5505
rect 1480 5504 1517 5536
rect 1793 5532 1857 5544
rect 1897 5506 1924 5684
rect 1756 5504 1924 5506
rect 1480 5490 1924 5504
rect 1948 5527 1976 6473
rect 1948 5497 1993 5527
rect 1480 5478 1927 5490
rect 1523 5476 1556 5478
rect 890 5458 1028 5467
rect 684 5457 721 5458
rect 414 5404 455 5405
rect 188 5383 240 5401
rect 306 5397 455 5404
rect 306 5377 365 5397
rect 385 5377 424 5397
rect 444 5377 455 5397
rect 306 5369 455 5377
rect 522 5400 679 5407
rect 522 5380 642 5400
rect 662 5380 679 5400
rect 522 5370 679 5380
rect 522 5369 557 5370
rect 522 5348 553 5369
rect 740 5348 776 5458
rect 795 5457 832 5458
rect 891 5457 928 5458
rect 851 5398 941 5404
rect 851 5378 860 5398
rect 880 5396 941 5398
rect 880 5378 905 5396
rect 851 5376 905 5378
rect 925 5376 941 5396
rect 851 5370 941 5376
rect 365 5347 402 5348
rect 364 5338 402 5347
rect 192 5320 232 5330
rect 192 5302 202 5320
rect 220 5302 232 5320
rect 364 5318 373 5338
rect 393 5318 402 5338
rect 364 5310 402 5318
rect 468 5342 553 5348
rect 583 5347 620 5348
rect 468 5322 476 5342
rect 496 5322 553 5342
rect 468 5314 553 5322
rect 582 5338 620 5347
rect 582 5318 591 5338
rect 611 5318 620 5338
rect 468 5313 504 5314
rect 582 5310 620 5318
rect 686 5342 830 5348
rect 686 5322 694 5342
rect 714 5322 747 5342
rect 767 5322 802 5342
rect 822 5322 830 5342
rect 686 5314 830 5322
rect 686 5313 722 5314
rect 794 5313 830 5314
rect 896 5347 933 5348
rect 896 5346 934 5347
rect 896 5338 960 5346
rect 896 5318 905 5338
rect 925 5324 960 5338
rect 980 5324 983 5344
rect 925 5319 983 5324
rect 925 5318 960 5319
rect 192 5246 232 5302
rect 365 5281 402 5310
rect 366 5279 402 5281
rect 366 5257 557 5279
rect 583 5278 620 5310
rect 896 5306 960 5318
rect 1000 5280 1027 5458
rect 1885 5433 1927 5478
rect 1948 5479 1959 5497
rect 1981 5479 1993 5497
rect 1948 5473 1993 5479
rect 1949 5472 1993 5473
rect 859 5278 1027 5280
rect 583 5268 1027 5278
rect 1168 5374 1355 5398
rect 1386 5379 1779 5399
rect 1799 5379 1802 5399
rect 1386 5374 1802 5379
rect 1168 5303 1205 5374
rect 1386 5373 1727 5374
rect 1320 5313 1351 5314
rect 1168 5283 1177 5303
rect 1197 5283 1205 5303
rect 1168 5273 1205 5283
rect 1264 5303 1351 5313
rect 1264 5283 1273 5303
rect 1293 5283 1351 5303
rect 1264 5274 1351 5283
rect 1264 5273 1301 5274
rect 189 5241 232 5246
rect 580 5252 1027 5268
rect 580 5246 608 5252
rect 859 5251 1027 5252
rect 189 5238 339 5241
rect 580 5238 607 5246
rect 189 5236 607 5238
rect 189 5218 198 5236
rect 216 5218 607 5236
rect 1320 5223 1351 5274
rect 1386 5303 1423 5373
rect 1689 5372 1726 5373
rect 1538 5313 1574 5314
rect 1386 5283 1395 5303
rect 1415 5283 1423 5303
rect 1386 5273 1423 5283
rect 1482 5303 1630 5313
rect 1730 5310 1826 5312
rect 1482 5283 1491 5303
rect 1511 5283 1601 5303
rect 1621 5283 1630 5303
rect 1482 5274 1630 5283
rect 1688 5303 1826 5310
rect 1688 5283 1697 5303
rect 1717 5283 1826 5303
rect 1688 5274 1826 5283
rect 1482 5273 1519 5274
rect 1212 5220 1253 5221
rect 189 5215 607 5218
rect 189 5209 232 5215
rect 192 5206 232 5209
rect 1107 5213 1253 5220
rect 589 5197 629 5198
rect 300 5180 629 5197
rect 1107 5193 1163 5213
rect 1183 5193 1222 5213
rect 1242 5193 1253 5213
rect 1107 5185 1253 5193
rect 1320 5216 1477 5223
rect 1320 5196 1440 5216
rect 1460 5196 1477 5216
rect 1320 5186 1477 5196
rect 1320 5185 1355 5186
rect 184 5137 227 5148
rect 184 5119 196 5137
rect 214 5119 227 5137
rect 184 5093 227 5119
rect 300 5093 327 5180
rect 589 5171 629 5180
rect 184 5072 327 5093
rect 371 5145 405 5161
rect 589 5151 982 5171
rect 1002 5151 1005 5171
rect 1320 5164 1351 5185
rect 1538 5164 1574 5274
rect 1593 5273 1630 5274
rect 1689 5273 1726 5274
rect 1649 5214 1739 5220
rect 1649 5194 1658 5214
rect 1678 5212 1739 5214
rect 1678 5194 1703 5212
rect 1649 5192 1703 5194
rect 1723 5192 1739 5212
rect 1649 5186 1739 5192
rect 1163 5163 1200 5164
rect 589 5146 1005 5151
rect 1162 5154 1200 5163
rect 589 5145 930 5146
rect 371 5075 408 5145
rect 523 5085 554 5086
rect 184 5070 321 5072
rect 184 5028 227 5070
rect 371 5055 380 5075
rect 400 5055 408 5075
rect 371 5045 408 5055
rect 467 5075 554 5085
rect 467 5055 476 5075
rect 496 5055 554 5075
rect 467 5046 554 5055
rect 467 5045 504 5046
rect 182 5018 227 5028
rect 182 5000 191 5018
rect 209 5000 227 5018
rect 182 4994 227 5000
rect 523 4995 554 5046
rect 589 5075 626 5145
rect 892 5144 929 5145
rect 1162 5134 1171 5154
rect 1191 5134 1200 5154
rect 1162 5126 1200 5134
rect 1266 5158 1351 5164
rect 1381 5163 1418 5164
rect 1266 5138 1274 5158
rect 1294 5138 1351 5158
rect 1266 5130 1351 5138
rect 1380 5154 1418 5163
rect 1380 5134 1389 5154
rect 1409 5134 1418 5154
rect 1266 5129 1302 5130
rect 1380 5126 1418 5134
rect 1484 5158 1628 5164
rect 1484 5138 1492 5158
rect 1512 5155 1600 5158
rect 1512 5138 1547 5155
rect 1484 5137 1547 5138
rect 1566 5138 1600 5155
rect 1620 5138 1628 5158
rect 1566 5137 1628 5138
rect 1484 5130 1628 5137
rect 1484 5129 1520 5130
rect 1592 5129 1628 5130
rect 1694 5163 1731 5164
rect 1694 5162 1732 5163
rect 1754 5162 1781 5166
rect 1694 5160 1781 5162
rect 1694 5154 1758 5160
rect 1694 5134 1703 5154
rect 1723 5140 1758 5154
rect 1778 5140 1781 5160
rect 1723 5135 1781 5140
rect 1723 5134 1758 5135
rect 1163 5097 1200 5126
rect 1164 5095 1200 5097
rect 741 5085 777 5086
rect 589 5055 598 5075
rect 618 5055 626 5075
rect 589 5045 626 5055
rect 685 5075 833 5085
rect 933 5082 1029 5084
rect 685 5055 694 5075
rect 714 5055 804 5075
rect 824 5055 833 5075
rect 685 5046 833 5055
rect 891 5075 1029 5082
rect 891 5055 900 5075
rect 920 5055 1029 5075
rect 1164 5073 1355 5095
rect 1381 5094 1418 5126
rect 1694 5122 1758 5134
rect 1798 5096 1825 5274
rect 1657 5094 1825 5096
rect 1381 5068 1825 5094
rect 891 5046 1029 5055
rect 685 5045 722 5046
rect 182 4991 219 4994
rect 415 4992 456 4993
rect 307 4985 456 4992
rect 307 4965 366 4985
rect 386 4965 425 4985
rect 445 4965 456 4985
rect 307 4957 456 4965
rect 523 4988 680 4995
rect 523 4968 643 4988
rect 663 4968 680 4988
rect 523 4958 680 4968
rect 523 4957 558 4958
rect 523 4936 554 4957
rect 741 4936 777 5046
rect 796 5045 833 5046
rect 892 5045 929 5046
rect 852 4986 942 4992
rect 852 4966 861 4986
rect 881 4984 942 4986
rect 881 4966 906 4984
rect 852 4964 906 4966
rect 926 4964 942 4984
rect 852 4958 942 4964
rect 366 4935 403 4936
rect 179 4927 216 4929
rect 179 4919 221 4927
rect 179 4901 189 4919
rect 207 4901 221 4919
rect 179 4892 221 4901
rect 365 4926 403 4935
rect 365 4906 374 4926
rect 394 4906 403 4926
rect 365 4898 403 4906
rect 469 4930 554 4936
rect 584 4935 621 4936
rect 469 4910 477 4930
rect 497 4910 554 4930
rect 469 4902 554 4910
rect 583 4926 621 4935
rect 583 4906 592 4926
rect 612 4906 621 4926
rect 469 4901 505 4902
rect 583 4898 621 4906
rect 687 4934 831 4936
rect 687 4930 739 4934
rect 687 4910 695 4930
rect 715 4914 739 4930
rect 759 4930 831 4934
rect 759 4914 803 4930
rect 715 4910 803 4914
rect 823 4910 831 4930
rect 687 4902 831 4910
rect 687 4901 723 4902
rect 795 4901 831 4902
rect 897 4935 934 4936
rect 897 4934 935 4935
rect 897 4926 961 4934
rect 897 4906 906 4926
rect 926 4912 961 4926
rect 981 4912 984 4932
rect 926 4907 984 4912
rect 926 4906 961 4907
rect 180 4867 221 4892
rect 366 4867 403 4898
rect 584 4867 621 4898
rect 897 4894 961 4906
rect 1001 4868 1028 5046
rect 180 4833 223 4867
rect 362 4841 429 4867
rect 584 4866 664 4867
rect 860 4866 1028 4868
rect 584 4840 1028 4866
rect 180 4822 227 4833
rect 584 4823 619 4840
rect 860 4839 1028 4840
rect 1491 4844 1531 5068
rect 1657 5067 1825 5068
rect 1889 5100 1922 5433
rect 2224 5420 2263 7235
rect 2399 7241 2843 7266
rect 2399 7060 2426 7241
rect 2568 7240 2843 7241
rect 2466 7200 2530 7212
rect 2806 7208 2843 7240
rect 2869 7239 3060 7261
rect 3361 7255 3470 7275
rect 3490 7255 3499 7275
rect 3361 7248 3499 7255
rect 3557 7275 3705 7284
rect 3557 7255 3566 7275
rect 3586 7255 3676 7275
rect 3696 7255 3705 7275
rect 3361 7246 3457 7248
rect 3557 7245 3705 7255
rect 3764 7275 3801 7285
rect 3764 7255 3772 7275
rect 3792 7255 3801 7275
rect 3613 7244 3649 7245
rect 3024 7237 3060 7239
rect 3024 7208 3061 7237
rect 2466 7199 2501 7200
rect 2443 7194 2501 7199
rect 2443 7174 2446 7194
rect 2466 7180 2501 7194
rect 2521 7180 2530 7200
rect 2466 7172 2530 7180
rect 2492 7171 2530 7172
rect 2493 7170 2530 7171
rect 2596 7204 2632 7205
rect 2704 7204 2740 7205
rect 2596 7196 2740 7204
rect 2596 7176 2604 7196
rect 2624 7194 2712 7196
rect 2624 7176 2657 7194
rect 2596 7172 2657 7176
rect 2680 7176 2712 7194
rect 2732 7176 2740 7196
rect 2680 7172 2740 7176
rect 2596 7170 2740 7172
rect 2806 7200 2844 7208
rect 2922 7204 2958 7205
rect 2806 7180 2815 7200
rect 2835 7180 2844 7200
rect 2806 7171 2844 7180
rect 2873 7196 2958 7204
rect 2873 7176 2930 7196
rect 2950 7176 2958 7196
rect 2806 7170 2843 7171
rect 2873 7170 2958 7176
rect 3024 7200 3062 7208
rect 3024 7180 3033 7200
rect 3053 7180 3062 7200
rect 3764 7188 3801 7255
rect 3836 7284 3867 7335
rect 4149 7323 4167 7341
rect 4185 7323 4201 7341
rect 3886 7284 3923 7285
rect 3836 7275 3923 7284
rect 3836 7255 3894 7275
rect 3914 7255 3923 7275
rect 3836 7245 3923 7255
rect 3982 7275 4019 7285
rect 3982 7255 3990 7275
rect 4010 7255 4019 7275
rect 3836 7244 3867 7245
rect 3461 7185 3498 7186
rect 3764 7185 3803 7188
rect 3460 7184 3803 7185
rect 3982 7184 4019 7255
rect 3024 7171 3062 7180
rect 3385 7179 3803 7184
rect 3024 7170 3061 7171
rect 2485 7142 2575 7148
rect 2485 7122 2501 7142
rect 2521 7140 2575 7142
rect 2521 7122 2546 7140
rect 2485 7120 2546 7122
rect 2566 7120 2575 7140
rect 2485 7114 2575 7120
rect 2498 7060 2535 7061
rect 2594 7060 2631 7061
rect 2650 7060 2686 7170
rect 2873 7149 2904 7170
rect 3385 7159 3388 7179
rect 3408 7159 3803 7179
rect 3832 7160 4019 7184
rect 2869 7148 2904 7149
rect 2747 7138 2904 7148
rect 2747 7118 2764 7138
rect 2784 7118 2904 7138
rect 2747 7111 2904 7118
rect 2971 7141 3120 7149
rect 2971 7121 2982 7141
rect 3002 7121 3041 7141
rect 3061 7121 3120 7141
rect 2971 7114 3120 7121
rect 3764 7134 3803 7159
rect 4149 7134 4201 7323
rect 4593 7351 4603 7369
rect 4621 7351 4633 7369
rect 4765 7367 4774 7387
rect 4794 7367 4803 7387
rect 4765 7359 4803 7367
rect 4869 7391 4954 7397
rect 4984 7396 5021 7397
rect 4869 7371 4877 7391
rect 4897 7371 4954 7391
rect 4869 7363 4954 7371
rect 4983 7387 5021 7396
rect 4983 7367 4992 7387
rect 5012 7367 5021 7387
rect 4869 7362 4905 7363
rect 4983 7359 5021 7367
rect 5087 7391 5231 7397
rect 5087 7371 5095 7391
rect 5115 7371 5148 7391
rect 5168 7371 5203 7391
rect 5223 7371 5231 7391
rect 5087 7363 5231 7371
rect 5087 7362 5123 7363
rect 5195 7362 5231 7363
rect 5297 7396 5334 7397
rect 5297 7395 5335 7396
rect 5297 7387 5361 7395
rect 5297 7367 5306 7387
rect 5326 7373 5361 7387
rect 5381 7373 5384 7393
rect 5326 7368 5384 7373
rect 5326 7367 5361 7368
rect 4593 7295 4633 7351
rect 4766 7330 4803 7359
rect 4767 7328 4803 7330
rect 4767 7306 4958 7328
rect 4984 7327 5021 7359
rect 5297 7355 5361 7367
rect 5401 7329 5428 7507
rect 6286 7482 6328 7527
rect 5260 7327 5428 7329
rect 4984 7317 5428 7327
rect 5569 7423 5756 7447
rect 5787 7428 6180 7448
rect 6200 7428 6203 7448
rect 5787 7423 6203 7428
rect 5569 7352 5606 7423
rect 5787 7422 6128 7423
rect 5721 7362 5752 7363
rect 5569 7332 5578 7352
rect 5598 7332 5606 7352
rect 5569 7322 5606 7332
rect 5665 7352 5752 7362
rect 5665 7332 5674 7352
rect 5694 7332 5752 7352
rect 5665 7323 5752 7332
rect 5665 7322 5702 7323
rect 4590 7290 4633 7295
rect 4981 7301 5428 7317
rect 4981 7295 5009 7301
rect 5260 7300 5428 7301
rect 4590 7287 4740 7290
rect 4981 7287 5008 7295
rect 4590 7285 5008 7287
rect 4590 7267 4599 7285
rect 4617 7267 5008 7285
rect 5721 7272 5752 7323
rect 5787 7352 5824 7422
rect 6090 7421 6127 7422
rect 5939 7362 5975 7363
rect 5787 7332 5796 7352
rect 5816 7332 5824 7352
rect 5787 7322 5824 7332
rect 5883 7352 6031 7362
rect 6131 7359 6227 7361
rect 5883 7332 5892 7352
rect 5912 7332 6002 7352
rect 6022 7332 6031 7352
rect 5883 7323 6031 7332
rect 6089 7352 6227 7359
rect 6089 7332 6098 7352
rect 6118 7332 6227 7352
rect 6089 7323 6227 7332
rect 5883 7322 5920 7323
rect 5613 7269 5654 7270
rect 4590 7264 5008 7267
rect 4590 7258 4633 7264
rect 4593 7255 4633 7258
rect 5508 7262 5654 7269
rect 4990 7246 5030 7247
rect 4701 7229 5030 7246
rect 5508 7242 5564 7262
rect 5584 7242 5623 7262
rect 5643 7242 5654 7262
rect 5508 7234 5654 7242
rect 5721 7265 5878 7272
rect 5721 7245 5841 7265
rect 5861 7245 5878 7265
rect 5721 7235 5878 7245
rect 5721 7234 5756 7235
rect 4585 7186 4628 7197
rect 4585 7168 4597 7186
rect 4615 7168 4628 7186
rect 4585 7142 4628 7168
rect 4701 7142 4728 7229
rect 4990 7220 5030 7229
rect 3764 7116 4203 7134
rect 2971 7113 3012 7114
rect 2705 7060 2742 7061
rect 2398 7051 2536 7060
rect 2398 7031 2507 7051
rect 2527 7031 2536 7051
rect 2398 7024 2536 7031
rect 2594 7051 2742 7060
rect 2594 7031 2603 7051
rect 2623 7031 2713 7051
rect 2733 7031 2742 7051
rect 2398 7022 2494 7024
rect 2594 7021 2742 7031
rect 2801 7051 2838 7061
rect 2801 7031 2809 7051
rect 2829 7031 2838 7051
rect 2650 7020 2686 7021
rect 2498 6961 2535 6962
rect 2801 6961 2838 7031
rect 2873 7060 2904 7111
rect 3764 7098 4164 7116
rect 4182 7098 4203 7116
rect 3764 7092 4203 7098
rect 3770 7088 4203 7092
rect 4585 7121 4728 7142
rect 4772 7194 4806 7210
rect 4990 7200 5383 7220
rect 5403 7200 5406 7220
rect 5721 7213 5752 7234
rect 5939 7213 5975 7323
rect 5994 7322 6031 7323
rect 6090 7322 6127 7323
rect 6050 7263 6140 7269
rect 6050 7243 6059 7263
rect 6079 7261 6140 7263
rect 6079 7243 6104 7261
rect 6050 7241 6104 7243
rect 6124 7241 6140 7261
rect 6050 7235 6140 7241
rect 5564 7212 5601 7213
rect 4990 7195 5406 7200
rect 5563 7203 5601 7212
rect 4990 7194 5331 7195
rect 4772 7124 4809 7194
rect 4924 7134 4955 7135
rect 4585 7119 4722 7121
rect 4149 7086 4201 7088
rect 4585 7077 4628 7119
rect 4772 7104 4781 7124
rect 4801 7104 4809 7124
rect 4772 7094 4809 7104
rect 4868 7124 4955 7134
rect 4868 7104 4877 7124
rect 4897 7104 4955 7124
rect 4868 7095 4955 7104
rect 4868 7094 4905 7095
rect 4583 7067 4628 7077
rect 2923 7060 2960 7061
rect 2873 7051 2960 7060
rect 2873 7031 2931 7051
rect 2951 7031 2960 7051
rect 2873 7021 2960 7031
rect 3019 7051 3056 7061
rect 3019 7031 3027 7051
rect 3047 7031 3056 7051
rect 4583 7049 4592 7067
rect 4610 7049 4628 7067
rect 4583 7043 4628 7049
rect 4924 7044 4955 7095
rect 4990 7124 5027 7194
rect 5293 7193 5330 7194
rect 5563 7183 5572 7203
rect 5592 7183 5601 7203
rect 5563 7175 5601 7183
rect 5667 7207 5752 7213
rect 5782 7212 5819 7213
rect 5667 7187 5675 7207
rect 5695 7187 5752 7207
rect 5667 7179 5752 7187
rect 5781 7203 5819 7212
rect 5781 7183 5790 7203
rect 5810 7183 5819 7203
rect 5667 7178 5703 7179
rect 5781 7175 5819 7183
rect 5885 7207 6029 7213
rect 5885 7187 5893 7207
rect 5913 7204 6001 7207
rect 5913 7187 5948 7204
rect 5885 7186 5948 7187
rect 5967 7187 6001 7204
rect 6021 7187 6029 7207
rect 5967 7186 6029 7187
rect 5885 7179 6029 7186
rect 5885 7178 5921 7179
rect 5993 7178 6029 7179
rect 6095 7212 6132 7213
rect 6095 7211 6133 7212
rect 6155 7211 6182 7215
rect 6095 7209 6182 7211
rect 6095 7203 6159 7209
rect 6095 7183 6104 7203
rect 6124 7189 6159 7203
rect 6179 7189 6182 7209
rect 6124 7184 6182 7189
rect 6124 7183 6159 7184
rect 5564 7146 5601 7175
rect 5565 7144 5601 7146
rect 5142 7134 5178 7135
rect 4990 7104 4999 7124
rect 5019 7104 5027 7124
rect 4990 7094 5027 7104
rect 5086 7124 5234 7134
rect 5334 7131 5430 7133
rect 5086 7104 5095 7124
rect 5115 7104 5205 7124
rect 5225 7104 5234 7124
rect 5086 7095 5234 7104
rect 5292 7124 5430 7131
rect 5292 7104 5301 7124
rect 5321 7104 5430 7124
rect 5565 7122 5756 7144
rect 5782 7143 5819 7175
rect 6095 7171 6159 7183
rect 6199 7145 6226 7323
rect 6058 7143 6226 7145
rect 5782 7117 6226 7143
rect 5292 7095 5430 7104
rect 5086 7094 5123 7095
rect 4583 7040 4620 7043
rect 4816 7041 4857 7042
rect 2873 7020 2904 7021
rect 2497 6960 2838 6961
rect 3019 6960 3056 7031
rect 4708 7034 4857 7041
rect 4152 7021 4189 7026
rect 2422 6955 2838 6960
rect 2422 6935 2425 6955
rect 2445 6935 2838 6955
rect 2869 6936 3056 6960
rect 4143 7017 4190 7021
rect 4143 6999 4162 7017
rect 4180 6999 4190 7017
rect 4708 7014 4767 7034
rect 4787 7014 4826 7034
rect 4846 7014 4857 7034
rect 4708 7006 4857 7014
rect 4924 7037 5081 7044
rect 4924 7017 5044 7037
rect 5064 7017 5081 7037
rect 4924 7007 5081 7017
rect 4924 7006 4959 7007
rect 4143 6951 4190 6999
rect 4924 6985 4955 7006
rect 5142 6985 5178 7095
rect 5197 7094 5234 7095
rect 5293 7094 5330 7095
rect 5253 7035 5343 7041
rect 5253 7015 5262 7035
rect 5282 7033 5343 7035
rect 5282 7015 5307 7033
rect 5253 7013 5307 7015
rect 5327 7013 5343 7033
rect 5253 7007 5343 7013
rect 4767 6984 4804 6985
rect 3767 6948 4190 6951
rect 2642 6934 2707 6935
rect 3745 6918 4190 6948
rect 4579 6976 4617 6978
rect 4579 6968 4622 6976
rect 4579 6950 4590 6968
rect 4608 6950 4622 6968
rect 4579 6923 4622 6950
rect 4766 6975 4804 6984
rect 4766 6955 4775 6975
rect 4795 6955 4804 6975
rect 4766 6947 4804 6955
rect 4870 6979 4955 6985
rect 4985 6984 5022 6985
rect 4870 6959 4878 6979
rect 4898 6959 4955 6979
rect 4870 6951 4955 6959
rect 4984 6975 5022 6984
rect 4984 6955 4993 6975
rect 5013 6955 5022 6975
rect 4870 6950 4906 6951
rect 4984 6947 5022 6955
rect 5088 6983 5232 6985
rect 5088 6979 5140 6983
rect 5088 6959 5096 6979
rect 5116 6963 5140 6979
rect 5160 6979 5232 6983
rect 5160 6963 5204 6979
rect 5116 6959 5204 6963
rect 5224 6959 5232 6979
rect 5088 6951 5232 6959
rect 5088 6950 5124 6951
rect 5196 6950 5232 6951
rect 5298 6984 5335 6985
rect 5298 6983 5336 6984
rect 5298 6975 5362 6983
rect 5298 6955 5307 6975
rect 5327 6961 5362 6975
rect 5382 6961 5385 6981
rect 5327 6956 5385 6961
rect 5327 6955 5362 6956
rect 2838 6902 2878 6910
rect 2838 6880 2846 6902
rect 2870 6880 2878 6902
rect 2443 6651 2480 6657
rect 2443 6632 2451 6651
rect 2472 6632 2480 6651
rect 2443 6624 2480 6632
rect 2447 6291 2480 6624
rect 2544 6656 2712 6657
rect 2838 6656 2878 6880
rect 3341 6884 3509 6885
rect 3745 6884 3786 6918
rect 4143 6897 4190 6918
rect 3341 6874 3786 6884
rect 3858 6882 4001 6883
rect 3341 6858 3785 6874
rect 3341 6856 3509 6858
rect 3705 6857 3785 6858
rect 3858 6857 4003 6882
rect 4145 6857 4190 6897
rect 3341 6678 3368 6856
rect 3408 6818 3472 6830
rect 3748 6826 3785 6857
rect 3966 6826 4003 6857
rect 4148 6850 4190 6857
rect 4580 6916 4622 6923
rect 4767 6916 4804 6947
rect 4985 6916 5022 6947
rect 5298 6943 5362 6955
rect 5402 6917 5429 7095
rect 4580 6876 4625 6916
rect 4767 6891 4912 6916
rect 4985 6915 5065 6916
rect 5261 6915 5429 6917
rect 4985 6899 5429 6915
rect 4769 6890 4912 6891
rect 4984 6889 5429 6899
rect 4580 6855 4627 6876
rect 4984 6855 5025 6889
rect 5261 6888 5429 6889
rect 5892 6893 5932 7117
rect 6058 7116 6226 7117
rect 6290 7149 6323 7482
rect 6928 7481 6955 7659
rect 6995 7621 7059 7633
rect 7335 7629 7372 7661
rect 7398 7660 7589 7682
rect 7724 7680 7833 7700
rect 7853 7680 7862 7700
rect 7724 7673 7862 7680
rect 7920 7700 8068 7709
rect 7920 7680 7929 7700
rect 7949 7680 8039 7700
rect 8059 7680 8068 7700
rect 7724 7671 7820 7673
rect 7920 7670 8068 7680
rect 8127 7700 8164 7710
rect 8127 7680 8135 7700
rect 8155 7680 8164 7700
rect 7976 7669 8012 7670
rect 7553 7658 7589 7660
rect 7553 7629 7590 7658
rect 6995 7620 7030 7621
rect 6972 7615 7030 7620
rect 6972 7595 6975 7615
rect 6995 7601 7030 7615
rect 7050 7601 7059 7621
rect 6995 7593 7059 7601
rect 7021 7592 7059 7593
rect 7022 7591 7059 7592
rect 7125 7625 7161 7626
rect 7233 7625 7269 7626
rect 7125 7617 7269 7625
rect 7125 7597 7133 7617
rect 7153 7616 7241 7617
rect 7153 7597 7188 7616
rect 7209 7597 7241 7616
rect 7261 7597 7269 7617
rect 7125 7591 7269 7597
rect 7335 7621 7373 7629
rect 7451 7625 7487 7626
rect 7335 7601 7344 7621
rect 7364 7601 7373 7621
rect 7335 7592 7373 7601
rect 7402 7617 7487 7625
rect 7402 7597 7459 7617
rect 7479 7597 7487 7617
rect 7335 7591 7372 7592
rect 7402 7591 7487 7597
rect 7553 7621 7591 7629
rect 7553 7601 7562 7621
rect 7582 7601 7591 7621
rect 7824 7610 7861 7611
rect 8127 7610 8164 7680
rect 8199 7709 8230 7760
rect 8526 7755 8571 7761
rect 8526 7737 8544 7755
rect 8562 7737 8571 7755
rect 10045 7754 10054 7774
rect 10074 7754 10082 7774
rect 10045 7744 10082 7754
rect 10141 7774 10228 7784
rect 10141 7754 10150 7774
rect 10170 7754 10228 7774
rect 10141 7745 10228 7754
rect 10141 7744 10178 7745
rect 8526 7727 8571 7737
rect 8249 7709 8286 7710
rect 8199 7700 8286 7709
rect 8199 7680 8257 7700
rect 8277 7680 8286 7700
rect 8199 7670 8286 7680
rect 8345 7700 8382 7710
rect 8345 7680 8353 7700
rect 8373 7680 8382 7700
rect 8526 7685 8569 7727
rect 8966 7715 9018 7717
rect 8432 7683 8569 7685
rect 8199 7669 8230 7670
rect 8345 7610 8382 7680
rect 7823 7609 8164 7610
rect 7553 7592 7591 7601
rect 7748 7604 8164 7609
rect 7553 7591 7590 7592
rect 7014 7563 7104 7569
rect 7014 7543 7030 7563
rect 7050 7561 7104 7563
rect 7050 7543 7075 7561
rect 7014 7541 7075 7543
rect 7095 7541 7104 7561
rect 7014 7535 7104 7541
rect 7027 7481 7064 7482
rect 7123 7481 7160 7482
rect 7179 7481 7215 7591
rect 7402 7570 7433 7591
rect 7748 7584 7751 7604
rect 7771 7584 8164 7604
rect 8348 7594 8382 7610
rect 8426 7662 8569 7683
rect 8964 7711 9397 7715
rect 8964 7705 9403 7711
rect 8964 7687 8985 7705
rect 9003 7687 9403 7705
rect 10197 7694 10228 7745
rect 10263 7774 10300 7844
rect 10566 7843 10603 7844
rect 10415 7784 10451 7785
rect 10263 7754 10272 7774
rect 10292 7754 10300 7774
rect 10263 7744 10300 7754
rect 10359 7774 10507 7784
rect 10607 7781 10703 7783
rect 10359 7754 10368 7774
rect 10388 7754 10478 7774
rect 10498 7754 10507 7774
rect 10359 7745 10507 7754
rect 10565 7774 10703 7781
rect 10565 7754 10574 7774
rect 10594 7754 10703 7774
rect 10565 7745 10703 7754
rect 10359 7744 10396 7745
rect 10089 7691 10130 7692
rect 8964 7669 9403 7687
rect 8124 7575 8164 7584
rect 8426 7575 8453 7662
rect 8526 7636 8569 7662
rect 8526 7618 8539 7636
rect 8557 7618 8569 7636
rect 8526 7607 8569 7618
rect 7398 7569 7433 7570
rect 7276 7559 7433 7569
rect 7276 7539 7293 7559
rect 7313 7539 7433 7559
rect 7276 7532 7433 7539
rect 7500 7562 7649 7570
rect 7500 7542 7511 7562
rect 7531 7542 7570 7562
rect 7590 7542 7649 7562
rect 8124 7558 8453 7575
rect 8124 7557 8164 7558
rect 7500 7535 7649 7542
rect 8521 7546 8561 7549
rect 8521 7540 8564 7546
rect 8146 7537 8564 7540
rect 7500 7534 7541 7535
rect 7234 7481 7271 7482
rect 6927 7472 7065 7481
rect 6790 7462 6826 7468
rect 6790 7444 6795 7462
rect 6817 7444 6826 7462
rect 6790 7440 6826 7444
rect 6927 7452 7036 7472
rect 7056 7452 7065 7472
rect 6927 7445 7065 7452
rect 7123 7472 7271 7481
rect 7123 7452 7132 7472
rect 7152 7452 7242 7472
rect 7262 7452 7271 7472
rect 6927 7443 7023 7445
rect 7123 7442 7271 7452
rect 7330 7472 7367 7482
rect 7330 7452 7338 7472
rect 7358 7452 7367 7472
rect 7179 7441 7215 7442
rect 6793 7281 6826 7440
rect 7027 7382 7064 7383
rect 7330 7382 7367 7452
rect 7402 7481 7433 7532
rect 8146 7519 8537 7537
rect 8555 7519 8564 7537
rect 8146 7517 8564 7519
rect 8146 7509 8173 7517
rect 8414 7514 8564 7517
rect 7726 7503 7894 7504
rect 8145 7503 8173 7509
rect 7726 7487 8173 7503
rect 8521 7509 8564 7514
rect 7452 7481 7489 7482
rect 7402 7472 7489 7481
rect 7402 7452 7460 7472
rect 7480 7452 7489 7472
rect 7402 7442 7489 7452
rect 7548 7472 7585 7482
rect 7548 7452 7556 7472
rect 7576 7452 7585 7472
rect 7402 7441 7433 7442
rect 7026 7381 7367 7382
rect 7548 7381 7585 7452
rect 6951 7376 7367 7381
rect 6951 7356 6954 7376
rect 6974 7356 7367 7376
rect 7398 7357 7585 7381
rect 7726 7477 8170 7487
rect 7726 7475 7894 7477
rect 7726 7297 7753 7475
rect 7793 7437 7857 7449
rect 8133 7445 8170 7477
rect 8196 7476 8387 7498
rect 8351 7474 8387 7476
rect 8351 7445 8388 7474
rect 8521 7453 8561 7509
rect 7793 7436 7828 7437
rect 7770 7431 7828 7436
rect 7770 7411 7773 7431
rect 7793 7417 7828 7431
rect 7848 7417 7857 7437
rect 7793 7409 7857 7417
rect 7819 7408 7857 7409
rect 7820 7407 7857 7408
rect 7923 7441 7959 7442
rect 8031 7441 8067 7442
rect 7923 7433 8067 7441
rect 7923 7413 7931 7433
rect 7951 7413 7986 7433
rect 8006 7413 8039 7433
rect 8059 7413 8067 7433
rect 7923 7407 8067 7413
rect 8133 7437 8171 7445
rect 8249 7441 8285 7442
rect 8133 7417 8142 7437
rect 8162 7417 8171 7437
rect 8133 7408 8171 7417
rect 8200 7433 8285 7441
rect 8200 7413 8257 7433
rect 8277 7413 8285 7433
rect 8133 7407 8170 7408
rect 8200 7407 8285 7413
rect 8351 7437 8389 7445
rect 8351 7417 8360 7437
rect 8380 7417 8389 7437
rect 8521 7435 8533 7453
rect 8551 7435 8561 7453
rect 8966 7480 9018 7669
rect 9364 7644 9403 7669
rect 9981 7684 10130 7691
rect 9981 7664 10040 7684
rect 10060 7664 10099 7684
rect 10119 7664 10130 7684
rect 9981 7656 10130 7664
rect 10197 7687 10354 7694
rect 10197 7667 10317 7687
rect 10337 7667 10354 7687
rect 10197 7657 10354 7667
rect 10197 7656 10232 7657
rect 9148 7619 9335 7643
rect 9364 7624 9759 7644
rect 9779 7624 9782 7644
rect 10197 7635 10228 7656
rect 10415 7635 10451 7745
rect 10470 7744 10507 7745
rect 10566 7744 10603 7745
rect 10526 7685 10616 7691
rect 10526 7665 10535 7685
rect 10555 7683 10616 7685
rect 10555 7665 10580 7683
rect 10526 7663 10580 7665
rect 10600 7663 10616 7683
rect 10526 7657 10616 7663
rect 10040 7634 10077 7635
rect 9364 7619 9782 7624
rect 10039 7625 10077 7634
rect 9148 7548 9185 7619
rect 9364 7618 9707 7619
rect 9364 7615 9403 7618
rect 9669 7617 9706 7618
rect 9300 7558 9331 7559
rect 9148 7528 9157 7548
rect 9177 7528 9185 7548
rect 9148 7518 9185 7528
rect 9244 7548 9331 7558
rect 9244 7528 9253 7548
rect 9273 7528 9331 7548
rect 9244 7519 9331 7528
rect 9244 7518 9281 7519
rect 8966 7462 8982 7480
rect 9000 7462 9018 7480
rect 9300 7468 9331 7519
rect 9366 7548 9403 7615
rect 10039 7605 10048 7625
rect 10068 7605 10077 7625
rect 10039 7597 10077 7605
rect 10143 7629 10228 7635
rect 10258 7634 10295 7635
rect 10143 7609 10151 7629
rect 10171 7609 10228 7629
rect 10143 7601 10228 7609
rect 10257 7625 10295 7634
rect 10257 7605 10266 7625
rect 10286 7605 10295 7625
rect 10143 7600 10179 7601
rect 10257 7597 10295 7605
rect 10361 7630 10505 7635
rect 10361 7629 10423 7630
rect 10361 7609 10369 7629
rect 10389 7611 10423 7629
rect 10444 7629 10505 7630
rect 10444 7611 10477 7629
rect 10389 7609 10477 7611
rect 10497 7609 10505 7629
rect 10361 7601 10505 7609
rect 10361 7600 10397 7601
rect 10469 7600 10505 7601
rect 10571 7634 10608 7635
rect 10571 7633 10609 7634
rect 10571 7625 10635 7633
rect 10571 7605 10580 7625
rect 10600 7611 10635 7625
rect 10655 7611 10658 7631
rect 10600 7606 10658 7611
rect 10600 7605 10635 7606
rect 10040 7568 10077 7597
rect 10041 7566 10077 7568
rect 9518 7558 9554 7559
rect 9366 7528 9375 7548
rect 9395 7528 9403 7548
rect 9366 7518 9403 7528
rect 9462 7548 9610 7558
rect 9710 7555 9806 7557
rect 9462 7528 9471 7548
rect 9491 7528 9581 7548
rect 9601 7528 9610 7548
rect 9462 7519 9610 7528
rect 9668 7548 9806 7555
rect 9668 7528 9677 7548
rect 9697 7528 9806 7548
rect 10041 7544 10232 7566
rect 10258 7565 10295 7597
rect 10571 7593 10635 7605
rect 10675 7567 10702 7745
rect 10534 7565 10702 7567
rect 10258 7551 10702 7565
rect 11305 7699 11473 7700
rect 11599 7699 11639 7923
rect 12102 7927 12270 7928
rect 12505 7927 12545 7960
rect 12901 7927 12948 7960
rect 13339 7959 13380 7984
rect 13525 7959 13562 7990
rect 13743 7959 13780 7990
rect 14056 7986 14120 7998
rect 14160 7960 14187 8138
rect 13339 7932 13388 7959
rect 13524 7933 13573 7959
rect 13742 7958 13823 7959
rect 14019 7958 14187 7960
rect 13742 7933 14187 7958
rect 13743 7932 14187 7933
rect 12102 7926 12546 7927
rect 12102 7901 12547 7926
rect 12102 7899 12270 7901
rect 12466 7900 12547 7901
rect 12716 7900 12765 7926
rect 12901 7900 12950 7927
rect 12102 7721 12129 7899
rect 12169 7861 12233 7873
rect 12509 7869 12546 7900
rect 12727 7869 12764 7900
rect 12909 7875 12950 7900
rect 13341 7899 13388 7932
rect 13744 7899 13784 7932
rect 14019 7931 14187 7932
rect 14650 7936 14690 8160
rect 14816 8159 14984 8160
rect 15587 8294 16031 8308
rect 15587 8292 15755 8294
rect 15587 8114 15614 8292
rect 15654 8254 15718 8266
rect 15994 8262 16031 8294
rect 16057 8293 16248 8315
rect 16483 8311 16592 8331
rect 16612 8311 16621 8331
rect 16483 8304 16621 8311
rect 16679 8331 16827 8340
rect 16679 8311 16688 8331
rect 16708 8311 16798 8331
rect 16818 8311 16827 8331
rect 16483 8302 16579 8304
rect 16679 8301 16827 8311
rect 16886 8331 16923 8341
rect 16886 8311 16894 8331
rect 16914 8311 16923 8331
rect 16735 8300 16771 8301
rect 16212 8291 16248 8293
rect 16212 8262 16249 8291
rect 15654 8253 15689 8254
rect 15631 8248 15689 8253
rect 15631 8228 15634 8248
rect 15654 8234 15689 8248
rect 15709 8234 15718 8254
rect 15654 8226 15718 8234
rect 15680 8225 15718 8226
rect 15681 8224 15718 8225
rect 15784 8258 15820 8259
rect 15892 8258 15928 8259
rect 15784 8252 15928 8258
rect 15784 8250 15845 8252
rect 15784 8230 15792 8250
rect 15812 8235 15845 8250
rect 15864 8250 15928 8252
rect 15864 8235 15900 8250
rect 15812 8230 15900 8235
rect 15920 8230 15928 8250
rect 15784 8224 15928 8230
rect 15994 8254 16032 8262
rect 16110 8258 16146 8259
rect 15994 8234 16003 8254
rect 16023 8234 16032 8254
rect 15994 8225 16032 8234
rect 16061 8250 16146 8258
rect 16061 8230 16118 8250
rect 16138 8230 16146 8250
rect 15994 8224 16031 8225
rect 16061 8224 16146 8230
rect 16212 8254 16250 8262
rect 16212 8234 16221 8254
rect 16241 8234 16250 8254
rect 16886 8244 16923 8311
rect 16958 8340 16989 8391
rect 17271 8379 17289 8397
rect 17307 8379 17323 8397
rect 17789 8404 17827 8413
rect 17008 8340 17045 8341
rect 16958 8331 17045 8340
rect 16958 8311 17016 8331
rect 17036 8311 17045 8331
rect 16958 8301 17045 8311
rect 17104 8331 17141 8341
rect 17104 8311 17112 8331
rect 17132 8311 17141 8331
rect 16958 8300 16989 8301
rect 16583 8241 16620 8242
rect 16886 8241 16925 8244
rect 16582 8240 16925 8241
rect 17104 8240 17141 8311
rect 16212 8225 16250 8234
rect 16507 8235 16925 8240
rect 16212 8224 16249 8225
rect 15673 8196 15763 8202
rect 15673 8176 15689 8196
rect 15709 8194 15763 8196
rect 15709 8176 15734 8194
rect 15673 8174 15734 8176
rect 15754 8174 15763 8194
rect 15673 8168 15763 8174
rect 15686 8114 15723 8115
rect 15782 8114 15819 8115
rect 15838 8114 15874 8224
rect 16061 8203 16092 8224
rect 16507 8215 16510 8235
rect 16530 8215 16925 8235
rect 16954 8216 17141 8240
rect 16057 8202 16092 8203
rect 15935 8192 16092 8202
rect 15935 8172 15952 8192
rect 15972 8172 16092 8192
rect 15935 8165 16092 8172
rect 16159 8195 16308 8203
rect 16159 8175 16170 8195
rect 16190 8175 16229 8195
rect 16249 8175 16308 8195
rect 16159 8168 16308 8175
rect 16886 8190 16925 8215
rect 17271 8190 17323 8379
rect 17617 8386 17657 8396
rect 17617 8368 17627 8386
rect 17645 8368 17657 8386
rect 17789 8384 17798 8404
rect 17818 8384 17827 8404
rect 17789 8376 17827 8384
rect 17893 8408 17978 8414
rect 18008 8413 18045 8414
rect 17893 8388 17901 8408
rect 17921 8388 17978 8408
rect 17893 8380 17978 8388
rect 18007 8404 18045 8413
rect 18007 8384 18016 8404
rect 18036 8384 18045 8404
rect 17893 8379 17929 8380
rect 18007 8376 18045 8384
rect 18111 8408 18255 8414
rect 18111 8388 18119 8408
rect 18139 8388 18172 8408
rect 18192 8388 18227 8408
rect 18247 8388 18255 8408
rect 18111 8380 18255 8388
rect 18111 8379 18147 8380
rect 18219 8379 18255 8380
rect 18321 8413 18358 8414
rect 18321 8412 18359 8413
rect 18321 8404 18385 8412
rect 18321 8384 18330 8404
rect 18350 8390 18385 8404
rect 18405 8390 18408 8410
rect 18350 8385 18408 8390
rect 18350 8384 18385 8385
rect 17617 8312 17657 8368
rect 17790 8347 17827 8376
rect 17791 8345 17827 8347
rect 17791 8323 17982 8345
rect 18008 8344 18045 8376
rect 18321 8372 18385 8384
rect 18425 8346 18452 8524
rect 18284 8344 18452 8346
rect 18008 8334 18452 8344
rect 18593 8440 18780 8464
rect 18811 8445 19204 8465
rect 19224 8445 19227 8465
rect 18811 8440 19227 8445
rect 18593 8369 18630 8440
rect 18811 8439 19152 8440
rect 18745 8379 18776 8380
rect 18593 8349 18602 8369
rect 18622 8349 18630 8369
rect 18593 8339 18630 8349
rect 18689 8369 18776 8379
rect 18689 8349 18698 8369
rect 18718 8349 18776 8369
rect 18689 8340 18776 8349
rect 18689 8339 18726 8340
rect 17614 8307 17657 8312
rect 18005 8318 18452 8334
rect 18005 8312 18033 8318
rect 18284 8317 18452 8318
rect 17614 8304 17764 8307
rect 18005 8304 18032 8312
rect 17614 8302 18032 8304
rect 17614 8284 17623 8302
rect 17641 8284 18032 8302
rect 18745 8289 18776 8340
rect 18811 8369 18848 8439
rect 19114 8438 19151 8439
rect 18963 8379 18999 8380
rect 18811 8349 18820 8369
rect 18840 8349 18848 8369
rect 18811 8339 18848 8349
rect 18907 8369 19055 8379
rect 19155 8376 19251 8378
rect 18907 8349 18916 8369
rect 18936 8349 19026 8369
rect 19046 8349 19055 8369
rect 18907 8340 19055 8349
rect 19113 8369 19251 8376
rect 19113 8349 19122 8369
rect 19142 8349 19251 8369
rect 19113 8340 19251 8349
rect 18907 8339 18944 8340
rect 18637 8286 18678 8287
rect 17614 8281 18032 8284
rect 17614 8275 17657 8281
rect 17617 8272 17657 8275
rect 18529 8279 18678 8286
rect 18014 8263 18054 8264
rect 17725 8246 18054 8263
rect 18529 8259 18588 8279
rect 18608 8259 18647 8279
rect 18667 8259 18678 8279
rect 18529 8251 18678 8259
rect 18745 8282 18902 8289
rect 18745 8262 18865 8282
rect 18885 8262 18902 8282
rect 18745 8252 18902 8262
rect 18745 8251 18780 8252
rect 17609 8203 17652 8214
rect 16886 8172 17325 8190
rect 16159 8167 16200 8168
rect 15893 8114 15930 8115
rect 15586 8105 15724 8114
rect 15586 8085 15695 8105
rect 15715 8085 15724 8105
rect 15586 8078 15724 8085
rect 15782 8105 15930 8114
rect 15782 8085 15791 8105
rect 15811 8085 15901 8105
rect 15921 8085 15930 8105
rect 15586 8076 15682 8078
rect 15782 8075 15930 8085
rect 15989 8105 16026 8115
rect 15989 8085 15997 8105
rect 16017 8085 16026 8105
rect 15838 8074 15874 8075
rect 15686 8015 15723 8016
rect 15989 8015 16026 8085
rect 16061 8114 16092 8165
rect 16886 8154 17286 8172
rect 17304 8154 17325 8172
rect 16886 8148 17325 8154
rect 16892 8144 17325 8148
rect 17609 8185 17621 8203
rect 17639 8185 17652 8203
rect 17609 8159 17652 8185
rect 17725 8159 17752 8246
rect 18014 8237 18054 8246
rect 17271 8142 17323 8144
rect 17609 8138 17752 8159
rect 17796 8211 17830 8227
rect 18014 8217 18407 8237
rect 18427 8217 18430 8237
rect 18745 8230 18776 8251
rect 18963 8230 18999 8340
rect 19018 8339 19055 8340
rect 19114 8339 19151 8340
rect 19074 8280 19164 8286
rect 19074 8260 19083 8280
rect 19103 8278 19164 8280
rect 19103 8260 19128 8278
rect 19074 8258 19128 8260
rect 19148 8258 19164 8278
rect 19074 8252 19164 8258
rect 18588 8229 18625 8230
rect 18014 8212 18430 8217
rect 18587 8220 18625 8229
rect 18014 8211 18355 8212
rect 17796 8141 17833 8211
rect 17948 8151 17979 8152
rect 17609 8136 17746 8138
rect 16111 8114 16148 8115
rect 16061 8105 16148 8114
rect 16061 8085 16119 8105
rect 16139 8085 16148 8105
rect 16061 8075 16148 8085
rect 16207 8105 16244 8115
rect 16207 8085 16215 8105
rect 16235 8085 16244 8105
rect 17609 8094 17652 8136
rect 17796 8121 17805 8141
rect 17825 8121 17833 8141
rect 17796 8111 17833 8121
rect 17892 8141 17979 8151
rect 17892 8121 17901 8141
rect 17921 8121 17979 8141
rect 17892 8112 17979 8121
rect 17892 8111 17929 8112
rect 16061 8074 16092 8075
rect 15685 8014 16026 8015
rect 16207 8014 16244 8085
rect 17607 8084 17652 8094
rect 17274 8077 17311 8082
rect 17265 8073 17312 8077
rect 17265 8055 17284 8073
rect 17302 8055 17312 8073
rect 17607 8066 17616 8084
rect 17634 8066 17652 8084
rect 17607 8060 17652 8066
rect 17948 8061 17979 8112
rect 18014 8141 18051 8211
rect 18317 8210 18354 8211
rect 18587 8200 18596 8220
rect 18616 8200 18625 8220
rect 18587 8192 18625 8200
rect 18691 8224 18776 8230
rect 18806 8229 18843 8230
rect 18691 8204 18699 8224
rect 18719 8204 18776 8224
rect 18691 8196 18776 8204
rect 18805 8220 18843 8229
rect 18805 8200 18814 8220
rect 18834 8200 18843 8220
rect 18691 8195 18727 8196
rect 18805 8192 18843 8200
rect 18909 8224 19053 8230
rect 18909 8204 18917 8224
rect 18937 8205 18969 8224
rect 18990 8205 19025 8224
rect 18937 8204 19025 8205
rect 19045 8204 19053 8224
rect 18909 8196 19053 8204
rect 18909 8195 18945 8196
rect 19017 8195 19053 8196
rect 19119 8229 19156 8230
rect 19119 8228 19157 8229
rect 19119 8220 19183 8228
rect 19119 8200 19128 8220
rect 19148 8206 19183 8220
rect 19203 8206 19206 8226
rect 19148 8201 19206 8206
rect 19148 8200 19183 8201
rect 18588 8163 18625 8192
rect 18589 8161 18625 8163
rect 18166 8151 18202 8152
rect 18014 8121 18023 8141
rect 18043 8121 18051 8141
rect 18014 8111 18051 8121
rect 18110 8141 18258 8151
rect 18358 8148 18454 8150
rect 18110 8121 18119 8141
rect 18139 8121 18229 8141
rect 18249 8121 18258 8141
rect 18110 8112 18258 8121
rect 18316 8141 18454 8148
rect 18316 8121 18325 8141
rect 18345 8121 18454 8141
rect 18589 8139 18780 8161
rect 18806 8160 18843 8192
rect 19119 8188 19183 8200
rect 19223 8162 19250 8340
rect 19855 8339 19888 8672
rect 19952 8704 20120 8705
rect 20246 8704 20286 8928
rect 20749 8932 20917 8933
rect 21150 8932 21195 8953
rect 20749 8906 21195 8932
rect 20749 8904 20917 8906
rect 21113 8905 21195 8906
rect 21330 8905 21411 8931
rect 21555 8918 22036 8953
rect 24610 8941 24618 8963
rect 24642 8941 24650 8963
rect 20749 8726 20776 8904
rect 20816 8866 20880 8878
rect 21156 8874 21193 8905
rect 21374 8874 21411 8905
rect 21558 8899 21597 8918
rect 21556 8880 21597 8899
rect 20816 8865 20851 8866
rect 20793 8860 20851 8865
rect 20793 8840 20796 8860
rect 20816 8846 20851 8860
rect 20871 8846 20880 8866
rect 20816 8838 20880 8846
rect 20842 8837 20880 8838
rect 20843 8836 20880 8837
rect 20946 8870 20982 8871
rect 21054 8870 21090 8871
rect 20946 8862 21090 8870
rect 20946 8842 20954 8862
rect 20974 8858 21062 8862
rect 20974 8842 21018 8858
rect 20946 8838 21018 8842
rect 21038 8842 21062 8858
rect 21082 8842 21090 8862
rect 21038 8838 21090 8842
rect 20946 8836 21090 8838
rect 21156 8866 21194 8874
rect 21272 8870 21308 8871
rect 21156 8846 21165 8866
rect 21185 8846 21194 8866
rect 21156 8837 21194 8846
rect 21223 8862 21308 8870
rect 21223 8842 21280 8862
rect 21300 8842 21308 8862
rect 21156 8836 21193 8837
rect 21223 8836 21308 8842
rect 21374 8866 21412 8874
rect 21374 8846 21383 8866
rect 21403 8846 21412 8866
rect 21374 8837 21412 8846
rect 21556 8871 21598 8880
rect 21556 8853 21570 8871
rect 21588 8853 21598 8871
rect 21556 8845 21598 8853
rect 21561 8843 21598 8845
rect 21374 8836 21411 8837
rect 20835 8808 20925 8814
rect 20835 8788 20851 8808
rect 20871 8806 20925 8808
rect 20871 8788 20896 8806
rect 20835 8786 20896 8788
rect 20916 8786 20925 8806
rect 20835 8780 20925 8786
rect 20848 8726 20885 8727
rect 20944 8726 20981 8727
rect 21000 8726 21036 8836
rect 21223 8815 21254 8836
rect 21988 8822 22035 8918
rect 21219 8814 21254 8815
rect 21097 8804 21254 8814
rect 21097 8784 21114 8804
rect 21134 8784 21254 8804
rect 21097 8777 21254 8784
rect 21321 8807 21470 8815
rect 21321 8787 21332 8807
rect 21352 8787 21391 8807
rect 21411 8787 21470 8807
rect 21988 8804 21998 8822
rect 22016 8804 22035 8822
rect 21988 8800 22035 8804
rect 21989 8795 22026 8800
rect 21321 8780 21470 8787
rect 21321 8779 21362 8780
rect 21558 8778 21595 8781
rect 21055 8726 21092 8727
rect 20748 8717 20886 8726
rect 19952 8678 20396 8704
rect 19952 8676 20120 8678
rect 19952 8498 19979 8676
rect 20019 8638 20083 8650
rect 20359 8646 20396 8678
rect 20422 8677 20613 8699
rect 20748 8697 20857 8717
rect 20877 8697 20886 8717
rect 20748 8690 20886 8697
rect 20944 8717 21092 8726
rect 20944 8697 20953 8717
rect 20973 8697 21063 8717
rect 21083 8697 21092 8717
rect 20748 8688 20844 8690
rect 20944 8687 21092 8697
rect 21151 8717 21188 8727
rect 21151 8697 21159 8717
rect 21179 8697 21188 8717
rect 21000 8686 21036 8687
rect 20577 8675 20613 8677
rect 20577 8646 20614 8675
rect 20019 8637 20054 8638
rect 19996 8632 20054 8637
rect 19996 8612 19999 8632
rect 20019 8618 20054 8632
rect 20074 8618 20083 8638
rect 20019 8612 20083 8618
rect 19996 8610 20083 8612
rect 19996 8606 20023 8610
rect 20045 8609 20083 8610
rect 20046 8608 20083 8609
rect 20149 8642 20185 8643
rect 20257 8642 20293 8643
rect 20149 8635 20293 8642
rect 20149 8634 20211 8635
rect 20149 8614 20157 8634
rect 20177 8617 20211 8634
rect 20230 8634 20293 8635
rect 20230 8617 20265 8634
rect 20177 8614 20265 8617
rect 20285 8614 20293 8634
rect 20149 8608 20293 8614
rect 20359 8638 20397 8646
rect 20475 8642 20511 8643
rect 20359 8618 20368 8638
rect 20388 8618 20397 8638
rect 20359 8609 20397 8618
rect 20426 8634 20511 8642
rect 20426 8614 20483 8634
rect 20503 8614 20511 8634
rect 20359 8608 20396 8609
rect 20426 8608 20511 8614
rect 20577 8638 20615 8646
rect 20577 8618 20586 8638
rect 20606 8618 20615 8638
rect 20848 8627 20885 8628
rect 21151 8627 21188 8697
rect 21223 8726 21254 8777
rect 21550 8772 21595 8778
rect 21550 8754 21568 8772
rect 21586 8754 21595 8772
rect 21550 8744 21595 8754
rect 21273 8726 21310 8727
rect 21223 8717 21310 8726
rect 21223 8697 21281 8717
rect 21301 8697 21310 8717
rect 21223 8687 21310 8697
rect 21369 8717 21406 8727
rect 21369 8697 21377 8717
rect 21397 8697 21406 8717
rect 21550 8702 21593 8744
rect 21977 8733 22029 8735
rect 21456 8700 21593 8702
rect 21223 8686 21254 8687
rect 21369 8627 21406 8697
rect 20847 8626 21188 8627
rect 20577 8609 20615 8618
rect 20772 8621 21188 8626
rect 20577 8608 20614 8609
rect 20038 8580 20128 8586
rect 20038 8560 20054 8580
rect 20074 8578 20128 8580
rect 20074 8560 20099 8578
rect 20038 8558 20099 8560
rect 20119 8558 20128 8578
rect 20038 8552 20128 8558
rect 20051 8498 20088 8499
rect 20147 8498 20184 8499
rect 20203 8498 20239 8608
rect 20426 8587 20457 8608
rect 20772 8601 20775 8621
rect 20795 8601 21188 8621
rect 21372 8611 21406 8627
rect 21450 8679 21593 8700
rect 21975 8729 22408 8733
rect 21975 8723 22414 8729
rect 21975 8705 21996 8723
rect 22014 8705 22414 8723
rect 21975 8687 22414 8705
rect 21148 8592 21188 8601
rect 21450 8592 21477 8679
rect 21550 8653 21593 8679
rect 21550 8635 21563 8653
rect 21581 8635 21593 8653
rect 21550 8624 21593 8635
rect 20422 8586 20457 8587
rect 20300 8576 20457 8586
rect 20300 8556 20317 8576
rect 20337 8556 20457 8576
rect 20300 8549 20457 8556
rect 20524 8579 20670 8587
rect 20524 8559 20535 8579
rect 20555 8559 20594 8579
rect 20614 8559 20670 8579
rect 21148 8575 21477 8592
rect 21148 8574 21188 8575
rect 20524 8552 20670 8559
rect 21545 8563 21585 8566
rect 21545 8557 21588 8563
rect 21170 8554 21588 8557
rect 20524 8551 20565 8552
rect 20258 8498 20295 8499
rect 19951 8489 20089 8498
rect 19951 8469 20060 8489
rect 20080 8469 20089 8489
rect 19951 8462 20089 8469
rect 20147 8489 20295 8498
rect 20147 8469 20156 8489
rect 20176 8469 20266 8489
rect 20286 8469 20295 8489
rect 19951 8460 20047 8462
rect 20147 8459 20295 8469
rect 20354 8489 20391 8499
rect 20354 8469 20362 8489
rect 20382 8469 20391 8489
rect 20203 8458 20239 8459
rect 20051 8399 20088 8400
rect 20354 8399 20391 8469
rect 20426 8498 20457 8549
rect 21170 8536 21561 8554
rect 21579 8536 21588 8554
rect 21170 8534 21588 8536
rect 21170 8526 21197 8534
rect 21438 8531 21588 8534
rect 20750 8520 20918 8521
rect 21169 8520 21197 8526
rect 20750 8504 21197 8520
rect 21545 8526 21588 8531
rect 20476 8498 20513 8499
rect 20426 8489 20513 8498
rect 20426 8469 20484 8489
rect 20504 8469 20513 8489
rect 20426 8459 20513 8469
rect 20572 8489 20609 8499
rect 20572 8469 20580 8489
rect 20600 8469 20609 8489
rect 20426 8458 20457 8459
rect 20050 8398 20391 8399
rect 20572 8398 20609 8469
rect 19975 8393 20391 8398
rect 19975 8373 19978 8393
rect 19998 8373 20391 8393
rect 20422 8374 20609 8398
rect 20750 8494 21194 8504
rect 20750 8492 20918 8494
rect 19850 8294 19892 8339
rect 20750 8314 20777 8492
rect 20817 8454 20881 8466
rect 21157 8462 21194 8494
rect 21220 8493 21411 8515
rect 21375 8491 21411 8493
rect 21375 8462 21412 8491
rect 21545 8470 21585 8526
rect 20817 8453 20852 8454
rect 20794 8448 20852 8453
rect 20794 8428 20797 8448
rect 20817 8434 20852 8448
rect 20872 8434 20881 8454
rect 20817 8426 20881 8434
rect 20843 8425 20881 8426
rect 20844 8424 20881 8425
rect 20947 8458 20983 8459
rect 21055 8458 21091 8459
rect 20947 8450 21091 8458
rect 20947 8430 20955 8450
rect 20975 8430 21010 8450
rect 21030 8430 21063 8450
rect 21083 8430 21091 8450
rect 20947 8424 21091 8430
rect 21157 8454 21195 8462
rect 21273 8458 21309 8459
rect 21157 8434 21166 8454
rect 21186 8434 21195 8454
rect 21157 8425 21195 8434
rect 21224 8450 21309 8458
rect 21224 8430 21281 8450
rect 21301 8430 21309 8450
rect 21157 8424 21194 8425
rect 21224 8424 21309 8430
rect 21375 8454 21413 8462
rect 21375 8434 21384 8454
rect 21404 8434 21413 8454
rect 21545 8452 21557 8470
rect 21575 8452 21585 8470
rect 21977 8498 22029 8687
rect 22375 8662 22414 8687
rect 24215 8712 24252 8718
rect 24215 8693 24223 8712
rect 24244 8693 24252 8712
rect 24215 8685 24252 8693
rect 22159 8637 22346 8661
rect 22375 8642 22770 8662
rect 22790 8642 22793 8662
rect 22375 8637 22793 8642
rect 22159 8566 22196 8637
rect 22375 8636 22718 8637
rect 22375 8633 22414 8636
rect 22680 8635 22717 8636
rect 22311 8576 22342 8577
rect 22159 8546 22168 8566
rect 22188 8546 22196 8566
rect 22159 8536 22196 8546
rect 22255 8566 22342 8576
rect 22255 8546 22264 8566
rect 22284 8546 22342 8566
rect 22255 8537 22342 8546
rect 22255 8536 22292 8537
rect 21977 8480 21993 8498
rect 22011 8480 22029 8498
rect 22311 8486 22342 8537
rect 22377 8566 22414 8633
rect 22529 8576 22565 8577
rect 22377 8546 22386 8566
rect 22406 8546 22414 8566
rect 22377 8536 22414 8546
rect 22473 8566 22621 8576
rect 22721 8573 22817 8575
rect 22473 8546 22482 8566
rect 22502 8546 22592 8566
rect 22612 8546 22621 8566
rect 22473 8537 22621 8546
rect 22679 8566 22817 8573
rect 22679 8546 22688 8566
rect 22708 8546 22817 8566
rect 22679 8537 22817 8546
rect 22473 8536 22510 8537
rect 22203 8483 22244 8484
rect 21977 8462 22029 8480
rect 22095 8476 22244 8483
rect 21545 8442 21585 8452
rect 22095 8456 22154 8476
rect 22174 8456 22213 8476
rect 22233 8456 22244 8476
rect 22095 8448 22244 8456
rect 22311 8479 22468 8486
rect 22311 8459 22431 8479
rect 22451 8459 22468 8479
rect 22311 8449 22468 8459
rect 22311 8448 22346 8449
rect 21375 8425 21413 8434
rect 22311 8427 22342 8448
rect 22529 8427 22565 8537
rect 22584 8536 22621 8537
rect 22680 8536 22717 8537
rect 22640 8477 22730 8483
rect 22640 8457 22649 8477
rect 22669 8475 22730 8477
rect 22669 8457 22694 8475
rect 22640 8455 22694 8457
rect 22714 8455 22730 8475
rect 22640 8449 22730 8455
rect 22154 8426 22191 8427
rect 21375 8424 21412 8425
rect 20836 8396 20926 8402
rect 20836 8376 20852 8396
rect 20872 8394 20926 8396
rect 20872 8376 20897 8394
rect 20836 8374 20897 8376
rect 20917 8374 20926 8394
rect 20836 8368 20926 8374
rect 20849 8314 20886 8315
rect 20945 8314 20982 8315
rect 21001 8314 21037 8424
rect 21224 8403 21255 8424
rect 22153 8417 22191 8426
rect 21220 8402 21255 8403
rect 21098 8392 21255 8402
rect 21098 8372 21115 8392
rect 21135 8372 21255 8392
rect 21098 8365 21255 8372
rect 21322 8395 21471 8403
rect 21322 8375 21333 8395
rect 21353 8375 21392 8395
rect 21412 8375 21471 8395
rect 21981 8399 22021 8409
rect 21322 8368 21471 8375
rect 21537 8371 21589 8389
rect 21322 8367 21363 8368
rect 21056 8314 21093 8315
rect 20749 8305 20887 8314
rect 20221 8294 20254 8296
rect 19850 8282 20297 8294
rect 19082 8160 19250 8162
rect 18806 8134 19250 8160
rect 18316 8112 18454 8121
rect 18110 8111 18147 8112
rect 17607 8057 17644 8060
rect 17840 8058 17881 8059
rect 15610 8009 16026 8014
rect 15610 7989 15613 8009
rect 15633 7989 16026 8009
rect 16057 7990 16244 8014
rect 16869 8012 16909 8017
rect 17265 8012 17312 8055
rect 17732 8051 17881 8058
rect 17732 8031 17791 8051
rect 17811 8031 17850 8051
rect 17870 8031 17881 8051
rect 17732 8023 17881 8031
rect 17948 8054 18105 8061
rect 17948 8034 18068 8054
rect 18088 8034 18105 8054
rect 17948 8024 18105 8034
rect 17948 8023 17983 8024
rect 16869 7973 17312 8012
rect 17948 8002 17979 8023
rect 18166 8002 18202 8112
rect 18221 8111 18258 8112
rect 18317 8111 18354 8112
rect 18277 8052 18367 8058
rect 18277 8032 18286 8052
rect 18306 8050 18367 8052
rect 18306 8032 18331 8050
rect 18277 8030 18331 8032
rect 18351 8030 18367 8050
rect 18277 8024 18367 8030
rect 17791 8001 17828 8002
rect 14650 7914 14658 7936
rect 14682 7914 14690 7936
rect 14650 7906 14690 7914
rect 15963 7958 16003 7966
rect 15963 7936 15971 7958
rect 15995 7936 16003 7958
rect 12169 7860 12204 7861
rect 12146 7855 12204 7860
rect 12146 7835 12149 7855
rect 12169 7841 12204 7855
rect 12224 7841 12233 7861
rect 12169 7833 12233 7841
rect 12195 7832 12233 7833
rect 12196 7831 12233 7832
rect 12299 7865 12335 7866
rect 12407 7865 12443 7866
rect 12299 7857 12443 7865
rect 12299 7837 12307 7857
rect 12327 7853 12415 7857
rect 12327 7837 12371 7853
rect 12299 7833 12371 7837
rect 12391 7837 12415 7853
rect 12435 7837 12443 7857
rect 12391 7833 12443 7837
rect 12299 7831 12443 7833
rect 12509 7861 12547 7869
rect 12625 7865 12661 7866
rect 12509 7841 12518 7861
rect 12538 7841 12547 7861
rect 12509 7832 12547 7841
rect 12576 7857 12661 7865
rect 12576 7837 12633 7857
rect 12653 7837 12661 7857
rect 12509 7831 12546 7832
rect 12576 7831 12661 7837
rect 12727 7861 12765 7869
rect 12727 7841 12736 7861
rect 12756 7841 12765 7861
rect 12727 7832 12765 7841
rect 12909 7866 12951 7875
rect 12909 7848 12923 7866
rect 12941 7848 12951 7866
rect 12909 7840 12951 7848
rect 12914 7838 12951 7840
rect 13341 7860 13784 7899
rect 12727 7831 12764 7832
rect 12188 7803 12278 7809
rect 12188 7783 12204 7803
rect 12224 7801 12278 7803
rect 12224 7783 12249 7801
rect 12188 7781 12249 7783
rect 12269 7781 12278 7801
rect 12188 7775 12278 7781
rect 12201 7721 12238 7722
rect 12297 7721 12334 7722
rect 12353 7721 12389 7831
rect 12576 7810 12607 7831
rect 13341 7817 13388 7860
rect 13744 7855 13784 7860
rect 14409 7858 14596 7882
rect 14627 7863 15020 7883
rect 15040 7863 15043 7883
rect 14627 7858 15043 7863
rect 12572 7809 12607 7810
rect 12450 7799 12607 7809
rect 12450 7779 12467 7799
rect 12487 7779 12607 7799
rect 12450 7772 12607 7779
rect 12674 7802 12823 7810
rect 12674 7782 12685 7802
rect 12705 7782 12744 7802
rect 12764 7782 12823 7802
rect 13341 7799 13351 7817
rect 13369 7799 13388 7817
rect 13341 7795 13388 7799
rect 13342 7790 13379 7795
rect 12674 7775 12823 7782
rect 14409 7787 14446 7858
rect 14627 7857 14968 7858
rect 14561 7797 14592 7798
rect 12674 7774 12715 7775
rect 12911 7773 12948 7776
rect 12408 7721 12445 7722
rect 12101 7712 12239 7721
rect 11305 7673 11749 7699
rect 11305 7671 11473 7673
rect 10258 7539 10705 7551
rect 10301 7537 10334 7539
rect 9668 7519 9806 7528
rect 9462 7518 9499 7519
rect 9192 7465 9233 7466
rect 8966 7444 9018 7462
rect 9084 7458 9233 7465
rect 8521 7425 8561 7435
rect 9084 7438 9143 7458
rect 9163 7438 9202 7458
rect 9222 7438 9233 7458
rect 9084 7430 9233 7438
rect 9300 7461 9457 7468
rect 9300 7441 9420 7461
rect 9440 7441 9457 7461
rect 9300 7431 9457 7441
rect 9300 7430 9335 7431
rect 8351 7408 8389 7417
rect 9300 7409 9331 7430
rect 9518 7409 9554 7519
rect 9573 7518 9610 7519
rect 9669 7518 9706 7519
rect 9629 7459 9719 7465
rect 9629 7439 9638 7459
rect 9658 7457 9719 7459
rect 9658 7439 9683 7457
rect 9629 7437 9683 7439
rect 9703 7437 9719 7457
rect 9629 7431 9719 7437
rect 9143 7408 9180 7409
rect 8351 7407 8388 7408
rect 7812 7379 7902 7385
rect 7812 7359 7828 7379
rect 7848 7377 7902 7379
rect 7848 7359 7873 7377
rect 7812 7357 7873 7359
rect 7893 7357 7902 7377
rect 7812 7351 7902 7357
rect 7825 7297 7862 7298
rect 7921 7297 7958 7298
rect 7977 7297 8013 7407
rect 8200 7386 8231 7407
rect 9142 7399 9180 7408
rect 8196 7385 8231 7386
rect 8074 7375 8231 7385
rect 8074 7355 8091 7375
rect 8111 7355 8231 7375
rect 8074 7348 8231 7355
rect 8298 7378 8447 7386
rect 8298 7358 8309 7378
rect 8329 7358 8368 7378
rect 8388 7358 8447 7378
rect 8970 7381 9010 7391
rect 8298 7351 8447 7358
rect 8513 7354 8565 7372
rect 8298 7350 8339 7351
rect 8032 7297 8069 7298
rect 7725 7288 7863 7297
rect 6792 7280 6829 7281
rect 6763 7279 6931 7280
rect 7057 7279 7097 7281
rect 6588 7270 6627 7276
rect 6588 7248 6596 7270
rect 6620 7248 6627 7270
rect 6290 7141 6327 7149
rect 6290 7122 6298 7141
rect 6319 7122 6327 7141
rect 6290 7116 6327 7122
rect 5892 6871 5900 6893
rect 5924 6871 5932 6893
rect 5892 6863 5932 6871
rect 3408 6817 3443 6818
rect 3385 6812 3443 6817
rect 3385 6792 3388 6812
rect 3408 6798 3443 6812
rect 3463 6798 3472 6818
rect 3408 6790 3472 6798
rect 3434 6789 3472 6790
rect 3435 6788 3472 6789
rect 3538 6822 3574 6823
rect 3646 6822 3682 6823
rect 3538 6814 3682 6822
rect 3538 6794 3546 6814
rect 3566 6810 3654 6814
rect 3566 6794 3610 6810
rect 3538 6790 3610 6794
rect 3630 6794 3654 6810
rect 3674 6794 3682 6814
rect 3630 6790 3682 6794
rect 3538 6788 3682 6790
rect 3748 6818 3786 6826
rect 3864 6822 3900 6823
rect 3748 6798 3757 6818
rect 3777 6798 3786 6818
rect 3748 6789 3786 6798
rect 3815 6814 3900 6822
rect 3815 6794 3872 6814
rect 3892 6794 3900 6814
rect 3748 6788 3785 6789
rect 3815 6788 3900 6794
rect 3966 6818 4004 6826
rect 3966 6798 3975 6818
rect 3995 6798 4004 6818
rect 3966 6789 4004 6798
rect 4148 6823 4191 6850
rect 4148 6805 4162 6823
rect 4180 6805 4191 6823
rect 4148 6797 4191 6805
rect 4153 6795 4191 6797
rect 4580 6825 5025 6855
rect 6063 6838 6128 6839
rect 4580 6822 5003 6825
rect 3966 6788 4003 6789
rect 3427 6760 3517 6766
rect 3427 6740 3443 6760
rect 3463 6758 3517 6760
rect 3463 6740 3488 6758
rect 3427 6738 3488 6740
rect 3508 6738 3517 6758
rect 3427 6732 3517 6738
rect 3440 6678 3477 6679
rect 3536 6678 3573 6679
rect 3592 6678 3628 6788
rect 3815 6767 3846 6788
rect 4580 6774 4627 6822
rect 3811 6766 3846 6767
rect 3689 6756 3846 6766
rect 3689 6736 3706 6756
rect 3726 6736 3846 6756
rect 3689 6729 3846 6736
rect 3913 6759 4062 6767
rect 3913 6739 3924 6759
rect 3944 6739 3983 6759
rect 4003 6739 4062 6759
rect 4580 6756 4590 6774
rect 4608 6756 4627 6774
rect 4580 6752 4627 6756
rect 5714 6813 5901 6837
rect 5932 6818 6325 6838
rect 6345 6818 6348 6838
rect 5932 6813 6348 6818
rect 4581 6747 4618 6752
rect 3913 6732 4062 6739
rect 5714 6742 5751 6813
rect 5932 6812 6273 6813
rect 5866 6752 5897 6753
rect 3913 6731 3954 6732
rect 4150 6730 4187 6733
rect 3647 6678 3684 6679
rect 3340 6669 3478 6678
rect 2544 6630 2988 6656
rect 2544 6628 2712 6630
rect 2544 6450 2571 6628
rect 2611 6590 2675 6602
rect 2951 6598 2988 6630
rect 3014 6629 3205 6651
rect 3340 6649 3449 6669
rect 3469 6649 3478 6669
rect 3340 6642 3478 6649
rect 3536 6669 3684 6678
rect 3536 6649 3545 6669
rect 3565 6649 3655 6669
rect 3675 6649 3684 6669
rect 3340 6640 3436 6642
rect 3536 6639 3684 6649
rect 3743 6669 3780 6679
rect 3743 6649 3751 6669
rect 3771 6649 3780 6669
rect 3592 6638 3628 6639
rect 3169 6627 3205 6629
rect 3169 6598 3206 6627
rect 2611 6589 2646 6590
rect 2588 6584 2646 6589
rect 2588 6564 2591 6584
rect 2611 6570 2646 6584
rect 2666 6570 2675 6590
rect 2611 6564 2675 6570
rect 2588 6562 2675 6564
rect 2588 6558 2615 6562
rect 2637 6561 2675 6562
rect 2638 6560 2675 6561
rect 2741 6594 2777 6595
rect 2849 6594 2885 6595
rect 2741 6587 2885 6594
rect 2741 6586 2803 6587
rect 2741 6566 2749 6586
rect 2769 6569 2803 6586
rect 2822 6586 2885 6587
rect 2822 6569 2857 6586
rect 2769 6566 2857 6569
rect 2877 6566 2885 6586
rect 2741 6560 2885 6566
rect 2951 6590 2989 6598
rect 3067 6594 3103 6595
rect 2951 6570 2960 6590
rect 2980 6570 2989 6590
rect 2951 6561 2989 6570
rect 3018 6586 3103 6594
rect 3018 6566 3075 6586
rect 3095 6566 3103 6586
rect 2951 6560 2988 6561
rect 3018 6560 3103 6566
rect 3169 6590 3207 6598
rect 3169 6570 3178 6590
rect 3198 6570 3207 6590
rect 3440 6579 3477 6580
rect 3743 6579 3780 6649
rect 3815 6678 3846 6729
rect 4142 6724 4187 6730
rect 4142 6706 4160 6724
rect 4178 6706 4187 6724
rect 5714 6722 5723 6742
rect 5743 6722 5751 6742
rect 5714 6712 5751 6722
rect 5810 6742 5897 6752
rect 5810 6722 5819 6742
rect 5839 6722 5897 6742
rect 5810 6713 5897 6722
rect 5810 6712 5847 6713
rect 4142 6696 4187 6706
rect 3865 6678 3902 6679
rect 3815 6669 3902 6678
rect 3815 6649 3873 6669
rect 3893 6649 3902 6669
rect 3815 6639 3902 6649
rect 3961 6669 3998 6679
rect 3961 6649 3969 6669
rect 3989 6649 3998 6669
rect 4142 6654 4185 6696
rect 4569 6685 4621 6687
rect 4048 6652 4185 6654
rect 3815 6638 3846 6639
rect 3961 6579 3998 6649
rect 3439 6578 3780 6579
rect 3169 6561 3207 6570
rect 3364 6573 3780 6578
rect 3169 6560 3206 6561
rect 2630 6532 2720 6538
rect 2630 6512 2646 6532
rect 2666 6530 2720 6532
rect 2666 6512 2691 6530
rect 2630 6510 2691 6512
rect 2711 6510 2720 6530
rect 2630 6504 2720 6510
rect 2643 6450 2680 6451
rect 2739 6450 2776 6451
rect 2795 6450 2831 6560
rect 3018 6539 3049 6560
rect 3364 6553 3367 6573
rect 3387 6553 3780 6573
rect 3964 6563 3998 6579
rect 4042 6631 4185 6652
rect 4567 6681 5000 6685
rect 4567 6675 5006 6681
rect 4567 6657 4588 6675
rect 4606 6657 5006 6675
rect 5866 6662 5897 6713
rect 5932 6742 5969 6812
rect 6235 6811 6272 6812
rect 6084 6752 6120 6753
rect 5932 6722 5941 6742
rect 5961 6722 5969 6742
rect 5932 6712 5969 6722
rect 6028 6742 6176 6752
rect 6276 6749 6372 6751
rect 6028 6722 6037 6742
rect 6057 6722 6147 6742
rect 6167 6722 6176 6742
rect 6028 6713 6176 6722
rect 6234 6742 6372 6749
rect 6234 6722 6243 6742
rect 6263 6722 6372 6742
rect 6234 6713 6372 6722
rect 6028 6712 6065 6713
rect 5758 6659 5799 6660
rect 4567 6639 5006 6657
rect 3740 6544 3780 6553
rect 4042 6544 4069 6631
rect 4142 6605 4185 6631
rect 4142 6587 4155 6605
rect 4173 6587 4185 6605
rect 4142 6576 4185 6587
rect 3014 6538 3049 6539
rect 2892 6528 3049 6538
rect 2892 6508 2909 6528
rect 2929 6508 3049 6528
rect 2892 6501 3049 6508
rect 3116 6531 3262 6539
rect 3116 6511 3127 6531
rect 3147 6511 3186 6531
rect 3206 6511 3262 6531
rect 3740 6527 4069 6544
rect 3740 6526 3780 6527
rect 3116 6504 3262 6511
rect 4137 6515 4177 6518
rect 4137 6509 4180 6515
rect 3762 6506 4180 6509
rect 3116 6503 3157 6504
rect 2850 6450 2887 6451
rect 2543 6441 2681 6450
rect 2543 6421 2652 6441
rect 2672 6421 2681 6441
rect 2543 6414 2681 6421
rect 2739 6441 2887 6450
rect 2739 6421 2748 6441
rect 2768 6421 2858 6441
rect 2878 6421 2887 6441
rect 2543 6412 2639 6414
rect 2739 6411 2887 6421
rect 2946 6441 2983 6451
rect 2946 6421 2954 6441
rect 2974 6421 2983 6441
rect 2795 6410 2831 6411
rect 2643 6351 2680 6352
rect 2946 6351 2983 6421
rect 3018 6450 3049 6501
rect 3762 6488 4153 6506
rect 4171 6488 4180 6506
rect 3762 6486 4180 6488
rect 3762 6478 3789 6486
rect 4030 6483 4180 6486
rect 3342 6472 3510 6473
rect 3761 6472 3789 6478
rect 3342 6456 3789 6472
rect 4137 6478 4180 6483
rect 3068 6450 3105 6451
rect 3018 6441 3105 6450
rect 3018 6421 3076 6441
rect 3096 6421 3105 6441
rect 3018 6411 3105 6421
rect 3164 6441 3201 6451
rect 3164 6421 3172 6441
rect 3192 6421 3201 6441
rect 3018 6410 3049 6411
rect 2642 6350 2983 6351
rect 3164 6350 3201 6421
rect 2567 6345 2983 6350
rect 2567 6325 2570 6345
rect 2590 6325 2983 6345
rect 3014 6326 3201 6350
rect 3342 6446 3786 6456
rect 3342 6444 3510 6446
rect 2442 6246 2484 6291
rect 3342 6266 3369 6444
rect 3409 6406 3473 6418
rect 3749 6414 3786 6446
rect 3812 6445 4003 6467
rect 3967 6443 4003 6445
rect 3967 6414 4004 6443
rect 4137 6422 4177 6478
rect 3409 6405 3444 6406
rect 3386 6400 3444 6405
rect 3386 6380 3389 6400
rect 3409 6386 3444 6400
rect 3464 6386 3473 6406
rect 3409 6378 3473 6386
rect 3435 6377 3473 6378
rect 3436 6376 3473 6377
rect 3539 6410 3575 6411
rect 3647 6410 3683 6411
rect 3539 6402 3683 6410
rect 3539 6382 3547 6402
rect 3567 6382 3602 6402
rect 3622 6382 3655 6402
rect 3675 6382 3683 6402
rect 3539 6376 3683 6382
rect 3749 6406 3787 6414
rect 3865 6410 3901 6411
rect 3749 6386 3758 6406
rect 3778 6386 3787 6406
rect 3749 6377 3787 6386
rect 3816 6402 3901 6410
rect 3816 6382 3873 6402
rect 3893 6382 3901 6402
rect 3749 6376 3786 6377
rect 3816 6376 3901 6382
rect 3967 6406 4005 6414
rect 3967 6386 3976 6406
rect 3996 6386 4005 6406
rect 4137 6404 4149 6422
rect 4167 6404 4177 6422
rect 4569 6450 4621 6639
rect 4967 6614 5006 6639
rect 5650 6652 5799 6659
rect 5650 6632 5709 6652
rect 5729 6632 5768 6652
rect 5788 6632 5799 6652
rect 5650 6624 5799 6632
rect 5866 6655 6023 6662
rect 5866 6635 5986 6655
rect 6006 6635 6023 6655
rect 5866 6625 6023 6635
rect 5866 6624 5901 6625
rect 4751 6589 4938 6613
rect 4967 6594 5362 6614
rect 5382 6594 5385 6614
rect 5866 6603 5897 6624
rect 6084 6603 6120 6713
rect 6139 6712 6176 6713
rect 6235 6712 6272 6713
rect 6195 6653 6285 6659
rect 6195 6633 6204 6653
rect 6224 6651 6285 6653
rect 6224 6633 6249 6651
rect 6195 6631 6249 6633
rect 6269 6631 6285 6651
rect 6195 6625 6285 6631
rect 5709 6602 5746 6603
rect 4967 6589 5385 6594
rect 5708 6593 5746 6602
rect 4751 6518 4788 6589
rect 4967 6588 5310 6589
rect 4967 6585 5006 6588
rect 5272 6587 5309 6588
rect 4903 6528 4934 6529
rect 4751 6498 4760 6518
rect 4780 6498 4788 6518
rect 4751 6488 4788 6498
rect 4847 6518 4934 6528
rect 4847 6498 4856 6518
rect 4876 6498 4934 6518
rect 4847 6489 4934 6498
rect 4847 6488 4884 6489
rect 4569 6432 4585 6450
rect 4603 6432 4621 6450
rect 4903 6438 4934 6489
rect 4969 6518 5006 6585
rect 5708 6573 5717 6593
rect 5737 6573 5746 6593
rect 5708 6565 5746 6573
rect 5812 6597 5897 6603
rect 5927 6602 5964 6603
rect 5812 6577 5820 6597
rect 5840 6577 5897 6597
rect 5812 6569 5897 6577
rect 5926 6593 5964 6602
rect 5926 6573 5935 6593
rect 5955 6573 5964 6593
rect 5812 6568 5848 6569
rect 5926 6565 5964 6573
rect 6030 6597 6174 6603
rect 6030 6577 6038 6597
rect 6058 6596 6146 6597
rect 6058 6578 6093 6596
rect 6111 6578 6146 6596
rect 6058 6577 6146 6578
rect 6166 6577 6174 6597
rect 6030 6569 6174 6577
rect 6030 6568 6066 6569
rect 6138 6568 6174 6569
rect 6240 6602 6277 6603
rect 6240 6601 6278 6602
rect 6240 6593 6304 6601
rect 6240 6573 6249 6593
rect 6269 6579 6304 6593
rect 6324 6579 6327 6599
rect 6269 6574 6327 6579
rect 6269 6573 6304 6574
rect 5709 6536 5746 6565
rect 5710 6534 5746 6536
rect 5121 6528 5157 6529
rect 4969 6498 4978 6518
rect 4998 6498 5006 6518
rect 4969 6488 5006 6498
rect 5065 6518 5213 6528
rect 5313 6525 5409 6527
rect 5065 6498 5074 6518
rect 5094 6498 5184 6518
rect 5204 6498 5213 6518
rect 5065 6489 5213 6498
rect 5271 6518 5409 6525
rect 5271 6498 5280 6518
rect 5300 6498 5409 6518
rect 5710 6512 5901 6534
rect 5927 6533 5964 6565
rect 6240 6561 6304 6573
rect 6344 6537 6371 6713
rect 6290 6535 6371 6537
rect 6203 6533 6371 6535
rect 5927 6507 6371 6533
rect 6037 6505 6077 6507
rect 6203 6506 6371 6507
rect 5271 6489 5409 6498
rect 6312 6504 6371 6506
rect 5065 6488 5102 6489
rect 4795 6435 4836 6436
rect 4569 6414 4621 6432
rect 4687 6428 4836 6435
rect 4137 6394 4177 6404
rect 4687 6408 4746 6428
rect 4766 6408 4805 6428
rect 4825 6408 4836 6428
rect 4687 6400 4836 6408
rect 4903 6431 5060 6438
rect 4903 6411 5023 6431
rect 5043 6411 5060 6431
rect 4903 6401 5060 6411
rect 4903 6400 4938 6401
rect 3967 6377 4005 6386
rect 4903 6379 4934 6400
rect 5121 6379 5157 6489
rect 5176 6488 5213 6489
rect 5272 6488 5309 6489
rect 5232 6429 5322 6435
rect 5232 6409 5241 6429
rect 5261 6427 5322 6429
rect 5261 6409 5286 6427
rect 5232 6407 5286 6409
rect 5306 6407 5322 6427
rect 5232 6401 5322 6407
rect 4746 6378 4783 6379
rect 3967 6376 4004 6377
rect 3428 6348 3518 6354
rect 3428 6328 3444 6348
rect 3464 6346 3518 6348
rect 3464 6328 3489 6346
rect 3428 6326 3489 6328
rect 3509 6326 3518 6346
rect 3428 6320 3518 6326
rect 3441 6266 3478 6267
rect 3537 6266 3574 6267
rect 3593 6266 3629 6376
rect 3816 6355 3847 6376
rect 4745 6369 4783 6378
rect 3812 6354 3847 6355
rect 3690 6344 3847 6354
rect 3690 6324 3707 6344
rect 3727 6324 3847 6344
rect 3690 6317 3847 6324
rect 3914 6347 4063 6355
rect 3914 6327 3925 6347
rect 3945 6327 3984 6347
rect 4004 6327 4063 6347
rect 4573 6351 4613 6361
rect 3914 6320 4063 6327
rect 4129 6323 4181 6341
rect 3914 6319 3955 6320
rect 3648 6266 3685 6267
rect 3341 6257 3479 6266
rect 2813 6246 2846 6248
rect 2442 6234 2889 6246
rect 2445 6220 2889 6234
rect 2445 6218 2613 6220
rect 2445 6040 2472 6218
rect 2512 6180 2576 6192
rect 2852 6188 2889 6220
rect 2915 6219 3106 6241
rect 3341 6237 3450 6257
rect 3470 6237 3479 6257
rect 3341 6230 3479 6237
rect 3537 6257 3685 6266
rect 3537 6237 3546 6257
rect 3566 6237 3656 6257
rect 3676 6237 3685 6257
rect 3341 6228 3437 6230
rect 3537 6227 3685 6237
rect 3744 6257 3781 6267
rect 3744 6237 3752 6257
rect 3772 6237 3781 6257
rect 3593 6226 3629 6227
rect 3070 6217 3106 6219
rect 3070 6188 3107 6217
rect 2512 6179 2547 6180
rect 2489 6174 2547 6179
rect 2489 6154 2492 6174
rect 2512 6160 2547 6174
rect 2567 6160 2576 6180
rect 2512 6152 2576 6160
rect 2538 6151 2576 6152
rect 2539 6150 2576 6151
rect 2642 6184 2678 6185
rect 2750 6184 2786 6185
rect 2642 6176 2786 6184
rect 2642 6156 2650 6176
rect 2670 6174 2758 6176
rect 2670 6156 2703 6174
rect 2642 6155 2703 6156
rect 2724 6156 2758 6174
rect 2778 6156 2786 6176
rect 2724 6155 2786 6156
rect 2642 6150 2786 6155
rect 2852 6180 2890 6188
rect 2968 6184 3004 6185
rect 2852 6160 2861 6180
rect 2881 6160 2890 6180
rect 2852 6151 2890 6160
rect 2919 6176 3004 6184
rect 2919 6156 2976 6176
rect 2996 6156 3004 6176
rect 2852 6150 2889 6151
rect 2919 6150 3004 6156
rect 3070 6180 3108 6188
rect 3070 6160 3079 6180
rect 3099 6160 3108 6180
rect 3744 6170 3781 6237
rect 3816 6266 3847 6317
rect 4129 6305 4147 6323
rect 4165 6305 4181 6323
rect 3866 6266 3903 6267
rect 3816 6257 3903 6266
rect 3816 6237 3874 6257
rect 3894 6237 3903 6257
rect 3816 6227 3903 6237
rect 3962 6257 3999 6267
rect 3962 6237 3970 6257
rect 3990 6237 3999 6257
rect 3816 6226 3847 6227
rect 3441 6167 3478 6168
rect 3744 6167 3783 6170
rect 3440 6166 3783 6167
rect 3962 6166 3999 6237
rect 3070 6151 3108 6160
rect 3365 6161 3783 6166
rect 3070 6150 3107 6151
rect 2531 6122 2621 6128
rect 2531 6102 2547 6122
rect 2567 6120 2621 6122
rect 2567 6102 2592 6120
rect 2531 6100 2592 6102
rect 2612 6100 2621 6120
rect 2531 6094 2621 6100
rect 2544 6040 2581 6041
rect 2640 6040 2677 6041
rect 2696 6040 2732 6150
rect 2919 6129 2950 6150
rect 3365 6141 3368 6161
rect 3388 6141 3783 6161
rect 3812 6142 3999 6166
rect 2915 6128 2950 6129
rect 2793 6118 2950 6128
rect 2793 6098 2810 6118
rect 2830 6098 2950 6118
rect 2793 6091 2950 6098
rect 3017 6121 3166 6129
rect 3017 6101 3028 6121
rect 3048 6101 3087 6121
rect 3107 6101 3166 6121
rect 3017 6094 3166 6101
rect 3744 6116 3783 6141
rect 4129 6116 4181 6305
rect 4573 6333 4583 6351
rect 4601 6333 4613 6351
rect 4745 6349 4754 6369
rect 4774 6349 4783 6369
rect 4745 6341 4783 6349
rect 4849 6373 4934 6379
rect 4964 6378 5001 6379
rect 4849 6353 4857 6373
rect 4877 6353 4934 6373
rect 4849 6345 4934 6353
rect 4963 6369 5001 6378
rect 4963 6349 4972 6369
rect 4992 6349 5001 6369
rect 4849 6344 4885 6345
rect 4963 6341 5001 6349
rect 5067 6373 5211 6379
rect 5067 6353 5075 6373
rect 5095 6353 5128 6373
rect 5148 6353 5183 6373
rect 5203 6353 5211 6373
rect 5067 6345 5211 6353
rect 5067 6344 5103 6345
rect 5175 6344 5211 6345
rect 5277 6378 5314 6379
rect 5277 6377 5315 6378
rect 5277 6369 5341 6377
rect 5277 6349 5286 6369
rect 5306 6355 5341 6369
rect 5361 6355 5364 6375
rect 5306 6350 5364 6355
rect 5306 6349 5341 6350
rect 4573 6277 4613 6333
rect 4746 6312 4783 6341
rect 4747 6310 4783 6312
rect 4747 6288 4938 6310
rect 4964 6309 5001 6341
rect 5277 6337 5341 6349
rect 5381 6311 5408 6489
rect 6312 6486 6341 6504
rect 5240 6309 5408 6311
rect 4964 6299 5408 6309
rect 5549 6405 5736 6429
rect 5767 6410 6160 6430
rect 6180 6410 6183 6430
rect 5767 6405 6183 6410
rect 5549 6334 5586 6405
rect 5767 6404 6108 6405
rect 5701 6344 5732 6345
rect 5549 6314 5558 6334
rect 5578 6314 5586 6334
rect 5549 6304 5586 6314
rect 5645 6334 5732 6344
rect 5645 6314 5654 6334
rect 5674 6314 5732 6334
rect 5645 6305 5732 6314
rect 5645 6304 5682 6305
rect 4570 6272 4613 6277
rect 4961 6283 5408 6299
rect 4961 6277 4989 6283
rect 5240 6282 5408 6283
rect 4570 6269 4720 6272
rect 4961 6269 4988 6277
rect 4570 6267 4988 6269
rect 4570 6249 4579 6267
rect 4597 6249 4988 6267
rect 5701 6254 5732 6305
rect 5767 6334 5804 6404
rect 6070 6403 6107 6404
rect 5919 6344 5955 6345
rect 5767 6314 5776 6334
rect 5796 6314 5804 6334
rect 5767 6304 5804 6314
rect 5863 6334 6011 6344
rect 6111 6341 6207 6343
rect 5863 6314 5872 6334
rect 5892 6314 5982 6334
rect 6002 6314 6011 6334
rect 5863 6305 6011 6314
rect 6069 6334 6207 6341
rect 6069 6314 6078 6334
rect 6098 6314 6207 6334
rect 6069 6305 6207 6314
rect 5863 6304 5900 6305
rect 5593 6251 5634 6252
rect 4570 6246 4988 6249
rect 4570 6240 4613 6246
rect 4573 6237 4613 6240
rect 5485 6244 5634 6251
rect 4970 6228 5010 6229
rect 4681 6211 5010 6228
rect 5485 6224 5544 6244
rect 5564 6224 5603 6244
rect 5623 6224 5634 6244
rect 5485 6216 5634 6224
rect 5701 6247 5858 6254
rect 5701 6227 5821 6247
rect 5841 6227 5858 6247
rect 5701 6217 5858 6227
rect 5701 6216 5736 6217
rect 4565 6168 4608 6179
rect 4565 6150 4577 6168
rect 4595 6150 4608 6168
rect 4565 6124 4608 6150
rect 4681 6124 4708 6211
rect 4970 6202 5010 6211
rect 3744 6098 4183 6116
rect 3017 6093 3058 6094
rect 2751 6040 2788 6041
rect 2444 6031 2582 6040
rect 2444 6011 2553 6031
rect 2573 6011 2582 6031
rect 2444 6004 2582 6011
rect 2640 6031 2788 6040
rect 2640 6011 2649 6031
rect 2669 6011 2759 6031
rect 2779 6011 2788 6031
rect 2444 6002 2540 6004
rect 2640 6001 2788 6011
rect 2847 6031 2884 6041
rect 2847 6011 2855 6031
rect 2875 6011 2884 6031
rect 2696 6000 2732 6001
rect 2544 5941 2581 5942
rect 2847 5941 2884 6011
rect 2919 6040 2950 6091
rect 3744 6080 4144 6098
rect 4162 6080 4183 6098
rect 3744 6074 4183 6080
rect 3750 6070 4183 6074
rect 4565 6103 4708 6124
rect 4752 6176 4786 6192
rect 4970 6182 5363 6202
rect 5383 6182 5386 6202
rect 5701 6195 5732 6216
rect 5919 6195 5955 6305
rect 5974 6304 6011 6305
rect 6070 6304 6107 6305
rect 6030 6245 6120 6251
rect 6030 6225 6039 6245
rect 6059 6243 6120 6245
rect 6059 6225 6084 6243
rect 6030 6223 6084 6225
rect 6104 6223 6120 6243
rect 6030 6217 6120 6223
rect 5544 6194 5581 6195
rect 4970 6177 5386 6182
rect 5543 6185 5581 6194
rect 4970 6176 5311 6177
rect 4752 6106 4789 6176
rect 4904 6116 4935 6117
rect 4565 6101 4702 6103
rect 4129 6068 4181 6070
rect 4565 6059 4608 6101
rect 4752 6086 4761 6106
rect 4781 6086 4789 6106
rect 4752 6076 4789 6086
rect 4848 6106 4935 6116
rect 4848 6086 4857 6106
rect 4877 6086 4935 6106
rect 4848 6077 4935 6086
rect 4848 6076 4885 6077
rect 4563 6049 4608 6059
rect 2969 6040 3006 6041
rect 2919 6031 3006 6040
rect 2919 6011 2977 6031
rect 2997 6011 3006 6031
rect 2919 6001 3006 6011
rect 3065 6031 3102 6041
rect 3065 6011 3073 6031
rect 3093 6011 3102 6031
rect 4563 6031 4572 6049
rect 4590 6031 4608 6049
rect 4563 6025 4608 6031
rect 4904 6026 4935 6077
rect 4970 6106 5007 6176
rect 5273 6175 5310 6176
rect 5543 6165 5552 6185
rect 5572 6165 5581 6185
rect 5543 6157 5581 6165
rect 5647 6189 5732 6195
rect 5762 6194 5799 6195
rect 5647 6169 5655 6189
rect 5675 6169 5732 6189
rect 5647 6161 5732 6169
rect 5761 6185 5799 6194
rect 5761 6165 5770 6185
rect 5790 6165 5799 6185
rect 5647 6160 5683 6161
rect 5761 6157 5799 6165
rect 5865 6189 6009 6195
rect 5865 6169 5873 6189
rect 5893 6170 5925 6189
rect 5946 6170 5981 6189
rect 5893 6169 5981 6170
rect 6001 6169 6009 6189
rect 5865 6161 6009 6169
rect 5865 6160 5901 6161
rect 5973 6160 6009 6161
rect 6075 6194 6112 6195
rect 6075 6193 6113 6194
rect 6075 6185 6139 6193
rect 6075 6165 6084 6185
rect 6104 6171 6139 6185
rect 6159 6171 6162 6191
rect 6104 6166 6162 6171
rect 6104 6165 6139 6166
rect 5544 6128 5581 6157
rect 5545 6126 5581 6128
rect 5122 6116 5158 6117
rect 4970 6086 4979 6106
rect 4999 6086 5007 6106
rect 4970 6076 5007 6086
rect 5066 6106 5214 6116
rect 5314 6113 5410 6115
rect 5066 6086 5075 6106
rect 5095 6086 5185 6106
rect 5205 6086 5214 6106
rect 5066 6077 5214 6086
rect 5272 6106 5410 6113
rect 5272 6086 5281 6106
rect 5301 6086 5410 6106
rect 5545 6104 5736 6126
rect 5762 6125 5799 6157
rect 6075 6153 6139 6165
rect 6179 6127 6206 6305
rect 6038 6125 6206 6127
rect 5762 6099 6206 6125
rect 5272 6077 5410 6086
rect 5066 6076 5103 6077
rect 4563 6022 4600 6025
rect 4796 6023 4837 6024
rect 2919 6000 2950 6001
rect 2543 5940 2884 5941
rect 3065 5940 3102 6011
rect 4688 6016 4837 6023
rect 4132 6003 4169 6008
rect 4123 5999 4170 6003
rect 4123 5981 4142 5999
rect 4160 5981 4170 5999
rect 4688 5996 4747 6016
rect 4767 5996 4806 6016
rect 4826 5996 4837 6016
rect 4688 5988 4837 5996
rect 4904 6019 5061 6026
rect 4904 5999 5024 6019
rect 5044 5999 5061 6019
rect 4904 5989 5061 5999
rect 4904 5988 4939 5989
rect 2468 5935 2884 5940
rect 2468 5915 2471 5935
rect 2491 5915 2884 5935
rect 2915 5916 3102 5940
rect 3727 5938 3767 5943
rect 4123 5938 4170 5981
rect 4904 5967 4935 5988
rect 5122 5967 5158 6077
rect 5177 6076 5214 6077
rect 5273 6076 5310 6077
rect 5233 6017 5323 6023
rect 5233 5997 5242 6017
rect 5262 6015 5323 6017
rect 5262 5997 5287 6015
rect 5233 5995 5287 5997
rect 5307 5995 5323 6015
rect 5233 5989 5323 5995
rect 4747 5966 4784 5967
rect 3727 5899 4170 5938
rect 4560 5958 4597 5960
rect 4560 5950 4602 5958
rect 4560 5932 4570 5950
rect 4588 5932 4602 5950
rect 4560 5923 4602 5932
rect 4746 5957 4784 5966
rect 4746 5937 4755 5957
rect 4775 5937 4784 5957
rect 4746 5929 4784 5937
rect 4850 5961 4935 5967
rect 4965 5966 5002 5967
rect 4850 5941 4858 5961
rect 4878 5941 4935 5961
rect 4850 5933 4935 5941
rect 4964 5957 5002 5966
rect 4964 5937 4973 5957
rect 4993 5937 5002 5957
rect 4850 5932 4886 5933
rect 4964 5929 5002 5937
rect 5068 5965 5212 5967
rect 5068 5961 5120 5965
rect 5068 5941 5076 5961
rect 5096 5945 5120 5961
rect 5140 5961 5212 5965
rect 5140 5945 5184 5961
rect 5096 5941 5184 5945
rect 5204 5941 5212 5961
rect 5068 5933 5212 5941
rect 5068 5932 5104 5933
rect 5176 5932 5212 5933
rect 5278 5966 5315 5967
rect 5278 5965 5316 5966
rect 5278 5957 5342 5965
rect 5278 5937 5287 5957
rect 5307 5943 5342 5957
rect 5362 5943 5365 5963
rect 5307 5938 5365 5943
rect 5307 5937 5342 5938
rect 2821 5884 2861 5892
rect 2821 5862 2829 5884
rect 2853 5862 2861 5884
rect 2527 5638 2695 5639
rect 2821 5638 2861 5862
rect 3324 5866 3492 5867
rect 3727 5866 3767 5899
rect 4123 5866 4170 5899
rect 4561 5898 4602 5923
rect 4747 5898 4784 5929
rect 4965 5898 5002 5929
rect 5278 5925 5342 5937
rect 5382 5899 5409 6077
rect 4561 5871 4610 5898
rect 4746 5872 4795 5898
rect 4964 5897 5045 5898
rect 5241 5897 5409 5899
rect 4964 5872 5409 5897
rect 4965 5871 5409 5872
rect 3324 5865 3768 5866
rect 3324 5840 3769 5865
rect 3324 5838 3492 5840
rect 3688 5839 3769 5840
rect 3938 5839 3987 5865
rect 4123 5839 4172 5866
rect 3324 5660 3351 5838
rect 3391 5800 3455 5812
rect 3731 5808 3768 5839
rect 3949 5808 3986 5839
rect 4131 5814 4172 5839
rect 4563 5838 4610 5871
rect 4966 5838 5006 5871
rect 5241 5870 5409 5871
rect 5872 5875 5912 6099
rect 6038 6098 6206 6099
rect 5872 5853 5880 5875
rect 5904 5853 5912 5875
rect 5872 5845 5912 5853
rect 3391 5799 3426 5800
rect 3368 5794 3426 5799
rect 3368 5774 3371 5794
rect 3391 5780 3426 5794
rect 3446 5780 3455 5800
rect 3391 5772 3455 5780
rect 3417 5771 3455 5772
rect 3418 5770 3455 5771
rect 3521 5804 3557 5805
rect 3629 5804 3665 5805
rect 3521 5796 3665 5804
rect 3521 5776 3529 5796
rect 3549 5792 3637 5796
rect 3549 5776 3593 5792
rect 3521 5772 3593 5776
rect 3613 5776 3637 5792
rect 3657 5776 3665 5796
rect 3613 5772 3665 5776
rect 3521 5770 3665 5772
rect 3731 5800 3769 5808
rect 3847 5804 3883 5805
rect 3731 5780 3740 5800
rect 3760 5780 3769 5800
rect 3731 5771 3769 5780
rect 3798 5796 3883 5804
rect 3798 5776 3855 5796
rect 3875 5776 3883 5796
rect 3731 5770 3768 5771
rect 3798 5770 3883 5776
rect 3949 5800 3987 5808
rect 3949 5780 3958 5800
rect 3978 5780 3987 5800
rect 3949 5771 3987 5780
rect 4131 5805 4173 5814
rect 4131 5787 4145 5805
rect 4163 5787 4173 5805
rect 4131 5779 4173 5787
rect 4136 5777 4173 5779
rect 4563 5799 5006 5838
rect 3949 5770 3986 5771
rect 3410 5742 3500 5748
rect 3410 5722 3426 5742
rect 3446 5740 3500 5742
rect 3446 5722 3471 5740
rect 3410 5720 3471 5722
rect 3491 5720 3500 5740
rect 3410 5714 3500 5720
rect 3423 5660 3460 5661
rect 3519 5660 3556 5661
rect 3575 5660 3611 5770
rect 3798 5749 3829 5770
rect 4563 5756 4610 5799
rect 4966 5794 5006 5799
rect 5631 5797 5818 5821
rect 5849 5802 6242 5822
rect 6262 5802 6265 5822
rect 5849 5797 6265 5802
rect 3794 5748 3829 5749
rect 3672 5738 3829 5748
rect 3672 5718 3689 5738
rect 3709 5718 3829 5738
rect 3672 5711 3829 5718
rect 3896 5741 4045 5749
rect 3896 5721 3907 5741
rect 3927 5721 3966 5741
rect 3986 5721 4045 5741
rect 4563 5738 4573 5756
rect 4591 5738 4610 5756
rect 4563 5734 4610 5738
rect 4564 5729 4601 5734
rect 3896 5714 4045 5721
rect 5631 5726 5668 5797
rect 5849 5796 6190 5797
rect 5783 5736 5814 5737
rect 3896 5713 3937 5714
rect 4133 5712 4170 5715
rect 3630 5660 3667 5661
rect 3323 5651 3461 5660
rect 2527 5612 2971 5638
rect 2527 5610 2695 5612
rect 2527 5432 2554 5610
rect 2594 5572 2658 5584
rect 2934 5580 2971 5612
rect 2997 5611 3188 5633
rect 3323 5631 3432 5651
rect 3452 5631 3461 5651
rect 3323 5624 3461 5631
rect 3519 5651 3667 5660
rect 3519 5631 3528 5651
rect 3548 5631 3638 5651
rect 3658 5631 3667 5651
rect 3323 5622 3419 5624
rect 3519 5621 3667 5631
rect 3726 5651 3763 5661
rect 3726 5631 3734 5651
rect 3754 5631 3763 5651
rect 3575 5620 3611 5621
rect 3152 5609 3188 5611
rect 3152 5580 3189 5609
rect 2594 5571 2629 5572
rect 2571 5566 2629 5571
rect 2571 5546 2574 5566
rect 2594 5552 2629 5566
rect 2649 5552 2658 5572
rect 2594 5544 2658 5552
rect 2620 5543 2658 5544
rect 2621 5542 2658 5543
rect 2724 5576 2760 5577
rect 2832 5576 2868 5577
rect 2724 5568 2868 5576
rect 2724 5548 2732 5568
rect 2752 5567 2840 5568
rect 2752 5548 2787 5567
rect 2808 5548 2840 5567
rect 2860 5548 2868 5568
rect 2724 5542 2868 5548
rect 2934 5572 2972 5580
rect 3050 5576 3086 5577
rect 2934 5552 2943 5572
rect 2963 5552 2972 5572
rect 2934 5543 2972 5552
rect 3001 5568 3086 5576
rect 3001 5548 3058 5568
rect 3078 5548 3086 5568
rect 2934 5542 2971 5543
rect 3001 5542 3086 5548
rect 3152 5572 3190 5580
rect 3152 5552 3161 5572
rect 3181 5552 3190 5572
rect 3423 5561 3460 5562
rect 3726 5561 3763 5631
rect 3798 5660 3829 5711
rect 4125 5706 4170 5712
rect 4125 5688 4143 5706
rect 4161 5688 4170 5706
rect 5631 5706 5640 5726
rect 5660 5706 5668 5726
rect 5631 5696 5668 5706
rect 5727 5726 5814 5736
rect 5727 5706 5736 5726
rect 5756 5706 5814 5726
rect 5727 5697 5814 5706
rect 5727 5696 5764 5697
rect 4125 5678 4170 5688
rect 3848 5660 3885 5661
rect 3798 5651 3885 5660
rect 3798 5631 3856 5651
rect 3876 5631 3885 5651
rect 3798 5621 3885 5631
rect 3944 5651 3981 5661
rect 3944 5631 3952 5651
rect 3972 5631 3981 5651
rect 4125 5636 4168 5678
rect 4552 5667 4604 5669
rect 4031 5634 4168 5636
rect 3798 5620 3829 5621
rect 3944 5561 3981 5631
rect 3422 5560 3763 5561
rect 3152 5543 3190 5552
rect 3347 5555 3763 5560
rect 3152 5542 3189 5543
rect 2613 5514 2703 5520
rect 2613 5494 2629 5514
rect 2649 5512 2703 5514
rect 2649 5494 2674 5512
rect 2613 5492 2674 5494
rect 2694 5492 2703 5512
rect 2613 5486 2703 5492
rect 2626 5432 2663 5433
rect 2722 5432 2759 5433
rect 2778 5432 2814 5542
rect 3001 5521 3032 5542
rect 3347 5535 3350 5555
rect 3370 5535 3763 5555
rect 3947 5545 3981 5561
rect 4025 5613 4168 5634
rect 4550 5663 4983 5667
rect 4550 5657 4989 5663
rect 4550 5639 4571 5657
rect 4589 5639 4989 5657
rect 5783 5646 5814 5697
rect 5849 5726 5886 5796
rect 6152 5795 6189 5796
rect 6001 5736 6037 5737
rect 5849 5706 5858 5726
rect 5878 5706 5886 5726
rect 5849 5696 5886 5706
rect 5945 5726 6093 5736
rect 6193 5733 6289 5735
rect 5945 5706 5954 5726
rect 5974 5706 6064 5726
rect 6084 5706 6093 5726
rect 5945 5697 6093 5706
rect 6151 5726 6289 5733
rect 6151 5706 6160 5726
rect 6180 5706 6289 5726
rect 6151 5697 6289 5706
rect 5945 5696 5982 5697
rect 5675 5643 5716 5644
rect 4550 5621 4989 5639
rect 3723 5526 3763 5535
rect 4025 5526 4052 5613
rect 4125 5587 4168 5613
rect 4125 5569 4138 5587
rect 4156 5569 4168 5587
rect 4125 5558 4168 5569
rect 2997 5520 3032 5521
rect 2875 5510 3032 5520
rect 2875 5490 2892 5510
rect 2912 5490 3032 5510
rect 2875 5483 3032 5490
rect 3099 5513 3248 5521
rect 3099 5493 3110 5513
rect 3130 5493 3169 5513
rect 3189 5493 3248 5513
rect 3723 5509 4052 5526
rect 3723 5508 3763 5509
rect 3099 5486 3248 5493
rect 4120 5497 4160 5500
rect 4120 5491 4163 5497
rect 3745 5488 4163 5491
rect 3099 5485 3140 5486
rect 2833 5432 2870 5433
rect 2526 5423 2664 5432
rect 2224 5248 2264 5420
rect 2526 5403 2635 5423
rect 2655 5403 2664 5423
rect 2526 5396 2664 5403
rect 2722 5423 2870 5432
rect 2722 5403 2731 5423
rect 2751 5403 2841 5423
rect 2861 5403 2870 5423
rect 2526 5394 2622 5396
rect 2722 5393 2870 5403
rect 2929 5423 2966 5433
rect 2929 5403 2937 5423
rect 2957 5403 2966 5423
rect 2778 5392 2814 5393
rect 2626 5333 2663 5334
rect 2929 5333 2966 5403
rect 3001 5432 3032 5483
rect 3745 5470 4136 5488
rect 4154 5470 4163 5488
rect 3745 5468 4163 5470
rect 3745 5460 3772 5468
rect 4013 5465 4163 5468
rect 3325 5454 3493 5455
rect 3744 5454 3772 5460
rect 3325 5438 3772 5454
rect 4120 5460 4163 5465
rect 3051 5432 3088 5433
rect 3001 5423 3088 5432
rect 3001 5403 3059 5423
rect 3079 5403 3088 5423
rect 3001 5393 3088 5403
rect 3147 5423 3184 5433
rect 3147 5403 3155 5423
rect 3175 5403 3184 5423
rect 3001 5392 3032 5393
rect 2625 5332 2966 5333
rect 3147 5332 3184 5403
rect 2550 5327 2966 5332
rect 2550 5307 2553 5327
rect 2573 5307 2966 5327
rect 2997 5308 3184 5332
rect 3325 5428 3769 5438
rect 3325 5426 3493 5428
rect 3325 5248 3352 5426
rect 3392 5388 3456 5400
rect 3732 5396 3769 5428
rect 3795 5427 3986 5449
rect 3950 5425 3986 5427
rect 3950 5396 3987 5425
rect 4120 5404 4160 5460
rect 3392 5387 3427 5388
rect 3369 5382 3427 5387
rect 3369 5362 3372 5382
rect 3392 5368 3427 5382
rect 3447 5368 3456 5388
rect 3392 5360 3456 5368
rect 3418 5359 3456 5360
rect 3419 5358 3456 5359
rect 3522 5392 3558 5393
rect 3630 5392 3666 5393
rect 3522 5384 3666 5392
rect 3522 5364 3530 5384
rect 3550 5364 3585 5384
rect 3605 5364 3638 5384
rect 3658 5364 3666 5384
rect 3522 5358 3666 5364
rect 3732 5388 3770 5396
rect 3848 5392 3884 5393
rect 3732 5368 3741 5388
rect 3761 5368 3770 5388
rect 3732 5359 3770 5368
rect 3799 5384 3884 5392
rect 3799 5364 3856 5384
rect 3876 5364 3884 5384
rect 3732 5358 3769 5359
rect 3799 5358 3884 5364
rect 3950 5388 3988 5396
rect 3950 5368 3959 5388
rect 3979 5368 3988 5388
rect 4120 5386 4132 5404
rect 4150 5386 4160 5404
rect 4552 5432 4604 5621
rect 4950 5596 4989 5621
rect 5567 5636 5716 5643
rect 5567 5616 5626 5636
rect 5646 5616 5685 5636
rect 5705 5616 5716 5636
rect 5567 5608 5716 5616
rect 5783 5639 5940 5646
rect 5783 5619 5903 5639
rect 5923 5619 5940 5639
rect 5783 5609 5940 5619
rect 5783 5608 5818 5609
rect 4734 5571 4921 5595
rect 4950 5576 5345 5596
rect 5365 5576 5368 5596
rect 5783 5587 5814 5608
rect 6001 5587 6037 5697
rect 6056 5696 6093 5697
rect 6152 5696 6189 5697
rect 6112 5637 6202 5643
rect 6112 5617 6121 5637
rect 6141 5635 6202 5637
rect 6141 5617 6166 5635
rect 6112 5615 6166 5617
rect 6186 5615 6202 5635
rect 6112 5609 6202 5615
rect 5626 5586 5663 5587
rect 4950 5571 5368 5576
rect 5625 5577 5663 5586
rect 4734 5500 4771 5571
rect 4950 5570 5293 5571
rect 4950 5567 4989 5570
rect 5255 5569 5292 5570
rect 4886 5510 4917 5511
rect 4734 5480 4743 5500
rect 4763 5480 4771 5500
rect 4734 5470 4771 5480
rect 4830 5500 4917 5510
rect 4830 5480 4839 5500
rect 4859 5480 4917 5500
rect 4830 5471 4917 5480
rect 4830 5470 4867 5471
rect 4552 5414 4568 5432
rect 4586 5414 4604 5432
rect 4886 5420 4917 5471
rect 4952 5500 4989 5567
rect 5625 5557 5634 5577
rect 5654 5557 5663 5577
rect 5625 5549 5663 5557
rect 5729 5581 5814 5587
rect 5844 5586 5881 5587
rect 5729 5561 5737 5581
rect 5757 5561 5814 5581
rect 5729 5553 5814 5561
rect 5843 5577 5881 5586
rect 5843 5557 5852 5577
rect 5872 5557 5881 5577
rect 5729 5552 5765 5553
rect 5843 5549 5881 5557
rect 5947 5581 6091 5587
rect 5947 5561 5955 5581
rect 5975 5576 6063 5581
rect 5975 5561 6011 5576
rect 5947 5559 6011 5561
rect 6030 5561 6063 5576
rect 6083 5561 6091 5581
rect 6030 5559 6091 5561
rect 5947 5553 6091 5559
rect 5947 5552 5983 5553
rect 6055 5552 6091 5553
rect 6157 5586 6194 5587
rect 6157 5585 6195 5586
rect 6157 5577 6221 5585
rect 6157 5557 6166 5577
rect 6186 5563 6221 5577
rect 6241 5563 6244 5583
rect 6186 5558 6244 5563
rect 6186 5557 6221 5558
rect 5626 5520 5663 5549
rect 5627 5518 5663 5520
rect 5104 5510 5140 5511
rect 4952 5480 4961 5500
rect 4981 5480 4989 5500
rect 4952 5470 4989 5480
rect 5048 5500 5196 5510
rect 5296 5507 5392 5509
rect 5048 5480 5057 5500
rect 5077 5480 5167 5500
rect 5187 5480 5196 5500
rect 5048 5471 5196 5480
rect 5254 5500 5392 5507
rect 5254 5480 5263 5500
rect 5283 5480 5392 5500
rect 5627 5496 5818 5518
rect 5844 5517 5881 5549
rect 6157 5545 6221 5557
rect 6261 5519 6288 5697
rect 6120 5517 6288 5519
rect 5844 5503 6288 5517
rect 6312 5540 6340 6486
rect 6312 5510 6357 5540
rect 5844 5491 6291 5503
rect 5887 5489 5920 5491
rect 5254 5471 5392 5480
rect 5048 5470 5085 5471
rect 4778 5417 4819 5418
rect 4552 5396 4604 5414
rect 4670 5410 4819 5417
rect 4120 5376 4160 5386
rect 4670 5390 4729 5410
rect 4749 5390 4788 5410
rect 4808 5390 4819 5410
rect 4670 5382 4819 5390
rect 4886 5413 5043 5420
rect 4886 5393 5006 5413
rect 5026 5393 5043 5413
rect 4886 5383 5043 5393
rect 4886 5382 4921 5383
rect 3950 5359 3988 5368
rect 4886 5361 4917 5382
rect 5104 5361 5140 5471
rect 5159 5470 5196 5471
rect 5255 5470 5292 5471
rect 5215 5411 5305 5417
rect 5215 5391 5224 5411
rect 5244 5409 5305 5411
rect 5244 5391 5269 5409
rect 5215 5389 5269 5391
rect 5289 5389 5305 5409
rect 5215 5383 5305 5389
rect 4729 5360 4766 5361
rect 3950 5358 3987 5359
rect 3411 5330 3501 5336
rect 3411 5310 3427 5330
rect 3447 5328 3501 5330
rect 3447 5310 3472 5328
rect 3411 5308 3472 5310
rect 3492 5308 3501 5328
rect 3411 5302 3501 5308
rect 3424 5248 3461 5249
rect 3520 5248 3557 5249
rect 3576 5248 3612 5358
rect 3799 5337 3830 5358
rect 4728 5351 4766 5360
rect 3795 5336 3830 5337
rect 3673 5326 3830 5336
rect 3673 5306 3690 5326
rect 3710 5306 3830 5326
rect 3673 5299 3830 5306
rect 3897 5329 4046 5337
rect 3897 5309 3908 5329
rect 3928 5309 3967 5329
rect 3987 5309 4046 5329
rect 4556 5333 4596 5343
rect 3897 5302 4046 5309
rect 4112 5305 4164 5323
rect 3897 5301 3938 5302
rect 3631 5248 3668 5249
rect 2225 5233 2264 5248
rect 3324 5239 3462 5248
rect 2225 5232 2391 5233
rect 2517 5232 2557 5234
rect 2225 5206 2667 5232
rect 2225 5204 2391 5206
rect 1889 5092 1926 5100
rect 1889 5073 1897 5092
rect 1918 5073 1926 5092
rect 1889 5067 1926 5073
rect 2225 5026 2250 5204
rect 2290 5166 2354 5178
rect 2630 5174 2667 5206
rect 2693 5205 2884 5227
rect 3324 5219 3433 5239
rect 3453 5219 3462 5239
rect 3324 5212 3462 5219
rect 3520 5239 3668 5248
rect 3520 5219 3529 5239
rect 3549 5219 3639 5239
rect 3659 5219 3668 5239
rect 3324 5210 3420 5212
rect 3520 5209 3668 5219
rect 3727 5239 3764 5249
rect 3727 5219 3735 5239
rect 3755 5219 3764 5239
rect 3576 5208 3612 5209
rect 2848 5203 2884 5205
rect 2848 5174 2885 5203
rect 2290 5165 2325 5166
rect 2267 5160 2325 5165
rect 2267 5140 2270 5160
rect 2290 5146 2325 5160
rect 2345 5146 2354 5166
rect 2290 5138 2354 5146
rect 2316 5137 2354 5138
rect 2317 5136 2354 5137
rect 2420 5170 2456 5171
rect 2528 5170 2564 5171
rect 2420 5165 2564 5170
rect 2420 5162 2482 5165
rect 2420 5142 2428 5162
rect 2448 5142 2482 5162
rect 2420 5139 2482 5142
rect 2508 5162 2564 5165
rect 2508 5142 2536 5162
rect 2556 5142 2564 5162
rect 2508 5139 2564 5142
rect 2420 5136 2564 5139
rect 2630 5166 2668 5174
rect 2746 5170 2782 5171
rect 2630 5146 2639 5166
rect 2659 5146 2668 5166
rect 2630 5137 2668 5146
rect 2697 5162 2782 5170
rect 2697 5142 2754 5162
rect 2774 5142 2782 5162
rect 2630 5136 2667 5137
rect 2697 5136 2782 5142
rect 2848 5166 2886 5174
rect 2848 5146 2857 5166
rect 2877 5146 2886 5166
rect 3727 5152 3764 5219
rect 3799 5248 3830 5299
rect 4112 5287 4130 5305
rect 4148 5287 4164 5305
rect 3849 5248 3886 5249
rect 3799 5239 3886 5248
rect 3799 5219 3857 5239
rect 3877 5219 3886 5239
rect 3799 5209 3886 5219
rect 3945 5239 3982 5249
rect 3945 5219 3953 5239
rect 3973 5219 3982 5239
rect 3799 5208 3830 5209
rect 3424 5149 3461 5150
rect 3727 5149 3766 5152
rect 3423 5148 3766 5149
rect 3945 5148 3982 5219
rect 2848 5137 2886 5146
rect 3348 5143 3766 5148
rect 2848 5136 2885 5137
rect 2309 5108 2399 5114
rect 2309 5088 2325 5108
rect 2345 5106 2399 5108
rect 2345 5088 2370 5106
rect 2309 5086 2370 5088
rect 2390 5086 2399 5106
rect 2309 5080 2399 5086
rect 2322 5026 2359 5027
rect 2418 5026 2455 5027
rect 2474 5026 2510 5136
rect 2697 5115 2728 5136
rect 3348 5123 3351 5143
rect 3371 5123 3766 5143
rect 3795 5124 3982 5148
rect 2693 5114 2728 5115
rect 2571 5104 2728 5114
rect 2571 5084 2588 5104
rect 2608 5084 2728 5104
rect 2571 5077 2728 5084
rect 2795 5107 2944 5115
rect 2795 5087 2806 5107
rect 2826 5087 2865 5107
rect 2885 5087 2944 5107
rect 2795 5080 2944 5087
rect 3727 5098 3766 5123
rect 4112 5098 4164 5287
rect 4556 5315 4566 5333
rect 4584 5315 4596 5333
rect 4728 5331 4737 5351
rect 4757 5331 4766 5351
rect 4728 5323 4766 5331
rect 4832 5355 4917 5361
rect 4947 5360 4984 5361
rect 4832 5335 4840 5355
rect 4860 5335 4917 5355
rect 4832 5327 4917 5335
rect 4946 5351 4984 5360
rect 4946 5331 4955 5351
rect 4975 5331 4984 5351
rect 4832 5326 4868 5327
rect 4946 5323 4984 5331
rect 5050 5355 5194 5361
rect 5050 5335 5058 5355
rect 5078 5335 5111 5355
rect 5131 5335 5166 5355
rect 5186 5335 5194 5355
rect 5050 5327 5194 5335
rect 5050 5326 5086 5327
rect 5158 5326 5194 5327
rect 5260 5360 5297 5361
rect 5260 5359 5298 5360
rect 5260 5351 5324 5359
rect 5260 5331 5269 5351
rect 5289 5337 5324 5351
rect 5344 5337 5347 5357
rect 5289 5332 5347 5337
rect 5289 5331 5324 5332
rect 4556 5259 4596 5315
rect 4729 5294 4766 5323
rect 4730 5292 4766 5294
rect 4730 5270 4921 5292
rect 4947 5291 4984 5323
rect 5260 5319 5324 5331
rect 5364 5293 5391 5471
rect 6249 5446 6291 5491
rect 6312 5492 6323 5510
rect 6345 5492 6357 5510
rect 6312 5486 6357 5492
rect 6313 5485 6357 5486
rect 5223 5291 5391 5293
rect 4947 5281 5391 5291
rect 5532 5387 5719 5411
rect 5750 5392 6143 5412
rect 6163 5392 6166 5412
rect 5750 5387 6166 5392
rect 5532 5316 5569 5387
rect 5750 5386 6091 5387
rect 5684 5326 5715 5327
rect 5532 5296 5541 5316
rect 5561 5296 5569 5316
rect 5532 5286 5569 5296
rect 5628 5316 5715 5326
rect 5628 5296 5637 5316
rect 5657 5296 5715 5316
rect 5628 5287 5715 5296
rect 5628 5286 5665 5287
rect 4553 5254 4596 5259
rect 4944 5265 5391 5281
rect 4944 5259 4972 5265
rect 5223 5264 5391 5265
rect 4553 5251 4703 5254
rect 4944 5251 4971 5259
rect 4553 5249 4971 5251
rect 4553 5231 4562 5249
rect 4580 5231 4971 5249
rect 5684 5236 5715 5287
rect 5750 5316 5787 5386
rect 6053 5385 6090 5386
rect 5902 5326 5938 5327
rect 5750 5296 5759 5316
rect 5779 5296 5787 5316
rect 5750 5286 5787 5296
rect 5846 5316 5994 5326
rect 6094 5323 6190 5325
rect 5846 5296 5855 5316
rect 5875 5296 5965 5316
rect 5985 5296 5994 5316
rect 5846 5287 5994 5296
rect 6052 5316 6190 5323
rect 6052 5296 6061 5316
rect 6081 5296 6190 5316
rect 6052 5287 6190 5296
rect 5846 5286 5883 5287
rect 5576 5233 5617 5234
rect 4553 5228 4971 5231
rect 4553 5222 4596 5228
rect 4556 5219 4596 5222
rect 5471 5226 5617 5233
rect 4953 5210 4993 5211
rect 4664 5193 4993 5210
rect 5471 5206 5527 5226
rect 5547 5206 5586 5226
rect 5606 5206 5617 5226
rect 5471 5198 5617 5206
rect 5684 5229 5841 5236
rect 5684 5209 5804 5229
rect 5824 5209 5841 5229
rect 5684 5199 5841 5209
rect 5684 5198 5719 5199
rect 4548 5150 4591 5161
rect 4548 5132 4560 5150
rect 4578 5132 4591 5150
rect 4548 5106 4591 5132
rect 4664 5106 4691 5193
rect 4953 5184 4993 5193
rect 3727 5080 4166 5098
rect 2795 5079 2836 5080
rect 2529 5026 2566 5027
rect 2225 5017 2360 5026
rect 2225 4997 2331 5017
rect 2351 4997 2360 5017
rect 2225 4990 2360 4997
rect 2418 5017 2566 5026
rect 2418 4997 2427 5017
rect 2447 4997 2537 5017
rect 2557 4997 2566 5017
rect 2225 4988 2318 4990
rect 2418 4987 2566 4997
rect 2625 5017 2662 5027
rect 2625 4997 2633 5017
rect 2653 4997 2662 5017
rect 2474 4986 2510 4987
rect 2322 4927 2359 4928
rect 2625 4927 2662 4997
rect 2697 5026 2728 5077
rect 3727 5062 4127 5080
rect 4145 5062 4166 5080
rect 3727 5056 4166 5062
rect 3733 5052 4166 5056
rect 4548 5085 4691 5106
rect 4735 5158 4769 5174
rect 4953 5164 5346 5184
rect 5366 5164 5369 5184
rect 5684 5177 5715 5198
rect 5902 5177 5938 5287
rect 5957 5286 5994 5287
rect 6053 5286 6090 5287
rect 6013 5227 6103 5233
rect 6013 5207 6022 5227
rect 6042 5225 6103 5227
rect 6042 5207 6067 5225
rect 6013 5205 6067 5207
rect 6087 5205 6103 5225
rect 6013 5199 6103 5205
rect 5527 5176 5564 5177
rect 4953 5159 5369 5164
rect 5526 5167 5564 5176
rect 4953 5158 5294 5159
rect 4735 5088 4772 5158
rect 4887 5098 4918 5099
rect 4548 5083 4685 5085
rect 4112 5050 4164 5052
rect 4548 5041 4591 5083
rect 4735 5068 4744 5088
rect 4764 5068 4772 5088
rect 4735 5058 4772 5068
rect 4831 5088 4918 5098
rect 4831 5068 4840 5088
rect 4860 5068 4918 5088
rect 4831 5059 4918 5068
rect 4831 5058 4868 5059
rect 4546 5031 4591 5041
rect 2747 5026 2784 5027
rect 2697 5017 2784 5026
rect 2697 4997 2755 5017
rect 2775 4997 2784 5017
rect 2697 4987 2784 4997
rect 2843 5017 2880 5027
rect 2843 4997 2851 5017
rect 2871 4997 2880 5017
rect 4546 5013 4555 5031
rect 4573 5013 4591 5031
rect 4546 5007 4591 5013
rect 4887 5008 4918 5059
rect 4953 5088 4990 5158
rect 5256 5157 5293 5158
rect 5526 5147 5535 5167
rect 5555 5147 5564 5167
rect 5526 5139 5564 5147
rect 5630 5171 5715 5177
rect 5745 5176 5782 5177
rect 5630 5151 5638 5171
rect 5658 5151 5715 5171
rect 5630 5143 5715 5151
rect 5744 5167 5782 5176
rect 5744 5147 5753 5167
rect 5773 5147 5782 5167
rect 5630 5142 5666 5143
rect 5744 5139 5782 5147
rect 5848 5171 5992 5177
rect 5848 5151 5856 5171
rect 5876 5168 5964 5171
rect 5876 5151 5911 5168
rect 5848 5150 5911 5151
rect 5930 5151 5964 5168
rect 5984 5151 5992 5171
rect 5930 5150 5992 5151
rect 5848 5143 5992 5150
rect 5848 5142 5884 5143
rect 5956 5142 5992 5143
rect 6058 5176 6095 5177
rect 6058 5175 6096 5176
rect 6118 5175 6145 5179
rect 6058 5173 6145 5175
rect 6058 5167 6122 5173
rect 6058 5147 6067 5167
rect 6087 5153 6122 5167
rect 6142 5153 6145 5173
rect 6087 5148 6145 5153
rect 6087 5147 6122 5148
rect 5527 5110 5564 5139
rect 5528 5108 5564 5110
rect 5105 5098 5141 5099
rect 4953 5068 4962 5088
rect 4982 5068 4990 5088
rect 4953 5058 4990 5068
rect 5049 5088 5197 5098
rect 5297 5095 5393 5097
rect 5049 5068 5058 5088
rect 5078 5068 5168 5088
rect 5188 5068 5197 5088
rect 5049 5059 5197 5068
rect 5255 5088 5393 5095
rect 5255 5068 5264 5088
rect 5284 5068 5393 5088
rect 5528 5086 5719 5108
rect 5745 5107 5782 5139
rect 6058 5135 6122 5147
rect 6162 5109 6189 5287
rect 6021 5107 6189 5109
rect 5745 5081 6189 5107
rect 5255 5059 5393 5068
rect 5049 5058 5086 5059
rect 4546 5004 4583 5007
rect 4779 5005 4820 5006
rect 2697 4986 2728 4987
rect 2321 4926 2662 4927
rect 2843 4926 2880 4997
rect 4671 4998 4820 5005
rect 4115 4985 4152 4990
rect 2246 4921 2662 4926
rect 2246 4901 2249 4921
rect 2269 4901 2662 4921
rect 2693 4902 2880 4926
rect 4106 4981 4153 4985
rect 4106 4963 4125 4981
rect 4143 4963 4153 4981
rect 4671 4978 4730 4998
rect 4750 4978 4789 4998
rect 4809 4978 4820 4998
rect 4671 4970 4820 4978
rect 4887 5001 5044 5008
rect 4887 4981 5007 5001
rect 5027 4981 5044 5001
rect 4887 4971 5044 4981
rect 4887 4970 4922 4971
rect 3714 4904 3752 4905
rect 4106 4904 4153 4963
rect 4887 4949 4918 4970
rect 5105 4949 5141 5059
rect 5160 5058 5197 5059
rect 5256 5058 5293 5059
rect 5216 4999 5306 5005
rect 5216 4979 5225 4999
rect 5245 4997 5306 4999
rect 5245 4979 5270 4997
rect 5216 4977 5270 4979
rect 5290 4977 5306 4997
rect 5216 4971 5306 4977
rect 4730 4948 4767 4949
rect 4543 4940 4580 4942
rect 4543 4932 4585 4940
rect 4543 4914 4553 4932
rect 4571 4914 4585 4932
rect 4543 4905 4585 4914
rect 4729 4939 4767 4948
rect 4729 4919 4738 4939
rect 4758 4919 4767 4939
rect 4729 4911 4767 4919
rect 4833 4943 4918 4949
rect 4948 4948 4985 4949
rect 4833 4923 4841 4943
rect 4861 4923 4918 4943
rect 4833 4915 4918 4923
rect 4947 4939 4985 4948
rect 4947 4919 4956 4939
rect 4976 4919 4985 4939
rect 4833 4914 4869 4915
rect 4947 4911 4985 4919
rect 5051 4947 5195 4949
rect 5051 4943 5103 4947
rect 5051 4923 5059 4943
rect 5079 4927 5103 4943
rect 5123 4943 5195 4947
rect 5123 4927 5167 4943
rect 5079 4923 5167 4927
rect 5187 4923 5195 4943
rect 5051 4915 5195 4923
rect 5051 4914 5087 4915
rect 5159 4914 5195 4915
rect 5261 4948 5298 4949
rect 5261 4947 5299 4948
rect 5261 4939 5325 4947
rect 5261 4919 5270 4939
rect 5290 4925 5325 4939
rect 5345 4925 5348 4945
rect 5290 4920 5348 4925
rect 5290 4919 5325 4920
rect 2466 4900 2531 4901
rect 581 4822 619 4823
rect 180 4784 619 4822
rect 1491 4822 1499 4844
rect 1523 4822 1531 4844
rect 1491 4814 1531 4822
rect 2802 4866 2842 4874
rect 2802 4844 2810 4866
rect 2834 4844 2842 4866
rect 3714 4866 4153 4904
rect 3714 4865 3752 4866
rect 1802 4787 1867 4788
rect 180 4725 227 4784
rect 581 4783 619 4784
rect 180 4707 190 4725
rect 208 4707 227 4725
rect 180 4703 227 4707
rect 1453 4762 1640 4786
rect 1671 4767 2064 4787
rect 2084 4767 2087 4787
rect 1671 4762 2087 4767
rect 181 4698 218 4703
rect 1453 4691 1490 4762
rect 1671 4761 2012 4762
rect 1605 4701 1636 4702
rect 1453 4671 1462 4691
rect 1482 4671 1490 4691
rect 1453 4661 1490 4671
rect 1549 4691 1636 4701
rect 1549 4671 1558 4691
rect 1578 4671 1636 4691
rect 1549 4662 1636 4671
rect 1549 4661 1586 4662
rect 169 4636 221 4638
rect 167 4632 600 4636
rect 167 4626 606 4632
rect 167 4608 188 4626
rect 206 4608 606 4626
rect 1605 4611 1636 4662
rect 1671 4691 1708 4761
rect 1974 4760 2011 4761
rect 1823 4701 1859 4702
rect 1671 4671 1680 4691
rect 1700 4671 1708 4691
rect 1671 4661 1708 4671
rect 1767 4691 1915 4701
rect 2015 4698 2111 4700
rect 1767 4671 1776 4691
rect 1796 4671 1886 4691
rect 1906 4671 1915 4691
rect 1767 4662 1915 4671
rect 1973 4691 2111 4698
rect 1973 4671 1982 4691
rect 2002 4671 2111 4691
rect 1973 4662 2111 4671
rect 1767 4661 1804 4662
rect 1497 4608 1538 4609
rect 167 4590 606 4608
rect 169 4401 221 4590
rect 567 4565 606 4590
rect 1389 4601 1538 4608
rect 1389 4581 1448 4601
rect 1468 4581 1507 4601
rect 1527 4581 1538 4601
rect 1389 4573 1538 4581
rect 1605 4604 1762 4611
rect 1605 4584 1725 4604
rect 1745 4584 1762 4604
rect 1605 4574 1762 4584
rect 1605 4573 1640 4574
rect 351 4540 538 4564
rect 567 4545 962 4565
rect 982 4545 985 4565
rect 1605 4552 1636 4573
rect 1823 4552 1859 4662
rect 1878 4661 1915 4662
rect 1974 4661 2011 4662
rect 1934 4602 2024 4608
rect 1934 4582 1943 4602
rect 1963 4600 2024 4602
rect 1963 4582 1988 4600
rect 1934 4580 1988 4582
rect 2008 4580 2024 4600
rect 1934 4574 2024 4580
rect 1448 4551 1485 4552
rect 567 4540 985 4545
rect 1447 4542 1485 4551
rect 351 4469 388 4540
rect 567 4539 910 4540
rect 567 4536 606 4539
rect 872 4538 909 4539
rect 503 4479 534 4480
rect 351 4449 360 4469
rect 380 4449 388 4469
rect 351 4439 388 4449
rect 447 4469 534 4479
rect 447 4449 456 4469
rect 476 4449 534 4469
rect 447 4440 534 4449
rect 447 4439 484 4440
rect 169 4383 185 4401
rect 203 4383 221 4401
rect 503 4389 534 4440
rect 569 4469 606 4536
rect 1447 4522 1456 4542
rect 1476 4522 1485 4542
rect 1447 4514 1485 4522
rect 1551 4546 1636 4552
rect 1666 4551 1703 4552
rect 1551 4526 1559 4546
rect 1579 4526 1636 4546
rect 1551 4518 1636 4526
rect 1665 4542 1703 4551
rect 1665 4522 1674 4542
rect 1694 4522 1703 4542
rect 1551 4517 1587 4518
rect 1665 4514 1703 4522
rect 1769 4546 1913 4552
rect 1769 4526 1777 4546
rect 1797 4540 1885 4546
rect 1797 4526 1826 4540
rect 1769 4518 1826 4526
rect 1769 4517 1805 4518
rect 1849 4526 1885 4540
rect 1905 4526 1913 4546
rect 1849 4518 1913 4526
rect 1877 4517 1913 4518
rect 1979 4551 2016 4552
rect 1979 4550 2017 4551
rect 1979 4542 2043 4550
rect 1979 4522 1988 4542
rect 2008 4528 2043 4542
rect 2063 4528 2066 4548
rect 2008 4523 2066 4528
rect 2008 4522 2043 4523
rect 1448 4485 1485 4514
rect 1449 4483 1485 4485
rect 721 4479 757 4480
rect 569 4449 578 4469
rect 598 4449 606 4469
rect 569 4439 606 4449
rect 665 4469 813 4479
rect 913 4476 1009 4478
rect 665 4449 674 4469
rect 694 4449 784 4469
rect 804 4449 813 4469
rect 665 4440 813 4449
rect 871 4469 1009 4476
rect 871 4449 880 4469
rect 900 4449 1009 4469
rect 1449 4461 1640 4483
rect 1666 4482 1703 4514
rect 1979 4510 2043 4522
rect 2083 4484 2110 4662
rect 2407 4615 2444 4621
rect 2407 4596 2415 4615
rect 2436 4596 2444 4615
rect 2407 4588 2444 4596
rect 1942 4482 2110 4484
rect 1666 4456 2110 4482
rect 1776 4454 1816 4456
rect 1942 4455 2110 4456
rect 871 4440 1009 4449
rect 2069 4450 2110 4455
rect 665 4439 702 4440
rect 395 4386 436 4387
rect 169 4365 221 4383
rect 287 4379 436 4386
rect 287 4359 346 4379
rect 366 4359 405 4379
rect 425 4359 436 4379
rect 287 4351 436 4359
rect 503 4382 660 4389
rect 503 4362 623 4382
rect 643 4362 660 4382
rect 503 4352 660 4362
rect 503 4351 538 4352
rect 503 4330 534 4351
rect 721 4330 757 4440
rect 776 4439 813 4440
rect 872 4439 909 4440
rect 832 4380 922 4386
rect 832 4360 841 4380
rect 861 4378 922 4380
rect 861 4360 886 4378
rect 832 4358 886 4360
rect 906 4358 922 4378
rect 832 4352 922 4358
rect 346 4329 383 4330
rect 345 4320 383 4329
rect 173 4302 213 4312
rect 173 4284 183 4302
rect 201 4284 213 4302
rect 345 4300 354 4320
rect 374 4300 383 4320
rect 345 4292 383 4300
rect 449 4324 534 4330
rect 564 4329 601 4330
rect 449 4304 457 4324
rect 477 4304 534 4324
rect 449 4296 534 4304
rect 563 4320 601 4329
rect 563 4300 572 4320
rect 592 4300 601 4320
rect 449 4295 485 4296
rect 563 4292 601 4300
rect 667 4324 811 4330
rect 667 4304 675 4324
rect 695 4304 728 4324
rect 748 4304 783 4324
rect 803 4304 811 4324
rect 667 4296 811 4304
rect 667 4295 703 4296
rect 775 4295 811 4296
rect 877 4329 914 4330
rect 877 4328 915 4329
rect 877 4320 941 4328
rect 877 4300 886 4320
rect 906 4306 941 4320
rect 961 4306 964 4326
rect 906 4301 964 4306
rect 906 4300 941 4301
rect 173 4228 213 4284
rect 346 4263 383 4292
rect 347 4261 383 4263
rect 347 4239 538 4261
rect 564 4260 601 4292
rect 877 4288 941 4300
rect 981 4262 1008 4440
rect 840 4260 1008 4262
rect 564 4250 1008 4260
rect 1149 4356 1336 4380
rect 1367 4361 1760 4381
rect 1780 4361 1783 4381
rect 1367 4356 1783 4361
rect 1149 4285 1186 4356
rect 1367 4355 1708 4356
rect 1301 4295 1332 4296
rect 1149 4265 1158 4285
rect 1178 4265 1186 4285
rect 1149 4255 1186 4265
rect 1245 4285 1332 4295
rect 1245 4265 1254 4285
rect 1274 4265 1332 4285
rect 1245 4256 1332 4265
rect 1245 4255 1282 4256
rect 170 4223 213 4228
rect 561 4234 1008 4250
rect 561 4228 589 4234
rect 840 4233 1008 4234
rect 170 4220 320 4223
rect 561 4220 588 4228
rect 170 4218 588 4220
rect 170 4200 179 4218
rect 197 4200 588 4218
rect 1301 4205 1332 4256
rect 1367 4285 1404 4355
rect 1670 4354 1707 4355
rect 1519 4295 1555 4296
rect 1367 4265 1376 4285
rect 1396 4265 1404 4285
rect 1367 4255 1404 4265
rect 1463 4285 1611 4295
rect 1711 4292 1807 4294
rect 1463 4265 1472 4285
rect 1492 4265 1582 4285
rect 1602 4265 1611 4285
rect 1463 4256 1611 4265
rect 1669 4285 1807 4292
rect 1669 4265 1678 4285
rect 1698 4265 1807 4285
rect 2069 4268 2109 4450
rect 1669 4256 1807 4265
rect 1463 4255 1500 4256
rect 1193 4202 1234 4203
rect 170 4197 588 4200
rect 170 4191 213 4197
rect 173 4188 213 4191
rect 1085 4195 1234 4202
rect 570 4179 610 4180
rect 281 4162 610 4179
rect 1085 4175 1144 4195
rect 1164 4175 1203 4195
rect 1223 4175 1234 4195
rect 1085 4167 1234 4175
rect 1301 4198 1458 4205
rect 1301 4178 1421 4198
rect 1441 4178 1458 4198
rect 1301 4168 1458 4178
rect 1301 4167 1336 4168
rect 165 4119 208 4130
rect 165 4101 177 4119
rect 195 4101 208 4119
rect 165 4075 208 4101
rect 281 4075 308 4162
rect 570 4153 610 4162
rect 165 4054 308 4075
rect 352 4127 386 4143
rect 570 4133 963 4153
rect 983 4133 986 4153
rect 1301 4146 1332 4167
rect 1519 4146 1555 4256
rect 1574 4255 1611 4256
rect 1670 4255 1707 4256
rect 1630 4196 1720 4202
rect 1630 4176 1639 4196
rect 1659 4194 1720 4196
rect 1659 4176 1684 4194
rect 1630 4174 1684 4176
rect 1704 4174 1720 4194
rect 1630 4168 1720 4174
rect 1144 4145 1181 4146
rect 570 4128 986 4133
rect 1143 4136 1181 4145
rect 570 4127 911 4128
rect 352 4057 389 4127
rect 504 4067 535 4068
rect 165 4052 302 4054
rect 165 4010 208 4052
rect 352 4037 361 4057
rect 381 4037 389 4057
rect 352 4027 389 4037
rect 448 4057 535 4067
rect 448 4037 457 4057
rect 477 4037 535 4057
rect 448 4028 535 4037
rect 448 4027 485 4028
rect 163 4000 208 4010
rect 163 3982 172 4000
rect 190 3982 208 4000
rect 163 3976 208 3982
rect 504 3977 535 4028
rect 570 4057 607 4127
rect 873 4126 910 4127
rect 1143 4116 1152 4136
rect 1172 4116 1181 4136
rect 1143 4108 1181 4116
rect 1247 4140 1332 4146
rect 1362 4145 1399 4146
rect 1247 4120 1255 4140
rect 1275 4120 1332 4140
rect 1247 4112 1332 4120
rect 1361 4136 1399 4145
rect 1361 4116 1370 4136
rect 1390 4116 1399 4136
rect 1247 4111 1283 4112
rect 1361 4108 1399 4116
rect 1465 4140 1609 4146
rect 1465 4120 1473 4140
rect 1493 4121 1525 4140
rect 1546 4121 1581 4140
rect 1493 4120 1581 4121
rect 1601 4120 1609 4140
rect 1465 4112 1609 4120
rect 1465 4111 1501 4112
rect 1573 4111 1609 4112
rect 1675 4145 1712 4146
rect 1675 4144 1713 4145
rect 1675 4136 1739 4144
rect 1675 4116 1684 4136
rect 1704 4122 1739 4136
rect 1759 4122 1762 4142
rect 1704 4117 1762 4122
rect 1704 4116 1739 4117
rect 1144 4079 1181 4108
rect 1145 4077 1181 4079
rect 722 4067 758 4068
rect 570 4037 579 4057
rect 599 4037 607 4057
rect 570 4027 607 4037
rect 666 4057 814 4067
rect 914 4064 1010 4066
rect 666 4037 675 4057
rect 695 4037 785 4057
rect 805 4037 814 4057
rect 666 4028 814 4037
rect 872 4057 1010 4064
rect 872 4037 881 4057
rect 901 4037 1010 4057
rect 1145 4055 1336 4077
rect 1362 4076 1399 4108
rect 1675 4104 1739 4116
rect 1779 4078 1806 4256
rect 1638 4076 1806 4078
rect 1362 4050 1806 4076
rect 872 4028 1010 4037
rect 666 4027 703 4028
rect 163 3973 200 3976
rect 396 3974 437 3975
rect 288 3967 437 3974
rect 288 3947 347 3967
rect 367 3947 406 3967
rect 426 3947 437 3967
rect 288 3939 437 3947
rect 504 3970 661 3977
rect 504 3950 624 3970
rect 644 3950 661 3970
rect 504 3940 661 3950
rect 504 3939 539 3940
rect 504 3918 535 3939
rect 722 3918 758 4028
rect 777 4027 814 4028
rect 873 4027 910 4028
rect 833 3968 923 3974
rect 833 3948 842 3968
rect 862 3966 923 3968
rect 862 3948 887 3966
rect 833 3946 887 3948
rect 907 3946 923 3966
rect 833 3940 923 3946
rect 347 3917 384 3918
rect 160 3909 197 3911
rect 160 3901 202 3909
rect 160 3883 170 3901
rect 188 3883 202 3901
rect 160 3874 202 3883
rect 346 3908 384 3917
rect 346 3888 355 3908
rect 375 3888 384 3908
rect 346 3880 384 3888
rect 450 3912 535 3918
rect 565 3917 602 3918
rect 450 3892 458 3912
rect 478 3892 535 3912
rect 450 3884 535 3892
rect 564 3908 602 3917
rect 564 3888 573 3908
rect 593 3888 602 3908
rect 450 3883 486 3884
rect 564 3880 602 3888
rect 668 3916 812 3918
rect 668 3912 720 3916
rect 668 3892 676 3912
rect 696 3896 720 3912
rect 740 3912 812 3916
rect 740 3896 784 3912
rect 696 3892 784 3896
rect 804 3892 812 3912
rect 668 3884 812 3892
rect 668 3883 704 3884
rect 776 3883 812 3884
rect 878 3917 915 3918
rect 878 3916 916 3917
rect 878 3908 942 3916
rect 878 3888 887 3908
rect 907 3894 942 3908
rect 962 3894 965 3914
rect 907 3889 965 3894
rect 907 3888 942 3889
rect 161 3849 202 3874
rect 347 3849 384 3880
rect 565 3849 602 3880
rect 878 3876 942 3888
rect 982 3850 1009 4028
rect 161 3822 210 3849
rect 346 3823 395 3849
rect 564 3848 645 3849
rect 841 3848 1009 3850
rect 564 3823 1009 3848
rect 565 3822 1009 3823
rect 163 3789 210 3822
rect 566 3789 606 3822
rect 841 3821 1009 3822
rect 1472 3826 1512 4050
rect 1638 4049 1806 4050
rect 1472 3804 1480 3826
rect 1504 3804 1512 3826
rect 1472 3796 1512 3804
rect 163 3750 606 3789
rect 163 3707 210 3750
rect 566 3745 606 3750
rect 1231 3748 1418 3772
rect 1449 3753 1842 3773
rect 1862 3753 1865 3773
rect 1449 3748 1865 3753
rect 163 3689 173 3707
rect 191 3689 210 3707
rect 163 3685 210 3689
rect 164 3680 201 3685
rect 1231 3677 1268 3748
rect 1449 3747 1790 3748
rect 1383 3687 1414 3688
rect 1231 3657 1240 3677
rect 1260 3657 1268 3677
rect 1231 3647 1268 3657
rect 1327 3677 1414 3687
rect 1327 3657 1336 3677
rect 1356 3657 1414 3677
rect 1327 3648 1414 3657
rect 1327 3647 1364 3648
rect 152 3618 204 3620
rect 150 3614 583 3618
rect 150 3608 589 3614
rect 150 3590 171 3608
rect 189 3590 589 3608
rect 1383 3597 1414 3648
rect 1449 3677 1486 3747
rect 1752 3746 1789 3747
rect 1601 3687 1637 3688
rect 1449 3657 1458 3677
rect 1478 3657 1486 3677
rect 1449 3647 1486 3657
rect 1545 3677 1693 3687
rect 1793 3684 1889 3686
rect 1545 3657 1554 3677
rect 1574 3657 1664 3677
rect 1684 3657 1693 3677
rect 1545 3648 1693 3657
rect 1751 3677 1889 3684
rect 1751 3657 1760 3677
rect 1780 3657 1889 3677
rect 1751 3648 1889 3657
rect 1545 3647 1582 3648
rect 1275 3594 1316 3595
rect 150 3572 589 3590
rect 152 3383 204 3572
rect 550 3547 589 3572
rect 1167 3587 1316 3594
rect 1167 3567 1226 3587
rect 1246 3567 1285 3587
rect 1305 3567 1316 3587
rect 1167 3559 1316 3567
rect 1383 3590 1540 3597
rect 1383 3570 1503 3590
rect 1523 3570 1540 3590
rect 1383 3560 1540 3570
rect 1383 3559 1418 3560
rect 334 3522 521 3546
rect 550 3527 945 3547
rect 965 3527 968 3547
rect 1383 3538 1414 3559
rect 1601 3538 1637 3648
rect 1656 3647 1693 3648
rect 1752 3647 1789 3648
rect 1712 3588 1802 3594
rect 1712 3568 1721 3588
rect 1741 3586 1802 3588
rect 1741 3568 1766 3586
rect 1712 3566 1766 3568
rect 1786 3566 1802 3586
rect 1712 3560 1802 3566
rect 1226 3537 1263 3538
rect 550 3522 968 3527
rect 1225 3528 1263 3537
rect 334 3451 371 3522
rect 550 3521 893 3522
rect 550 3518 589 3521
rect 855 3520 892 3521
rect 486 3461 517 3462
rect 334 3431 343 3451
rect 363 3431 371 3451
rect 334 3421 371 3431
rect 430 3451 517 3461
rect 430 3431 439 3451
rect 459 3431 517 3451
rect 430 3422 517 3431
rect 430 3421 467 3422
rect 152 3365 168 3383
rect 186 3365 204 3383
rect 486 3371 517 3422
rect 552 3451 589 3518
rect 1225 3508 1234 3528
rect 1254 3508 1263 3528
rect 1225 3500 1263 3508
rect 1329 3532 1414 3538
rect 1444 3537 1481 3538
rect 1329 3512 1337 3532
rect 1357 3512 1414 3532
rect 1329 3504 1414 3512
rect 1443 3528 1481 3537
rect 1443 3508 1452 3528
rect 1472 3508 1481 3528
rect 1329 3503 1365 3504
rect 1443 3500 1481 3508
rect 1547 3533 1691 3538
rect 1547 3532 1609 3533
rect 1547 3512 1555 3532
rect 1575 3514 1609 3532
rect 1630 3532 1691 3533
rect 1630 3514 1663 3532
rect 1575 3512 1663 3514
rect 1683 3512 1691 3532
rect 1547 3504 1691 3512
rect 1547 3503 1583 3504
rect 1655 3503 1691 3504
rect 1757 3537 1794 3538
rect 1757 3536 1795 3537
rect 1757 3528 1821 3536
rect 1757 3508 1766 3528
rect 1786 3514 1821 3528
rect 1841 3514 1844 3534
rect 1786 3509 1844 3514
rect 1786 3508 1821 3509
rect 1226 3471 1263 3500
rect 1227 3469 1263 3471
rect 704 3461 740 3462
rect 552 3431 561 3451
rect 581 3431 589 3451
rect 552 3421 589 3431
rect 648 3451 796 3461
rect 896 3458 992 3460
rect 648 3431 657 3451
rect 677 3431 767 3451
rect 787 3431 796 3451
rect 648 3422 796 3431
rect 854 3451 992 3458
rect 854 3431 863 3451
rect 883 3431 992 3451
rect 1227 3447 1418 3469
rect 1444 3468 1481 3500
rect 1757 3496 1821 3508
rect 1861 3470 1888 3648
rect 1720 3468 1888 3470
rect 1444 3454 1888 3468
rect 1444 3442 1891 3454
rect 1487 3440 1520 3442
rect 854 3422 992 3431
rect 648 3421 685 3422
rect 378 3368 419 3369
rect 152 3347 204 3365
rect 270 3361 419 3368
rect 270 3341 329 3361
rect 349 3341 388 3361
rect 408 3341 419 3361
rect 270 3333 419 3341
rect 486 3364 643 3371
rect 486 3344 606 3364
rect 626 3344 643 3364
rect 486 3334 643 3344
rect 486 3333 521 3334
rect 486 3312 517 3333
rect 704 3312 740 3422
rect 759 3421 796 3422
rect 855 3421 892 3422
rect 815 3362 905 3368
rect 815 3342 824 3362
rect 844 3360 905 3362
rect 844 3342 869 3360
rect 815 3340 869 3342
rect 889 3340 905 3360
rect 815 3334 905 3340
rect 329 3311 366 3312
rect 328 3302 366 3311
rect 156 3284 196 3294
rect 156 3266 166 3284
rect 184 3266 196 3284
rect 328 3282 337 3302
rect 357 3282 366 3302
rect 328 3274 366 3282
rect 432 3306 517 3312
rect 547 3311 584 3312
rect 432 3286 440 3306
rect 460 3286 517 3306
rect 432 3278 517 3286
rect 546 3302 584 3311
rect 546 3282 555 3302
rect 575 3282 584 3302
rect 432 3277 468 3278
rect 546 3274 584 3282
rect 650 3306 794 3312
rect 650 3286 658 3306
rect 678 3286 711 3306
rect 731 3286 766 3306
rect 786 3286 794 3306
rect 650 3278 794 3286
rect 650 3277 686 3278
rect 758 3277 794 3278
rect 860 3311 897 3312
rect 860 3310 898 3311
rect 860 3302 924 3310
rect 860 3282 869 3302
rect 889 3288 924 3302
rect 944 3288 947 3308
rect 889 3283 947 3288
rect 889 3282 924 3283
rect 156 3210 196 3266
rect 329 3245 366 3274
rect 330 3243 366 3245
rect 330 3221 521 3243
rect 547 3242 584 3274
rect 860 3270 924 3282
rect 964 3244 991 3422
rect 1849 3397 1891 3442
rect 823 3242 991 3244
rect 547 3232 991 3242
rect 1132 3338 1319 3362
rect 1350 3343 1743 3363
rect 1763 3343 1766 3363
rect 1350 3338 1766 3343
rect 1132 3267 1169 3338
rect 1350 3337 1691 3338
rect 1284 3277 1315 3278
rect 1132 3247 1141 3267
rect 1161 3247 1169 3267
rect 1132 3237 1169 3247
rect 1228 3267 1315 3277
rect 1228 3247 1237 3267
rect 1257 3247 1315 3267
rect 1228 3238 1315 3247
rect 1228 3237 1265 3238
rect 153 3205 196 3210
rect 544 3216 991 3232
rect 544 3210 572 3216
rect 823 3215 991 3216
rect 153 3202 303 3205
rect 544 3202 571 3210
rect 153 3200 571 3202
rect 153 3182 162 3200
rect 180 3182 571 3200
rect 1284 3187 1315 3238
rect 1350 3267 1387 3337
rect 1653 3336 1690 3337
rect 1502 3277 1538 3278
rect 1350 3247 1359 3267
rect 1379 3247 1387 3267
rect 1350 3237 1387 3247
rect 1446 3267 1594 3277
rect 1694 3274 1790 3276
rect 1446 3247 1455 3267
rect 1475 3247 1565 3267
rect 1585 3247 1594 3267
rect 1446 3238 1594 3247
rect 1652 3267 1790 3274
rect 1652 3247 1661 3267
rect 1681 3247 1790 3267
rect 1652 3238 1790 3247
rect 1446 3237 1483 3238
rect 1176 3184 1217 3185
rect 153 3179 571 3182
rect 153 3173 196 3179
rect 156 3170 196 3173
rect 1071 3177 1217 3184
rect 553 3161 593 3162
rect 264 3144 593 3161
rect 1071 3157 1127 3177
rect 1147 3157 1186 3177
rect 1206 3157 1217 3177
rect 1071 3149 1217 3157
rect 1284 3180 1441 3187
rect 1284 3160 1404 3180
rect 1424 3160 1441 3180
rect 1284 3150 1441 3160
rect 1284 3149 1319 3150
rect 148 3101 191 3112
rect 148 3083 160 3101
rect 178 3083 191 3101
rect 148 3057 191 3083
rect 264 3057 291 3144
rect 553 3135 593 3144
rect 148 3036 291 3057
rect 335 3109 369 3125
rect 553 3115 946 3135
rect 966 3115 969 3135
rect 1284 3128 1315 3149
rect 1502 3128 1538 3238
rect 1557 3237 1594 3238
rect 1653 3237 1690 3238
rect 1613 3178 1703 3184
rect 1613 3158 1622 3178
rect 1642 3176 1703 3178
rect 1642 3158 1667 3176
rect 1613 3156 1667 3158
rect 1687 3156 1703 3176
rect 1613 3150 1703 3156
rect 1127 3127 1164 3128
rect 553 3110 969 3115
rect 1126 3118 1164 3127
rect 553 3109 894 3110
rect 335 3039 372 3109
rect 487 3049 518 3050
rect 148 3034 285 3036
rect 148 2992 191 3034
rect 335 3019 344 3039
rect 364 3019 372 3039
rect 335 3009 372 3019
rect 431 3039 518 3049
rect 431 3019 440 3039
rect 460 3019 518 3039
rect 431 3010 518 3019
rect 431 3009 468 3010
rect 146 2982 191 2992
rect 146 2964 155 2982
rect 173 2964 191 2982
rect 146 2958 191 2964
rect 487 2959 518 3010
rect 553 3039 590 3109
rect 856 3108 893 3109
rect 1126 3098 1135 3118
rect 1155 3098 1164 3118
rect 1126 3090 1164 3098
rect 1230 3122 1315 3128
rect 1345 3127 1382 3128
rect 1230 3102 1238 3122
rect 1258 3102 1315 3122
rect 1230 3094 1315 3102
rect 1344 3118 1382 3127
rect 1344 3098 1353 3118
rect 1373 3098 1382 3118
rect 1230 3093 1266 3094
rect 1344 3090 1382 3098
rect 1448 3122 1592 3128
rect 1448 3102 1456 3122
rect 1476 3119 1564 3122
rect 1476 3102 1511 3119
rect 1448 3101 1511 3102
rect 1530 3102 1564 3119
rect 1584 3102 1592 3122
rect 1530 3101 1592 3102
rect 1448 3094 1592 3101
rect 1448 3093 1484 3094
rect 1556 3093 1592 3094
rect 1658 3127 1695 3128
rect 1658 3126 1696 3127
rect 1718 3126 1745 3130
rect 1658 3124 1745 3126
rect 1658 3118 1722 3124
rect 1658 3098 1667 3118
rect 1687 3104 1722 3118
rect 1742 3104 1745 3124
rect 1687 3099 1745 3104
rect 1687 3098 1722 3099
rect 1127 3061 1164 3090
rect 1128 3059 1164 3061
rect 705 3049 741 3050
rect 553 3019 562 3039
rect 582 3019 590 3039
rect 553 3009 590 3019
rect 649 3039 797 3049
rect 897 3046 993 3048
rect 649 3019 658 3039
rect 678 3019 768 3039
rect 788 3019 797 3039
rect 649 3010 797 3019
rect 855 3039 993 3046
rect 855 3019 864 3039
rect 884 3019 993 3039
rect 1128 3037 1319 3059
rect 1345 3058 1382 3090
rect 1658 3086 1722 3098
rect 1762 3060 1789 3238
rect 1621 3058 1789 3060
rect 1345 3032 1789 3058
rect 855 3010 993 3019
rect 649 3009 686 3010
rect 146 2955 183 2958
rect 379 2956 420 2957
rect 271 2949 420 2956
rect 271 2929 330 2949
rect 350 2929 389 2949
rect 409 2929 420 2949
rect 271 2921 420 2929
rect 487 2952 644 2959
rect 487 2932 607 2952
rect 627 2932 644 2952
rect 487 2922 644 2932
rect 487 2921 522 2922
rect 487 2900 518 2921
rect 705 2900 741 3010
rect 760 3009 797 3010
rect 856 3009 893 3010
rect 816 2950 906 2956
rect 816 2930 825 2950
rect 845 2948 906 2950
rect 845 2930 870 2948
rect 816 2928 870 2930
rect 890 2928 906 2948
rect 816 2922 906 2928
rect 330 2899 367 2900
rect 142 2891 180 2893
rect 142 2883 185 2891
rect 142 2865 153 2883
rect 171 2865 185 2883
rect 142 2838 185 2865
rect 329 2890 367 2899
rect 329 2870 338 2890
rect 358 2870 367 2890
rect 329 2862 367 2870
rect 433 2894 518 2900
rect 548 2899 585 2900
rect 433 2874 441 2894
rect 461 2874 518 2894
rect 433 2866 518 2874
rect 547 2890 585 2899
rect 547 2870 556 2890
rect 576 2870 585 2890
rect 433 2865 469 2866
rect 547 2862 585 2870
rect 651 2898 795 2900
rect 651 2894 703 2898
rect 651 2874 659 2894
rect 679 2878 703 2894
rect 723 2894 795 2898
rect 723 2878 767 2894
rect 679 2874 767 2878
rect 787 2874 795 2894
rect 651 2866 795 2874
rect 651 2865 687 2866
rect 759 2865 795 2866
rect 861 2899 898 2900
rect 861 2898 899 2899
rect 861 2890 925 2898
rect 861 2870 870 2890
rect 890 2876 925 2890
rect 945 2876 948 2896
rect 890 2871 948 2876
rect 890 2870 925 2871
rect 143 2831 185 2838
rect 330 2831 367 2862
rect 548 2831 585 2862
rect 861 2858 925 2870
rect 965 2832 992 3010
rect 143 2791 188 2831
rect 330 2806 475 2831
rect 548 2830 628 2831
rect 824 2830 992 2832
rect 548 2814 992 2830
rect 332 2805 475 2806
rect 547 2804 992 2814
rect 143 2770 190 2791
rect 547 2770 588 2804
rect 824 2803 992 2804
rect 1455 2808 1495 3032
rect 1621 3031 1789 3032
rect 1853 3064 1886 3397
rect 1853 3056 1890 3064
rect 1853 3037 1861 3056
rect 1882 3037 1890 3056
rect 1853 3031 1890 3037
rect 1455 2786 1463 2808
rect 1487 2786 1495 2808
rect 1455 2778 1495 2786
rect 143 2740 588 2770
rect 1626 2753 1691 2754
rect 143 2737 566 2740
rect 143 2689 190 2737
rect 143 2671 153 2689
rect 171 2671 190 2689
rect 143 2667 190 2671
rect 1277 2728 1464 2752
rect 1495 2733 1888 2753
rect 1908 2733 1911 2753
rect 1495 2728 1911 2733
rect 144 2662 181 2667
rect 1277 2657 1314 2728
rect 1495 2727 1836 2728
rect 1429 2667 1460 2668
rect 1277 2637 1286 2657
rect 1306 2637 1314 2657
rect 1277 2627 1314 2637
rect 1373 2657 1460 2667
rect 1373 2637 1382 2657
rect 1402 2637 1460 2657
rect 1373 2628 1460 2637
rect 1373 2627 1410 2628
rect 132 2600 184 2602
rect 130 2596 563 2600
rect 130 2590 569 2596
rect 130 2572 151 2590
rect 169 2572 569 2590
rect 1429 2577 1460 2628
rect 1495 2657 1532 2727
rect 1798 2726 1835 2727
rect 1647 2667 1683 2668
rect 1495 2637 1504 2657
rect 1524 2637 1532 2657
rect 1495 2627 1532 2637
rect 1591 2657 1739 2667
rect 1839 2664 1935 2666
rect 1591 2637 1600 2657
rect 1620 2637 1710 2657
rect 1730 2637 1739 2657
rect 1591 2628 1739 2637
rect 1797 2657 1935 2664
rect 1797 2637 1806 2657
rect 1826 2637 1935 2657
rect 1797 2628 1935 2637
rect 1591 2627 1628 2628
rect 1321 2574 1362 2575
rect 130 2554 569 2572
rect 132 2365 184 2554
rect 530 2529 569 2554
rect 1213 2567 1362 2574
rect 1213 2547 1272 2567
rect 1292 2547 1331 2567
rect 1351 2547 1362 2567
rect 1213 2539 1362 2547
rect 1429 2570 1586 2577
rect 1429 2550 1549 2570
rect 1569 2550 1586 2570
rect 1429 2540 1586 2550
rect 1429 2539 1464 2540
rect 314 2504 501 2528
rect 530 2509 925 2529
rect 945 2509 948 2529
rect 1429 2518 1460 2539
rect 1647 2518 1683 2628
rect 1702 2627 1739 2628
rect 1798 2627 1835 2628
rect 1758 2568 1848 2574
rect 1758 2548 1767 2568
rect 1787 2566 1848 2568
rect 1787 2548 1812 2566
rect 1758 2546 1812 2548
rect 1832 2546 1848 2566
rect 1758 2540 1848 2546
rect 1272 2517 1309 2518
rect 530 2504 948 2509
rect 1271 2508 1309 2517
rect 314 2433 351 2504
rect 530 2503 873 2504
rect 530 2500 569 2503
rect 835 2502 872 2503
rect 466 2443 497 2444
rect 314 2413 323 2433
rect 343 2413 351 2433
rect 314 2403 351 2413
rect 410 2433 497 2443
rect 410 2413 419 2433
rect 439 2413 497 2433
rect 410 2404 497 2413
rect 410 2403 447 2404
rect 132 2347 148 2365
rect 166 2347 184 2365
rect 466 2353 497 2404
rect 532 2433 569 2500
rect 1271 2488 1280 2508
rect 1300 2488 1309 2508
rect 1271 2480 1309 2488
rect 1375 2512 1460 2518
rect 1490 2517 1527 2518
rect 1375 2492 1383 2512
rect 1403 2492 1460 2512
rect 1375 2484 1460 2492
rect 1489 2508 1527 2517
rect 1489 2488 1498 2508
rect 1518 2488 1527 2508
rect 1375 2483 1411 2484
rect 1489 2480 1527 2488
rect 1593 2516 1737 2518
rect 1593 2512 1653 2516
rect 1593 2492 1601 2512
rect 1621 2494 1653 2512
rect 1676 2512 1737 2516
rect 1676 2494 1709 2512
rect 1621 2492 1709 2494
rect 1729 2492 1737 2512
rect 1593 2484 1737 2492
rect 1593 2483 1629 2484
rect 1701 2483 1737 2484
rect 1803 2517 1840 2518
rect 1803 2516 1841 2517
rect 1803 2508 1867 2516
rect 1803 2488 1812 2508
rect 1832 2494 1867 2508
rect 1887 2494 1890 2514
rect 1832 2489 1890 2494
rect 1832 2488 1867 2489
rect 1272 2451 1309 2480
rect 1273 2449 1309 2451
rect 684 2443 720 2444
rect 532 2413 541 2433
rect 561 2413 569 2433
rect 532 2403 569 2413
rect 628 2433 776 2443
rect 876 2440 972 2442
rect 628 2413 637 2433
rect 657 2413 747 2433
rect 767 2413 776 2433
rect 628 2404 776 2413
rect 834 2433 972 2440
rect 834 2413 843 2433
rect 863 2413 972 2433
rect 1273 2427 1464 2449
rect 1490 2448 1527 2480
rect 1803 2476 1867 2488
rect 1490 2447 1765 2448
rect 1907 2447 1934 2628
rect 1490 2422 1934 2447
rect 2070 2453 2109 4268
rect 2411 4255 2444 4588
rect 2508 4620 2676 4621
rect 2802 4620 2842 4844
rect 3305 4848 3473 4849
rect 3714 4848 3749 4865
rect 4106 4855 4153 4866
rect 3305 4822 3749 4848
rect 3305 4820 3473 4822
rect 3669 4821 3749 4822
rect 3904 4821 3971 4847
rect 4110 4821 4153 4855
rect 3305 4642 3332 4820
rect 3372 4782 3436 4794
rect 3712 4790 3749 4821
rect 3930 4790 3967 4821
rect 4112 4796 4153 4821
rect 4544 4880 4585 4905
rect 4730 4880 4767 4911
rect 4948 4880 4985 4911
rect 5261 4907 5325 4919
rect 5365 4881 5392 5059
rect 4544 4846 4587 4880
rect 4726 4854 4793 4880
rect 4948 4879 5028 4880
rect 5224 4879 5392 4881
rect 4948 4853 5392 4879
rect 4544 4835 4591 4846
rect 4948 4836 4983 4853
rect 5224 4852 5392 4853
rect 5855 4857 5895 5081
rect 6021 5080 6189 5081
rect 6253 5113 6286 5446
rect 6588 5433 6627 7248
rect 6763 7254 7207 7279
rect 6763 7073 6790 7254
rect 6932 7253 7207 7254
rect 6830 7213 6894 7225
rect 7170 7221 7207 7253
rect 7233 7252 7424 7274
rect 7725 7268 7834 7288
rect 7854 7268 7863 7288
rect 7725 7261 7863 7268
rect 7921 7288 8069 7297
rect 7921 7268 7930 7288
rect 7950 7268 8040 7288
rect 8060 7268 8069 7288
rect 7725 7259 7821 7261
rect 7921 7258 8069 7268
rect 8128 7288 8165 7298
rect 8128 7268 8136 7288
rect 8156 7268 8165 7288
rect 7977 7257 8013 7258
rect 7388 7250 7424 7252
rect 7388 7221 7425 7250
rect 6830 7212 6865 7213
rect 6807 7207 6865 7212
rect 6807 7187 6810 7207
rect 6830 7193 6865 7207
rect 6885 7193 6894 7213
rect 6830 7185 6894 7193
rect 6856 7184 6894 7185
rect 6857 7183 6894 7184
rect 6960 7217 6996 7218
rect 7068 7217 7104 7218
rect 6960 7209 7104 7217
rect 6960 7189 6968 7209
rect 6988 7207 7076 7209
rect 6988 7189 7021 7207
rect 6960 7185 7021 7189
rect 7044 7189 7076 7207
rect 7096 7189 7104 7209
rect 7044 7185 7104 7189
rect 6960 7183 7104 7185
rect 7170 7213 7208 7221
rect 7286 7217 7322 7218
rect 7170 7193 7179 7213
rect 7199 7193 7208 7213
rect 7170 7184 7208 7193
rect 7237 7209 7322 7217
rect 7237 7189 7294 7209
rect 7314 7189 7322 7209
rect 7170 7183 7207 7184
rect 7237 7183 7322 7189
rect 7388 7213 7426 7221
rect 7388 7193 7397 7213
rect 7417 7193 7426 7213
rect 8128 7201 8165 7268
rect 8200 7297 8231 7348
rect 8513 7336 8531 7354
rect 8549 7336 8565 7354
rect 8250 7297 8287 7298
rect 8200 7288 8287 7297
rect 8200 7268 8258 7288
rect 8278 7268 8287 7288
rect 8200 7258 8287 7268
rect 8346 7288 8383 7298
rect 8346 7268 8354 7288
rect 8374 7268 8383 7288
rect 8200 7257 8231 7258
rect 7825 7198 7862 7199
rect 8128 7198 8167 7201
rect 7824 7197 8167 7198
rect 8346 7197 8383 7268
rect 7388 7184 7426 7193
rect 7749 7192 8167 7197
rect 7388 7183 7425 7184
rect 6849 7155 6939 7161
rect 6849 7135 6865 7155
rect 6885 7153 6939 7155
rect 6885 7135 6910 7153
rect 6849 7133 6910 7135
rect 6930 7133 6939 7153
rect 6849 7127 6939 7133
rect 6862 7073 6899 7074
rect 6958 7073 6995 7074
rect 7014 7073 7050 7183
rect 7237 7162 7268 7183
rect 7749 7172 7752 7192
rect 7772 7172 8167 7192
rect 8196 7173 8383 7197
rect 7233 7161 7268 7162
rect 7111 7151 7268 7161
rect 7111 7131 7128 7151
rect 7148 7131 7268 7151
rect 7111 7124 7268 7131
rect 7335 7154 7484 7162
rect 7335 7134 7346 7154
rect 7366 7134 7405 7154
rect 7425 7134 7484 7154
rect 7335 7127 7484 7134
rect 8128 7147 8167 7172
rect 8513 7147 8565 7336
rect 8970 7363 8980 7381
rect 8998 7363 9010 7381
rect 9142 7379 9151 7399
rect 9171 7379 9180 7399
rect 9142 7371 9180 7379
rect 9246 7403 9331 7409
rect 9361 7408 9398 7409
rect 9246 7383 9254 7403
rect 9274 7383 9331 7403
rect 9246 7375 9331 7383
rect 9360 7399 9398 7408
rect 9360 7379 9369 7399
rect 9389 7379 9398 7399
rect 9246 7374 9282 7375
rect 9360 7371 9398 7379
rect 9464 7403 9608 7409
rect 9464 7383 9472 7403
rect 9492 7383 9525 7403
rect 9545 7383 9580 7403
rect 9600 7383 9608 7403
rect 9464 7375 9608 7383
rect 9464 7374 9500 7375
rect 9572 7374 9608 7375
rect 9674 7408 9711 7409
rect 9674 7407 9712 7408
rect 9674 7399 9738 7407
rect 9674 7379 9683 7399
rect 9703 7385 9738 7399
rect 9758 7385 9761 7405
rect 9703 7380 9761 7385
rect 9703 7379 9738 7380
rect 8970 7307 9010 7363
rect 9143 7342 9180 7371
rect 9144 7340 9180 7342
rect 9144 7318 9335 7340
rect 9361 7339 9398 7371
rect 9674 7367 9738 7379
rect 9778 7341 9805 7519
rect 10663 7494 10705 7539
rect 9637 7339 9805 7341
rect 9361 7329 9805 7339
rect 9946 7435 10133 7459
rect 10164 7440 10557 7460
rect 10577 7440 10580 7460
rect 10164 7435 10580 7440
rect 9946 7364 9983 7435
rect 10164 7434 10505 7435
rect 10098 7374 10129 7375
rect 9946 7344 9955 7364
rect 9975 7344 9983 7364
rect 9946 7334 9983 7344
rect 10042 7364 10129 7374
rect 10042 7344 10051 7364
rect 10071 7344 10129 7364
rect 10042 7335 10129 7344
rect 10042 7334 10079 7335
rect 8967 7302 9010 7307
rect 9358 7313 9805 7329
rect 9358 7307 9386 7313
rect 9637 7312 9805 7313
rect 8967 7299 9117 7302
rect 9358 7299 9385 7307
rect 8967 7297 9385 7299
rect 8967 7279 8976 7297
rect 8994 7279 9385 7297
rect 10098 7284 10129 7335
rect 10164 7364 10201 7434
rect 10467 7433 10504 7434
rect 10316 7374 10352 7375
rect 10164 7344 10173 7364
rect 10193 7344 10201 7364
rect 10164 7334 10201 7344
rect 10260 7364 10408 7374
rect 10508 7371 10604 7373
rect 10260 7344 10269 7364
rect 10289 7344 10379 7364
rect 10399 7344 10408 7364
rect 10260 7335 10408 7344
rect 10466 7364 10604 7371
rect 10466 7344 10475 7364
rect 10495 7344 10604 7364
rect 10466 7335 10604 7344
rect 10260 7334 10297 7335
rect 9990 7281 10031 7282
rect 8967 7276 9385 7279
rect 8967 7270 9010 7276
rect 8970 7267 9010 7270
rect 9885 7274 10031 7281
rect 9367 7258 9407 7259
rect 9078 7241 9407 7258
rect 9885 7254 9941 7274
rect 9961 7254 10000 7274
rect 10020 7254 10031 7274
rect 9885 7246 10031 7254
rect 10098 7277 10255 7284
rect 10098 7257 10218 7277
rect 10238 7257 10255 7277
rect 10098 7247 10255 7257
rect 10098 7246 10133 7247
rect 8962 7198 9005 7209
rect 8962 7180 8974 7198
rect 8992 7180 9005 7198
rect 8962 7154 9005 7180
rect 9078 7154 9105 7241
rect 9367 7232 9407 7241
rect 8128 7129 8567 7147
rect 7335 7126 7376 7127
rect 7069 7073 7106 7074
rect 6762 7064 6900 7073
rect 6762 7044 6871 7064
rect 6891 7044 6900 7064
rect 6762 7037 6900 7044
rect 6958 7064 7106 7073
rect 6958 7044 6967 7064
rect 6987 7044 7077 7064
rect 7097 7044 7106 7064
rect 6762 7035 6858 7037
rect 6958 7034 7106 7044
rect 7165 7064 7202 7074
rect 7165 7044 7173 7064
rect 7193 7044 7202 7064
rect 7014 7033 7050 7034
rect 6862 6974 6899 6975
rect 7165 6974 7202 7044
rect 7237 7073 7268 7124
rect 8128 7111 8528 7129
rect 8546 7111 8567 7129
rect 8128 7105 8567 7111
rect 8134 7101 8567 7105
rect 8962 7133 9105 7154
rect 9149 7206 9183 7222
rect 9367 7212 9760 7232
rect 9780 7212 9783 7232
rect 10098 7225 10129 7246
rect 10316 7225 10352 7335
rect 10371 7334 10408 7335
rect 10467 7334 10504 7335
rect 10427 7275 10517 7281
rect 10427 7255 10436 7275
rect 10456 7273 10517 7275
rect 10456 7255 10481 7273
rect 10427 7253 10481 7255
rect 10501 7253 10517 7273
rect 10427 7247 10517 7253
rect 9941 7224 9978 7225
rect 9367 7207 9783 7212
rect 9940 7215 9978 7224
rect 9367 7206 9708 7207
rect 9149 7136 9186 7206
rect 9301 7146 9332 7147
rect 8962 7131 9099 7133
rect 8513 7099 8565 7101
rect 8962 7089 9005 7131
rect 9149 7116 9158 7136
rect 9178 7116 9186 7136
rect 9149 7106 9186 7116
rect 9245 7136 9332 7146
rect 9245 7116 9254 7136
rect 9274 7116 9332 7136
rect 9245 7107 9332 7116
rect 9245 7106 9282 7107
rect 8960 7079 9005 7089
rect 7287 7073 7324 7074
rect 7237 7064 7324 7073
rect 7237 7044 7295 7064
rect 7315 7044 7324 7064
rect 7237 7034 7324 7044
rect 7383 7064 7420 7074
rect 7383 7044 7391 7064
rect 7411 7044 7420 7064
rect 8960 7061 8969 7079
rect 8987 7061 9005 7079
rect 8960 7055 9005 7061
rect 9301 7056 9332 7107
rect 9367 7136 9404 7206
rect 9670 7205 9707 7206
rect 9940 7195 9949 7215
rect 9969 7195 9978 7215
rect 9940 7187 9978 7195
rect 10044 7219 10129 7225
rect 10159 7224 10196 7225
rect 10044 7199 10052 7219
rect 10072 7199 10129 7219
rect 10044 7191 10129 7199
rect 10158 7215 10196 7224
rect 10158 7195 10167 7215
rect 10187 7195 10196 7215
rect 10044 7190 10080 7191
rect 10158 7187 10196 7195
rect 10262 7219 10406 7225
rect 10262 7199 10270 7219
rect 10290 7216 10378 7219
rect 10290 7199 10325 7216
rect 10262 7198 10325 7199
rect 10344 7199 10378 7216
rect 10398 7199 10406 7219
rect 10344 7198 10406 7199
rect 10262 7191 10406 7198
rect 10262 7190 10298 7191
rect 10370 7190 10406 7191
rect 10472 7224 10509 7225
rect 10472 7223 10510 7224
rect 10532 7223 10559 7227
rect 10472 7221 10559 7223
rect 10472 7215 10536 7221
rect 10472 7195 10481 7215
rect 10501 7201 10536 7215
rect 10556 7201 10559 7221
rect 10501 7196 10559 7201
rect 10501 7195 10536 7196
rect 9941 7158 9978 7187
rect 9942 7156 9978 7158
rect 9519 7146 9555 7147
rect 9367 7116 9376 7136
rect 9396 7116 9404 7136
rect 9367 7106 9404 7116
rect 9463 7136 9611 7146
rect 9711 7143 9807 7145
rect 9463 7116 9472 7136
rect 9492 7116 9582 7136
rect 9602 7116 9611 7136
rect 9463 7107 9611 7116
rect 9669 7136 9807 7143
rect 9669 7116 9678 7136
rect 9698 7116 9807 7136
rect 9942 7134 10133 7156
rect 10159 7155 10196 7187
rect 10472 7183 10536 7195
rect 10576 7157 10603 7335
rect 10435 7155 10603 7157
rect 10159 7129 10603 7155
rect 9669 7107 9807 7116
rect 9463 7106 9500 7107
rect 8960 7052 8997 7055
rect 9193 7053 9234 7054
rect 7237 7033 7268 7034
rect 6861 6973 7202 6974
rect 7383 6973 7420 7044
rect 9085 7046 9234 7053
rect 8516 7034 8553 7039
rect 6786 6968 7202 6973
rect 6786 6948 6789 6968
rect 6809 6948 7202 6968
rect 7233 6949 7420 6973
rect 8507 7030 8554 7034
rect 8507 7012 8526 7030
rect 8544 7012 8554 7030
rect 9085 7026 9144 7046
rect 9164 7026 9203 7046
rect 9223 7026 9234 7046
rect 9085 7018 9234 7026
rect 9301 7049 9458 7056
rect 9301 7029 9421 7049
rect 9441 7029 9458 7049
rect 9301 7019 9458 7029
rect 9301 7018 9336 7019
rect 8507 6964 8554 7012
rect 9301 6997 9332 7018
rect 9519 6997 9555 7107
rect 9574 7106 9611 7107
rect 9670 7106 9707 7107
rect 9630 7047 9720 7053
rect 9630 7027 9639 7047
rect 9659 7045 9720 7047
rect 9659 7027 9684 7045
rect 9630 7025 9684 7027
rect 9704 7025 9720 7045
rect 9630 7019 9720 7025
rect 9144 6996 9181 6997
rect 8131 6961 8554 6964
rect 7006 6947 7071 6948
rect 8109 6931 8554 6961
rect 8956 6988 8994 6990
rect 8956 6980 8999 6988
rect 8956 6962 8967 6980
rect 8985 6962 8999 6980
rect 8956 6935 8999 6962
rect 9143 6987 9181 6996
rect 9143 6967 9152 6987
rect 9172 6967 9181 6987
rect 9143 6959 9181 6967
rect 9247 6991 9332 6997
rect 9362 6996 9399 6997
rect 9247 6971 9255 6991
rect 9275 6971 9332 6991
rect 9247 6963 9332 6971
rect 9361 6987 9399 6996
rect 9361 6967 9370 6987
rect 9390 6967 9399 6987
rect 9247 6962 9283 6963
rect 9361 6959 9399 6967
rect 9465 6995 9609 6997
rect 9465 6991 9517 6995
rect 9465 6971 9473 6991
rect 9493 6975 9517 6991
rect 9537 6991 9609 6995
rect 9537 6975 9581 6991
rect 9493 6971 9581 6975
rect 9601 6971 9609 6991
rect 9465 6963 9609 6971
rect 9465 6962 9501 6963
rect 9573 6962 9609 6963
rect 9675 6996 9712 6997
rect 9675 6995 9713 6996
rect 9675 6987 9739 6995
rect 9675 6967 9684 6987
rect 9704 6973 9739 6987
rect 9759 6973 9762 6993
rect 9704 6968 9762 6973
rect 9704 6967 9739 6968
rect 7202 6915 7242 6923
rect 7202 6893 7210 6915
rect 7234 6893 7242 6915
rect 6807 6664 6844 6670
rect 6807 6645 6815 6664
rect 6836 6645 6844 6664
rect 6807 6637 6844 6645
rect 6811 6304 6844 6637
rect 6908 6669 7076 6670
rect 7202 6669 7242 6893
rect 7705 6897 7873 6898
rect 8109 6897 8150 6931
rect 8507 6910 8554 6931
rect 7705 6887 8150 6897
rect 8222 6895 8365 6896
rect 7705 6871 8149 6887
rect 7705 6869 7873 6871
rect 8069 6870 8149 6871
rect 8222 6870 8367 6895
rect 8509 6870 8554 6910
rect 7705 6691 7732 6869
rect 7772 6831 7836 6843
rect 8112 6839 8149 6870
rect 8330 6839 8367 6870
rect 8512 6863 8554 6870
rect 8957 6928 8999 6935
rect 9144 6928 9181 6959
rect 9362 6928 9399 6959
rect 9675 6955 9739 6967
rect 9779 6929 9806 7107
rect 8957 6888 9002 6928
rect 9144 6903 9289 6928
rect 9362 6927 9442 6928
rect 9638 6927 9806 6929
rect 9362 6911 9806 6927
rect 9146 6902 9289 6903
rect 9361 6901 9806 6911
rect 8957 6867 9004 6888
rect 9361 6867 9402 6901
rect 9638 6900 9806 6901
rect 10269 6905 10309 7129
rect 10435 7128 10603 7129
rect 10667 7161 10700 7494
rect 11305 7493 11332 7671
rect 11372 7633 11436 7645
rect 11712 7641 11749 7673
rect 11775 7672 11966 7694
rect 12101 7692 12210 7712
rect 12230 7692 12239 7712
rect 12101 7685 12239 7692
rect 12297 7712 12445 7721
rect 12297 7692 12306 7712
rect 12326 7692 12416 7712
rect 12436 7692 12445 7712
rect 12101 7683 12197 7685
rect 12297 7682 12445 7692
rect 12504 7712 12541 7722
rect 12504 7692 12512 7712
rect 12532 7692 12541 7712
rect 12353 7681 12389 7682
rect 11930 7670 11966 7672
rect 11930 7641 11967 7670
rect 11372 7632 11407 7633
rect 11349 7627 11407 7632
rect 11349 7607 11352 7627
rect 11372 7613 11407 7627
rect 11427 7613 11436 7633
rect 11372 7605 11436 7613
rect 11398 7604 11436 7605
rect 11399 7603 11436 7604
rect 11502 7637 11538 7638
rect 11610 7637 11646 7638
rect 11502 7629 11646 7637
rect 11502 7609 11510 7629
rect 11530 7628 11618 7629
rect 11530 7609 11565 7628
rect 11586 7609 11618 7628
rect 11638 7609 11646 7629
rect 11502 7603 11646 7609
rect 11712 7633 11750 7641
rect 11828 7637 11864 7638
rect 11712 7613 11721 7633
rect 11741 7613 11750 7633
rect 11712 7604 11750 7613
rect 11779 7629 11864 7637
rect 11779 7609 11836 7629
rect 11856 7609 11864 7629
rect 11712 7603 11749 7604
rect 11779 7603 11864 7609
rect 11930 7633 11968 7641
rect 11930 7613 11939 7633
rect 11959 7613 11968 7633
rect 12201 7622 12238 7623
rect 12504 7622 12541 7692
rect 12576 7721 12607 7772
rect 12903 7767 12948 7773
rect 12903 7749 12921 7767
rect 12939 7749 12948 7767
rect 14409 7767 14418 7787
rect 14438 7767 14446 7787
rect 14409 7757 14446 7767
rect 14505 7787 14592 7797
rect 14505 7767 14514 7787
rect 14534 7767 14592 7787
rect 14505 7758 14592 7767
rect 14505 7757 14542 7758
rect 12903 7739 12948 7749
rect 12626 7721 12663 7722
rect 12576 7712 12663 7721
rect 12576 7692 12634 7712
rect 12654 7692 12663 7712
rect 12576 7682 12663 7692
rect 12722 7712 12759 7722
rect 12722 7692 12730 7712
rect 12750 7692 12759 7712
rect 12903 7697 12946 7739
rect 13330 7728 13382 7730
rect 12809 7695 12946 7697
rect 12576 7681 12607 7682
rect 12722 7622 12759 7692
rect 12200 7621 12541 7622
rect 11930 7604 11968 7613
rect 12125 7616 12541 7621
rect 11930 7603 11967 7604
rect 11391 7575 11481 7581
rect 11391 7555 11407 7575
rect 11427 7573 11481 7575
rect 11427 7555 11452 7573
rect 11391 7553 11452 7555
rect 11472 7553 11481 7573
rect 11391 7547 11481 7553
rect 11404 7493 11441 7494
rect 11500 7493 11537 7494
rect 11556 7493 11592 7603
rect 11779 7582 11810 7603
rect 12125 7596 12128 7616
rect 12148 7596 12541 7616
rect 12725 7606 12759 7622
rect 12803 7674 12946 7695
rect 13328 7724 13761 7728
rect 13328 7718 13767 7724
rect 13328 7700 13349 7718
rect 13367 7700 13767 7718
rect 14561 7707 14592 7758
rect 14627 7787 14664 7857
rect 14930 7856 14967 7857
rect 14779 7797 14815 7798
rect 14627 7767 14636 7787
rect 14656 7767 14664 7787
rect 14627 7757 14664 7767
rect 14723 7787 14871 7797
rect 14971 7794 15067 7796
rect 14723 7767 14732 7787
rect 14752 7767 14842 7787
rect 14862 7767 14871 7787
rect 14723 7758 14871 7767
rect 14929 7787 15067 7794
rect 14929 7767 14938 7787
rect 14958 7767 15067 7787
rect 14929 7758 15067 7767
rect 14723 7757 14760 7758
rect 14453 7704 14494 7705
rect 13328 7682 13767 7700
rect 12501 7587 12541 7596
rect 12803 7587 12830 7674
rect 12903 7648 12946 7674
rect 12903 7630 12916 7648
rect 12934 7630 12946 7648
rect 12903 7619 12946 7630
rect 11775 7581 11810 7582
rect 11653 7571 11810 7581
rect 11653 7551 11670 7571
rect 11690 7551 11810 7571
rect 11653 7544 11810 7551
rect 11877 7574 12026 7582
rect 11877 7554 11888 7574
rect 11908 7554 11947 7574
rect 11967 7554 12026 7574
rect 12501 7570 12830 7587
rect 12501 7569 12541 7570
rect 11877 7547 12026 7554
rect 12898 7558 12938 7561
rect 12898 7552 12941 7558
rect 12523 7549 12941 7552
rect 11877 7546 11918 7547
rect 11611 7493 11648 7494
rect 11304 7484 11442 7493
rect 11167 7474 11203 7480
rect 11167 7456 11172 7474
rect 11194 7456 11203 7474
rect 11167 7452 11203 7456
rect 11304 7464 11413 7484
rect 11433 7464 11442 7484
rect 11304 7457 11442 7464
rect 11500 7484 11648 7493
rect 11500 7464 11509 7484
rect 11529 7464 11619 7484
rect 11639 7464 11648 7484
rect 11304 7455 11400 7457
rect 11500 7454 11648 7464
rect 11707 7484 11744 7494
rect 11707 7464 11715 7484
rect 11735 7464 11744 7484
rect 11556 7453 11592 7454
rect 11170 7293 11203 7452
rect 11404 7394 11441 7395
rect 11707 7394 11744 7464
rect 11779 7493 11810 7544
rect 12523 7531 12914 7549
rect 12932 7531 12941 7549
rect 12523 7529 12941 7531
rect 12523 7521 12550 7529
rect 12791 7526 12941 7529
rect 12103 7515 12271 7516
rect 12522 7515 12550 7521
rect 12103 7499 12550 7515
rect 12898 7521 12941 7526
rect 11829 7493 11866 7494
rect 11779 7484 11866 7493
rect 11779 7464 11837 7484
rect 11857 7464 11866 7484
rect 11779 7454 11866 7464
rect 11925 7484 11962 7494
rect 11925 7464 11933 7484
rect 11953 7464 11962 7484
rect 11779 7453 11810 7454
rect 11403 7393 11744 7394
rect 11925 7393 11962 7464
rect 11328 7388 11744 7393
rect 11328 7368 11331 7388
rect 11351 7368 11744 7388
rect 11775 7369 11962 7393
rect 12103 7489 12547 7499
rect 12103 7487 12271 7489
rect 12103 7309 12130 7487
rect 12170 7449 12234 7461
rect 12510 7457 12547 7489
rect 12573 7488 12764 7510
rect 12728 7486 12764 7488
rect 12728 7457 12765 7486
rect 12898 7465 12938 7521
rect 12170 7448 12205 7449
rect 12147 7443 12205 7448
rect 12147 7423 12150 7443
rect 12170 7429 12205 7443
rect 12225 7429 12234 7449
rect 12170 7421 12234 7429
rect 12196 7420 12234 7421
rect 12197 7419 12234 7420
rect 12300 7453 12336 7454
rect 12408 7453 12444 7454
rect 12300 7445 12444 7453
rect 12300 7425 12308 7445
rect 12328 7425 12363 7445
rect 12383 7425 12416 7445
rect 12436 7425 12444 7445
rect 12300 7419 12444 7425
rect 12510 7449 12548 7457
rect 12626 7453 12662 7454
rect 12510 7429 12519 7449
rect 12539 7429 12548 7449
rect 12510 7420 12548 7429
rect 12577 7445 12662 7453
rect 12577 7425 12634 7445
rect 12654 7425 12662 7445
rect 12510 7419 12547 7420
rect 12577 7419 12662 7425
rect 12728 7449 12766 7457
rect 12728 7429 12737 7449
rect 12757 7429 12766 7449
rect 12898 7447 12910 7465
rect 12928 7447 12938 7465
rect 13330 7493 13382 7682
rect 13728 7657 13767 7682
rect 14345 7697 14494 7704
rect 14345 7677 14404 7697
rect 14424 7677 14463 7697
rect 14483 7677 14494 7697
rect 14345 7669 14494 7677
rect 14561 7700 14718 7707
rect 14561 7680 14681 7700
rect 14701 7680 14718 7700
rect 14561 7670 14718 7680
rect 14561 7669 14596 7670
rect 13512 7632 13699 7656
rect 13728 7637 14123 7657
rect 14143 7637 14146 7657
rect 14561 7648 14592 7669
rect 14779 7648 14815 7758
rect 14834 7757 14871 7758
rect 14930 7757 14967 7758
rect 14890 7698 14980 7704
rect 14890 7678 14899 7698
rect 14919 7696 14980 7698
rect 14919 7678 14944 7696
rect 14890 7676 14944 7678
rect 14964 7676 14980 7696
rect 14890 7670 14980 7676
rect 14404 7647 14441 7648
rect 13728 7632 14146 7637
rect 14403 7638 14441 7647
rect 13512 7561 13549 7632
rect 13728 7631 14071 7632
rect 13728 7628 13767 7631
rect 14033 7630 14070 7631
rect 13664 7571 13695 7572
rect 13512 7541 13521 7561
rect 13541 7541 13549 7561
rect 13512 7531 13549 7541
rect 13608 7561 13695 7571
rect 13608 7541 13617 7561
rect 13637 7541 13695 7561
rect 13608 7532 13695 7541
rect 13608 7531 13645 7532
rect 13330 7475 13346 7493
rect 13364 7475 13382 7493
rect 13664 7481 13695 7532
rect 13730 7561 13767 7628
rect 14403 7618 14412 7638
rect 14432 7618 14441 7638
rect 14403 7610 14441 7618
rect 14507 7642 14592 7648
rect 14622 7647 14659 7648
rect 14507 7622 14515 7642
rect 14535 7622 14592 7642
rect 14507 7614 14592 7622
rect 14621 7638 14659 7647
rect 14621 7618 14630 7638
rect 14650 7618 14659 7638
rect 14507 7613 14543 7614
rect 14621 7610 14659 7618
rect 14725 7643 14869 7648
rect 14725 7642 14787 7643
rect 14725 7622 14733 7642
rect 14753 7624 14787 7642
rect 14808 7642 14869 7643
rect 14808 7624 14841 7642
rect 14753 7622 14841 7624
rect 14861 7622 14869 7642
rect 14725 7614 14869 7622
rect 14725 7613 14761 7614
rect 14833 7613 14869 7614
rect 14935 7647 14972 7648
rect 14935 7646 14973 7647
rect 14935 7638 14999 7646
rect 14935 7618 14944 7638
rect 14964 7624 14999 7638
rect 15019 7624 15022 7644
rect 14964 7619 15022 7624
rect 14964 7618 14999 7619
rect 14404 7581 14441 7610
rect 14405 7579 14441 7581
rect 13882 7571 13918 7572
rect 13730 7541 13739 7561
rect 13759 7541 13767 7561
rect 13730 7531 13767 7541
rect 13826 7561 13974 7571
rect 14074 7568 14170 7570
rect 13826 7541 13835 7561
rect 13855 7541 13945 7561
rect 13965 7541 13974 7561
rect 13826 7532 13974 7541
rect 14032 7561 14170 7568
rect 14032 7541 14041 7561
rect 14061 7541 14170 7561
rect 14405 7557 14596 7579
rect 14622 7578 14659 7610
rect 14935 7606 14999 7618
rect 15039 7580 15066 7758
rect 14898 7578 15066 7580
rect 14622 7564 15066 7578
rect 15669 7712 15837 7713
rect 15963 7712 16003 7936
rect 16466 7940 16634 7941
rect 16869 7940 16909 7973
rect 17265 7940 17312 7973
rect 17604 7993 17641 7995
rect 17604 7985 17646 7993
rect 17604 7967 17614 7985
rect 17632 7967 17646 7985
rect 17604 7958 17646 7967
rect 17790 7992 17828 8001
rect 17790 7972 17799 7992
rect 17819 7972 17828 7992
rect 17790 7964 17828 7972
rect 17894 7996 17979 8002
rect 18009 8001 18046 8002
rect 17894 7976 17902 7996
rect 17922 7976 17979 7996
rect 17894 7968 17979 7976
rect 18008 7992 18046 8001
rect 18008 7972 18017 7992
rect 18037 7972 18046 7992
rect 17894 7967 17930 7968
rect 18008 7964 18046 7972
rect 18112 8000 18256 8002
rect 18112 7996 18164 8000
rect 18112 7976 18120 7996
rect 18140 7980 18164 7996
rect 18184 7996 18256 8000
rect 18184 7980 18228 7996
rect 18140 7976 18228 7980
rect 18248 7976 18256 7996
rect 18112 7968 18256 7976
rect 18112 7967 18148 7968
rect 18220 7967 18256 7968
rect 18322 8001 18359 8002
rect 18322 8000 18360 8001
rect 18322 7992 18386 8000
rect 18322 7972 18331 7992
rect 18351 7978 18386 7992
rect 18406 7978 18409 7998
rect 18351 7973 18409 7978
rect 18351 7972 18386 7973
rect 16466 7939 16910 7940
rect 16466 7914 16911 7939
rect 16466 7912 16634 7914
rect 16830 7913 16911 7914
rect 17080 7913 17129 7939
rect 17265 7913 17314 7940
rect 16466 7734 16493 7912
rect 16533 7874 16597 7886
rect 16873 7882 16910 7913
rect 17091 7882 17128 7913
rect 17273 7888 17314 7913
rect 17605 7933 17646 7958
rect 17791 7933 17828 7964
rect 18009 7933 18046 7964
rect 18322 7960 18386 7972
rect 18426 7934 18453 8112
rect 17605 7906 17654 7933
rect 17790 7907 17839 7933
rect 18008 7932 18089 7933
rect 18285 7932 18453 7934
rect 18008 7907 18453 7932
rect 18009 7906 18453 7907
rect 16533 7873 16568 7874
rect 16510 7868 16568 7873
rect 16510 7848 16513 7868
rect 16533 7854 16568 7868
rect 16588 7854 16597 7874
rect 16533 7846 16597 7854
rect 16559 7845 16597 7846
rect 16560 7844 16597 7845
rect 16663 7878 16699 7879
rect 16771 7878 16807 7879
rect 16663 7870 16807 7878
rect 16663 7850 16671 7870
rect 16691 7866 16779 7870
rect 16691 7850 16735 7866
rect 16663 7846 16735 7850
rect 16755 7850 16779 7866
rect 16799 7850 16807 7870
rect 16755 7846 16807 7850
rect 16663 7844 16807 7846
rect 16873 7874 16911 7882
rect 16989 7878 17025 7879
rect 16873 7854 16882 7874
rect 16902 7854 16911 7874
rect 16873 7845 16911 7854
rect 16940 7870 17025 7878
rect 16940 7850 16997 7870
rect 17017 7850 17025 7870
rect 16873 7844 16910 7845
rect 16940 7844 17025 7850
rect 17091 7874 17129 7882
rect 17091 7854 17100 7874
rect 17120 7854 17129 7874
rect 17091 7845 17129 7854
rect 17273 7879 17315 7888
rect 17273 7861 17287 7879
rect 17305 7861 17315 7879
rect 17273 7853 17315 7861
rect 17278 7851 17315 7853
rect 17607 7873 17654 7906
rect 18010 7873 18050 7906
rect 18285 7905 18453 7906
rect 18916 7910 18956 8134
rect 19082 8133 19250 8134
rect 19853 8268 20297 8282
rect 19853 8266 20021 8268
rect 19853 8088 19880 8266
rect 19920 8228 19984 8240
rect 20260 8236 20297 8268
rect 20323 8267 20514 8289
rect 20749 8285 20858 8305
rect 20878 8285 20887 8305
rect 20749 8278 20887 8285
rect 20945 8305 21093 8314
rect 20945 8285 20954 8305
rect 20974 8285 21064 8305
rect 21084 8285 21093 8305
rect 20749 8276 20845 8278
rect 20945 8275 21093 8285
rect 21152 8305 21189 8315
rect 21152 8285 21160 8305
rect 21180 8285 21189 8305
rect 21001 8274 21037 8275
rect 20478 8265 20514 8267
rect 20478 8236 20515 8265
rect 19920 8227 19955 8228
rect 19897 8222 19955 8227
rect 19897 8202 19900 8222
rect 19920 8208 19955 8222
rect 19975 8208 19984 8228
rect 19920 8200 19984 8208
rect 19946 8199 19984 8200
rect 19947 8198 19984 8199
rect 20050 8232 20086 8233
rect 20158 8232 20194 8233
rect 20050 8226 20194 8232
rect 20050 8224 20111 8226
rect 20050 8204 20058 8224
rect 20078 8209 20111 8224
rect 20130 8224 20194 8226
rect 20130 8209 20166 8224
rect 20078 8204 20166 8209
rect 20186 8204 20194 8224
rect 20050 8198 20194 8204
rect 20260 8228 20298 8236
rect 20376 8232 20412 8233
rect 20260 8208 20269 8228
rect 20289 8208 20298 8228
rect 20260 8199 20298 8208
rect 20327 8224 20412 8232
rect 20327 8204 20384 8224
rect 20404 8204 20412 8224
rect 20260 8198 20297 8199
rect 20327 8198 20412 8204
rect 20478 8228 20516 8236
rect 20478 8208 20487 8228
rect 20507 8208 20516 8228
rect 21152 8218 21189 8285
rect 21224 8314 21255 8365
rect 21537 8353 21555 8371
rect 21573 8353 21589 8371
rect 21274 8314 21311 8315
rect 21224 8305 21311 8314
rect 21224 8285 21282 8305
rect 21302 8285 21311 8305
rect 21224 8275 21311 8285
rect 21370 8305 21407 8315
rect 21370 8285 21378 8305
rect 21398 8285 21407 8305
rect 21224 8274 21255 8275
rect 20849 8215 20886 8216
rect 21152 8215 21191 8218
rect 20848 8214 21191 8215
rect 21370 8214 21407 8285
rect 20478 8199 20516 8208
rect 20773 8209 21191 8214
rect 20478 8198 20515 8199
rect 19939 8170 20029 8176
rect 19939 8150 19955 8170
rect 19975 8168 20029 8170
rect 19975 8150 20000 8168
rect 19939 8148 20000 8150
rect 20020 8148 20029 8168
rect 19939 8142 20029 8148
rect 19952 8088 19989 8089
rect 20048 8088 20085 8089
rect 20104 8088 20140 8198
rect 20327 8177 20358 8198
rect 20773 8189 20776 8209
rect 20796 8189 21191 8209
rect 21220 8190 21407 8214
rect 20323 8176 20358 8177
rect 20201 8166 20358 8176
rect 20201 8146 20218 8166
rect 20238 8146 20358 8166
rect 20201 8139 20358 8146
rect 20425 8169 20574 8177
rect 20425 8149 20436 8169
rect 20456 8149 20495 8169
rect 20515 8149 20574 8169
rect 20425 8142 20574 8149
rect 21152 8164 21191 8189
rect 21537 8164 21589 8353
rect 21981 8381 21991 8399
rect 22009 8381 22021 8399
rect 22153 8397 22162 8417
rect 22182 8397 22191 8417
rect 22153 8389 22191 8397
rect 22257 8421 22342 8427
rect 22372 8426 22409 8427
rect 22257 8401 22265 8421
rect 22285 8401 22342 8421
rect 22257 8393 22342 8401
rect 22371 8417 22409 8426
rect 22371 8397 22380 8417
rect 22400 8397 22409 8417
rect 22257 8392 22293 8393
rect 22371 8389 22409 8397
rect 22475 8421 22619 8427
rect 22475 8401 22483 8421
rect 22503 8401 22536 8421
rect 22556 8401 22591 8421
rect 22611 8401 22619 8421
rect 22475 8393 22619 8401
rect 22475 8392 22511 8393
rect 22583 8392 22619 8393
rect 22685 8426 22722 8427
rect 22685 8425 22723 8426
rect 22685 8417 22749 8425
rect 22685 8397 22694 8417
rect 22714 8403 22749 8417
rect 22769 8403 22772 8423
rect 22714 8398 22772 8403
rect 22714 8397 22749 8398
rect 21981 8325 22021 8381
rect 22154 8360 22191 8389
rect 22155 8358 22191 8360
rect 22155 8336 22346 8358
rect 22372 8357 22409 8389
rect 22685 8385 22749 8397
rect 22789 8359 22816 8537
rect 22648 8357 22816 8359
rect 22372 8347 22816 8357
rect 22957 8453 23144 8477
rect 23175 8458 23568 8478
rect 23588 8458 23591 8478
rect 23175 8453 23591 8458
rect 22957 8382 22994 8453
rect 23175 8452 23516 8453
rect 23109 8392 23140 8393
rect 22957 8362 22966 8382
rect 22986 8362 22994 8382
rect 22957 8352 22994 8362
rect 23053 8382 23140 8392
rect 23053 8362 23062 8382
rect 23082 8362 23140 8382
rect 23053 8353 23140 8362
rect 23053 8352 23090 8353
rect 21978 8320 22021 8325
rect 22369 8331 22816 8347
rect 22369 8325 22397 8331
rect 22648 8330 22816 8331
rect 21978 8317 22128 8320
rect 22369 8317 22396 8325
rect 21978 8315 22396 8317
rect 21978 8297 21987 8315
rect 22005 8297 22396 8315
rect 23109 8302 23140 8353
rect 23175 8382 23212 8452
rect 23478 8451 23515 8452
rect 23327 8392 23363 8393
rect 23175 8362 23184 8382
rect 23204 8362 23212 8382
rect 23175 8352 23212 8362
rect 23271 8382 23419 8392
rect 23519 8389 23615 8391
rect 23271 8362 23280 8382
rect 23300 8362 23390 8382
rect 23410 8362 23419 8382
rect 23271 8353 23419 8362
rect 23477 8382 23615 8389
rect 23477 8362 23486 8382
rect 23506 8362 23615 8382
rect 23477 8353 23615 8362
rect 23271 8352 23308 8353
rect 23001 8299 23042 8300
rect 21978 8294 22396 8297
rect 21978 8288 22021 8294
rect 21981 8285 22021 8288
rect 22893 8292 23042 8299
rect 22378 8276 22418 8277
rect 22089 8259 22418 8276
rect 22893 8272 22952 8292
rect 22972 8272 23011 8292
rect 23031 8272 23042 8292
rect 22893 8264 23042 8272
rect 23109 8295 23266 8302
rect 23109 8275 23229 8295
rect 23249 8275 23266 8295
rect 23109 8265 23266 8275
rect 23109 8264 23144 8265
rect 21973 8216 22016 8227
rect 21973 8198 21985 8216
rect 22003 8198 22016 8216
rect 21973 8172 22016 8198
rect 22089 8172 22116 8259
rect 22378 8250 22418 8259
rect 21152 8146 21591 8164
rect 20425 8141 20466 8142
rect 20159 8088 20196 8089
rect 19852 8079 19990 8088
rect 19852 8059 19961 8079
rect 19981 8059 19990 8079
rect 19852 8052 19990 8059
rect 20048 8079 20196 8088
rect 20048 8059 20057 8079
rect 20077 8059 20167 8079
rect 20187 8059 20196 8079
rect 19852 8050 19948 8052
rect 20048 8049 20196 8059
rect 20255 8079 20292 8089
rect 20255 8059 20263 8079
rect 20283 8059 20292 8079
rect 20104 8048 20140 8049
rect 19952 7989 19989 7990
rect 20255 7989 20292 8059
rect 20327 8088 20358 8139
rect 21152 8128 21552 8146
rect 21570 8128 21591 8146
rect 21152 8122 21591 8128
rect 21158 8118 21591 8122
rect 21973 8151 22116 8172
rect 22160 8224 22194 8240
rect 22378 8230 22771 8250
rect 22791 8230 22794 8250
rect 23109 8243 23140 8264
rect 23327 8243 23363 8353
rect 23382 8352 23419 8353
rect 23478 8352 23515 8353
rect 23438 8293 23528 8299
rect 23438 8273 23447 8293
rect 23467 8291 23528 8293
rect 23467 8273 23492 8291
rect 23438 8271 23492 8273
rect 23512 8271 23528 8291
rect 23438 8265 23528 8271
rect 22952 8242 22989 8243
rect 22378 8225 22794 8230
rect 22951 8233 22989 8242
rect 22378 8224 22719 8225
rect 22160 8154 22197 8224
rect 22312 8164 22343 8165
rect 21973 8149 22110 8151
rect 21537 8116 21589 8118
rect 21973 8107 22016 8149
rect 22160 8134 22169 8154
rect 22189 8134 22197 8154
rect 22160 8124 22197 8134
rect 22256 8154 22343 8164
rect 22256 8134 22265 8154
rect 22285 8134 22343 8154
rect 22256 8125 22343 8134
rect 22256 8124 22293 8125
rect 21971 8097 22016 8107
rect 20377 8088 20414 8089
rect 20327 8079 20414 8088
rect 20327 8059 20385 8079
rect 20405 8059 20414 8079
rect 20327 8049 20414 8059
rect 20473 8079 20510 8089
rect 20473 8059 20481 8079
rect 20501 8059 20510 8079
rect 21971 8079 21980 8097
rect 21998 8079 22016 8097
rect 21971 8073 22016 8079
rect 22312 8074 22343 8125
rect 22378 8154 22415 8224
rect 22681 8223 22718 8224
rect 22951 8213 22960 8233
rect 22980 8213 22989 8233
rect 22951 8205 22989 8213
rect 23055 8237 23140 8243
rect 23170 8242 23207 8243
rect 23055 8217 23063 8237
rect 23083 8217 23140 8237
rect 23055 8209 23140 8217
rect 23169 8233 23207 8242
rect 23169 8213 23178 8233
rect 23198 8213 23207 8233
rect 23055 8208 23091 8209
rect 23169 8205 23207 8213
rect 23273 8237 23417 8243
rect 23273 8217 23281 8237
rect 23301 8218 23333 8237
rect 23354 8218 23389 8237
rect 23301 8217 23389 8218
rect 23409 8217 23417 8237
rect 23273 8209 23417 8217
rect 23273 8208 23309 8209
rect 23381 8208 23417 8209
rect 23483 8242 23520 8243
rect 23483 8241 23521 8242
rect 23483 8233 23547 8241
rect 23483 8213 23492 8233
rect 23512 8219 23547 8233
rect 23567 8219 23570 8239
rect 23512 8214 23570 8219
rect 23512 8213 23547 8214
rect 22952 8176 22989 8205
rect 22953 8174 22989 8176
rect 22530 8164 22566 8165
rect 22378 8134 22387 8154
rect 22407 8134 22415 8154
rect 22378 8124 22415 8134
rect 22474 8154 22622 8164
rect 22722 8161 22818 8163
rect 22474 8134 22483 8154
rect 22503 8134 22593 8154
rect 22613 8134 22622 8154
rect 22474 8125 22622 8134
rect 22680 8154 22818 8161
rect 22680 8134 22689 8154
rect 22709 8134 22818 8154
rect 22953 8152 23144 8174
rect 23170 8173 23207 8205
rect 23483 8201 23547 8213
rect 23587 8175 23614 8353
rect 24219 8352 24252 8685
rect 24316 8717 24484 8718
rect 24610 8717 24650 8941
rect 25113 8945 25281 8946
rect 25517 8945 25566 8980
rect 25113 8919 25566 8945
rect 25113 8917 25281 8919
rect 25477 8918 25559 8919
rect 25699 8918 25777 8944
rect 25917 8922 25964 8980
rect 26365 8976 26412 8981
rect 25113 8739 25140 8917
rect 25180 8879 25244 8891
rect 25520 8887 25557 8918
rect 25738 8887 25775 8918
rect 25917 8909 25965 8922
rect 25180 8878 25215 8879
rect 25157 8873 25215 8878
rect 25157 8853 25160 8873
rect 25180 8859 25215 8873
rect 25235 8859 25244 8879
rect 25180 8851 25244 8859
rect 25206 8850 25244 8851
rect 25207 8849 25244 8850
rect 25310 8883 25346 8884
rect 25418 8883 25454 8884
rect 25310 8875 25454 8883
rect 25310 8855 25318 8875
rect 25338 8871 25426 8875
rect 25338 8855 25382 8871
rect 25310 8851 25382 8855
rect 25402 8855 25426 8871
rect 25446 8855 25454 8875
rect 25402 8851 25454 8855
rect 25310 8849 25454 8851
rect 25520 8879 25558 8887
rect 25636 8883 25672 8884
rect 25520 8859 25529 8879
rect 25549 8859 25558 8879
rect 25520 8850 25558 8859
rect 25587 8875 25672 8883
rect 25587 8855 25644 8875
rect 25664 8855 25672 8875
rect 25520 8849 25557 8850
rect 25587 8849 25672 8855
rect 25738 8879 25776 8887
rect 25738 8859 25747 8879
rect 25767 8859 25776 8879
rect 25738 8850 25776 8859
rect 25920 8884 25965 8909
rect 25920 8866 25934 8884
rect 25952 8866 25965 8884
rect 25920 8858 25965 8866
rect 25925 8856 25965 8858
rect 26365 8914 26413 8976
rect 28987 8975 29027 8983
rect 28987 8953 28995 8975
rect 29019 8953 29027 8975
rect 29891 8978 30347 9013
rect 33351 8988 33391 8996
rect 25738 8849 25775 8850
rect 25199 8821 25289 8827
rect 25199 8801 25215 8821
rect 25235 8819 25289 8821
rect 25235 8801 25260 8819
rect 25199 8799 25260 8801
rect 25280 8799 25289 8819
rect 25199 8793 25289 8799
rect 25212 8739 25249 8740
rect 25308 8739 25345 8740
rect 25364 8739 25400 8849
rect 25587 8828 25618 8849
rect 26365 8834 26412 8914
rect 25583 8827 25618 8828
rect 25461 8817 25618 8827
rect 25461 8797 25478 8817
rect 25498 8797 25618 8817
rect 25461 8790 25618 8797
rect 25685 8820 25834 8828
rect 25685 8800 25696 8820
rect 25716 8800 25755 8820
rect 25775 8800 25834 8820
rect 26365 8816 26375 8834
rect 26393 8816 26412 8834
rect 26365 8812 26412 8816
rect 26366 8807 26403 8812
rect 25685 8793 25834 8800
rect 25685 8792 25726 8793
rect 25922 8791 25959 8794
rect 25419 8739 25456 8740
rect 25112 8730 25250 8739
rect 24316 8691 24760 8717
rect 24316 8689 24484 8691
rect 24316 8511 24343 8689
rect 24383 8651 24447 8663
rect 24723 8659 24760 8691
rect 24786 8690 24977 8712
rect 25112 8710 25221 8730
rect 25241 8710 25250 8730
rect 25112 8703 25250 8710
rect 25308 8730 25456 8739
rect 25308 8710 25317 8730
rect 25337 8710 25427 8730
rect 25447 8710 25456 8730
rect 25112 8701 25208 8703
rect 25308 8700 25456 8710
rect 25515 8730 25552 8740
rect 25515 8710 25523 8730
rect 25543 8710 25552 8730
rect 25364 8699 25400 8700
rect 24941 8688 24977 8690
rect 24941 8659 24978 8688
rect 24383 8650 24418 8651
rect 24360 8645 24418 8650
rect 24360 8625 24363 8645
rect 24383 8631 24418 8645
rect 24438 8631 24447 8651
rect 24383 8625 24447 8631
rect 24360 8623 24447 8625
rect 24360 8619 24387 8623
rect 24409 8622 24447 8623
rect 24410 8621 24447 8622
rect 24513 8655 24549 8656
rect 24621 8655 24657 8656
rect 24513 8648 24657 8655
rect 24513 8647 24575 8648
rect 24513 8627 24521 8647
rect 24541 8630 24575 8647
rect 24594 8647 24657 8648
rect 24594 8630 24629 8647
rect 24541 8627 24629 8630
rect 24649 8627 24657 8647
rect 24513 8621 24657 8627
rect 24723 8651 24761 8659
rect 24839 8655 24875 8656
rect 24723 8631 24732 8651
rect 24752 8631 24761 8651
rect 24723 8622 24761 8631
rect 24790 8647 24875 8655
rect 24790 8627 24847 8647
rect 24867 8627 24875 8647
rect 24723 8621 24760 8622
rect 24790 8621 24875 8627
rect 24941 8651 24979 8659
rect 24941 8631 24950 8651
rect 24970 8631 24979 8651
rect 25212 8640 25249 8641
rect 25515 8640 25552 8710
rect 25587 8739 25618 8790
rect 25914 8785 25959 8791
rect 25914 8767 25932 8785
rect 25950 8767 25959 8785
rect 25914 8757 25959 8767
rect 25637 8739 25674 8740
rect 25587 8730 25674 8739
rect 25587 8710 25645 8730
rect 25665 8710 25674 8730
rect 25587 8700 25674 8710
rect 25733 8730 25770 8740
rect 25733 8710 25741 8730
rect 25761 8710 25770 8730
rect 25914 8715 25957 8757
rect 26354 8745 26406 8747
rect 25820 8713 25957 8715
rect 25587 8699 25618 8700
rect 25733 8640 25770 8710
rect 25211 8639 25552 8640
rect 24941 8622 24979 8631
rect 25136 8634 25552 8639
rect 24941 8621 24978 8622
rect 24402 8593 24492 8599
rect 24402 8573 24418 8593
rect 24438 8591 24492 8593
rect 24438 8573 24463 8591
rect 24402 8571 24463 8573
rect 24483 8571 24492 8591
rect 24402 8565 24492 8571
rect 24415 8511 24452 8512
rect 24511 8511 24548 8512
rect 24567 8511 24603 8621
rect 24790 8600 24821 8621
rect 25136 8614 25139 8634
rect 25159 8614 25552 8634
rect 25736 8624 25770 8640
rect 25814 8692 25957 8713
rect 26352 8741 26785 8745
rect 26352 8735 26791 8741
rect 26352 8717 26373 8735
rect 26391 8717 26791 8735
rect 26352 8699 26791 8717
rect 25512 8605 25552 8614
rect 25814 8605 25841 8692
rect 25914 8666 25957 8692
rect 25914 8648 25927 8666
rect 25945 8648 25957 8666
rect 25914 8637 25957 8648
rect 24786 8599 24821 8600
rect 24664 8589 24821 8599
rect 24664 8569 24681 8589
rect 24701 8569 24821 8589
rect 24664 8562 24821 8569
rect 24888 8592 25034 8600
rect 24888 8572 24899 8592
rect 24919 8572 24958 8592
rect 24978 8572 25034 8592
rect 25512 8588 25841 8605
rect 25512 8587 25552 8588
rect 24888 8565 25034 8572
rect 25909 8576 25949 8579
rect 25909 8570 25952 8576
rect 25534 8567 25952 8570
rect 24888 8564 24929 8565
rect 24622 8511 24659 8512
rect 24315 8502 24453 8511
rect 24315 8482 24424 8502
rect 24444 8482 24453 8502
rect 24315 8475 24453 8482
rect 24511 8502 24659 8511
rect 24511 8482 24520 8502
rect 24540 8482 24630 8502
rect 24650 8482 24659 8502
rect 24315 8473 24411 8475
rect 24511 8472 24659 8482
rect 24718 8502 24755 8512
rect 24718 8482 24726 8502
rect 24746 8482 24755 8502
rect 24567 8471 24603 8472
rect 24415 8412 24452 8413
rect 24718 8412 24755 8482
rect 24790 8511 24821 8562
rect 25534 8549 25925 8567
rect 25943 8549 25952 8567
rect 25534 8547 25952 8549
rect 25534 8539 25561 8547
rect 25802 8544 25952 8547
rect 25114 8533 25282 8534
rect 25533 8533 25561 8539
rect 25114 8517 25561 8533
rect 25909 8539 25952 8544
rect 24840 8511 24877 8512
rect 24790 8502 24877 8511
rect 24790 8482 24848 8502
rect 24868 8482 24877 8502
rect 24790 8472 24877 8482
rect 24936 8502 24973 8512
rect 24936 8482 24944 8502
rect 24964 8482 24973 8502
rect 24790 8471 24821 8472
rect 24414 8411 24755 8412
rect 24936 8411 24973 8482
rect 24339 8406 24755 8411
rect 24339 8386 24342 8406
rect 24362 8386 24755 8406
rect 24786 8387 24973 8411
rect 25114 8507 25558 8517
rect 25114 8505 25282 8507
rect 24214 8307 24256 8352
rect 25114 8327 25141 8505
rect 25181 8467 25245 8479
rect 25521 8475 25558 8507
rect 25584 8506 25775 8528
rect 25739 8504 25775 8506
rect 25739 8475 25776 8504
rect 25909 8483 25949 8539
rect 25181 8466 25216 8467
rect 25158 8461 25216 8466
rect 25158 8441 25161 8461
rect 25181 8447 25216 8461
rect 25236 8447 25245 8467
rect 25181 8439 25245 8447
rect 25207 8438 25245 8439
rect 25208 8437 25245 8438
rect 25311 8471 25347 8472
rect 25419 8471 25455 8472
rect 25311 8463 25455 8471
rect 25311 8443 25319 8463
rect 25339 8443 25374 8463
rect 25394 8443 25427 8463
rect 25447 8443 25455 8463
rect 25311 8437 25455 8443
rect 25521 8467 25559 8475
rect 25637 8471 25673 8472
rect 25521 8447 25530 8467
rect 25550 8447 25559 8467
rect 25521 8438 25559 8447
rect 25588 8463 25673 8471
rect 25588 8443 25645 8463
rect 25665 8443 25673 8463
rect 25521 8437 25558 8438
rect 25588 8437 25673 8443
rect 25739 8467 25777 8475
rect 25739 8447 25748 8467
rect 25768 8447 25777 8467
rect 25909 8465 25921 8483
rect 25939 8465 25949 8483
rect 26354 8510 26406 8699
rect 26752 8674 26791 8699
rect 28592 8724 28629 8730
rect 28592 8705 28600 8724
rect 28621 8705 28629 8724
rect 28592 8697 28629 8705
rect 26536 8649 26723 8673
rect 26752 8654 27147 8674
rect 27167 8654 27170 8674
rect 26752 8649 27170 8654
rect 26536 8578 26573 8649
rect 26752 8648 27095 8649
rect 26752 8645 26791 8648
rect 27057 8647 27094 8648
rect 26688 8588 26719 8589
rect 26536 8558 26545 8578
rect 26565 8558 26573 8578
rect 26536 8548 26573 8558
rect 26632 8578 26719 8588
rect 26632 8558 26641 8578
rect 26661 8558 26719 8578
rect 26632 8549 26719 8558
rect 26632 8548 26669 8549
rect 26354 8492 26370 8510
rect 26388 8492 26406 8510
rect 26688 8498 26719 8549
rect 26754 8578 26791 8645
rect 26906 8588 26942 8589
rect 26754 8558 26763 8578
rect 26783 8558 26791 8578
rect 26754 8548 26791 8558
rect 26850 8578 26998 8588
rect 27098 8585 27194 8587
rect 26850 8558 26859 8578
rect 26879 8558 26969 8578
rect 26989 8558 26998 8578
rect 26850 8549 26998 8558
rect 27056 8578 27194 8585
rect 27056 8558 27065 8578
rect 27085 8558 27194 8578
rect 27056 8549 27194 8558
rect 26850 8548 26887 8549
rect 26580 8495 26621 8496
rect 26354 8474 26406 8492
rect 26472 8488 26621 8495
rect 25909 8455 25949 8465
rect 26472 8468 26531 8488
rect 26551 8468 26590 8488
rect 26610 8468 26621 8488
rect 26472 8460 26621 8468
rect 26688 8491 26845 8498
rect 26688 8471 26808 8491
rect 26828 8471 26845 8491
rect 26688 8461 26845 8471
rect 26688 8460 26723 8461
rect 25739 8438 25777 8447
rect 26688 8439 26719 8460
rect 26906 8439 26942 8549
rect 26961 8548 26998 8549
rect 27057 8548 27094 8549
rect 27017 8489 27107 8495
rect 27017 8469 27026 8489
rect 27046 8487 27107 8489
rect 27046 8469 27071 8487
rect 27017 8467 27071 8469
rect 27091 8467 27107 8487
rect 27017 8461 27107 8467
rect 26531 8438 26568 8439
rect 25739 8437 25776 8438
rect 25200 8409 25290 8415
rect 25200 8389 25216 8409
rect 25236 8407 25290 8409
rect 25236 8389 25261 8407
rect 25200 8387 25261 8389
rect 25281 8387 25290 8407
rect 25200 8381 25290 8387
rect 25213 8327 25250 8328
rect 25309 8327 25346 8328
rect 25365 8327 25401 8437
rect 25588 8416 25619 8437
rect 26530 8429 26568 8438
rect 25584 8415 25619 8416
rect 25462 8405 25619 8415
rect 25462 8385 25479 8405
rect 25499 8385 25619 8405
rect 25462 8378 25619 8385
rect 25686 8408 25835 8416
rect 25686 8388 25697 8408
rect 25717 8388 25756 8408
rect 25776 8388 25835 8408
rect 26358 8411 26398 8421
rect 25686 8381 25835 8388
rect 25901 8384 25953 8402
rect 25686 8380 25727 8381
rect 25420 8327 25457 8328
rect 25113 8318 25251 8327
rect 24585 8307 24618 8309
rect 24214 8295 24661 8307
rect 23446 8173 23614 8175
rect 23170 8147 23614 8173
rect 22680 8125 22818 8134
rect 22474 8124 22511 8125
rect 21971 8070 22008 8073
rect 22204 8071 22245 8072
rect 20327 8048 20358 8049
rect 19951 7988 20292 7989
rect 20473 7988 20510 8059
rect 22096 8064 22245 8071
rect 21540 8051 21577 8056
rect 21531 8047 21578 8051
rect 21531 8029 21550 8047
rect 21568 8029 21578 8047
rect 22096 8044 22155 8064
rect 22175 8044 22214 8064
rect 22234 8044 22245 8064
rect 22096 8036 22245 8044
rect 22312 8067 22469 8074
rect 22312 8047 22432 8067
rect 22452 8047 22469 8067
rect 22312 8037 22469 8047
rect 22312 8036 22347 8037
rect 19876 7983 20292 7988
rect 19876 7963 19879 7983
rect 19899 7963 20292 7983
rect 20323 7964 20510 7988
rect 21135 7986 21175 7991
rect 21531 7986 21578 8029
rect 22312 8015 22343 8036
rect 22530 8015 22566 8125
rect 22585 8124 22622 8125
rect 22681 8124 22718 8125
rect 22641 8065 22731 8071
rect 22641 8045 22650 8065
rect 22670 8063 22731 8065
rect 22670 8045 22695 8063
rect 22641 8043 22695 8045
rect 22715 8043 22731 8063
rect 22641 8037 22731 8043
rect 22155 8014 22192 8015
rect 21135 7947 21578 7986
rect 21968 8006 22005 8008
rect 21968 7998 22010 8006
rect 21968 7980 21978 7998
rect 21996 7980 22010 7998
rect 21968 7971 22010 7980
rect 22154 8005 22192 8014
rect 22154 7985 22163 8005
rect 22183 7985 22192 8005
rect 22154 7977 22192 7985
rect 22258 8009 22343 8015
rect 22373 8014 22410 8015
rect 22258 7989 22266 8009
rect 22286 7989 22343 8009
rect 22258 7981 22343 7989
rect 22372 8005 22410 8014
rect 22372 7985 22381 8005
rect 22401 7985 22410 8005
rect 22258 7980 22294 7981
rect 22372 7977 22410 7985
rect 22476 8013 22620 8015
rect 22476 8009 22528 8013
rect 22476 7989 22484 8009
rect 22504 7993 22528 8009
rect 22548 8009 22620 8013
rect 22548 7993 22592 8009
rect 22504 7989 22592 7993
rect 22612 7989 22620 8009
rect 22476 7981 22620 7989
rect 22476 7980 22512 7981
rect 22584 7980 22620 7981
rect 22686 8014 22723 8015
rect 22686 8013 22724 8014
rect 22686 8005 22750 8013
rect 22686 7985 22695 8005
rect 22715 7991 22750 8005
rect 22770 7991 22773 8011
rect 22715 7986 22773 7991
rect 22715 7985 22750 7986
rect 18916 7888 18924 7910
rect 18948 7888 18956 7910
rect 18916 7880 18956 7888
rect 20229 7932 20269 7940
rect 20229 7910 20237 7932
rect 20261 7910 20269 7932
rect 17091 7844 17128 7845
rect 16552 7816 16642 7822
rect 16552 7796 16568 7816
rect 16588 7814 16642 7816
rect 16588 7796 16613 7814
rect 16552 7794 16613 7796
rect 16633 7794 16642 7814
rect 16552 7788 16642 7794
rect 16565 7734 16602 7735
rect 16661 7734 16698 7735
rect 16717 7734 16753 7844
rect 16940 7823 16971 7844
rect 17607 7834 18050 7873
rect 16936 7822 16971 7823
rect 16814 7812 16971 7822
rect 16814 7792 16831 7812
rect 16851 7792 16971 7812
rect 16814 7785 16971 7792
rect 17038 7815 17187 7823
rect 17038 7795 17049 7815
rect 17069 7795 17108 7815
rect 17128 7795 17187 7815
rect 17038 7788 17187 7795
rect 17607 7791 17654 7834
rect 18010 7829 18050 7834
rect 18675 7832 18862 7856
rect 18893 7837 19286 7857
rect 19306 7837 19309 7857
rect 18893 7832 19309 7837
rect 17038 7787 17079 7788
rect 17275 7786 17312 7789
rect 16772 7734 16809 7735
rect 16465 7725 16603 7734
rect 15669 7686 16113 7712
rect 15669 7684 15837 7686
rect 14622 7552 15069 7564
rect 14665 7550 14698 7552
rect 14032 7532 14170 7541
rect 13826 7531 13863 7532
rect 13556 7478 13597 7479
rect 13330 7457 13382 7475
rect 13448 7471 13597 7478
rect 12898 7437 12938 7447
rect 13448 7451 13507 7471
rect 13527 7451 13566 7471
rect 13586 7451 13597 7471
rect 13448 7443 13597 7451
rect 13664 7474 13821 7481
rect 13664 7454 13784 7474
rect 13804 7454 13821 7474
rect 13664 7444 13821 7454
rect 13664 7443 13699 7444
rect 12728 7420 12766 7429
rect 13664 7422 13695 7443
rect 13882 7422 13918 7532
rect 13937 7531 13974 7532
rect 14033 7531 14070 7532
rect 13993 7472 14083 7478
rect 13993 7452 14002 7472
rect 14022 7470 14083 7472
rect 14022 7452 14047 7470
rect 13993 7450 14047 7452
rect 14067 7450 14083 7470
rect 13993 7444 14083 7450
rect 13507 7421 13544 7422
rect 12728 7419 12765 7420
rect 12189 7391 12279 7397
rect 12189 7371 12205 7391
rect 12225 7389 12279 7391
rect 12225 7371 12250 7389
rect 12189 7369 12250 7371
rect 12270 7369 12279 7389
rect 12189 7363 12279 7369
rect 12202 7309 12239 7310
rect 12298 7309 12335 7310
rect 12354 7309 12390 7419
rect 12577 7398 12608 7419
rect 13506 7412 13544 7421
rect 12573 7397 12608 7398
rect 12451 7387 12608 7397
rect 12451 7367 12468 7387
rect 12488 7367 12608 7387
rect 12451 7360 12608 7367
rect 12675 7390 12824 7398
rect 12675 7370 12686 7390
rect 12706 7370 12745 7390
rect 12765 7370 12824 7390
rect 13334 7394 13374 7404
rect 12675 7363 12824 7370
rect 12890 7366 12942 7384
rect 12675 7362 12716 7363
rect 12409 7309 12446 7310
rect 12102 7300 12240 7309
rect 11169 7292 11206 7293
rect 11140 7291 11308 7292
rect 11434 7291 11474 7293
rect 10965 7282 11004 7288
rect 10965 7260 10973 7282
rect 10997 7260 11004 7282
rect 10667 7153 10704 7161
rect 10667 7134 10675 7153
rect 10696 7134 10704 7153
rect 10667 7128 10704 7134
rect 10269 6883 10277 6905
rect 10301 6883 10309 6905
rect 10269 6875 10309 6883
rect 7772 6830 7807 6831
rect 7749 6825 7807 6830
rect 7749 6805 7752 6825
rect 7772 6811 7807 6825
rect 7827 6811 7836 6831
rect 7772 6803 7836 6811
rect 7798 6802 7836 6803
rect 7799 6801 7836 6802
rect 7902 6835 7938 6836
rect 8010 6835 8046 6836
rect 7902 6827 8046 6835
rect 7902 6807 7910 6827
rect 7930 6823 8018 6827
rect 7930 6807 7974 6823
rect 7902 6803 7974 6807
rect 7994 6807 8018 6823
rect 8038 6807 8046 6827
rect 7994 6803 8046 6807
rect 7902 6801 8046 6803
rect 8112 6831 8150 6839
rect 8228 6835 8264 6836
rect 8112 6811 8121 6831
rect 8141 6811 8150 6831
rect 8112 6802 8150 6811
rect 8179 6827 8264 6835
rect 8179 6807 8236 6827
rect 8256 6807 8264 6827
rect 8112 6801 8149 6802
rect 8179 6801 8264 6807
rect 8330 6831 8368 6839
rect 8330 6811 8339 6831
rect 8359 6811 8368 6831
rect 8330 6802 8368 6811
rect 8512 6836 8555 6863
rect 8512 6818 8526 6836
rect 8544 6818 8555 6836
rect 8512 6810 8555 6818
rect 8517 6808 8555 6810
rect 8957 6837 9402 6867
rect 10440 6850 10505 6851
rect 8957 6834 9380 6837
rect 8330 6801 8367 6802
rect 7791 6773 7881 6779
rect 7791 6753 7807 6773
rect 7827 6771 7881 6773
rect 7827 6753 7852 6771
rect 7791 6751 7852 6753
rect 7872 6751 7881 6771
rect 7791 6745 7881 6751
rect 7804 6691 7841 6692
rect 7900 6691 7937 6692
rect 7956 6691 7992 6801
rect 8179 6780 8210 6801
rect 8957 6786 9004 6834
rect 8175 6779 8210 6780
rect 8053 6769 8210 6779
rect 8053 6749 8070 6769
rect 8090 6749 8210 6769
rect 8053 6742 8210 6749
rect 8277 6772 8426 6780
rect 8277 6752 8288 6772
rect 8308 6752 8347 6772
rect 8367 6752 8426 6772
rect 8957 6768 8967 6786
rect 8985 6768 9004 6786
rect 8957 6764 9004 6768
rect 10091 6825 10278 6849
rect 10309 6830 10702 6850
rect 10722 6830 10725 6850
rect 10309 6825 10725 6830
rect 8958 6759 8995 6764
rect 8277 6745 8426 6752
rect 10091 6754 10128 6825
rect 10309 6824 10650 6825
rect 10243 6764 10274 6765
rect 8277 6744 8318 6745
rect 8514 6743 8551 6746
rect 8011 6691 8048 6692
rect 7704 6682 7842 6691
rect 6908 6643 7352 6669
rect 6908 6641 7076 6643
rect 6908 6463 6935 6641
rect 6975 6603 7039 6615
rect 7315 6611 7352 6643
rect 7378 6642 7569 6664
rect 7704 6662 7813 6682
rect 7833 6662 7842 6682
rect 7704 6655 7842 6662
rect 7900 6682 8048 6691
rect 7900 6662 7909 6682
rect 7929 6662 8019 6682
rect 8039 6662 8048 6682
rect 7704 6653 7800 6655
rect 7900 6652 8048 6662
rect 8107 6682 8144 6692
rect 8107 6662 8115 6682
rect 8135 6662 8144 6682
rect 7956 6651 7992 6652
rect 7533 6640 7569 6642
rect 7533 6611 7570 6640
rect 6975 6602 7010 6603
rect 6952 6597 7010 6602
rect 6952 6577 6955 6597
rect 6975 6583 7010 6597
rect 7030 6583 7039 6603
rect 6975 6577 7039 6583
rect 6952 6575 7039 6577
rect 6952 6571 6979 6575
rect 7001 6574 7039 6575
rect 7002 6573 7039 6574
rect 7105 6607 7141 6608
rect 7213 6607 7249 6608
rect 7105 6600 7249 6607
rect 7105 6599 7167 6600
rect 7105 6579 7113 6599
rect 7133 6582 7167 6599
rect 7186 6599 7249 6600
rect 7186 6582 7221 6599
rect 7133 6579 7221 6582
rect 7241 6579 7249 6599
rect 7105 6573 7249 6579
rect 7315 6603 7353 6611
rect 7431 6607 7467 6608
rect 7315 6583 7324 6603
rect 7344 6583 7353 6603
rect 7315 6574 7353 6583
rect 7382 6599 7467 6607
rect 7382 6579 7439 6599
rect 7459 6579 7467 6599
rect 7315 6573 7352 6574
rect 7382 6573 7467 6579
rect 7533 6603 7571 6611
rect 7533 6583 7542 6603
rect 7562 6583 7571 6603
rect 7804 6592 7841 6593
rect 8107 6592 8144 6662
rect 8179 6691 8210 6742
rect 8506 6737 8551 6743
rect 8506 6719 8524 6737
rect 8542 6719 8551 6737
rect 10091 6734 10100 6754
rect 10120 6734 10128 6754
rect 10091 6724 10128 6734
rect 10187 6754 10274 6764
rect 10187 6734 10196 6754
rect 10216 6734 10274 6754
rect 10187 6725 10274 6734
rect 10187 6724 10224 6725
rect 8506 6709 8551 6719
rect 8229 6691 8266 6692
rect 8179 6682 8266 6691
rect 8179 6662 8237 6682
rect 8257 6662 8266 6682
rect 8179 6652 8266 6662
rect 8325 6682 8362 6692
rect 8325 6662 8333 6682
rect 8353 6662 8362 6682
rect 8506 6667 8549 6709
rect 8946 6697 8998 6699
rect 8412 6665 8549 6667
rect 8179 6651 8210 6652
rect 8325 6592 8362 6662
rect 7803 6591 8144 6592
rect 7533 6574 7571 6583
rect 7728 6586 8144 6591
rect 7533 6573 7570 6574
rect 6994 6545 7084 6551
rect 6994 6525 7010 6545
rect 7030 6543 7084 6545
rect 7030 6525 7055 6543
rect 6994 6523 7055 6525
rect 7075 6523 7084 6543
rect 6994 6517 7084 6523
rect 7007 6463 7044 6464
rect 7103 6463 7140 6464
rect 7159 6463 7195 6573
rect 7382 6552 7413 6573
rect 7728 6566 7731 6586
rect 7751 6566 8144 6586
rect 8328 6576 8362 6592
rect 8406 6644 8549 6665
rect 8944 6693 9377 6697
rect 8944 6687 9383 6693
rect 8944 6669 8965 6687
rect 8983 6669 9383 6687
rect 10243 6674 10274 6725
rect 10309 6754 10346 6824
rect 10612 6823 10649 6824
rect 10461 6764 10497 6765
rect 10309 6734 10318 6754
rect 10338 6734 10346 6754
rect 10309 6724 10346 6734
rect 10405 6754 10553 6764
rect 10653 6761 10749 6763
rect 10405 6734 10414 6754
rect 10434 6734 10524 6754
rect 10544 6734 10553 6754
rect 10405 6725 10553 6734
rect 10611 6754 10749 6761
rect 10611 6734 10620 6754
rect 10640 6734 10749 6754
rect 10611 6725 10749 6734
rect 10405 6724 10442 6725
rect 10135 6671 10176 6672
rect 8944 6651 9383 6669
rect 8104 6557 8144 6566
rect 8406 6557 8433 6644
rect 8506 6618 8549 6644
rect 8506 6600 8519 6618
rect 8537 6600 8549 6618
rect 8506 6589 8549 6600
rect 7378 6551 7413 6552
rect 7256 6541 7413 6551
rect 7256 6521 7273 6541
rect 7293 6521 7413 6541
rect 7256 6514 7413 6521
rect 7480 6544 7626 6552
rect 7480 6524 7491 6544
rect 7511 6524 7550 6544
rect 7570 6524 7626 6544
rect 8104 6540 8433 6557
rect 8104 6539 8144 6540
rect 7480 6517 7626 6524
rect 8501 6528 8541 6531
rect 8501 6522 8544 6528
rect 8126 6519 8544 6522
rect 7480 6516 7521 6517
rect 7214 6463 7251 6464
rect 6907 6454 7045 6463
rect 6907 6434 7016 6454
rect 7036 6434 7045 6454
rect 6907 6427 7045 6434
rect 7103 6454 7251 6463
rect 7103 6434 7112 6454
rect 7132 6434 7222 6454
rect 7242 6434 7251 6454
rect 6907 6425 7003 6427
rect 7103 6424 7251 6434
rect 7310 6454 7347 6464
rect 7310 6434 7318 6454
rect 7338 6434 7347 6454
rect 7159 6423 7195 6424
rect 7007 6364 7044 6365
rect 7310 6364 7347 6434
rect 7382 6463 7413 6514
rect 8126 6501 8517 6519
rect 8535 6501 8544 6519
rect 8126 6499 8544 6501
rect 8126 6491 8153 6499
rect 8394 6496 8544 6499
rect 7706 6485 7874 6486
rect 8125 6485 8153 6491
rect 7706 6469 8153 6485
rect 8501 6491 8544 6496
rect 7432 6463 7469 6464
rect 7382 6454 7469 6463
rect 7382 6434 7440 6454
rect 7460 6434 7469 6454
rect 7382 6424 7469 6434
rect 7528 6454 7565 6464
rect 7528 6434 7536 6454
rect 7556 6434 7565 6454
rect 7382 6423 7413 6424
rect 7006 6363 7347 6364
rect 7528 6363 7565 6434
rect 6931 6358 7347 6363
rect 6931 6338 6934 6358
rect 6954 6338 7347 6358
rect 7378 6339 7565 6363
rect 7706 6459 8150 6469
rect 7706 6457 7874 6459
rect 6806 6259 6848 6304
rect 7706 6279 7733 6457
rect 7773 6419 7837 6431
rect 8113 6427 8150 6459
rect 8176 6458 8367 6480
rect 8331 6456 8367 6458
rect 8331 6427 8368 6456
rect 8501 6435 8541 6491
rect 7773 6418 7808 6419
rect 7750 6413 7808 6418
rect 7750 6393 7753 6413
rect 7773 6399 7808 6413
rect 7828 6399 7837 6419
rect 7773 6391 7837 6399
rect 7799 6390 7837 6391
rect 7800 6389 7837 6390
rect 7903 6423 7939 6424
rect 8011 6423 8047 6424
rect 7903 6415 8047 6423
rect 7903 6395 7911 6415
rect 7931 6395 7966 6415
rect 7986 6395 8019 6415
rect 8039 6395 8047 6415
rect 7903 6389 8047 6395
rect 8113 6419 8151 6427
rect 8229 6423 8265 6424
rect 8113 6399 8122 6419
rect 8142 6399 8151 6419
rect 8113 6390 8151 6399
rect 8180 6415 8265 6423
rect 8180 6395 8237 6415
rect 8257 6395 8265 6415
rect 8113 6389 8150 6390
rect 8180 6389 8265 6395
rect 8331 6419 8369 6427
rect 8331 6399 8340 6419
rect 8360 6399 8369 6419
rect 8501 6417 8513 6435
rect 8531 6417 8541 6435
rect 8946 6462 8998 6651
rect 9344 6626 9383 6651
rect 10027 6664 10176 6671
rect 10027 6644 10086 6664
rect 10106 6644 10145 6664
rect 10165 6644 10176 6664
rect 10027 6636 10176 6644
rect 10243 6667 10400 6674
rect 10243 6647 10363 6667
rect 10383 6647 10400 6667
rect 10243 6637 10400 6647
rect 10243 6636 10278 6637
rect 9128 6601 9315 6625
rect 9344 6606 9739 6626
rect 9759 6606 9762 6626
rect 10243 6615 10274 6636
rect 10461 6615 10497 6725
rect 10516 6724 10553 6725
rect 10612 6724 10649 6725
rect 10572 6665 10662 6671
rect 10572 6645 10581 6665
rect 10601 6663 10662 6665
rect 10601 6645 10626 6663
rect 10572 6643 10626 6645
rect 10646 6643 10662 6663
rect 10572 6637 10662 6643
rect 10086 6614 10123 6615
rect 9344 6601 9762 6606
rect 10085 6605 10123 6614
rect 9128 6530 9165 6601
rect 9344 6600 9687 6601
rect 9344 6597 9383 6600
rect 9649 6599 9686 6600
rect 9280 6540 9311 6541
rect 9128 6510 9137 6530
rect 9157 6510 9165 6530
rect 9128 6500 9165 6510
rect 9224 6530 9311 6540
rect 9224 6510 9233 6530
rect 9253 6510 9311 6530
rect 9224 6501 9311 6510
rect 9224 6500 9261 6501
rect 8946 6444 8962 6462
rect 8980 6444 8998 6462
rect 9280 6450 9311 6501
rect 9346 6530 9383 6597
rect 10085 6585 10094 6605
rect 10114 6585 10123 6605
rect 10085 6577 10123 6585
rect 10189 6609 10274 6615
rect 10304 6614 10341 6615
rect 10189 6589 10197 6609
rect 10217 6589 10274 6609
rect 10189 6581 10274 6589
rect 10303 6605 10341 6614
rect 10303 6585 10312 6605
rect 10332 6585 10341 6605
rect 10189 6580 10225 6581
rect 10303 6577 10341 6585
rect 10407 6609 10551 6615
rect 10407 6589 10415 6609
rect 10435 6608 10523 6609
rect 10435 6590 10470 6608
rect 10488 6590 10523 6608
rect 10435 6589 10523 6590
rect 10543 6589 10551 6609
rect 10407 6581 10551 6589
rect 10407 6580 10443 6581
rect 10515 6580 10551 6581
rect 10617 6614 10654 6615
rect 10617 6613 10655 6614
rect 10617 6605 10681 6613
rect 10617 6585 10626 6605
rect 10646 6591 10681 6605
rect 10701 6591 10704 6611
rect 10646 6586 10704 6591
rect 10646 6585 10681 6586
rect 10086 6548 10123 6577
rect 10087 6546 10123 6548
rect 9498 6540 9534 6541
rect 9346 6510 9355 6530
rect 9375 6510 9383 6530
rect 9346 6500 9383 6510
rect 9442 6530 9590 6540
rect 9690 6537 9786 6539
rect 9442 6510 9451 6530
rect 9471 6510 9561 6530
rect 9581 6510 9590 6530
rect 9442 6501 9590 6510
rect 9648 6530 9786 6537
rect 9648 6510 9657 6530
rect 9677 6510 9786 6530
rect 10087 6524 10278 6546
rect 10304 6545 10341 6577
rect 10617 6573 10681 6585
rect 10721 6549 10748 6725
rect 10667 6547 10748 6549
rect 10580 6545 10748 6547
rect 10304 6519 10748 6545
rect 10414 6517 10454 6519
rect 10580 6518 10748 6519
rect 9648 6501 9786 6510
rect 10689 6516 10748 6518
rect 9442 6500 9479 6501
rect 9172 6447 9213 6448
rect 8946 6426 8998 6444
rect 9064 6440 9213 6447
rect 8501 6407 8541 6417
rect 9064 6420 9123 6440
rect 9143 6420 9182 6440
rect 9202 6420 9213 6440
rect 9064 6412 9213 6420
rect 9280 6443 9437 6450
rect 9280 6423 9400 6443
rect 9420 6423 9437 6443
rect 9280 6413 9437 6423
rect 9280 6412 9315 6413
rect 8331 6390 8369 6399
rect 9280 6391 9311 6412
rect 9498 6391 9534 6501
rect 9553 6500 9590 6501
rect 9649 6500 9686 6501
rect 9609 6441 9699 6447
rect 9609 6421 9618 6441
rect 9638 6439 9699 6441
rect 9638 6421 9663 6439
rect 9609 6419 9663 6421
rect 9683 6419 9699 6439
rect 9609 6413 9699 6419
rect 9123 6390 9160 6391
rect 8331 6389 8368 6390
rect 7792 6361 7882 6367
rect 7792 6341 7808 6361
rect 7828 6359 7882 6361
rect 7828 6341 7853 6359
rect 7792 6339 7853 6341
rect 7873 6339 7882 6359
rect 7792 6333 7882 6339
rect 7805 6279 7842 6280
rect 7901 6279 7938 6280
rect 7957 6279 7993 6389
rect 8180 6368 8211 6389
rect 9122 6381 9160 6390
rect 8176 6367 8211 6368
rect 8054 6357 8211 6367
rect 8054 6337 8071 6357
rect 8091 6337 8211 6357
rect 8054 6330 8211 6337
rect 8278 6360 8427 6368
rect 8278 6340 8289 6360
rect 8309 6340 8348 6360
rect 8368 6340 8427 6360
rect 8950 6363 8990 6373
rect 8278 6333 8427 6340
rect 8493 6336 8545 6354
rect 8278 6332 8319 6333
rect 8012 6279 8049 6280
rect 7705 6270 7843 6279
rect 7177 6259 7210 6261
rect 6806 6247 7253 6259
rect 6809 6233 7253 6247
rect 6809 6231 6977 6233
rect 6809 6053 6836 6231
rect 6876 6193 6940 6205
rect 7216 6201 7253 6233
rect 7279 6232 7470 6254
rect 7705 6250 7814 6270
rect 7834 6250 7843 6270
rect 7705 6243 7843 6250
rect 7901 6270 8049 6279
rect 7901 6250 7910 6270
rect 7930 6250 8020 6270
rect 8040 6250 8049 6270
rect 7705 6241 7801 6243
rect 7901 6240 8049 6250
rect 8108 6270 8145 6280
rect 8108 6250 8116 6270
rect 8136 6250 8145 6270
rect 7957 6239 7993 6240
rect 7434 6230 7470 6232
rect 7434 6201 7471 6230
rect 6876 6192 6911 6193
rect 6853 6187 6911 6192
rect 6853 6167 6856 6187
rect 6876 6173 6911 6187
rect 6931 6173 6940 6193
rect 6876 6165 6940 6173
rect 6902 6164 6940 6165
rect 6903 6163 6940 6164
rect 7006 6197 7042 6198
rect 7114 6197 7150 6198
rect 7006 6189 7150 6197
rect 7006 6169 7014 6189
rect 7034 6187 7122 6189
rect 7034 6169 7067 6187
rect 7006 6168 7067 6169
rect 7088 6169 7122 6187
rect 7142 6169 7150 6189
rect 7088 6168 7150 6169
rect 7006 6163 7150 6168
rect 7216 6193 7254 6201
rect 7332 6197 7368 6198
rect 7216 6173 7225 6193
rect 7245 6173 7254 6193
rect 7216 6164 7254 6173
rect 7283 6189 7368 6197
rect 7283 6169 7340 6189
rect 7360 6169 7368 6189
rect 7216 6163 7253 6164
rect 7283 6163 7368 6169
rect 7434 6193 7472 6201
rect 7434 6173 7443 6193
rect 7463 6173 7472 6193
rect 8108 6183 8145 6250
rect 8180 6279 8211 6330
rect 8493 6318 8511 6336
rect 8529 6318 8545 6336
rect 8230 6279 8267 6280
rect 8180 6270 8267 6279
rect 8180 6250 8238 6270
rect 8258 6250 8267 6270
rect 8180 6240 8267 6250
rect 8326 6270 8363 6280
rect 8326 6250 8334 6270
rect 8354 6250 8363 6270
rect 8180 6239 8211 6240
rect 7805 6180 7842 6181
rect 8108 6180 8147 6183
rect 7804 6179 8147 6180
rect 8326 6179 8363 6250
rect 7434 6164 7472 6173
rect 7729 6174 8147 6179
rect 7434 6163 7471 6164
rect 6895 6135 6985 6141
rect 6895 6115 6911 6135
rect 6931 6133 6985 6135
rect 6931 6115 6956 6133
rect 6895 6113 6956 6115
rect 6976 6113 6985 6133
rect 6895 6107 6985 6113
rect 6908 6053 6945 6054
rect 7004 6053 7041 6054
rect 7060 6053 7096 6163
rect 7283 6142 7314 6163
rect 7729 6154 7732 6174
rect 7752 6154 8147 6174
rect 8176 6155 8363 6179
rect 7279 6141 7314 6142
rect 7157 6131 7314 6141
rect 7157 6111 7174 6131
rect 7194 6111 7314 6131
rect 7157 6104 7314 6111
rect 7381 6134 7530 6142
rect 7381 6114 7392 6134
rect 7412 6114 7451 6134
rect 7471 6114 7530 6134
rect 7381 6107 7530 6114
rect 8108 6129 8147 6154
rect 8493 6129 8545 6318
rect 8950 6345 8960 6363
rect 8978 6345 8990 6363
rect 9122 6361 9131 6381
rect 9151 6361 9160 6381
rect 9122 6353 9160 6361
rect 9226 6385 9311 6391
rect 9341 6390 9378 6391
rect 9226 6365 9234 6385
rect 9254 6365 9311 6385
rect 9226 6357 9311 6365
rect 9340 6381 9378 6390
rect 9340 6361 9349 6381
rect 9369 6361 9378 6381
rect 9226 6356 9262 6357
rect 9340 6353 9378 6361
rect 9444 6385 9588 6391
rect 9444 6365 9452 6385
rect 9472 6365 9505 6385
rect 9525 6365 9560 6385
rect 9580 6365 9588 6385
rect 9444 6357 9588 6365
rect 9444 6356 9480 6357
rect 9552 6356 9588 6357
rect 9654 6390 9691 6391
rect 9654 6389 9692 6390
rect 9654 6381 9718 6389
rect 9654 6361 9663 6381
rect 9683 6367 9718 6381
rect 9738 6367 9741 6387
rect 9683 6362 9741 6367
rect 9683 6361 9718 6362
rect 8950 6289 8990 6345
rect 9123 6324 9160 6353
rect 9124 6322 9160 6324
rect 9124 6300 9315 6322
rect 9341 6321 9378 6353
rect 9654 6349 9718 6361
rect 9758 6323 9785 6501
rect 10689 6498 10718 6516
rect 9617 6321 9785 6323
rect 9341 6311 9785 6321
rect 9926 6417 10113 6441
rect 10144 6422 10537 6442
rect 10557 6422 10560 6442
rect 10144 6417 10560 6422
rect 9926 6346 9963 6417
rect 10144 6416 10485 6417
rect 10078 6356 10109 6357
rect 9926 6326 9935 6346
rect 9955 6326 9963 6346
rect 9926 6316 9963 6326
rect 10022 6346 10109 6356
rect 10022 6326 10031 6346
rect 10051 6326 10109 6346
rect 10022 6317 10109 6326
rect 10022 6316 10059 6317
rect 8947 6284 8990 6289
rect 9338 6295 9785 6311
rect 9338 6289 9366 6295
rect 9617 6294 9785 6295
rect 8947 6281 9097 6284
rect 9338 6281 9365 6289
rect 8947 6279 9365 6281
rect 8947 6261 8956 6279
rect 8974 6261 9365 6279
rect 10078 6266 10109 6317
rect 10144 6346 10181 6416
rect 10447 6415 10484 6416
rect 10296 6356 10332 6357
rect 10144 6326 10153 6346
rect 10173 6326 10181 6346
rect 10144 6316 10181 6326
rect 10240 6346 10388 6356
rect 10488 6353 10584 6355
rect 10240 6326 10249 6346
rect 10269 6326 10359 6346
rect 10379 6326 10388 6346
rect 10240 6317 10388 6326
rect 10446 6346 10584 6353
rect 10446 6326 10455 6346
rect 10475 6326 10584 6346
rect 10446 6317 10584 6326
rect 10240 6316 10277 6317
rect 9970 6263 10011 6264
rect 8947 6258 9365 6261
rect 8947 6252 8990 6258
rect 8950 6249 8990 6252
rect 9862 6256 10011 6263
rect 9347 6240 9387 6241
rect 9058 6223 9387 6240
rect 9862 6236 9921 6256
rect 9941 6236 9980 6256
rect 10000 6236 10011 6256
rect 9862 6228 10011 6236
rect 10078 6259 10235 6266
rect 10078 6239 10198 6259
rect 10218 6239 10235 6259
rect 10078 6229 10235 6239
rect 10078 6228 10113 6229
rect 8942 6180 8985 6191
rect 8942 6162 8954 6180
rect 8972 6162 8985 6180
rect 8942 6136 8985 6162
rect 9058 6136 9085 6223
rect 9347 6214 9387 6223
rect 8108 6111 8547 6129
rect 7381 6106 7422 6107
rect 7115 6053 7152 6054
rect 6808 6044 6946 6053
rect 6808 6024 6917 6044
rect 6937 6024 6946 6044
rect 6808 6017 6946 6024
rect 7004 6044 7152 6053
rect 7004 6024 7013 6044
rect 7033 6024 7123 6044
rect 7143 6024 7152 6044
rect 6808 6015 6904 6017
rect 7004 6014 7152 6024
rect 7211 6044 7248 6054
rect 7211 6024 7219 6044
rect 7239 6024 7248 6044
rect 7060 6013 7096 6014
rect 6908 5954 6945 5955
rect 7211 5954 7248 6024
rect 7283 6053 7314 6104
rect 8108 6093 8508 6111
rect 8526 6093 8547 6111
rect 8108 6087 8547 6093
rect 8114 6083 8547 6087
rect 8942 6115 9085 6136
rect 9129 6188 9163 6204
rect 9347 6194 9740 6214
rect 9760 6194 9763 6214
rect 10078 6207 10109 6228
rect 10296 6207 10332 6317
rect 10351 6316 10388 6317
rect 10447 6316 10484 6317
rect 10407 6257 10497 6263
rect 10407 6237 10416 6257
rect 10436 6255 10497 6257
rect 10436 6237 10461 6255
rect 10407 6235 10461 6237
rect 10481 6235 10497 6255
rect 10407 6229 10497 6235
rect 9921 6206 9958 6207
rect 9347 6189 9763 6194
rect 9920 6197 9958 6206
rect 9347 6188 9688 6189
rect 9129 6118 9166 6188
rect 9281 6128 9312 6129
rect 8942 6113 9079 6115
rect 8493 6081 8545 6083
rect 8942 6071 8985 6113
rect 9129 6098 9138 6118
rect 9158 6098 9166 6118
rect 9129 6088 9166 6098
rect 9225 6118 9312 6128
rect 9225 6098 9234 6118
rect 9254 6098 9312 6118
rect 9225 6089 9312 6098
rect 9225 6088 9262 6089
rect 8940 6061 8985 6071
rect 7333 6053 7370 6054
rect 7283 6044 7370 6053
rect 7283 6024 7341 6044
rect 7361 6024 7370 6044
rect 7283 6014 7370 6024
rect 7429 6044 7466 6054
rect 7429 6024 7437 6044
rect 7457 6024 7466 6044
rect 8940 6043 8949 6061
rect 8967 6043 8985 6061
rect 8940 6037 8985 6043
rect 9281 6038 9312 6089
rect 9347 6118 9384 6188
rect 9650 6187 9687 6188
rect 9920 6177 9929 6197
rect 9949 6177 9958 6197
rect 9920 6169 9958 6177
rect 10024 6201 10109 6207
rect 10139 6206 10176 6207
rect 10024 6181 10032 6201
rect 10052 6181 10109 6201
rect 10024 6173 10109 6181
rect 10138 6197 10176 6206
rect 10138 6177 10147 6197
rect 10167 6177 10176 6197
rect 10024 6172 10060 6173
rect 10138 6169 10176 6177
rect 10242 6201 10386 6207
rect 10242 6181 10250 6201
rect 10270 6182 10302 6201
rect 10323 6182 10358 6201
rect 10270 6181 10358 6182
rect 10378 6181 10386 6201
rect 10242 6173 10386 6181
rect 10242 6172 10278 6173
rect 10350 6172 10386 6173
rect 10452 6206 10489 6207
rect 10452 6205 10490 6206
rect 10452 6197 10516 6205
rect 10452 6177 10461 6197
rect 10481 6183 10516 6197
rect 10536 6183 10539 6203
rect 10481 6178 10539 6183
rect 10481 6177 10516 6178
rect 9921 6140 9958 6169
rect 9922 6138 9958 6140
rect 9499 6128 9535 6129
rect 9347 6098 9356 6118
rect 9376 6098 9384 6118
rect 9347 6088 9384 6098
rect 9443 6118 9591 6128
rect 9691 6125 9787 6127
rect 9443 6098 9452 6118
rect 9472 6098 9562 6118
rect 9582 6098 9591 6118
rect 9443 6089 9591 6098
rect 9649 6118 9787 6125
rect 9649 6098 9658 6118
rect 9678 6098 9787 6118
rect 9922 6116 10113 6138
rect 10139 6137 10176 6169
rect 10452 6165 10516 6177
rect 10556 6139 10583 6317
rect 10415 6137 10583 6139
rect 10139 6111 10583 6137
rect 9649 6089 9787 6098
rect 9443 6088 9480 6089
rect 8940 6034 8977 6037
rect 9173 6035 9214 6036
rect 7283 6013 7314 6014
rect 6907 5953 7248 5954
rect 7429 5953 7466 6024
rect 9065 6028 9214 6035
rect 8496 6016 8533 6021
rect 8487 6012 8534 6016
rect 8487 5994 8506 6012
rect 8524 5994 8534 6012
rect 9065 6008 9124 6028
rect 9144 6008 9183 6028
rect 9203 6008 9214 6028
rect 9065 6000 9214 6008
rect 9281 6031 9438 6038
rect 9281 6011 9401 6031
rect 9421 6011 9438 6031
rect 9281 6001 9438 6011
rect 9281 6000 9316 6001
rect 6832 5948 7248 5953
rect 6832 5928 6835 5948
rect 6855 5928 7248 5948
rect 7279 5929 7466 5953
rect 8091 5951 8131 5956
rect 8487 5951 8534 5994
rect 9281 5979 9312 6000
rect 9499 5979 9535 6089
rect 9554 6088 9591 6089
rect 9650 6088 9687 6089
rect 9610 6029 9700 6035
rect 9610 6009 9619 6029
rect 9639 6027 9700 6029
rect 9639 6009 9664 6027
rect 9610 6007 9664 6009
rect 9684 6007 9700 6027
rect 9610 6001 9700 6007
rect 9124 5978 9161 5979
rect 8091 5912 8534 5951
rect 8937 5970 8974 5972
rect 8937 5962 8979 5970
rect 8937 5944 8947 5962
rect 8965 5944 8979 5962
rect 8937 5935 8979 5944
rect 9123 5969 9161 5978
rect 9123 5949 9132 5969
rect 9152 5949 9161 5969
rect 9123 5941 9161 5949
rect 9227 5973 9312 5979
rect 9342 5978 9379 5979
rect 9227 5953 9235 5973
rect 9255 5953 9312 5973
rect 9227 5945 9312 5953
rect 9341 5969 9379 5978
rect 9341 5949 9350 5969
rect 9370 5949 9379 5969
rect 9227 5944 9263 5945
rect 9341 5941 9379 5949
rect 9445 5977 9589 5979
rect 9445 5973 9497 5977
rect 9445 5953 9453 5973
rect 9473 5957 9497 5973
rect 9517 5973 9589 5977
rect 9517 5957 9561 5973
rect 9473 5953 9561 5957
rect 9581 5953 9589 5973
rect 9445 5945 9589 5953
rect 9445 5944 9481 5945
rect 9553 5944 9589 5945
rect 9655 5978 9692 5979
rect 9655 5977 9693 5978
rect 9655 5969 9719 5977
rect 9655 5949 9664 5969
rect 9684 5955 9719 5969
rect 9739 5955 9742 5975
rect 9684 5950 9742 5955
rect 9684 5949 9719 5950
rect 7185 5897 7225 5905
rect 7185 5875 7193 5897
rect 7217 5875 7225 5897
rect 6891 5651 7059 5652
rect 7185 5651 7225 5875
rect 7688 5879 7856 5880
rect 8091 5879 8131 5912
rect 8487 5879 8534 5912
rect 8938 5910 8979 5935
rect 9124 5910 9161 5941
rect 9342 5910 9379 5941
rect 9655 5937 9719 5949
rect 9759 5911 9786 6089
rect 8938 5883 8987 5910
rect 9123 5884 9172 5910
rect 9341 5909 9422 5910
rect 9618 5909 9786 5911
rect 9341 5884 9786 5909
rect 9342 5883 9786 5884
rect 7688 5878 8132 5879
rect 7688 5853 8133 5878
rect 7688 5851 7856 5853
rect 8052 5852 8133 5853
rect 8302 5852 8351 5878
rect 8487 5852 8536 5879
rect 7688 5673 7715 5851
rect 7755 5813 7819 5825
rect 8095 5821 8132 5852
rect 8313 5821 8350 5852
rect 8495 5827 8536 5852
rect 8940 5850 8987 5883
rect 9343 5850 9383 5883
rect 9618 5882 9786 5883
rect 10249 5887 10289 6111
rect 10415 6110 10583 6111
rect 10249 5865 10257 5887
rect 10281 5865 10289 5887
rect 10249 5857 10289 5865
rect 7755 5812 7790 5813
rect 7732 5807 7790 5812
rect 7732 5787 7735 5807
rect 7755 5793 7790 5807
rect 7810 5793 7819 5813
rect 7755 5785 7819 5793
rect 7781 5784 7819 5785
rect 7782 5783 7819 5784
rect 7885 5817 7921 5818
rect 7993 5817 8029 5818
rect 7885 5809 8029 5817
rect 7885 5789 7893 5809
rect 7913 5805 8001 5809
rect 7913 5789 7957 5805
rect 7885 5785 7957 5789
rect 7977 5789 8001 5805
rect 8021 5789 8029 5809
rect 7977 5785 8029 5789
rect 7885 5783 8029 5785
rect 8095 5813 8133 5821
rect 8211 5817 8247 5818
rect 8095 5793 8104 5813
rect 8124 5793 8133 5813
rect 8095 5784 8133 5793
rect 8162 5809 8247 5817
rect 8162 5789 8219 5809
rect 8239 5789 8247 5809
rect 8095 5783 8132 5784
rect 8162 5783 8247 5789
rect 8313 5813 8351 5821
rect 8313 5793 8322 5813
rect 8342 5793 8351 5813
rect 8313 5784 8351 5793
rect 8495 5818 8537 5827
rect 8495 5800 8509 5818
rect 8527 5800 8537 5818
rect 8495 5792 8537 5800
rect 8500 5790 8537 5792
rect 8940 5811 9383 5850
rect 8313 5783 8350 5784
rect 7774 5755 7864 5761
rect 7774 5735 7790 5755
rect 7810 5753 7864 5755
rect 7810 5735 7835 5753
rect 7774 5733 7835 5735
rect 7855 5733 7864 5753
rect 7774 5727 7864 5733
rect 7787 5673 7824 5674
rect 7883 5673 7920 5674
rect 7939 5673 7975 5783
rect 8162 5762 8193 5783
rect 8940 5768 8987 5811
rect 9343 5806 9383 5811
rect 10008 5809 10195 5833
rect 10226 5814 10619 5834
rect 10639 5814 10642 5834
rect 10226 5809 10642 5814
rect 8158 5761 8193 5762
rect 8036 5751 8193 5761
rect 8036 5731 8053 5751
rect 8073 5731 8193 5751
rect 8036 5724 8193 5731
rect 8260 5754 8409 5762
rect 8260 5734 8271 5754
rect 8291 5734 8330 5754
rect 8350 5734 8409 5754
rect 8940 5750 8950 5768
rect 8968 5750 8987 5768
rect 8940 5746 8987 5750
rect 8941 5741 8978 5746
rect 8260 5727 8409 5734
rect 10008 5738 10045 5809
rect 10226 5808 10567 5809
rect 10160 5748 10191 5749
rect 8260 5726 8301 5727
rect 8497 5725 8534 5728
rect 7994 5673 8031 5674
rect 7687 5664 7825 5673
rect 6891 5625 7335 5651
rect 6891 5623 7059 5625
rect 6891 5445 6918 5623
rect 6958 5585 7022 5597
rect 7298 5593 7335 5625
rect 7361 5624 7552 5646
rect 7687 5644 7796 5664
rect 7816 5644 7825 5664
rect 7687 5637 7825 5644
rect 7883 5664 8031 5673
rect 7883 5644 7892 5664
rect 7912 5644 8002 5664
rect 8022 5644 8031 5664
rect 7687 5635 7783 5637
rect 7883 5634 8031 5644
rect 8090 5664 8127 5674
rect 8090 5644 8098 5664
rect 8118 5644 8127 5664
rect 7939 5633 7975 5634
rect 7516 5622 7552 5624
rect 7516 5593 7553 5622
rect 6958 5584 6993 5585
rect 6935 5579 6993 5584
rect 6935 5559 6938 5579
rect 6958 5565 6993 5579
rect 7013 5565 7022 5585
rect 6958 5557 7022 5565
rect 6984 5556 7022 5557
rect 6985 5555 7022 5556
rect 7088 5589 7124 5590
rect 7196 5589 7232 5590
rect 7088 5581 7232 5589
rect 7088 5561 7096 5581
rect 7116 5580 7204 5581
rect 7116 5561 7151 5580
rect 7172 5561 7204 5580
rect 7224 5561 7232 5581
rect 7088 5555 7232 5561
rect 7298 5585 7336 5593
rect 7414 5589 7450 5590
rect 7298 5565 7307 5585
rect 7327 5565 7336 5585
rect 7298 5556 7336 5565
rect 7365 5581 7450 5589
rect 7365 5561 7422 5581
rect 7442 5561 7450 5581
rect 7298 5555 7335 5556
rect 7365 5555 7450 5561
rect 7516 5585 7554 5593
rect 7516 5565 7525 5585
rect 7545 5565 7554 5585
rect 7787 5574 7824 5575
rect 8090 5574 8127 5644
rect 8162 5673 8193 5724
rect 8489 5719 8534 5725
rect 8489 5701 8507 5719
rect 8525 5701 8534 5719
rect 10008 5718 10017 5738
rect 10037 5718 10045 5738
rect 10008 5708 10045 5718
rect 10104 5738 10191 5748
rect 10104 5718 10113 5738
rect 10133 5718 10191 5738
rect 10104 5709 10191 5718
rect 10104 5708 10141 5709
rect 8489 5691 8534 5701
rect 8212 5673 8249 5674
rect 8162 5664 8249 5673
rect 8162 5644 8220 5664
rect 8240 5644 8249 5664
rect 8162 5634 8249 5644
rect 8308 5664 8345 5674
rect 8308 5644 8316 5664
rect 8336 5644 8345 5664
rect 8489 5649 8532 5691
rect 8929 5679 8981 5681
rect 8395 5647 8532 5649
rect 8162 5633 8193 5634
rect 8308 5574 8345 5644
rect 7786 5573 8127 5574
rect 7516 5556 7554 5565
rect 7711 5568 8127 5573
rect 7516 5555 7553 5556
rect 6977 5527 7067 5533
rect 6977 5507 6993 5527
rect 7013 5525 7067 5527
rect 7013 5507 7038 5525
rect 6977 5505 7038 5507
rect 7058 5505 7067 5525
rect 6977 5499 7067 5505
rect 6990 5445 7027 5446
rect 7086 5445 7123 5446
rect 7142 5445 7178 5555
rect 7365 5534 7396 5555
rect 7711 5548 7714 5568
rect 7734 5548 8127 5568
rect 8311 5558 8345 5574
rect 8389 5626 8532 5647
rect 8927 5675 9360 5679
rect 8927 5669 9366 5675
rect 8927 5651 8948 5669
rect 8966 5651 9366 5669
rect 10160 5658 10191 5709
rect 10226 5738 10263 5808
rect 10529 5807 10566 5808
rect 10378 5748 10414 5749
rect 10226 5718 10235 5738
rect 10255 5718 10263 5738
rect 10226 5708 10263 5718
rect 10322 5738 10470 5748
rect 10570 5745 10666 5747
rect 10322 5718 10331 5738
rect 10351 5718 10441 5738
rect 10461 5718 10470 5738
rect 10322 5709 10470 5718
rect 10528 5738 10666 5745
rect 10528 5718 10537 5738
rect 10557 5718 10666 5738
rect 10528 5709 10666 5718
rect 10322 5708 10359 5709
rect 10052 5655 10093 5656
rect 8927 5633 9366 5651
rect 8087 5539 8127 5548
rect 8389 5539 8416 5626
rect 8489 5600 8532 5626
rect 8489 5582 8502 5600
rect 8520 5582 8532 5600
rect 8489 5571 8532 5582
rect 7361 5533 7396 5534
rect 7239 5523 7396 5533
rect 7239 5503 7256 5523
rect 7276 5503 7396 5523
rect 7239 5496 7396 5503
rect 7463 5526 7612 5534
rect 7463 5506 7474 5526
rect 7494 5506 7533 5526
rect 7553 5506 7612 5526
rect 8087 5522 8416 5539
rect 8087 5521 8127 5522
rect 7463 5499 7612 5506
rect 8484 5510 8524 5513
rect 8484 5504 8527 5510
rect 8109 5501 8527 5504
rect 7463 5498 7504 5499
rect 7197 5445 7234 5446
rect 6890 5436 7028 5445
rect 6588 5261 6628 5433
rect 6890 5416 6999 5436
rect 7019 5416 7028 5436
rect 6890 5409 7028 5416
rect 7086 5436 7234 5445
rect 7086 5416 7095 5436
rect 7115 5416 7205 5436
rect 7225 5416 7234 5436
rect 6890 5407 6986 5409
rect 7086 5406 7234 5416
rect 7293 5436 7330 5446
rect 7293 5416 7301 5436
rect 7321 5416 7330 5436
rect 7142 5405 7178 5406
rect 6990 5346 7027 5347
rect 7293 5346 7330 5416
rect 7365 5445 7396 5496
rect 8109 5483 8500 5501
rect 8518 5483 8527 5501
rect 8109 5481 8527 5483
rect 8109 5473 8136 5481
rect 8377 5478 8527 5481
rect 7689 5467 7857 5468
rect 8108 5467 8136 5473
rect 7689 5451 8136 5467
rect 8484 5473 8527 5478
rect 7415 5445 7452 5446
rect 7365 5436 7452 5445
rect 7365 5416 7423 5436
rect 7443 5416 7452 5436
rect 7365 5406 7452 5416
rect 7511 5436 7548 5446
rect 7511 5416 7519 5436
rect 7539 5416 7548 5436
rect 7365 5405 7396 5406
rect 6989 5345 7330 5346
rect 7511 5345 7548 5416
rect 6914 5340 7330 5345
rect 6914 5320 6917 5340
rect 6937 5320 7330 5340
rect 7361 5321 7548 5345
rect 7689 5441 8133 5451
rect 7689 5439 7857 5441
rect 7689 5261 7716 5439
rect 7756 5401 7820 5413
rect 8096 5409 8133 5441
rect 8159 5440 8350 5462
rect 8314 5438 8350 5440
rect 8314 5409 8351 5438
rect 8484 5417 8524 5473
rect 7756 5400 7791 5401
rect 7733 5395 7791 5400
rect 7733 5375 7736 5395
rect 7756 5381 7791 5395
rect 7811 5381 7820 5401
rect 7756 5373 7820 5381
rect 7782 5372 7820 5373
rect 7783 5371 7820 5372
rect 7886 5405 7922 5406
rect 7994 5405 8030 5406
rect 7886 5397 8030 5405
rect 7886 5377 7894 5397
rect 7914 5377 7949 5397
rect 7969 5377 8002 5397
rect 8022 5377 8030 5397
rect 7886 5371 8030 5377
rect 8096 5401 8134 5409
rect 8212 5405 8248 5406
rect 8096 5381 8105 5401
rect 8125 5381 8134 5401
rect 8096 5372 8134 5381
rect 8163 5397 8248 5405
rect 8163 5377 8220 5397
rect 8240 5377 8248 5397
rect 8096 5371 8133 5372
rect 8163 5371 8248 5377
rect 8314 5401 8352 5409
rect 8314 5381 8323 5401
rect 8343 5381 8352 5401
rect 8484 5399 8496 5417
rect 8514 5399 8524 5417
rect 8929 5444 8981 5633
rect 9327 5608 9366 5633
rect 9944 5648 10093 5655
rect 9944 5628 10003 5648
rect 10023 5628 10062 5648
rect 10082 5628 10093 5648
rect 9944 5620 10093 5628
rect 10160 5651 10317 5658
rect 10160 5631 10280 5651
rect 10300 5631 10317 5651
rect 10160 5621 10317 5631
rect 10160 5620 10195 5621
rect 9111 5583 9298 5607
rect 9327 5588 9722 5608
rect 9742 5588 9745 5608
rect 10160 5599 10191 5620
rect 10378 5599 10414 5709
rect 10433 5708 10470 5709
rect 10529 5708 10566 5709
rect 10489 5649 10579 5655
rect 10489 5629 10498 5649
rect 10518 5647 10579 5649
rect 10518 5629 10543 5647
rect 10489 5627 10543 5629
rect 10563 5627 10579 5647
rect 10489 5621 10579 5627
rect 10003 5598 10040 5599
rect 9327 5583 9745 5588
rect 10002 5589 10040 5598
rect 9111 5512 9148 5583
rect 9327 5582 9670 5583
rect 9327 5579 9366 5582
rect 9632 5581 9669 5582
rect 9263 5522 9294 5523
rect 9111 5492 9120 5512
rect 9140 5492 9148 5512
rect 9111 5482 9148 5492
rect 9207 5512 9294 5522
rect 9207 5492 9216 5512
rect 9236 5492 9294 5512
rect 9207 5483 9294 5492
rect 9207 5482 9244 5483
rect 8929 5426 8945 5444
rect 8963 5426 8981 5444
rect 9263 5432 9294 5483
rect 9329 5512 9366 5579
rect 10002 5569 10011 5589
rect 10031 5569 10040 5589
rect 10002 5561 10040 5569
rect 10106 5593 10191 5599
rect 10221 5598 10258 5599
rect 10106 5573 10114 5593
rect 10134 5573 10191 5593
rect 10106 5565 10191 5573
rect 10220 5589 10258 5598
rect 10220 5569 10229 5589
rect 10249 5569 10258 5589
rect 10106 5564 10142 5565
rect 10220 5561 10258 5569
rect 10324 5593 10468 5599
rect 10324 5573 10332 5593
rect 10352 5588 10440 5593
rect 10352 5573 10388 5588
rect 10324 5571 10388 5573
rect 10407 5573 10440 5588
rect 10460 5573 10468 5593
rect 10407 5571 10468 5573
rect 10324 5565 10468 5571
rect 10324 5564 10360 5565
rect 10432 5564 10468 5565
rect 10534 5598 10571 5599
rect 10534 5597 10572 5598
rect 10534 5589 10598 5597
rect 10534 5569 10543 5589
rect 10563 5575 10598 5589
rect 10618 5575 10621 5595
rect 10563 5570 10621 5575
rect 10563 5569 10598 5570
rect 10003 5532 10040 5561
rect 10004 5530 10040 5532
rect 9481 5522 9517 5523
rect 9329 5492 9338 5512
rect 9358 5492 9366 5512
rect 9329 5482 9366 5492
rect 9425 5512 9573 5522
rect 9673 5519 9769 5521
rect 9425 5492 9434 5512
rect 9454 5492 9544 5512
rect 9564 5492 9573 5512
rect 9425 5483 9573 5492
rect 9631 5512 9769 5519
rect 9631 5492 9640 5512
rect 9660 5492 9769 5512
rect 10004 5508 10195 5530
rect 10221 5529 10258 5561
rect 10534 5557 10598 5569
rect 10638 5531 10665 5709
rect 10497 5529 10665 5531
rect 10221 5515 10665 5529
rect 10689 5552 10717 6498
rect 10689 5522 10734 5552
rect 10221 5503 10668 5515
rect 10264 5501 10297 5503
rect 9631 5483 9769 5492
rect 9425 5482 9462 5483
rect 9155 5429 9196 5430
rect 8929 5408 8981 5426
rect 9047 5422 9196 5429
rect 8484 5389 8524 5399
rect 9047 5402 9106 5422
rect 9126 5402 9165 5422
rect 9185 5402 9196 5422
rect 9047 5394 9196 5402
rect 9263 5425 9420 5432
rect 9263 5405 9383 5425
rect 9403 5405 9420 5425
rect 9263 5395 9420 5405
rect 9263 5394 9298 5395
rect 8314 5372 8352 5381
rect 9263 5373 9294 5394
rect 9481 5373 9517 5483
rect 9536 5482 9573 5483
rect 9632 5482 9669 5483
rect 9592 5423 9682 5429
rect 9592 5403 9601 5423
rect 9621 5421 9682 5423
rect 9621 5403 9646 5421
rect 9592 5401 9646 5403
rect 9666 5401 9682 5421
rect 9592 5395 9682 5401
rect 9106 5372 9143 5373
rect 8314 5371 8351 5372
rect 7775 5343 7865 5349
rect 7775 5323 7791 5343
rect 7811 5341 7865 5343
rect 7811 5323 7836 5341
rect 7775 5321 7836 5323
rect 7856 5321 7865 5341
rect 7775 5315 7865 5321
rect 7788 5261 7825 5262
rect 7884 5261 7921 5262
rect 7940 5261 7976 5371
rect 8163 5350 8194 5371
rect 9105 5363 9143 5372
rect 8159 5349 8194 5350
rect 8037 5339 8194 5349
rect 8037 5319 8054 5339
rect 8074 5319 8194 5339
rect 8037 5312 8194 5319
rect 8261 5342 8410 5350
rect 8261 5322 8272 5342
rect 8292 5322 8331 5342
rect 8351 5322 8410 5342
rect 8933 5345 8973 5355
rect 8261 5315 8410 5322
rect 8476 5318 8528 5336
rect 8261 5314 8302 5315
rect 7995 5261 8032 5262
rect 6589 5246 6628 5261
rect 7688 5252 7826 5261
rect 6589 5245 6755 5246
rect 6881 5245 6921 5247
rect 6589 5219 7031 5245
rect 6589 5217 6755 5219
rect 6253 5105 6290 5113
rect 6253 5086 6261 5105
rect 6282 5086 6290 5105
rect 6253 5080 6290 5086
rect 6589 5039 6614 5217
rect 6654 5179 6718 5191
rect 6994 5187 7031 5219
rect 7057 5218 7248 5240
rect 7688 5232 7797 5252
rect 7817 5232 7826 5252
rect 7688 5225 7826 5232
rect 7884 5252 8032 5261
rect 7884 5232 7893 5252
rect 7913 5232 8003 5252
rect 8023 5232 8032 5252
rect 7688 5223 7784 5225
rect 7884 5222 8032 5232
rect 8091 5252 8128 5262
rect 8091 5232 8099 5252
rect 8119 5232 8128 5252
rect 7940 5221 7976 5222
rect 7212 5216 7248 5218
rect 7212 5187 7249 5216
rect 6654 5178 6689 5179
rect 6631 5173 6689 5178
rect 6631 5153 6634 5173
rect 6654 5159 6689 5173
rect 6709 5159 6718 5179
rect 6654 5151 6718 5159
rect 6680 5150 6718 5151
rect 6681 5149 6718 5150
rect 6784 5183 6820 5184
rect 6892 5183 6928 5184
rect 6784 5178 6928 5183
rect 6784 5175 6846 5178
rect 6784 5155 6792 5175
rect 6812 5155 6846 5175
rect 6784 5152 6846 5155
rect 6872 5175 6928 5178
rect 6872 5155 6900 5175
rect 6920 5155 6928 5175
rect 6872 5152 6928 5155
rect 6784 5149 6928 5152
rect 6994 5179 7032 5187
rect 7110 5183 7146 5184
rect 6994 5159 7003 5179
rect 7023 5159 7032 5179
rect 6994 5150 7032 5159
rect 7061 5175 7146 5183
rect 7061 5155 7118 5175
rect 7138 5155 7146 5175
rect 6994 5149 7031 5150
rect 7061 5149 7146 5155
rect 7212 5179 7250 5187
rect 7212 5159 7221 5179
rect 7241 5159 7250 5179
rect 8091 5165 8128 5232
rect 8163 5261 8194 5312
rect 8476 5300 8494 5318
rect 8512 5300 8528 5318
rect 8213 5261 8250 5262
rect 8163 5252 8250 5261
rect 8163 5232 8221 5252
rect 8241 5232 8250 5252
rect 8163 5222 8250 5232
rect 8309 5252 8346 5262
rect 8309 5232 8317 5252
rect 8337 5232 8346 5252
rect 8163 5221 8194 5222
rect 7788 5162 7825 5163
rect 8091 5162 8130 5165
rect 7787 5161 8130 5162
rect 8309 5161 8346 5232
rect 7212 5150 7250 5159
rect 7712 5156 8130 5161
rect 7212 5149 7249 5150
rect 6673 5121 6763 5127
rect 6673 5101 6689 5121
rect 6709 5119 6763 5121
rect 6709 5101 6734 5119
rect 6673 5099 6734 5101
rect 6754 5099 6763 5119
rect 6673 5093 6763 5099
rect 6686 5039 6723 5040
rect 6782 5039 6819 5040
rect 6838 5039 6874 5149
rect 7061 5128 7092 5149
rect 7712 5136 7715 5156
rect 7735 5136 8130 5156
rect 8159 5137 8346 5161
rect 7057 5127 7092 5128
rect 6935 5117 7092 5127
rect 6935 5097 6952 5117
rect 6972 5097 7092 5117
rect 6935 5090 7092 5097
rect 7159 5120 7308 5128
rect 7159 5100 7170 5120
rect 7190 5100 7229 5120
rect 7249 5100 7308 5120
rect 7159 5093 7308 5100
rect 8091 5111 8130 5136
rect 8476 5111 8528 5300
rect 8933 5327 8943 5345
rect 8961 5327 8973 5345
rect 9105 5343 9114 5363
rect 9134 5343 9143 5363
rect 9105 5335 9143 5343
rect 9209 5367 9294 5373
rect 9324 5372 9361 5373
rect 9209 5347 9217 5367
rect 9237 5347 9294 5367
rect 9209 5339 9294 5347
rect 9323 5363 9361 5372
rect 9323 5343 9332 5363
rect 9352 5343 9361 5363
rect 9209 5338 9245 5339
rect 9323 5335 9361 5343
rect 9427 5367 9571 5373
rect 9427 5347 9435 5367
rect 9455 5347 9488 5367
rect 9508 5347 9543 5367
rect 9563 5347 9571 5367
rect 9427 5339 9571 5347
rect 9427 5338 9463 5339
rect 9535 5338 9571 5339
rect 9637 5372 9674 5373
rect 9637 5371 9675 5372
rect 9637 5363 9701 5371
rect 9637 5343 9646 5363
rect 9666 5349 9701 5363
rect 9721 5349 9724 5369
rect 9666 5344 9724 5349
rect 9666 5343 9701 5344
rect 8933 5271 8973 5327
rect 9106 5306 9143 5335
rect 9107 5304 9143 5306
rect 9107 5282 9298 5304
rect 9324 5303 9361 5335
rect 9637 5331 9701 5343
rect 9741 5305 9768 5483
rect 10626 5458 10668 5503
rect 10689 5504 10700 5522
rect 10722 5504 10734 5522
rect 10689 5498 10734 5504
rect 10690 5497 10734 5498
rect 9600 5303 9768 5305
rect 9324 5293 9768 5303
rect 9909 5399 10096 5423
rect 10127 5404 10520 5424
rect 10540 5404 10543 5424
rect 10127 5399 10543 5404
rect 9909 5328 9946 5399
rect 10127 5398 10468 5399
rect 10061 5338 10092 5339
rect 9909 5308 9918 5328
rect 9938 5308 9946 5328
rect 9909 5298 9946 5308
rect 10005 5328 10092 5338
rect 10005 5308 10014 5328
rect 10034 5308 10092 5328
rect 10005 5299 10092 5308
rect 10005 5298 10042 5299
rect 8930 5266 8973 5271
rect 9321 5277 9768 5293
rect 9321 5271 9349 5277
rect 9600 5276 9768 5277
rect 8930 5263 9080 5266
rect 9321 5263 9348 5271
rect 8930 5261 9348 5263
rect 8930 5243 8939 5261
rect 8957 5243 9348 5261
rect 10061 5248 10092 5299
rect 10127 5328 10164 5398
rect 10430 5397 10467 5398
rect 10279 5338 10315 5339
rect 10127 5308 10136 5328
rect 10156 5308 10164 5328
rect 10127 5298 10164 5308
rect 10223 5328 10371 5338
rect 10471 5335 10567 5337
rect 10223 5308 10232 5328
rect 10252 5308 10342 5328
rect 10362 5308 10371 5328
rect 10223 5299 10371 5308
rect 10429 5328 10567 5335
rect 10429 5308 10438 5328
rect 10458 5308 10567 5328
rect 10429 5299 10567 5308
rect 10223 5298 10260 5299
rect 9953 5245 9994 5246
rect 8930 5240 9348 5243
rect 8930 5234 8973 5240
rect 8933 5231 8973 5234
rect 9848 5238 9994 5245
rect 9330 5222 9370 5223
rect 9041 5205 9370 5222
rect 9848 5218 9904 5238
rect 9924 5218 9963 5238
rect 9983 5218 9994 5238
rect 9848 5210 9994 5218
rect 10061 5241 10218 5248
rect 10061 5221 10181 5241
rect 10201 5221 10218 5241
rect 10061 5211 10218 5221
rect 10061 5210 10096 5211
rect 8925 5162 8968 5173
rect 8925 5144 8937 5162
rect 8955 5144 8968 5162
rect 8925 5118 8968 5144
rect 9041 5118 9068 5205
rect 9330 5196 9370 5205
rect 8091 5093 8530 5111
rect 7159 5092 7200 5093
rect 6893 5039 6930 5040
rect 6589 5030 6724 5039
rect 6589 5010 6695 5030
rect 6715 5010 6724 5030
rect 6589 5003 6724 5010
rect 6782 5030 6930 5039
rect 6782 5010 6791 5030
rect 6811 5010 6901 5030
rect 6921 5010 6930 5030
rect 6589 5001 6682 5003
rect 6782 5000 6930 5010
rect 6989 5030 7026 5040
rect 6989 5010 6997 5030
rect 7017 5010 7026 5030
rect 6838 4999 6874 5000
rect 6686 4940 6723 4941
rect 6989 4940 7026 5010
rect 7061 5039 7092 5090
rect 8091 5075 8491 5093
rect 8509 5075 8530 5093
rect 8091 5069 8530 5075
rect 8097 5065 8530 5069
rect 8925 5097 9068 5118
rect 9112 5170 9146 5186
rect 9330 5176 9723 5196
rect 9743 5176 9746 5196
rect 10061 5189 10092 5210
rect 10279 5189 10315 5299
rect 10334 5298 10371 5299
rect 10430 5298 10467 5299
rect 10390 5239 10480 5245
rect 10390 5219 10399 5239
rect 10419 5237 10480 5239
rect 10419 5219 10444 5237
rect 10390 5217 10444 5219
rect 10464 5217 10480 5237
rect 10390 5211 10480 5217
rect 9904 5188 9941 5189
rect 9330 5171 9746 5176
rect 9903 5179 9941 5188
rect 9330 5170 9671 5171
rect 9112 5100 9149 5170
rect 9264 5110 9295 5111
rect 8925 5095 9062 5097
rect 8476 5063 8528 5065
rect 8925 5053 8968 5095
rect 9112 5080 9121 5100
rect 9141 5080 9149 5100
rect 9112 5070 9149 5080
rect 9208 5100 9295 5110
rect 9208 5080 9217 5100
rect 9237 5080 9295 5100
rect 9208 5071 9295 5080
rect 9208 5070 9245 5071
rect 8923 5043 8968 5053
rect 7111 5039 7148 5040
rect 7061 5030 7148 5039
rect 7061 5010 7119 5030
rect 7139 5010 7148 5030
rect 7061 5000 7148 5010
rect 7207 5030 7244 5040
rect 7207 5010 7215 5030
rect 7235 5010 7244 5030
rect 8923 5025 8932 5043
rect 8950 5025 8968 5043
rect 8923 5019 8968 5025
rect 9264 5020 9295 5071
rect 9330 5100 9367 5170
rect 9633 5169 9670 5170
rect 9903 5159 9912 5179
rect 9932 5159 9941 5179
rect 9903 5151 9941 5159
rect 10007 5183 10092 5189
rect 10122 5188 10159 5189
rect 10007 5163 10015 5183
rect 10035 5163 10092 5183
rect 10007 5155 10092 5163
rect 10121 5179 10159 5188
rect 10121 5159 10130 5179
rect 10150 5159 10159 5179
rect 10007 5154 10043 5155
rect 10121 5151 10159 5159
rect 10225 5183 10369 5189
rect 10225 5163 10233 5183
rect 10253 5180 10341 5183
rect 10253 5163 10288 5180
rect 10225 5162 10288 5163
rect 10307 5163 10341 5180
rect 10361 5163 10369 5183
rect 10307 5162 10369 5163
rect 10225 5155 10369 5162
rect 10225 5154 10261 5155
rect 10333 5154 10369 5155
rect 10435 5188 10472 5189
rect 10435 5187 10473 5188
rect 10495 5187 10522 5191
rect 10435 5185 10522 5187
rect 10435 5179 10499 5185
rect 10435 5159 10444 5179
rect 10464 5165 10499 5179
rect 10519 5165 10522 5185
rect 10464 5160 10522 5165
rect 10464 5159 10499 5160
rect 9904 5122 9941 5151
rect 9905 5120 9941 5122
rect 9482 5110 9518 5111
rect 9330 5080 9339 5100
rect 9359 5080 9367 5100
rect 9330 5070 9367 5080
rect 9426 5100 9574 5110
rect 9674 5107 9770 5109
rect 9426 5080 9435 5100
rect 9455 5080 9545 5100
rect 9565 5080 9574 5100
rect 9426 5071 9574 5080
rect 9632 5100 9770 5107
rect 9632 5080 9641 5100
rect 9661 5080 9770 5100
rect 9905 5098 10096 5120
rect 10122 5119 10159 5151
rect 10435 5147 10499 5159
rect 10539 5121 10566 5299
rect 10398 5119 10566 5121
rect 10122 5093 10566 5119
rect 9632 5071 9770 5080
rect 9426 5070 9463 5071
rect 8923 5016 8960 5019
rect 9156 5017 9197 5018
rect 7061 4999 7092 5000
rect 6685 4939 7026 4940
rect 7207 4939 7244 5010
rect 9048 5010 9197 5017
rect 8479 4998 8516 5003
rect 6610 4934 7026 4939
rect 6610 4914 6613 4934
rect 6633 4914 7026 4934
rect 7057 4915 7244 4939
rect 8470 4994 8517 4998
rect 8470 4976 8489 4994
rect 8507 4976 8517 4994
rect 9048 4990 9107 5010
rect 9127 4990 9166 5010
rect 9186 4990 9197 5010
rect 9048 4982 9197 4990
rect 9264 5013 9421 5020
rect 9264 4993 9384 5013
rect 9404 4993 9421 5013
rect 9264 4983 9421 4993
rect 9264 4982 9299 4983
rect 8078 4917 8116 4918
rect 8470 4917 8517 4976
rect 9264 4961 9295 4982
rect 9482 4961 9518 5071
rect 9537 5070 9574 5071
rect 9633 5070 9670 5071
rect 9593 5011 9683 5017
rect 9593 4991 9602 5011
rect 9622 5009 9683 5011
rect 9622 4991 9647 5009
rect 9593 4989 9647 4991
rect 9667 4989 9683 5009
rect 9593 4983 9683 4989
rect 9107 4960 9144 4961
rect 8920 4952 8957 4954
rect 8920 4944 8962 4952
rect 8920 4926 8930 4944
rect 8948 4926 8962 4944
rect 8920 4917 8962 4926
rect 9106 4951 9144 4960
rect 9106 4931 9115 4951
rect 9135 4931 9144 4951
rect 9106 4923 9144 4931
rect 9210 4955 9295 4961
rect 9325 4960 9362 4961
rect 9210 4935 9218 4955
rect 9238 4935 9295 4955
rect 9210 4927 9295 4935
rect 9324 4951 9362 4960
rect 9324 4931 9333 4951
rect 9353 4931 9362 4951
rect 9210 4926 9246 4927
rect 9324 4923 9362 4931
rect 9428 4959 9572 4961
rect 9428 4955 9480 4959
rect 9428 4935 9436 4955
rect 9456 4939 9480 4955
rect 9500 4955 9572 4959
rect 9500 4939 9544 4955
rect 9456 4935 9544 4939
rect 9564 4935 9572 4955
rect 9428 4927 9572 4935
rect 9428 4926 9464 4927
rect 9536 4926 9572 4927
rect 9638 4960 9675 4961
rect 9638 4959 9676 4960
rect 9638 4951 9702 4959
rect 9638 4931 9647 4951
rect 9667 4937 9702 4951
rect 9722 4937 9725 4957
rect 9667 4932 9725 4937
rect 9667 4931 9702 4932
rect 6830 4913 6895 4914
rect 4945 4835 4983 4836
rect 4544 4797 4983 4835
rect 5855 4835 5863 4857
rect 5887 4835 5895 4857
rect 5855 4827 5895 4835
rect 7166 4879 7206 4887
rect 7166 4857 7174 4879
rect 7198 4857 7206 4879
rect 8078 4879 8517 4917
rect 8078 4878 8116 4879
rect 6166 4800 6231 4801
rect 3372 4781 3407 4782
rect 3349 4776 3407 4781
rect 3349 4756 3352 4776
rect 3372 4762 3407 4776
rect 3427 4762 3436 4782
rect 3372 4754 3436 4762
rect 3398 4753 3436 4754
rect 3399 4752 3436 4753
rect 3502 4786 3538 4787
rect 3610 4786 3646 4787
rect 3502 4778 3646 4786
rect 3502 4758 3510 4778
rect 3530 4774 3618 4778
rect 3530 4758 3574 4774
rect 3502 4754 3574 4758
rect 3594 4758 3618 4774
rect 3638 4758 3646 4778
rect 3594 4754 3646 4758
rect 3502 4752 3646 4754
rect 3712 4782 3750 4790
rect 3828 4786 3864 4787
rect 3712 4762 3721 4782
rect 3741 4762 3750 4782
rect 3712 4753 3750 4762
rect 3779 4778 3864 4786
rect 3779 4758 3836 4778
rect 3856 4758 3864 4778
rect 3712 4752 3749 4753
rect 3779 4752 3864 4758
rect 3930 4782 3968 4790
rect 3930 4762 3939 4782
rect 3959 4762 3968 4782
rect 3930 4753 3968 4762
rect 4112 4787 4154 4796
rect 4112 4769 4126 4787
rect 4144 4769 4154 4787
rect 4112 4761 4154 4769
rect 4117 4759 4154 4761
rect 3930 4752 3967 4753
rect 3391 4724 3481 4730
rect 3391 4704 3407 4724
rect 3427 4722 3481 4724
rect 3427 4704 3452 4722
rect 3391 4702 3452 4704
rect 3472 4702 3481 4722
rect 3391 4696 3481 4702
rect 3404 4642 3441 4643
rect 3500 4642 3537 4643
rect 3556 4642 3592 4752
rect 3779 4731 3810 4752
rect 4544 4738 4591 4797
rect 4945 4796 4983 4797
rect 3775 4730 3810 4731
rect 3653 4720 3810 4730
rect 3653 4700 3670 4720
rect 3690 4700 3810 4720
rect 3653 4693 3810 4700
rect 3877 4723 4026 4731
rect 3877 4703 3888 4723
rect 3908 4703 3947 4723
rect 3967 4703 4026 4723
rect 4544 4720 4554 4738
rect 4572 4720 4591 4738
rect 4544 4716 4591 4720
rect 5817 4775 6004 4799
rect 6035 4780 6428 4800
rect 6448 4780 6451 4800
rect 6035 4775 6451 4780
rect 4545 4711 4582 4716
rect 3877 4696 4026 4703
rect 5817 4704 5854 4775
rect 6035 4774 6376 4775
rect 5969 4714 6000 4715
rect 3877 4695 3918 4696
rect 4114 4694 4151 4697
rect 3611 4642 3648 4643
rect 3304 4633 3442 4642
rect 2508 4594 2952 4620
rect 2508 4592 2676 4594
rect 2508 4414 2535 4592
rect 2575 4554 2639 4566
rect 2915 4562 2952 4594
rect 2978 4593 3169 4615
rect 3304 4613 3413 4633
rect 3433 4613 3442 4633
rect 3304 4606 3442 4613
rect 3500 4633 3648 4642
rect 3500 4613 3509 4633
rect 3529 4613 3619 4633
rect 3639 4613 3648 4633
rect 3304 4604 3400 4606
rect 3500 4603 3648 4613
rect 3707 4633 3744 4643
rect 3707 4613 3715 4633
rect 3735 4613 3744 4633
rect 3556 4602 3592 4603
rect 3133 4591 3169 4593
rect 3133 4562 3170 4591
rect 2575 4553 2610 4554
rect 2552 4548 2610 4553
rect 2552 4528 2555 4548
rect 2575 4534 2610 4548
rect 2630 4534 2639 4554
rect 2575 4528 2639 4534
rect 2552 4526 2639 4528
rect 2552 4522 2579 4526
rect 2601 4525 2639 4526
rect 2602 4524 2639 4525
rect 2705 4558 2741 4559
rect 2813 4558 2849 4559
rect 2705 4551 2849 4558
rect 2705 4550 2767 4551
rect 2705 4530 2713 4550
rect 2733 4533 2767 4550
rect 2786 4550 2849 4551
rect 2786 4533 2821 4550
rect 2733 4530 2821 4533
rect 2841 4530 2849 4550
rect 2705 4524 2849 4530
rect 2915 4554 2953 4562
rect 3031 4558 3067 4559
rect 2915 4534 2924 4554
rect 2944 4534 2953 4554
rect 2915 4525 2953 4534
rect 2982 4550 3067 4558
rect 2982 4530 3039 4550
rect 3059 4530 3067 4550
rect 2915 4524 2952 4525
rect 2982 4524 3067 4530
rect 3133 4554 3171 4562
rect 3133 4534 3142 4554
rect 3162 4534 3171 4554
rect 3404 4543 3441 4544
rect 3707 4543 3744 4613
rect 3779 4642 3810 4693
rect 4106 4688 4151 4694
rect 4106 4670 4124 4688
rect 4142 4670 4151 4688
rect 5817 4684 5826 4704
rect 5846 4684 5854 4704
rect 5817 4674 5854 4684
rect 5913 4704 6000 4714
rect 5913 4684 5922 4704
rect 5942 4684 6000 4704
rect 5913 4675 6000 4684
rect 5913 4674 5950 4675
rect 4106 4660 4151 4670
rect 3829 4642 3866 4643
rect 3779 4633 3866 4642
rect 3779 4613 3837 4633
rect 3857 4613 3866 4633
rect 3779 4603 3866 4613
rect 3925 4633 3962 4643
rect 3925 4613 3933 4633
rect 3953 4613 3962 4633
rect 4106 4618 4149 4660
rect 4533 4649 4585 4651
rect 4012 4616 4149 4618
rect 3779 4602 3810 4603
rect 3925 4543 3962 4613
rect 3403 4542 3744 4543
rect 3133 4525 3171 4534
rect 3328 4537 3744 4542
rect 3133 4524 3170 4525
rect 2594 4496 2684 4502
rect 2594 4476 2610 4496
rect 2630 4494 2684 4496
rect 2630 4476 2655 4494
rect 2594 4474 2655 4476
rect 2675 4474 2684 4494
rect 2594 4468 2684 4474
rect 2607 4414 2644 4415
rect 2703 4414 2740 4415
rect 2759 4414 2795 4524
rect 2982 4503 3013 4524
rect 3328 4517 3331 4537
rect 3351 4517 3744 4537
rect 3928 4527 3962 4543
rect 4006 4595 4149 4616
rect 4531 4645 4964 4649
rect 4531 4639 4970 4645
rect 4531 4621 4552 4639
rect 4570 4621 4970 4639
rect 5969 4624 6000 4675
rect 6035 4704 6072 4774
rect 6338 4773 6375 4774
rect 6187 4714 6223 4715
rect 6035 4684 6044 4704
rect 6064 4684 6072 4704
rect 6035 4674 6072 4684
rect 6131 4704 6279 4714
rect 6379 4711 6475 4713
rect 6131 4684 6140 4704
rect 6160 4684 6250 4704
rect 6270 4684 6279 4704
rect 6131 4675 6279 4684
rect 6337 4704 6475 4711
rect 6337 4684 6346 4704
rect 6366 4684 6475 4704
rect 6337 4675 6475 4684
rect 6131 4674 6168 4675
rect 5861 4621 5902 4622
rect 4531 4603 4970 4621
rect 3704 4508 3744 4517
rect 4006 4508 4033 4595
rect 4106 4569 4149 4595
rect 4106 4551 4119 4569
rect 4137 4551 4149 4569
rect 4106 4540 4149 4551
rect 2978 4502 3013 4503
rect 2856 4492 3013 4502
rect 2856 4472 2873 4492
rect 2893 4472 3013 4492
rect 2856 4465 3013 4472
rect 3080 4495 3226 4503
rect 3080 4475 3091 4495
rect 3111 4475 3150 4495
rect 3170 4475 3226 4495
rect 3704 4491 4033 4508
rect 3704 4490 3744 4491
rect 3080 4468 3226 4475
rect 4101 4479 4141 4482
rect 4101 4473 4144 4479
rect 3726 4470 4144 4473
rect 3080 4467 3121 4468
rect 2814 4414 2851 4415
rect 2507 4405 2645 4414
rect 2507 4385 2616 4405
rect 2636 4385 2645 4405
rect 2507 4378 2645 4385
rect 2703 4405 2851 4414
rect 2703 4385 2712 4405
rect 2732 4385 2822 4405
rect 2842 4385 2851 4405
rect 2507 4376 2603 4378
rect 2703 4375 2851 4385
rect 2910 4405 2947 4415
rect 2910 4385 2918 4405
rect 2938 4385 2947 4405
rect 2759 4374 2795 4375
rect 2607 4315 2644 4316
rect 2910 4315 2947 4385
rect 2982 4414 3013 4465
rect 3726 4452 4117 4470
rect 4135 4452 4144 4470
rect 3726 4450 4144 4452
rect 3726 4442 3753 4450
rect 3994 4447 4144 4450
rect 3306 4436 3474 4437
rect 3725 4436 3753 4442
rect 3306 4420 3753 4436
rect 4101 4442 4144 4447
rect 3032 4414 3069 4415
rect 2982 4405 3069 4414
rect 2982 4385 3040 4405
rect 3060 4385 3069 4405
rect 2982 4375 3069 4385
rect 3128 4405 3165 4415
rect 3128 4385 3136 4405
rect 3156 4385 3165 4405
rect 2982 4374 3013 4375
rect 2606 4314 2947 4315
rect 3128 4314 3165 4385
rect 2531 4309 2947 4314
rect 2531 4289 2534 4309
rect 2554 4289 2947 4309
rect 2978 4290 3165 4314
rect 3306 4410 3750 4420
rect 3306 4408 3474 4410
rect 2340 4215 2384 4216
rect 2340 4209 2385 4215
rect 2340 4191 2352 4209
rect 2374 4191 2385 4209
rect 2406 4210 2448 4255
rect 3306 4230 3333 4408
rect 3373 4370 3437 4382
rect 3713 4378 3750 4410
rect 3776 4409 3967 4431
rect 3931 4407 3967 4409
rect 3931 4378 3968 4407
rect 4101 4386 4141 4442
rect 3373 4369 3408 4370
rect 3350 4364 3408 4369
rect 3350 4344 3353 4364
rect 3373 4350 3408 4364
rect 3428 4350 3437 4370
rect 3373 4342 3437 4350
rect 3399 4341 3437 4342
rect 3400 4340 3437 4341
rect 3503 4374 3539 4375
rect 3611 4374 3647 4375
rect 3503 4366 3647 4374
rect 3503 4346 3511 4366
rect 3531 4346 3566 4366
rect 3586 4346 3619 4366
rect 3639 4346 3647 4366
rect 3503 4340 3647 4346
rect 3713 4370 3751 4378
rect 3829 4374 3865 4375
rect 3713 4350 3722 4370
rect 3742 4350 3751 4370
rect 3713 4341 3751 4350
rect 3780 4366 3865 4374
rect 3780 4346 3837 4366
rect 3857 4346 3865 4366
rect 3713 4340 3750 4341
rect 3780 4340 3865 4346
rect 3931 4370 3969 4378
rect 3931 4350 3940 4370
rect 3960 4350 3969 4370
rect 4101 4368 4113 4386
rect 4131 4368 4141 4386
rect 4533 4414 4585 4603
rect 4931 4578 4970 4603
rect 5753 4614 5902 4621
rect 5753 4594 5812 4614
rect 5832 4594 5871 4614
rect 5891 4594 5902 4614
rect 5753 4586 5902 4594
rect 5969 4617 6126 4624
rect 5969 4597 6089 4617
rect 6109 4597 6126 4617
rect 5969 4587 6126 4597
rect 5969 4586 6004 4587
rect 4715 4553 4902 4577
rect 4931 4558 5326 4578
rect 5346 4558 5349 4578
rect 5969 4565 6000 4586
rect 6187 4565 6223 4675
rect 6242 4674 6279 4675
rect 6338 4674 6375 4675
rect 6298 4615 6388 4621
rect 6298 4595 6307 4615
rect 6327 4613 6388 4615
rect 6327 4595 6352 4613
rect 6298 4593 6352 4595
rect 6372 4593 6388 4613
rect 6298 4587 6388 4593
rect 5812 4564 5849 4565
rect 4931 4553 5349 4558
rect 5811 4555 5849 4564
rect 4715 4482 4752 4553
rect 4931 4552 5274 4553
rect 4931 4549 4970 4552
rect 5236 4551 5273 4552
rect 4867 4492 4898 4493
rect 4715 4462 4724 4482
rect 4744 4462 4752 4482
rect 4715 4452 4752 4462
rect 4811 4482 4898 4492
rect 4811 4462 4820 4482
rect 4840 4462 4898 4482
rect 4811 4453 4898 4462
rect 4811 4452 4848 4453
rect 4533 4396 4549 4414
rect 4567 4396 4585 4414
rect 4867 4402 4898 4453
rect 4933 4482 4970 4549
rect 5811 4535 5820 4555
rect 5840 4535 5849 4555
rect 5811 4527 5849 4535
rect 5915 4559 6000 4565
rect 6030 4564 6067 4565
rect 5915 4539 5923 4559
rect 5943 4539 6000 4559
rect 5915 4531 6000 4539
rect 6029 4555 6067 4564
rect 6029 4535 6038 4555
rect 6058 4535 6067 4555
rect 5915 4530 5951 4531
rect 6029 4527 6067 4535
rect 6133 4559 6277 4565
rect 6133 4539 6141 4559
rect 6161 4553 6249 4559
rect 6161 4539 6190 4553
rect 6133 4531 6190 4539
rect 6133 4530 6169 4531
rect 6213 4539 6249 4553
rect 6269 4539 6277 4559
rect 6213 4531 6277 4539
rect 6241 4530 6277 4531
rect 6343 4564 6380 4565
rect 6343 4563 6381 4564
rect 6343 4555 6407 4563
rect 6343 4535 6352 4555
rect 6372 4541 6407 4555
rect 6427 4541 6430 4561
rect 6372 4536 6430 4541
rect 6372 4535 6407 4536
rect 5812 4498 5849 4527
rect 5813 4496 5849 4498
rect 5085 4492 5121 4493
rect 4933 4462 4942 4482
rect 4962 4462 4970 4482
rect 4933 4452 4970 4462
rect 5029 4482 5177 4492
rect 5277 4489 5373 4491
rect 5029 4462 5038 4482
rect 5058 4462 5148 4482
rect 5168 4462 5177 4482
rect 5029 4453 5177 4462
rect 5235 4482 5373 4489
rect 5235 4462 5244 4482
rect 5264 4462 5373 4482
rect 5813 4474 6004 4496
rect 6030 4495 6067 4527
rect 6343 4523 6407 4535
rect 6447 4497 6474 4675
rect 6771 4628 6808 4634
rect 6771 4609 6779 4628
rect 6800 4609 6808 4628
rect 6771 4601 6808 4609
rect 6306 4495 6474 4497
rect 6030 4469 6474 4495
rect 6140 4467 6180 4469
rect 6306 4468 6474 4469
rect 5235 4453 5373 4462
rect 6433 4463 6474 4468
rect 5029 4452 5066 4453
rect 4759 4399 4800 4400
rect 4533 4378 4585 4396
rect 4651 4392 4800 4399
rect 4101 4358 4141 4368
rect 4651 4372 4710 4392
rect 4730 4372 4769 4392
rect 4789 4372 4800 4392
rect 4651 4364 4800 4372
rect 4867 4395 5024 4402
rect 4867 4375 4987 4395
rect 5007 4375 5024 4395
rect 4867 4365 5024 4375
rect 4867 4364 4902 4365
rect 3931 4341 3969 4350
rect 4867 4343 4898 4364
rect 5085 4343 5121 4453
rect 5140 4452 5177 4453
rect 5236 4452 5273 4453
rect 5196 4393 5286 4399
rect 5196 4373 5205 4393
rect 5225 4391 5286 4393
rect 5225 4373 5250 4391
rect 5196 4371 5250 4373
rect 5270 4371 5286 4391
rect 5196 4365 5286 4371
rect 4710 4342 4747 4343
rect 3931 4340 3968 4341
rect 3392 4312 3482 4318
rect 3392 4292 3408 4312
rect 3428 4310 3482 4312
rect 3428 4292 3453 4310
rect 3392 4290 3453 4292
rect 3473 4290 3482 4310
rect 3392 4284 3482 4290
rect 3405 4230 3442 4231
rect 3501 4230 3538 4231
rect 3557 4230 3593 4340
rect 3780 4319 3811 4340
rect 4709 4333 4747 4342
rect 3776 4318 3811 4319
rect 3654 4308 3811 4318
rect 3654 4288 3671 4308
rect 3691 4288 3811 4308
rect 3654 4281 3811 4288
rect 3878 4311 4027 4319
rect 3878 4291 3889 4311
rect 3909 4291 3948 4311
rect 3968 4291 4027 4311
rect 4537 4315 4577 4325
rect 3878 4284 4027 4291
rect 4093 4287 4145 4305
rect 3878 4283 3919 4284
rect 3612 4230 3649 4231
rect 3305 4221 3443 4230
rect 2777 4210 2810 4212
rect 2406 4198 2853 4210
rect 2340 4161 2385 4191
rect 2357 3215 2385 4161
rect 2409 4184 2853 4198
rect 2409 4182 2577 4184
rect 2409 4004 2436 4182
rect 2476 4144 2540 4156
rect 2816 4152 2853 4184
rect 2879 4183 3070 4205
rect 3305 4201 3414 4221
rect 3434 4201 3443 4221
rect 3305 4194 3443 4201
rect 3501 4221 3649 4230
rect 3501 4201 3510 4221
rect 3530 4201 3620 4221
rect 3640 4201 3649 4221
rect 3305 4192 3401 4194
rect 3501 4191 3649 4201
rect 3708 4221 3745 4231
rect 3708 4201 3716 4221
rect 3736 4201 3745 4221
rect 3557 4190 3593 4191
rect 3034 4181 3070 4183
rect 3034 4152 3071 4181
rect 2476 4143 2511 4144
rect 2453 4138 2511 4143
rect 2453 4118 2456 4138
rect 2476 4124 2511 4138
rect 2531 4124 2540 4144
rect 2476 4116 2540 4124
rect 2502 4115 2540 4116
rect 2503 4114 2540 4115
rect 2606 4148 2642 4149
rect 2714 4148 2750 4149
rect 2606 4142 2750 4148
rect 2606 4140 2667 4142
rect 2606 4120 2614 4140
rect 2634 4125 2667 4140
rect 2686 4140 2750 4142
rect 2686 4125 2722 4140
rect 2634 4120 2722 4125
rect 2742 4120 2750 4140
rect 2606 4114 2750 4120
rect 2816 4144 2854 4152
rect 2932 4148 2968 4149
rect 2816 4124 2825 4144
rect 2845 4124 2854 4144
rect 2816 4115 2854 4124
rect 2883 4140 2968 4148
rect 2883 4120 2940 4140
rect 2960 4120 2968 4140
rect 2816 4114 2853 4115
rect 2883 4114 2968 4120
rect 3034 4144 3072 4152
rect 3034 4124 3043 4144
rect 3063 4124 3072 4144
rect 3708 4134 3745 4201
rect 3780 4230 3811 4281
rect 4093 4269 4111 4287
rect 4129 4269 4145 4287
rect 3830 4230 3867 4231
rect 3780 4221 3867 4230
rect 3780 4201 3838 4221
rect 3858 4201 3867 4221
rect 3780 4191 3867 4201
rect 3926 4221 3963 4231
rect 3926 4201 3934 4221
rect 3954 4201 3963 4221
rect 3780 4190 3811 4191
rect 3405 4131 3442 4132
rect 3708 4131 3747 4134
rect 3404 4130 3747 4131
rect 3926 4130 3963 4201
rect 3034 4115 3072 4124
rect 3329 4125 3747 4130
rect 3034 4114 3071 4115
rect 2495 4086 2585 4092
rect 2495 4066 2511 4086
rect 2531 4084 2585 4086
rect 2531 4066 2556 4084
rect 2495 4064 2556 4066
rect 2576 4064 2585 4084
rect 2495 4058 2585 4064
rect 2508 4004 2545 4005
rect 2604 4004 2641 4005
rect 2660 4004 2696 4114
rect 2883 4093 2914 4114
rect 3329 4105 3332 4125
rect 3352 4105 3747 4125
rect 3776 4106 3963 4130
rect 2879 4092 2914 4093
rect 2757 4082 2914 4092
rect 2757 4062 2774 4082
rect 2794 4062 2914 4082
rect 2757 4055 2914 4062
rect 2981 4085 3130 4093
rect 2981 4065 2992 4085
rect 3012 4065 3051 4085
rect 3071 4065 3130 4085
rect 2981 4058 3130 4065
rect 3708 4080 3747 4105
rect 4093 4080 4145 4269
rect 4537 4297 4547 4315
rect 4565 4297 4577 4315
rect 4709 4313 4718 4333
rect 4738 4313 4747 4333
rect 4709 4305 4747 4313
rect 4813 4337 4898 4343
rect 4928 4342 4965 4343
rect 4813 4317 4821 4337
rect 4841 4317 4898 4337
rect 4813 4309 4898 4317
rect 4927 4333 4965 4342
rect 4927 4313 4936 4333
rect 4956 4313 4965 4333
rect 4813 4308 4849 4309
rect 4927 4305 4965 4313
rect 5031 4337 5175 4343
rect 5031 4317 5039 4337
rect 5059 4317 5092 4337
rect 5112 4317 5147 4337
rect 5167 4317 5175 4337
rect 5031 4309 5175 4317
rect 5031 4308 5067 4309
rect 5139 4308 5175 4309
rect 5241 4342 5278 4343
rect 5241 4341 5279 4342
rect 5241 4333 5305 4341
rect 5241 4313 5250 4333
rect 5270 4319 5305 4333
rect 5325 4319 5328 4339
rect 5270 4314 5328 4319
rect 5270 4313 5305 4314
rect 4537 4241 4577 4297
rect 4710 4276 4747 4305
rect 4711 4274 4747 4276
rect 4711 4252 4902 4274
rect 4928 4273 4965 4305
rect 5241 4301 5305 4313
rect 5345 4275 5372 4453
rect 5204 4273 5372 4275
rect 4928 4263 5372 4273
rect 5513 4369 5700 4393
rect 5731 4374 6124 4394
rect 6144 4374 6147 4394
rect 5731 4369 6147 4374
rect 5513 4298 5550 4369
rect 5731 4368 6072 4369
rect 5665 4308 5696 4309
rect 5513 4278 5522 4298
rect 5542 4278 5550 4298
rect 5513 4268 5550 4278
rect 5609 4298 5696 4308
rect 5609 4278 5618 4298
rect 5638 4278 5696 4298
rect 5609 4269 5696 4278
rect 5609 4268 5646 4269
rect 4534 4236 4577 4241
rect 4925 4247 5372 4263
rect 4925 4241 4953 4247
rect 5204 4246 5372 4247
rect 4534 4233 4684 4236
rect 4925 4233 4952 4241
rect 4534 4231 4952 4233
rect 4534 4213 4543 4231
rect 4561 4213 4952 4231
rect 5665 4218 5696 4269
rect 5731 4298 5768 4368
rect 6034 4367 6071 4368
rect 5883 4308 5919 4309
rect 5731 4278 5740 4298
rect 5760 4278 5768 4298
rect 5731 4268 5768 4278
rect 5827 4298 5975 4308
rect 6075 4305 6171 4307
rect 5827 4278 5836 4298
rect 5856 4278 5946 4298
rect 5966 4278 5975 4298
rect 5827 4269 5975 4278
rect 6033 4298 6171 4305
rect 6033 4278 6042 4298
rect 6062 4278 6171 4298
rect 6433 4281 6473 4463
rect 6033 4269 6171 4278
rect 5827 4268 5864 4269
rect 5557 4215 5598 4216
rect 4534 4210 4952 4213
rect 4534 4204 4577 4210
rect 4537 4201 4577 4204
rect 5449 4208 5598 4215
rect 4934 4192 4974 4193
rect 4645 4175 4974 4192
rect 5449 4188 5508 4208
rect 5528 4188 5567 4208
rect 5587 4188 5598 4208
rect 5449 4180 5598 4188
rect 5665 4211 5822 4218
rect 5665 4191 5785 4211
rect 5805 4191 5822 4211
rect 5665 4181 5822 4191
rect 5665 4180 5700 4181
rect 4529 4132 4572 4143
rect 4529 4114 4541 4132
rect 4559 4114 4572 4132
rect 4529 4088 4572 4114
rect 4645 4088 4672 4175
rect 4934 4166 4974 4175
rect 3708 4062 4147 4080
rect 2981 4057 3022 4058
rect 2715 4004 2752 4005
rect 2408 3995 2546 4004
rect 2408 3975 2517 3995
rect 2537 3975 2546 3995
rect 2408 3968 2546 3975
rect 2604 3995 2752 4004
rect 2604 3975 2613 3995
rect 2633 3975 2723 3995
rect 2743 3975 2752 3995
rect 2408 3966 2504 3968
rect 2604 3965 2752 3975
rect 2811 3995 2848 4005
rect 2811 3975 2819 3995
rect 2839 3975 2848 3995
rect 2660 3964 2696 3965
rect 2508 3905 2545 3906
rect 2811 3905 2848 3975
rect 2883 4004 2914 4055
rect 3708 4044 4108 4062
rect 4126 4044 4147 4062
rect 3708 4038 4147 4044
rect 3714 4034 4147 4038
rect 4529 4067 4672 4088
rect 4716 4140 4750 4156
rect 4934 4146 5327 4166
rect 5347 4146 5350 4166
rect 5665 4159 5696 4180
rect 5883 4159 5919 4269
rect 5938 4268 5975 4269
rect 6034 4268 6071 4269
rect 5994 4209 6084 4215
rect 5994 4189 6003 4209
rect 6023 4207 6084 4209
rect 6023 4189 6048 4207
rect 5994 4187 6048 4189
rect 6068 4187 6084 4207
rect 5994 4181 6084 4187
rect 5508 4158 5545 4159
rect 4934 4141 5350 4146
rect 5507 4149 5545 4158
rect 4934 4140 5275 4141
rect 4716 4070 4753 4140
rect 4868 4080 4899 4081
rect 4529 4065 4666 4067
rect 4093 4032 4145 4034
rect 4529 4023 4572 4065
rect 4716 4050 4725 4070
rect 4745 4050 4753 4070
rect 4716 4040 4753 4050
rect 4812 4070 4899 4080
rect 4812 4050 4821 4070
rect 4841 4050 4899 4070
rect 4812 4041 4899 4050
rect 4812 4040 4849 4041
rect 4527 4013 4572 4023
rect 2933 4004 2970 4005
rect 2883 3995 2970 4004
rect 2883 3975 2941 3995
rect 2961 3975 2970 3995
rect 2883 3965 2970 3975
rect 3029 3995 3066 4005
rect 3029 3975 3037 3995
rect 3057 3975 3066 3995
rect 4527 3995 4536 4013
rect 4554 3995 4572 4013
rect 4527 3989 4572 3995
rect 4868 3990 4899 4041
rect 4934 4070 4971 4140
rect 5237 4139 5274 4140
rect 5507 4129 5516 4149
rect 5536 4129 5545 4149
rect 5507 4121 5545 4129
rect 5611 4153 5696 4159
rect 5726 4158 5763 4159
rect 5611 4133 5619 4153
rect 5639 4133 5696 4153
rect 5611 4125 5696 4133
rect 5725 4149 5763 4158
rect 5725 4129 5734 4149
rect 5754 4129 5763 4149
rect 5611 4124 5647 4125
rect 5725 4121 5763 4129
rect 5829 4153 5973 4159
rect 5829 4133 5837 4153
rect 5857 4134 5889 4153
rect 5910 4134 5945 4153
rect 5857 4133 5945 4134
rect 5965 4133 5973 4153
rect 5829 4125 5973 4133
rect 5829 4124 5865 4125
rect 5937 4124 5973 4125
rect 6039 4158 6076 4159
rect 6039 4157 6077 4158
rect 6039 4149 6103 4157
rect 6039 4129 6048 4149
rect 6068 4135 6103 4149
rect 6123 4135 6126 4155
rect 6068 4130 6126 4135
rect 6068 4129 6103 4130
rect 5508 4092 5545 4121
rect 5509 4090 5545 4092
rect 5086 4080 5122 4081
rect 4934 4050 4943 4070
rect 4963 4050 4971 4070
rect 4934 4040 4971 4050
rect 5030 4070 5178 4080
rect 5278 4077 5374 4079
rect 5030 4050 5039 4070
rect 5059 4050 5149 4070
rect 5169 4050 5178 4070
rect 5030 4041 5178 4050
rect 5236 4070 5374 4077
rect 5236 4050 5245 4070
rect 5265 4050 5374 4070
rect 5509 4068 5700 4090
rect 5726 4089 5763 4121
rect 6039 4117 6103 4129
rect 6143 4091 6170 4269
rect 6002 4089 6170 4091
rect 5726 4063 6170 4089
rect 5236 4041 5374 4050
rect 5030 4040 5067 4041
rect 4527 3986 4564 3989
rect 4760 3987 4801 3988
rect 2883 3964 2914 3965
rect 2507 3904 2848 3905
rect 3029 3904 3066 3975
rect 4652 3980 4801 3987
rect 4096 3967 4133 3972
rect 4087 3963 4134 3967
rect 4087 3945 4106 3963
rect 4124 3945 4134 3963
rect 4652 3960 4711 3980
rect 4731 3960 4770 3980
rect 4790 3960 4801 3980
rect 4652 3952 4801 3960
rect 4868 3983 5025 3990
rect 4868 3963 4988 3983
rect 5008 3963 5025 3983
rect 4868 3953 5025 3963
rect 4868 3952 4903 3953
rect 2432 3899 2848 3904
rect 2432 3879 2435 3899
rect 2455 3879 2848 3899
rect 2879 3880 3066 3904
rect 3691 3902 3731 3907
rect 4087 3902 4134 3945
rect 4868 3931 4899 3952
rect 5086 3931 5122 4041
rect 5141 4040 5178 4041
rect 5237 4040 5274 4041
rect 5197 3981 5287 3987
rect 5197 3961 5206 3981
rect 5226 3979 5287 3981
rect 5226 3961 5251 3979
rect 5197 3959 5251 3961
rect 5271 3959 5287 3979
rect 5197 3953 5287 3959
rect 4711 3930 4748 3931
rect 3691 3863 4134 3902
rect 4524 3922 4561 3924
rect 4524 3914 4566 3922
rect 4524 3896 4534 3914
rect 4552 3896 4566 3914
rect 4524 3887 4566 3896
rect 4710 3921 4748 3930
rect 4710 3901 4719 3921
rect 4739 3901 4748 3921
rect 4710 3893 4748 3901
rect 4814 3925 4899 3931
rect 4929 3930 4966 3931
rect 4814 3905 4822 3925
rect 4842 3905 4899 3925
rect 4814 3897 4899 3905
rect 4928 3921 4966 3930
rect 4928 3901 4937 3921
rect 4957 3901 4966 3921
rect 4814 3896 4850 3897
rect 4928 3893 4966 3901
rect 5032 3929 5176 3931
rect 5032 3925 5084 3929
rect 5032 3905 5040 3925
rect 5060 3909 5084 3925
rect 5104 3925 5176 3929
rect 5104 3909 5148 3925
rect 5060 3905 5148 3909
rect 5168 3905 5176 3925
rect 5032 3897 5176 3905
rect 5032 3896 5068 3897
rect 5140 3896 5176 3897
rect 5242 3930 5279 3931
rect 5242 3929 5280 3930
rect 5242 3921 5306 3929
rect 5242 3901 5251 3921
rect 5271 3907 5306 3921
rect 5326 3907 5329 3927
rect 5271 3902 5329 3907
rect 5271 3901 5306 3902
rect 2785 3848 2825 3856
rect 2785 3826 2793 3848
rect 2817 3826 2825 3848
rect 2491 3602 2659 3603
rect 2785 3602 2825 3826
rect 3288 3830 3456 3831
rect 3691 3830 3731 3863
rect 4087 3830 4134 3863
rect 4525 3862 4566 3887
rect 4711 3862 4748 3893
rect 4929 3862 4966 3893
rect 5242 3889 5306 3901
rect 5346 3863 5373 4041
rect 4525 3835 4574 3862
rect 4710 3836 4759 3862
rect 4928 3861 5009 3862
rect 5205 3861 5373 3863
rect 4928 3836 5373 3861
rect 4929 3835 5373 3836
rect 3288 3829 3732 3830
rect 3288 3804 3733 3829
rect 3288 3802 3456 3804
rect 3652 3803 3733 3804
rect 3902 3803 3951 3829
rect 4087 3803 4136 3830
rect 3288 3624 3315 3802
rect 3355 3764 3419 3776
rect 3695 3772 3732 3803
rect 3913 3772 3950 3803
rect 4095 3778 4136 3803
rect 4527 3802 4574 3835
rect 4930 3802 4970 3835
rect 5205 3834 5373 3835
rect 5836 3839 5876 4063
rect 6002 4062 6170 4063
rect 5836 3817 5844 3839
rect 5868 3817 5876 3839
rect 5836 3809 5876 3817
rect 3355 3763 3390 3764
rect 3332 3758 3390 3763
rect 3332 3738 3335 3758
rect 3355 3744 3390 3758
rect 3410 3744 3419 3764
rect 3355 3736 3419 3744
rect 3381 3735 3419 3736
rect 3382 3734 3419 3735
rect 3485 3768 3521 3769
rect 3593 3768 3629 3769
rect 3485 3760 3629 3768
rect 3485 3740 3493 3760
rect 3513 3756 3601 3760
rect 3513 3740 3557 3756
rect 3485 3736 3557 3740
rect 3577 3740 3601 3756
rect 3621 3740 3629 3760
rect 3577 3736 3629 3740
rect 3485 3734 3629 3736
rect 3695 3764 3733 3772
rect 3811 3768 3847 3769
rect 3695 3744 3704 3764
rect 3724 3744 3733 3764
rect 3695 3735 3733 3744
rect 3762 3760 3847 3768
rect 3762 3740 3819 3760
rect 3839 3740 3847 3760
rect 3695 3734 3732 3735
rect 3762 3734 3847 3740
rect 3913 3764 3951 3772
rect 3913 3744 3922 3764
rect 3942 3744 3951 3764
rect 3913 3735 3951 3744
rect 4095 3769 4137 3778
rect 4095 3751 4109 3769
rect 4127 3751 4137 3769
rect 4095 3743 4137 3751
rect 4100 3741 4137 3743
rect 4527 3763 4970 3802
rect 3913 3734 3950 3735
rect 3374 3706 3464 3712
rect 3374 3686 3390 3706
rect 3410 3704 3464 3706
rect 3410 3686 3435 3704
rect 3374 3684 3435 3686
rect 3455 3684 3464 3704
rect 3374 3678 3464 3684
rect 3387 3624 3424 3625
rect 3483 3624 3520 3625
rect 3539 3624 3575 3734
rect 3762 3713 3793 3734
rect 4527 3720 4574 3763
rect 4930 3758 4970 3763
rect 5595 3761 5782 3785
rect 5813 3766 6206 3786
rect 6226 3766 6229 3786
rect 5813 3761 6229 3766
rect 3758 3712 3793 3713
rect 3636 3702 3793 3712
rect 3636 3682 3653 3702
rect 3673 3682 3793 3702
rect 3636 3675 3793 3682
rect 3860 3705 4009 3713
rect 3860 3685 3871 3705
rect 3891 3685 3930 3705
rect 3950 3685 4009 3705
rect 4527 3702 4537 3720
rect 4555 3702 4574 3720
rect 4527 3698 4574 3702
rect 4528 3693 4565 3698
rect 3860 3678 4009 3685
rect 5595 3690 5632 3761
rect 5813 3760 6154 3761
rect 5747 3700 5778 3701
rect 3860 3677 3901 3678
rect 4097 3676 4134 3679
rect 3594 3624 3631 3625
rect 3287 3615 3425 3624
rect 2491 3576 2935 3602
rect 2491 3574 2659 3576
rect 2491 3396 2518 3574
rect 2558 3536 2622 3548
rect 2898 3544 2935 3576
rect 2961 3575 3152 3597
rect 3287 3595 3396 3615
rect 3416 3595 3425 3615
rect 3287 3588 3425 3595
rect 3483 3615 3631 3624
rect 3483 3595 3492 3615
rect 3512 3595 3602 3615
rect 3622 3595 3631 3615
rect 3287 3586 3383 3588
rect 3483 3585 3631 3595
rect 3690 3615 3727 3625
rect 3690 3595 3698 3615
rect 3718 3595 3727 3615
rect 3539 3584 3575 3585
rect 3116 3573 3152 3575
rect 3116 3544 3153 3573
rect 2558 3535 2593 3536
rect 2535 3530 2593 3535
rect 2535 3510 2538 3530
rect 2558 3516 2593 3530
rect 2613 3516 2622 3536
rect 2558 3508 2622 3516
rect 2584 3507 2622 3508
rect 2585 3506 2622 3507
rect 2688 3540 2724 3541
rect 2796 3540 2832 3541
rect 2688 3532 2832 3540
rect 2688 3512 2696 3532
rect 2716 3531 2804 3532
rect 2716 3512 2751 3531
rect 2772 3512 2804 3531
rect 2824 3512 2832 3532
rect 2688 3506 2832 3512
rect 2898 3536 2936 3544
rect 3014 3540 3050 3541
rect 2898 3516 2907 3536
rect 2927 3516 2936 3536
rect 2898 3507 2936 3516
rect 2965 3532 3050 3540
rect 2965 3512 3022 3532
rect 3042 3512 3050 3532
rect 2898 3506 2935 3507
rect 2965 3506 3050 3512
rect 3116 3536 3154 3544
rect 3116 3516 3125 3536
rect 3145 3516 3154 3536
rect 3387 3525 3424 3526
rect 3690 3525 3727 3595
rect 3762 3624 3793 3675
rect 4089 3670 4134 3676
rect 4089 3652 4107 3670
rect 4125 3652 4134 3670
rect 5595 3670 5604 3690
rect 5624 3670 5632 3690
rect 5595 3660 5632 3670
rect 5691 3690 5778 3700
rect 5691 3670 5700 3690
rect 5720 3670 5778 3690
rect 5691 3661 5778 3670
rect 5691 3660 5728 3661
rect 4089 3642 4134 3652
rect 3812 3624 3849 3625
rect 3762 3615 3849 3624
rect 3762 3595 3820 3615
rect 3840 3595 3849 3615
rect 3762 3585 3849 3595
rect 3908 3615 3945 3625
rect 3908 3595 3916 3615
rect 3936 3595 3945 3615
rect 4089 3600 4132 3642
rect 4516 3631 4568 3633
rect 3995 3598 4132 3600
rect 3762 3584 3793 3585
rect 3908 3525 3945 3595
rect 3386 3524 3727 3525
rect 3116 3507 3154 3516
rect 3311 3519 3727 3524
rect 3116 3506 3153 3507
rect 2577 3478 2667 3484
rect 2577 3458 2593 3478
rect 2613 3476 2667 3478
rect 2613 3458 2638 3476
rect 2577 3456 2638 3458
rect 2658 3456 2667 3476
rect 2577 3450 2667 3456
rect 2590 3396 2627 3397
rect 2686 3396 2723 3397
rect 2742 3396 2778 3506
rect 2965 3485 2996 3506
rect 3311 3499 3314 3519
rect 3334 3499 3727 3519
rect 3911 3509 3945 3525
rect 3989 3577 4132 3598
rect 4514 3627 4947 3631
rect 4514 3621 4953 3627
rect 4514 3603 4535 3621
rect 4553 3603 4953 3621
rect 5747 3610 5778 3661
rect 5813 3690 5850 3760
rect 6116 3759 6153 3760
rect 5965 3700 6001 3701
rect 5813 3670 5822 3690
rect 5842 3670 5850 3690
rect 5813 3660 5850 3670
rect 5909 3690 6057 3700
rect 6157 3697 6253 3699
rect 5909 3670 5918 3690
rect 5938 3670 6028 3690
rect 6048 3670 6057 3690
rect 5909 3661 6057 3670
rect 6115 3690 6253 3697
rect 6115 3670 6124 3690
rect 6144 3670 6253 3690
rect 6115 3661 6253 3670
rect 5909 3660 5946 3661
rect 5639 3607 5680 3608
rect 4514 3585 4953 3603
rect 3687 3490 3727 3499
rect 3989 3490 4016 3577
rect 4089 3551 4132 3577
rect 4089 3533 4102 3551
rect 4120 3533 4132 3551
rect 4089 3522 4132 3533
rect 2961 3484 2996 3485
rect 2839 3474 2996 3484
rect 2839 3454 2856 3474
rect 2876 3454 2996 3474
rect 2839 3447 2996 3454
rect 3063 3477 3212 3485
rect 3063 3457 3074 3477
rect 3094 3457 3133 3477
rect 3153 3457 3212 3477
rect 3687 3473 4016 3490
rect 3687 3472 3727 3473
rect 3063 3450 3212 3457
rect 4084 3461 4124 3464
rect 4084 3455 4127 3461
rect 3709 3452 4127 3455
rect 3063 3449 3104 3450
rect 2797 3396 2834 3397
rect 2490 3387 2628 3396
rect 2490 3367 2599 3387
rect 2619 3367 2628 3387
rect 2490 3360 2628 3367
rect 2686 3387 2834 3396
rect 2686 3367 2695 3387
rect 2715 3367 2805 3387
rect 2825 3367 2834 3387
rect 2490 3358 2586 3360
rect 2686 3357 2834 3367
rect 2893 3387 2930 3397
rect 2893 3367 2901 3387
rect 2921 3367 2930 3387
rect 2742 3356 2778 3357
rect 2590 3297 2627 3298
rect 2893 3297 2930 3367
rect 2965 3396 2996 3447
rect 3709 3434 4100 3452
rect 4118 3434 4127 3452
rect 3709 3432 4127 3434
rect 3709 3424 3736 3432
rect 3977 3429 4127 3432
rect 3289 3418 3457 3419
rect 3708 3418 3736 3424
rect 3289 3402 3736 3418
rect 4084 3424 4127 3429
rect 3015 3396 3052 3397
rect 2965 3387 3052 3396
rect 2965 3367 3023 3387
rect 3043 3367 3052 3387
rect 2965 3357 3052 3367
rect 3111 3387 3148 3397
rect 3111 3367 3119 3387
rect 3139 3367 3148 3387
rect 2965 3356 2996 3357
rect 2589 3296 2930 3297
rect 3111 3296 3148 3367
rect 2514 3291 2930 3296
rect 2514 3271 2517 3291
rect 2537 3271 2930 3291
rect 2961 3272 3148 3296
rect 3289 3392 3733 3402
rect 3289 3390 3457 3392
rect 2356 3197 2385 3215
rect 3289 3212 3316 3390
rect 3356 3352 3420 3364
rect 3696 3360 3733 3392
rect 3759 3391 3950 3413
rect 3914 3389 3950 3391
rect 3914 3360 3951 3389
rect 4084 3368 4124 3424
rect 3356 3351 3391 3352
rect 3333 3346 3391 3351
rect 3333 3326 3336 3346
rect 3356 3332 3391 3346
rect 3411 3332 3420 3352
rect 3356 3324 3420 3332
rect 3382 3323 3420 3324
rect 3383 3322 3420 3323
rect 3486 3356 3522 3357
rect 3594 3356 3630 3357
rect 3486 3348 3630 3356
rect 3486 3328 3494 3348
rect 3514 3328 3549 3348
rect 3569 3328 3602 3348
rect 3622 3328 3630 3348
rect 3486 3322 3630 3328
rect 3696 3352 3734 3360
rect 3812 3356 3848 3357
rect 3696 3332 3705 3352
rect 3725 3332 3734 3352
rect 3696 3323 3734 3332
rect 3763 3348 3848 3356
rect 3763 3328 3820 3348
rect 3840 3328 3848 3348
rect 3696 3322 3733 3323
rect 3763 3322 3848 3328
rect 3914 3352 3952 3360
rect 3914 3332 3923 3352
rect 3943 3332 3952 3352
rect 4084 3350 4096 3368
rect 4114 3350 4124 3368
rect 4516 3396 4568 3585
rect 4914 3560 4953 3585
rect 5531 3600 5680 3607
rect 5531 3580 5590 3600
rect 5610 3580 5649 3600
rect 5669 3580 5680 3600
rect 5531 3572 5680 3580
rect 5747 3603 5904 3610
rect 5747 3583 5867 3603
rect 5887 3583 5904 3603
rect 5747 3573 5904 3583
rect 5747 3572 5782 3573
rect 4698 3535 4885 3559
rect 4914 3540 5309 3560
rect 5329 3540 5332 3560
rect 5747 3551 5778 3572
rect 5965 3551 6001 3661
rect 6020 3660 6057 3661
rect 6116 3660 6153 3661
rect 6076 3601 6166 3607
rect 6076 3581 6085 3601
rect 6105 3599 6166 3601
rect 6105 3581 6130 3599
rect 6076 3579 6130 3581
rect 6150 3579 6166 3599
rect 6076 3573 6166 3579
rect 5590 3550 5627 3551
rect 4914 3535 5332 3540
rect 5589 3541 5627 3550
rect 4698 3464 4735 3535
rect 4914 3534 5257 3535
rect 4914 3531 4953 3534
rect 5219 3533 5256 3534
rect 4850 3474 4881 3475
rect 4698 3444 4707 3464
rect 4727 3444 4735 3464
rect 4698 3434 4735 3444
rect 4794 3464 4881 3474
rect 4794 3444 4803 3464
rect 4823 3444 4881 3464
rect 4794 3435 4881 3444
rect 4794 3434 4831 3435
rect 4516 3378 4532 3396
rect 4550 3378 4568 3396
rect 4850 3384 4881 3435
rect 4916 3464 4953 3531
rect 5589 3521 5598 3541
rect 5618 3521 5627 3541
rect 5589 3513 5627 3521
rect 5693 3545 5778 3551
rect 5808 3550 5845 3551
rect 5693 3525 5701 3545
rect 5721 3525 5778 3545
rect 5693 3517 5778 3525
rect 5807 3541 5845 3550
rect 5807 3521 5816 3541
rect 5836 3521 5845 3541
rect 5693 3516 5729 3517
rect 5807 3513 5845 3521
rect 5911 3546 6055 3551
rect 5911 3545 5973 3546
rect 5911 3525 5919 3545
rect 5939 3527 5973 3545
rect 5994 3545 6055 3546
rect 5994 3527 6027 3545
rect 5939 3525 6027 3527
rect 6047 3525 6055 3545
rect 5911 3517 6055 3525
rect 5911 3516 5947 3517
rect 6019 3516 6055 3517
rect 6121 3550 6158 3551
rect 6121 3549 6159 3550
rect 6121 3541 6185 3549
rect 6121 3521 6130 3541
rect 6150 3527 6185 3541
rect 6205 3527 6208 3547
rect 6150 3522 6208 3527
rect 6150 3521 6185 3522
rect 5590 3484 5627 3513
rect 5591 3482 5627 3484
rect 5068 3474 5104 3475
rect 4916 3444 4925 3464
rect 4945 3444 4953 3464
rect 4916 3434 4953 3444
rect 5012 3464 5160 3474
rect 5260 3471 5356 3473
rect 5012 3444 5021 3464
rect 5041 3444 5131 3464
rect 5151 3444 5160 3464
rect 5012 3435 5160 3444
rect 5218 3464 5356 3471
rect 5218 3444 5227 3464
rect 5247 3444 5356 3464
rect 5591 3460 5782 3482
rect 5808 3481 5845 3513
rect 6121 3509 6185 3521
rect 6225 3483 6252 3661
rect 6084 3481 6252 3483
rect 5808 3467 6252 3481
rect 5808 3455 6255 3467
rect 5851 3453 5884 3455
rect 5218 3435 5356 3444
rect 5012 3434 5049 3435
rect 4742 3381 4783 3382
rect 4516 3360 4568 3378
rect 4634 3374 4783 3381
rect 4084 3340 4124 3350
rect 4634 3354 4693 3374
rect 4713 3354 4752 3374
rect 4772 3354 4783 3374
rect 4634 3346 4783 3354
rect 4850 3377 5007 3384
rect 4850 3357 4970 3377
rect 4990 3357 5007 3377
rect 4850 3347 5007 3357
rect 4850 3346 4885 3347
rect 3914 3323 3952 3332
rect 4850 3325 4881 3346
rect 5068 3325 5104 3435
rect 5123 3434 5160 3435
rect 5219 3434 5256 3435
rect 5179 3375 5269 3381
rect 5179 3355 5188 3375
rect 5208 3373 5269 3375
rect 5208 3355 5233 3373
rect 5179 3353 5233 3355
rect 5253 3353 5269 3373
rect 5179 3347 5269 3353
rect 4693 3324 4730 3325
rect 3914 3322 3951 3323
rect 3375 3294 3465 3300
rect 3375 3274 3391 3294
rect 3411 3292 3465 3294
rect 3411 3274 3436 3292
rect 3375 3272 3436 3274
rect 3456 3272 3465 3292
rect 3375 3266 3465 3272
rect 3388 3212 3425 3213
rect 3484 3212 3521 3213
rect 3540 3212 3576 3322
rect 3763 3301 3794 3322
rect 4692 3315 4730 3324
rect 3759 3300 3794 3301
rect 3637 3290 3794 3300
rect 3637 3270 3654 3290
rect 3674 3270 3794 3290
rect 3637 3263 3794 3270
rect 3861 3293 4010 3301
rect 3861 3273 3872 3293
rect 3892 3273 3931 3293
rect 3951 3273 4010 3293
rect 4520 3297 4560 3307
rect 3861 3266 4010 3273
rect 4076 3269 4128 3287
rect 3861 3265 3902 3266
rect 3595 3212 3632 3213
rect 2326 3195 2385 3197
rect 3288 3203 3426 3212
rect 2326 3194 2494 3195
rect 2620 3194 2660 3196
rect 2326 3168 2770 3194
rect 2326 3166 2494 3168
rect 2326 3164 2407 3166
rect 2326 2988 2353 3164
rect 2393 3128 2457 3140
rect 2733 3136 2770 3168
rect 2796 3167 2987 3189
rect 3288 3183 3397 3203
rect 3417 3183 3426 3203
rect 3288 3176 3426 3183
rect 3484 3203 3632 3212
rect 3484 3183 3493 3203
rect 3513 3183 3603 3203
rect 3623 3183 3632 3203
rect 3288 3174 3384 3176
rect 3484 3173 3632 3183
rect 3691 3203 3728 3213
rect 3691 3183 3699 3203
rect 3719 3183 3728 3203
rect 3540 3172 3576 3173
rect 2951 3165 2987 3167
rect 2951 3136 2988 3165
rect 2393 3127 2428 3128
rect 2370 3122 2428 3127
rect 2370 3102 2373 3122
rect 2393 3108 2428 3122
rect 2448 3108 2457 3128
rect 2393 3100 2457 3108
rect 2419 3099 2457 3100
rect 2420 3098 2457 3099
rect 2523 3132 2559 3133
rect 2631 3132 2667 3133
rect 2523 3124 2667 3132
rect 2523 3104 2531 3124
rect 2551 3123 2639 3124
rect 2551 3105 2586 3123
rect 2604 3105 2639 3123
rect 2551 3104 2639 3105
rect 2659 3104 2667 3124
rect 2523 3098 2667 3104
rect 2733 3128 2771 3136
rect 2849 3132 2885 3133
rect 2733 3108 2742 3128
rect 2762 3108 2771 3128
rect 2733 3099 2771 3108
rect 2800 3124 2885 3132
rect 2800 3104 2857 3124
rect 2877 3104 2885 3124
rect 2733 3098 2770 3099
rect 2800 3098 2885 3104
rect 2951 3128 2989 3136
rect 2951 3108 2960 3128
rect 2980 3108 2989 3128
rect 3691 3116 3728 3183
rect 3763 3212 3794 3263
rect 4076 3251 4094 3269
rect 4112 3251 4128 3269
rect 3813 3212 3850 3213
rect 3763 3203 3850 3212
rect 3763 3183 3821 3203
rect 3841 3183 3850 3203
rect 3763 3173 3850 3183
rect 3909 3203 3946 3213
rect 3909 3183 3917 3203
rect 3937 3183 3946 3203
rect 3763 3172 3794 3173
rect 3388 3113 3425 3114
rect 3691 3113 3730 3116
rect 3387 3112 3730 3113
rect 3909 3112 3946 3183
rect 2951 3099 2989 3108
rect 3312 3107 3730 3112
rect 2951 3098 2988 3099
rect 2412 3070 2502 3076
rect 2412 3050 2428 3070
rect 2448 3068 2502 3070
rect 2448 3050 2473 3068
rect 2412 3048 2473 3050
rect 2493 3048 2502 3068
rect 2412 3042 2502 3048
rect 2425 2988 2462 2989
rect 2521 2988 2558 2989
rect 2577 2988 2613 3098
rect 2800 3077 2831 3098
rect 3312 3087 3315 3107
rect 3335 3087 3730 3107
rect 3759 3088 3946 3112
rect 2796 3076 2831 3077
rect 2674 3066 2831 3076
rect 2674 3046 2691 3066
rect 2711 3046 2831 3066
rect 2674 3039 2831 3046
rect 2898 3069 3047 3077
rect 2898 3049 2909 3069
rect 2929 3049 2968 3069
rect 2988 3049 3047 3069
rect 2898 3042 3047 3049
rect 3691 3062 3730 3087
rect 4076 3062 4128 3251
rect 4520 3279 4530 3297
rect 4548 3279 4560 3297
rect 4692 3295 4701 3315
rect 4721 3295 4730 3315
rect 4692 3287 4730 3295
rect 4796 3319 4881 3325
rect 4911 3324 4948 3325
rect 4796 3299 4804 3319
rect 4824 3299 4881 3319
rect 4796 3291 4881 3299
rect 4910 3315 4948 3324
rect 4910 3295 4919 3315
rect 4939 3295 4948 3315
rect 4796 3290 4832 3291
rect 4910 3287 4948 3295
rect 5014 3319 5158 3325
rect 5014 3299 5022 3319
rect 5042 3299 5075 3319
rect 5095 3299 5130 3319
rect 5150 3299 5158 3319
rect 5014 3291 5158 3299
rect 5014 3290 5050 3291
rect 5122 3290 5158 3291
rect 5224 3324 5261 3325
rect 5224 3323 5262 3324
rect 5224 3315 5288 3323
rect 5224 3295 5233 3315
rect 5253 3301 5288 3315
rect 5308 3301 5311 3321
rect 5253 3296 5311 3301
rect 5253 3295 5288 3296
rect 4520 3223 4560 3279
rect 4693 3258 4730 3287
rect 4694 3256 4730 3258
rect 4694 3234 4885 3256
rect 4911 3255 4948 3287
rect 5224 3283 5288 3295
rect 5328 3257 5355 3435
rect 6213 3410 6255 3455
rect 5187 3255 5355 3257
rect 4911 3245 5355 3255
rect 5496 3351 5683 3375
rect 5714 3356 6107 3376
rect 6127 3356 6130 3376
rect 5714 3351 6130 3356
rect 5496 3280 5533 3351
rect 5714 3350 6055 3351
rect 5648 3290 5679 3291
rect 5496 3260 5505 3280
rect 5525 3260 5533 3280
rect 5496 3250 5533 3260
rect 5592 3280 5679 3290
rect 5592 3260 5601 3280
rect 5621 3260 5679 3280
rect 5592 3251 5679 3260
rect 5592 3250 5629 3251
rect 4517 3218 4560 3223
rect 4908 3229 5355 3245
rect 4908 3223 4936 3229
rect 5187 3228 5355 3229
rect 4517 3215 4667 3218
rect 4908 3215 4935 3223
rect 4517 3213 4935 3215
rect 4517 3195 4526 3213
rect 4544 3195 4935 3213
rect 5648 3200 5679 3251
rect 5714 3280 5751 3350
rect 6017 3349 6054 3350
rect 5866 3290 5902 3291
rect 5714 3260 5723 3280
rect 5743 3260 5751 3280
rect 5714 3250 5751 3260
rect 5810 3280 5958 3290
rect 6058 3287 6154 3289
rect 5810 3260 5819 3280
rect 5839 3260 5929 3280
rect 5949 3260 5958 3280
rect 5810 3251 5958 3260
rect 6016 3280 6154 3287
rect 6016 3260 6025 3280
rect 6045 3260 6154 3280
rect 6016 3251 6154 3260
rect 5810 3250 5847 3251
rect 5540 3197 5581 3198
rect 4517 3192 4935 3195
rect 4517 3186 4560 3192
rect 4520 3183 4560 3186
rect 5435 3190 5581 3197
rect 4917 3174 4957 3175
rect 4628 3157 4957 3174
rect 5435 3170 5491 3190
rect 5511 3170 5550 3190
rect 5570 3170 5581 3190
rect 5435 3162 5581 3170
rect 5648 3193 5805 3200
rect 5648 3173 5768 3193
rect 5788 3173 5805 3193
rect 5648 3163 5805 3173
rect 5648 3162 5683 3163
rect 4512 3114 4555 3125
rect 4512 3096 4524 3114
rect 4542 3096 4555 3114
rect 4512 3070 4555 3096
rect 4628 3070 4655 3157
rect 4917 3148 4957 3157
rect 3691 3044 4130 3062
rect 2898 3041 2939 3042
rect 2632 2988 2669 2989
rect 2325 2979 2463 2988
rect 2325 2959 2434 2979
rect 2454 2959 2463 2979
rect 2325 2952 2463 2959
rect 2521 2979 2669 2988
rect 2521 2959 2530 2979
rect 2550 2959 2640 2979
rect 2660 2959 2669 2979
rect 2325 2950 2421 2952
rect 2521 2949 2669 2959
rect 2728 2979 2765 2989
rect 2728 2959 2736 2979
rect 2756 2959 2765 2979
rect 2577 2948 2613 2949
rect 2425 2889 2462 2890
rect 2728 2889 2765 2959
rect 2800 2988 2831 3039
rect 3691 3026 4091 3044
rect 4109 3026 4130 3044
rect 3691 3020 4130 3026
rect 3697 3016 4130 3020
rect 4512 3049 4655 3070
rect 4699 3122 4733 3138
rect 4917 3128 5310 3148
rect 5330 3128 5333 3148
rect 5648 3141 5679 3162
rect 5866 3141 5902 3251
rect 5921 3250 5958 3251
rect 6017 3250 6054 3251
rect 5977 3191 6067 3197
rect 5977 3171 5986 3191
rect 6006 3189 6067 3191
rect 6006 3171 6031 3189
rect 5977 3169 6031 3171
rect 6051 3169 6067 3189
rect 5977 3163 6067 3169
rect 5491 3140 5528 3141
rect 4917 3123 5333 3128
rect 5490 3131 5528 3140
rect 4917 3122 5258 3123
rect 4699 3052 4736 3122
rect 4851 3062 4882 3063
rect 4512 3047 4649 3049
rect 4076 3014 4128 3016
rect 4512 3005 4555 3047
rect 4699 3032 4708 3052
rect 4728 3032 4736 3052
rect 4699 3022 4736 3032
rect 4795 3052 4882 3062
rect 4795 3032 4804 3052
rect 4824 3032 4882 3052
rect 4795 3023 4882 3032
rect 4795 3022 4832 3023
rect 4510 2995 4555 3005
rect 2850 2988 2887 2989
rect 2800 2979 2887 2988
rect 2800 2959 2858 2979
rect 2878 2959 2887 2979
rect 2800 2949 2887 2959
rect 2946 2979 2983 2989
rect 2946 2959 2954 2979
rect 2974 2959 2983 2979
rect 4510 2977 4519 2995
rect 4537 2977 4555 2995
rect 4510 2971 4555 2977
rect 4851 2972 4882 3023
rect 4917 3052 4954 3122
rect 5220 3121 5257 3122
rect 5490 3111 5499 3131
rect 5519 3111 5528 3131
rect 5490 3103 5528 3111
rect 5594 3135 5679 3141
rect 5709 3140 5746 3141
rect 5594 3115 5602 3135
rect 5622 3115 5679 3135
rect 5594 3107 5679 3115
rect 5708 3131 5746 3140
rect 5708 3111 5717 3131
rect 5737 3111 5746 3131
rect 5594 3106 5630 3107
rect 5708 3103 5746 3111
rect 5812 3135 5956 3141
rect 5812 3115 5820 3135
rect 5840 3132 5928 3135
rect 5840 3115 5875 3132
rect 5812 3114 5875 3115
rect 5894 3115 5928 3132
rect 5948 3115 5956 3135
rect 5894 3114 5956 3115
rect 5812 3107 5956 3114
rect 5812 3106 5848 3107
rect 5920 3106 5956 3107
rect 6022 3140 6059 3141
rect 6022 3139 6060 3140
rect 6082 3139 6109 3143
rect 6022 3137 6109 3139
rect 6022 3131 6086 3137
rect 6022 3111 6031 3131
rect 6051 3117 6086 3131
rect 6106 3117 6109 3137
rect 6051 3112 6109 3117
rect 6051 3111 6086 3112
rect 5491 3074 5528 3103
rect 5492 3072 5528 3074
rect 5069 3062 5105 3063
rect 4917 3032 4926 3052
rect 4946 3032 4954 3052
rect 4917 3022 4954 3032
rect 5013 3052 5161 3062
rect 5261 3059 5357 3061
rect 5013 3032 5022 3052
rect 5042 3032 5132 3052
rect 5152 3032 5161 3052
rect 5013 3023 5161 3032
rect 5219 3052 5357 3059
rect 5219 3032 5228 3052
rect 5248 3032 5357 3052
rect 5492 3050 5683 3072
rect 5709 3071 5746 3103
rect 6022 3099 6086 3111
rect 6126 3073 6153 3251
rect 5985 3071 6153 3073
rect 5709 3045 6153 3071
rect 5219 3023 5357 3032
rect 5013 3022 5050 3023
rect 4510 2968 4547 2971
rect 4743 2969 4784 2970
rect 2800 2948 2831 2949
rect 2424 2888 2765 2889
rect 2946 2888 2983 2959
rect 4635 2962 4784 2969
rect 4079 2949 4116 2954
rect 2349 2883 2765 2888
rect 2349 2863 2352 2883
rect 2372 2863 2765 2883
rect 2796 2864 2983 2888
rect 4070 2945 4117 2949
rect 4070 2927 4089 2945
rect 4107 2927 4117 2945
rect 4635 2942 4694 2962
rect 4714 2942 4753 2962
rect 4773 2942 4784 2962
rect 4635 2934 4784 2942
rect 4851 2965 5008 2972
rect 4851 2945 4971 2965
rect 4991 2945 5008 2965
rect 4851 2935 5008 2945
rect 4851 2934 4886 2935
rect 4070 2879 4117 2927
rect 4851 2913 4882 2934
rect 5069 2913 5105 3023
rect 5124 3022 5161 3023
rect 5220 3022 5257 3023
rect 5180 2963 5270 2969
rect 5180 2943 5189 2963
rect 5209 2961 5270 2963
rect 5209 2943 5234 2961
rect 5180 2941 5234 2943
rect 5254 2941 5270 2961
rect 5180 2935 5270 2941
rect 4694 2912 4731 2913
rect 3694 2876 4117 2879
rect 2569 2862 2634 2863
rect 3672 2846 4117 2876
rect 4506 2904 4544 2906
rect 4506 2896 4549 2904
rect 4506 2878 4517 2896
rect 4535 2878 4549 2896
rect 4506 2851 4549 2878
rect 4693 2903 4731 2912
rect 4693 2883 4702 2903
rect 4722 2883 4731 2903
rect 4693 2875 4731 2883
rect 4797 2907 4882 2913
rect 4912 2912 4949 2913
rect 4797 2887 4805 2907
rect 4825 2887 4882 2907
rect 4797 2879 4882 2887
rect 4911 2903 4949 2912
rect 4911 2883 4920 2903
rect 4940 2883 4949 2903
rect 4797 2878 4833 2879
rect 4911 2875 4949 2883
rect 5015 2911 5159 2913
rect 5015 2907 5067 2911
rect 5015 2887 5023 2907
rect 5043 2891 5067 2907
rect 5087 2907 5159 2911
rect 5087 2891 5131 2907
rect 5043 2887 5131 2891
rect 5151 2887 5159 2907
rect 5015 2879 5159 2887
rect 5015 2878 5051 2879
rect 5123 2878 5159 2879
rect 5225 2912 5262 2913
rect 5225 2911 5263 2912
rect 5225 2903 5289 2911
rect 5225 2883 5234 2903
rect 5254 2889 5289 2903
rect 5309 2889 5312 2909
rect 5254 2884 5312 2889
rect 5254 2883 5289 2884
rect 2765 2830 2805 2838
rect 2765 2808 2773 2830
rect 2797 2808 2805 2830
rect 2370 2579 2407 2585
rect 2370 2560 2378 2579
rect 2399 2560 2407 2579
rect 2370 2552 2407 2560
rect 2070 2431 2077 2453
rect 2101 2431 2109 2453
rect 2070 2425 2109 2431
rect 1600 2420 1640 2422
rect 1766 2421 1934 2422
rect 1868 2420 1905 2421
rect 834 2404 972 2413
rect 628 2403 665 2404
rect 358 2350 399 2351
rect 132 2329 184 2347
rect 250 2343 399 2350
rect 250 2323 309 2343
rect 329 2323 368 2343
rect 388 2323 399 2343
rect 250 2315 399 2323
rect 466 2346 623 2353
rect 466 2326 586 2346
rect 606 2326 623 2346
rect 466 2316 623 2326
rect 466 2315 501 2316
rect 466 2294 497 2315
rect 684 2294 720 2404
rect 739 2403 776 2404
rect 835 2403 872 2404
rect 795 2344 885 2350
rect 795 2324 804 2344
rect 824 2342 885 2344
rect 824 2324 849 2342
rect 795 2322 849 2324
rect 869 2322 885 2342
rect 795 2316 885 2322
rect 309 2293 346 2294
rect 308 2284 346 2293
rect 136 2266 176 2276
rect 136 2248 146 2266
rect 164 2248 176 2266
rect 308 2264 317 2284
rect 337 2264 346 2284
rect 308 2256 346 2264
rect 412 2288 497 2294
rect 527 2293 564 2294
rect 412 2268 420 2288
rect 440 2268 497 2288
rect 412 2260 497 2268
rect 526 2284 564 2293
rect 526 2264 535 2284
rect 555 2264 564 2284
rect 412 2259 448 2260
rect 526 2256 564 2264
rect 630 2288 774 2294
rect 630 2268 638 2288
rect 658 2268 691 2288
rect 711 2268 746 2288
rect 766 2268 774 2288
rect 630 2260 774 2268
rect 630 2259 666 2260
rect 738 2259 774 2260
rect 840 2293 877 2294
rect 840 2292 878 2293
rect 840 2284 904 2292
rect 840 2264 849 2284
rect 869 2270 904 2284
rect 924 2270 927 2290
rect 869 2265 927 2270
rect 869 2264 904 2265
rect 136 2192 176 2248
rect 309 2227 346 2256
rect 310 2225 346 2227
rect 310 2203 501 2225
rect 527 2224 564 2256
rect 840 2252 904 2264
rect 944 2226 971 2404
rect 803 2224 971 2226
rect 527 2214 971 2224
rect 1112 2320 1299 2344
rect 1330 2325 1723 2345
rect 1743 2325 1746 2345
rect 1330 2320 1746 2325
rect 1112 2249 1149 2320
rect 1330 2319 1671 2320
rect 1264 2259 1295 2260
rect 1112 2229 1121 2249
rect 1141 2229 1149 2249
rect 1112 2219 1149 2229
rect 1208 2249 1295 2259
rect 1208 2229 1217 2249
rect 1237 2229 1295 2249
rect 1208 2220 1295 2229
rect 1208 2219 1245 2220
rect 133 2187 176 2192
rect 524 2198 971 2214
rect 524 2192 552 2198
rect 803 2197 971 2198
rect 133 2184 283 2187
rect 524 2184 551 2192
rect 133 2182 551 2184
rect 133 2164 142 2182
rect 160 2164 551 2182
rect 1264 2169 1295 2220
rect 1330 2249 1367 2319
rect 1633 2318 1670 2319
rect 1871 2261 1904 2420
rect 1482 2259 1518 2260
rect 1330 2229 1339 2249
rect 1359 2229 1367 2249
rect 1330 2219 1367 2229
rect 1426 2249 1574 2259
rect 1674 2256 1770 2258
rect 1426 2229 1435 2249
rect 1455 2229 1545 2249
rect 1565 2229 1574 2249
rect 1426 2220 1574 2229
rect 1632 2249 1770 2256
rect 1632 2229 1641 2249
rect 1661 2229 1770 2249
rect 1871 2257 1907 2261
rect 1871 2239 1880 2257
rect 1902 2239 1907 2257
rect 1871 2233 1907 2239
rect 1632 2220 1770 2229
rect 1426 2219 1463 2220
rect 1156 2166 1197 2167
rect 133 2161 551 2164
rect 133 2155 176 2161
rect 136 2152 176 2155
rect 1048 2159 1197 2166
rect 533 2143 573 2144
rect 244 2126 573 2143
rect 1048 2139 1107 2159
rect 1127 2139 1166 2159
rect 1186 2139 1197 2159
rect 1048 2131 1197 2139
rect 1264 2162 1421 2169
rect 1264 2142 1384 2162
rect 1404 2142 1421 2162
rect 1264 2132 1421 2142
rect 1264 2131 1299 2132
rect 128 2083 171 2094
rect 128 2065 140 2083
rect 158 2065 171 2083
rect 128 2039 171 2065
rect 244 2039 271 2126
rect 533 2117 573 2126
rect 128 2018 271 2039
rect 315 2091 349 2107
rect 533 2097 926 2117
rect 946 2097 949 2117
rect 1264 2110 1295 2131
rect 1482 2110 1518 2220
rect 1537 2219 1574 2220
rect 1633 2219 1670 2220
rect 1593 2160 1683 2166
rect 1593 2140 1602 2160
rect 1622 2158 1683 2160
rect 1622 2140 1647 2158
rect 1593 2138 1647 2140
rect 1667 2138 1683 2158
rect 1593 2132 1683 2138
rect 1107 2109 1144 2110
rect 533 2092 949 2097
rect 1106 2100 1144 2109
rect 533 2091 874 2092
rect 315 2021 352 2091
rect 467 2031 498 2032
rect 128 2016 265 2018
rect 128 1974 171 2016
rect 315 2001 324 2021
rect 344 2001 352 2021
rect 315 1991 352 2001
rect 411 2021 498 2031
rect 411 2001 420 2021
rect 440 2001 498 2021
rect 411 1992 498 2001
rect 411 1991 448 1992
rect 126 1964 171 1974
rect 126 1946 135 1964
rect 153 1946 171 1964
rect 126 1940 171 1946
rect 467 1941 498 1992
rect 533 2021 570 2091
rect 836 2090 873 2091
rect 1106 2080 1115 2100
rect 1135 2080 1144 2100
rect 1106 2072 1144 2080
rect 1210 2104 1295 2110
rect 1325 2109 1362 2110
rect 1210 2084 1218 2104
rect 1238 2084 1295 2104
rect 1210 2076 1295 2084
rect 1324 2100 1362 2109
rect 1324 2080 1333 2100
rect 1353 2080 1362 2100
rect 1210 2075 1246 2076
rect 1324 2072 1362 2080
rect 1428 2104 1572 2110
rect 1428 2084 1436 2104
rect 1456 2085 1488 2104
rect 1509 2085 1544 2104
rect 1456 2084 1544 2085
rect 1564 2084 1572 2104
rect 1428 2076 1572 2084
rect 1428 2075 1464 2076
rect 1536 2075 1572 2076
rect 1638 2109 1675 2110
rect 1638 2108 1676 2109
rect 1638 2100 1702 2108
rect 1638 2080 1647 2100
rect 1667 2086 1702 2100
rect 1722 2086 1725 2106
rect 1667 2081 1725 2086
rect 1667 2080 1702 2081
rect 1107 2043 1144 2072
rect 1108 2041 1144 2043
rect 685 2031 721 2032
rect 533 2001 542 2021
rect 562 2001 570 2021
rect 533 1991 570 2001
rect 629 2021 777 2031
rect 877 2028 973 2030
rect 629 2001 638 2021
rect 658 2001 748 2021
rect 768 2001 777 2021
rect 629 1992 777 2001
rect 835 2021 973 2028
rect 835 2001 844 2021
rect 864 2001 973 2021
rect 1108 2019 1299 2041
rect 1325 2040 1362 2072
rect 1638 2068 1702 2080
rect 1742 2042 1769 2220
rect 2374 2219 2407 2552
rect 2471 2584 2639 2585
rect 2765 2584 2805 2808
rect 3268 2812 3436 2813
rect 3672 2812 3713 2846
rect 4070 2825 4117 2846
rect 3268 2802 3713 2812
rect 3785 2810 3928 2811
rect 3268 2786 3712 2802
rect 3268 2784 3436 2786
rect 3632 2785 3712 2786
rect 3785 2785 3930 2810
rect 4072 2785 4117 2825
rect 3268 2606 3295 2784
rect 3335 2746 3399 2758
rect 3675 2754 3712 2785
rect 3893 2754 3930 2785
rect 4075 2778 4117 2785
rect 4507 2844 4549 2851
rect 4694 2844 4731 2875
rect 4912 2844 4949 2875
rect 5225 2871 5289 2883
rect 5329 2845 5356 3023
rect 4507 2804 4552 2844
rect 4694 2819 4839 2844
rect 4912 2843 4992 2844
rect 5188 2843 5356 2845
rect 4912 2827 5356 2843
rect 4696 2818 4839 2819
rect 4911 2817 5356 2827
rect 4507 2783 4554 2804
rect 4911 2783 4952 2817
rect 5188 2816 5356 2817
rect 5819 2821 5859 3045
rect 5985 3044 6153 3045
rect 6217 3077 6250 3410
rect 6217 3069 6254 3077
rect 6217 3050 6225 3069
rect 6246 3050 6254 3069
rect 6217 3044 6254 3050
rect 5819 2799 5827 2821
rect 5851 2799 5859 2821
rect 5819 2791 5859 2799
rect 3335 2745 3370 2746
rect 3312 2740 3370 2745
rect 3312 2720 3315 2740
rect 3335 2726 3370 2740
rect 3390 2726 3399 2746
rect 3335 2718 3399 2726
rect 3361 2717 3399 2718
rect 3362 2716 3399 2717
rect 3465 2750 3501 2751
rect 3573 2750 3609 2751
rect 3465 2742 3609 2750
rect 3465 2722 3473 2742
rect 3493 2738 3581 2742
rect 3493 2722 3537 2738
rect 3465 2718 3537 2722
rect 3557 2722 3581 2738
rect 3601 2722 3609 2742
rect 3557 2718 3609 2722
rect 3465 2716 3609 2718
rect 3675 2746 3713 2754
rect 3791 2750 3827 2751
rect 3675 2726 3684 2746
rect 3704 2726 3713 2746
rect 3675 2717 3713 2726
rect 3742 2742 3827 2750
rect 3742 2722 3799 2742
rect 3819 2722 3827 2742
rect 3675 2716 3712 2717
rect 3742 2716 3827 2722
rect 3893 2746 3931 2754
rect 3893 2726 3902 2746
rect 3922 2726 3931 2746
rect 3893 2717 3931 2726
rect 4075 2751 4118 2778
rect 4075 2733 4089 2751
rect 4107 2733 4118 2751
rect 4075 2725 4118 2733
rect 4080 2723 4118 2725
rect 4507 2753 4952 2783
rect 5990 2766 6055 2767
rect 4507 2750 4930 2753
rect 3893 2716 3930 2717
rect 3354 2688 3444 2694
rect 3354 2668 3370 2688
rect 3390 2686 3444 2688
rect 3390 2668 3415 2686
rect 3354 2666 3415 2668
rect 3435 2666 3444 2686
rect 3354 2660 3444 2666
rect 3367 2606 3404 2607
rect 3463 2606 3500 2607
rect 3519 2606 3555 2716
rect 3742 2695 3773 2716
rect 4507 2702 4554 2750
rect 3738 2694 3773 2695
rect 3616 2684 3773 2694
rect 3616 2664 3633 2684
rect 3653 2664 3773 2684
rect 3616 2657 3773 2664
rect 3840 2687 3989 2695
rect 3840 2667 3851 2687
rect 3871 2667 3910 2687
rect 3930 2667 3989 2687
rect 4507 2684 4517 2702
rect 4535 2684 4554 2702
rect 4507 2680 4554 2684
rect 5641 2741 5828 2765
rect 5859 2746 6252 2766
rect 6272 2746 6275 2766
rect 5859 2741 6275 2746
rect 4508 2675 4545 2680
rect 3840 2660 3989 2667
rect 5641 2670 5678 2741
rect 5859 2740 6200 2741
rect 5793 2680 5824 2681
rect 3840 2659 3881 2660
rect 4077 2658 4114 2661
rect 3574 2606 3611 2607
rect 3267 2597 3405 2606
rect 2471 2558 2915 2584
rect 2471 2556 2639 2558
rect 2471 2378 2498 2556
rect 2538 2518 2602 2530
rect 2878 2526 2915 2558
rect 2941 2557 3132 2579
rect 3267 2577 3376 2597
rect 3396 2577 3405 2597
rect 3267 2570 3405 2577
rect 3463 2597 3611 2606
rect 3463 2577 3472 2597
rect 3492 2577 3582 2597
rect 3602 2577 3611 2597
rect 3267 2568 3363 2570
rect 3463 2567 3611 2577
rect 3670 2597 3707 2607
rect 3670 2577 3678 2597
rect 3698 2577 3707 2597
rect 3519 2566 3555 2567
rect 3096 2555 3132 2557
rect 3096 2526 3133 2555
rect 2538 2517 2573 2518
rect 2515 2512 2573 2517
rect 2515 2492 2518 2512
rect 2538 2498 2573 2512
rect 2593 2498 2602 2518
rect 2538 2492 2602 2498
rect 2515 2490 2602 2492
rect 2515 2486 2542 2490
rect 2564 2489 2602 2490
rect 2565 2488 2602 2489
rect 2668 2522 2704 2523
rect 2776 2522 2812 2523
rect 2668 2515 2812 2522
rect 2668 2514 2730 2515
rect 2668 2494 2676 2514
rect 2696 2497 2730 2514
rect 2749 2514 2812 2515
rect 2749 2497 2784 2514
rect 2696 2494 2784 2497
rect 2804 2494 2812 2514
rect 2668 2488 2812 2494
rect 2878 2518 2916 2526
rect 2994 2522 3030 2523
rect 2878 2498 2887 2518
rect 2907 2498 2916 2518
rect 2878 2489 2916 2498
rect 2945 2514 3030 2522
rect 2945 2494 3002 2514
rect 3022 2494 3030 2514
rect 2878 2488 2915 2489
rect 2945 2488 3030 2494
rect 3096 2518 3134 2526
rect 3096 2498 3105 2518
rect 3125 2498 3134 2518
rect 3367 2507 3404 2508
rect 3670 2507 3707 2577
rect 3742 2606 3773 2657
rect 4069 2652 4114 2658
rect 4069 2634 4087 2652
rect 4105 2634 4114 2652
rect 5641 2650 5650 2670
rect 5670 2650 5678 2670
rect 5641 2640 5678 2650
rect 5737 2670 5824 2680
rect 5737 2650 5746 2670
rect 5766 2650 5824 2670
rect 5737 2641 5824 2650
rect 5737 2640 5774 2641
rect 4069 2624 4114 2634
rect 3792 2606 3829 2607
rect 3742 2597 3829 2606
rect 3742 2577 3800 2597
rect 3820 2577 3829 2597
rect 3742 2567 3829 2577
rect 3888 2597 3925 2607
rect 3888 2577 3896 2597
rect 3916 2577 3925 2597
rect 4069 2582 4112 2624
rect 4496 2613 4548 2615
rect 3975 2580 4112 2582
rect 3742 2566 3773 2567
rect 3888 2507 3925 2577
rect 3366 2506 3707 2507
rect 3096 2489 3134 2498
rect 3291 2501 3707 2506
rect 3096 2488 3133 2489
rect 2557 2460 2647 2466
rect 2557 2440 2573 2460
rect 2593 2458 2647 2460
rect 2593 2440 2618 2458
rect 2557 2438 2618 2440
rect 2638 2438 2647 2458
rect 2557 2432 2647 2438
rect 2570 2378 2607 2379
rect 2666 2378 2703 2379
rect 2722 2378 2758 2488
rect 2945 2467 2976 2488
rect 3291 2481 3294 2501
rect 3314 2481 3707 2501
rect 3891 2491 3925 2507
rect 3969 2559 4112 2580
rect 4494 2609 4927 2613
rect 4494 2603 4933 2609
rect 4494 2585 4515 2603
rect 4533 2585 4933 2603
rect 5793 2590 5824 2641
rect 5859 2670 5896 2740
rect 6162 2739 6199 2740
rect 6011 2680 6047 2681
rect 5859 2650 5868 2670
rect 5888 2650 5896 2670
rect 5859 2640 5896 2650
rect 5955 2670 6103 2680
rect 6203 2677 6299 2679
rect 5955 2650 5964 2670
rect 5984 2650 6074 2670
rect 6094 2650 6103 2670
rect 5955 2641 6103 2650
rect 6161 2670 6299 2677
rect 6161 2650 6170 2670
rect 6190 2650 6299 2670
rect 6161 2641 6299 2650
rect 5955 2640 5992 2641
rect 5685 2587 5726 2588
rect 4494 2567 4933 2585
rect 3667 2472 3707 2481
rect 3969 2472 3996 2559
rect 4069 2533 4112 2559
rect 4069 2515 4082 2533
rect 4100 2515 4112 2533
rect 4069 2504 4112 2515
rect 2941 2466 2976 2467
rect 2819 2456 2976 2466
rect 2819 2436 2836 2456
rect 2856 2436 2976 2456
rect 2819 2429 2976 2436
rect 3043 2459 3189 2467
rect 3043 2439 3054 2459
rect 3074 2439 3113 2459
rect 3133 2439 3189 2459
rect 3667 2455 3996 2472
rect 3667 2454 3707 2455
rect 3043 2432 3189 2439
rect 4064 2443 4104 2446
rect 4064 2437 4107 2443
rect 3689 2434 4107 2437
rect 3043 2431 3084 2432
rect 2777 2378 2814 2379
rect 2470 2369 2608 2378
rect 2470 2349 2579 2369
rect 2599 2349 2608 2369
rect 2470 2342 2608 2349
rect 2666 2369 2814 2378
rect 2666 2349 2675 2369
rect 2695 2349 2785 2369
rect 2805 2349 2814 2369
rect 2470 2340 2566 2342
rect 2666 2339 2814 2349
rect 2873 2369 2910 2379
rect 2873 2349 2881 2369
rect 2901 2349 2910 2369
rect 2722 2338 2758 2339
rect 2570 2279 2607 2280
rect 2873 2279 2910 2349
rect 2945 2378 2976 2429
rect 3689 2416 4080 2434
rect 4098 2416 4107 2434
rect 3689 2414 4107 2416
rect 3689 2406 3716 2414
rect 3957 2411 4107 2414
rect 3269 2400 3437 2401
rect 3688 2400 3716 2406
rect 3269 2384 3716 2400
rect 4064 2406 4107 2411
rect 2995 2378 3032 2379
rect 2945 2369 3032 2378
rect 2945 2349 3003 2369
rect 3023 2349 3032 2369
rect 2945 2339 3032 2349
rect 3091 2369 3128 2379
rect 3091 2349 3099 2369
rect 3119 2349 3128 2369
rect 2945 2338 2976 2339
rect 2569 2278 2910 2279
rect 3091 2278 3128 2349
rect 2494 2273 2910 2278
rect 2494 2253 2497 2273
rect 2517 2253 2910 2273
rect 2941 2254 3128 2278
rect 3269 2374 3713 2384
rect 3269 2372 3437 2374
rect 2369 2174 2411 2219
rect 3269 2194 3296 2372
rect 3336 2334 3400 2346
rect 3676 2342 3713 2374
rect 3739 2373 3930 2395
rect 3894 2371 3930 2373
rect 3894 2342 3931 2371
rect 4064 2350 4104 2406
rect 3336 2333 3371 2334
rect 3313 2328 3371 2333
rect 3313 2308 3316 2328
rect 3336 2314 3371 2328
rect 3391 2314 3400 2334
rect 3336 2306 3400 2314
rect 3362 2305 3400 2306
rect 3363 2304 3400 2305
rect 3466 2338 3502 2339
rect 3574 2338 3610 2339
rect 3466 2330 3610 2338
rect 3466 2310 3474 2330
rect 3494 2310 3529 2330
rect 3549 2310 3582 2330
rect 3602 2310 3610 2330
rect 3466 2304 3610 2310
rect 3676 2334 3714 2342
rect 3792 2338 3828 2339
rect 3676 2314 3685 2334
rect 3705 2314 3714 2334
rect 3676 2305 3714 2314
rect 3743 2330 3828 2338
rect 3743 2310 3800 2330
rect 3820 2310 3828 2330
rect 3676 2304 3713 2305
rect 3743 2304 3828 2310
rect 3894 2334 3932 2342
rect 3894 2314 3903 2334
rect 3923 2314 3932 2334
rect 4064 2332 4076 2350
rect 4094 2332 4104 2350
rect 4496 2378 4548 2567
rect 4894 2542 4933 2567
rect 5577 2580 5726 2587
rect 5577 2560 5636 2580
rect 5656 2560 5695 2580
rect 5715 2560 5726 2580
rect 5577 2552 5726 2560
rect 5793 2583 5950 2590
rect 5793 2563 5913 2583
rect 5933 2563 5950 2583
rect 5793 2553 5950 2563
rect 5793 2552 5828 2553
rect 4678 2517 4865 2541
rect 4894 2522 5289 2542
rect 5309 2522 5312 2542
rect 5793 2531 5824 2552
rect 6011 2531 6047 2641
rect 6066 2640 6103 2641
rect 6162 2640 6199 2641
rect 6122 2581 6212 2587
rect 6122 2561 6131 2581
rect 6151 2579 6212 2581
rect 6151 2561 6176 2579
rect 6122 2559 6176 2561
rect 6196 2559 6212 2579
rect 6122 2553 6212 2559
rect 5636 2530 5673 2531
rect 4894 2517 5312 2522
rect 5635 2521 5673 2530
rect 4678 2446 4715 2517
rect 4894 2516 5237 2517
rect 4894 2513 4933 2516
rect 5199 2515 5236 2516
rect 4830 2456 4861 2457
rect 4678 2426 4687 2446
rect 4707 2426 4715 2446
rect 4678 2416 4715 2426
rect 4774 2446 4861 2456
rect 4774 2426 4783 2446
rect 4803 2426 4861 2446
rect 4774 2417 4861 2426
rect 4774 2416 4811 2417
rect 4496 2360 4512 2378
rect 4530 2360 4548 2378
rect 4830 2366 4861 2417
rect 4896 2446 4933 2513
rect 5635 2501 5644 2521
rect 5664 2501 5673 2521
rect 5635 2493 5673 2501
rect 5739 2525 5824 2531
rect 5854 2530 5891 2531
rect 5739 2505 5747 2525
rect 5767 2505 5824 2525
rect 5739 2497 5824 2505
rect 5853 2521 5891 2530
rect 5853 2501 5862 2521
rect 5882 2501 5891 2521
rect 5739 2496 5775 2497
rect 5853 2493 5891 2501
rect 5957 2529 6101 2531
rect 5957 2525 6017 2529
rect 5957 2505 5965 2525
rect 5985 2507 6017 2525
rect 6040 2525 6101 2529
rect 6040 2507 6073 2525
rect 5985 2505 6073 2507
rect 6093 2505 6101 2525
rect 5957 2497 6101 2505
rect 5957 2496 5993 2497
rect 6065 2496 6101 2497
rect 6167 2530 6204 2531
rect 6167 2529 6205 2530
rect 6167 2521 6231 2529
rect 6167 2501 6176 2521
rect 6196 2507 6231 2521
rect 6251 2507 6254 2527
rect 6196 2502 6254 2507
rect 6196 2501 6231 2502
rect 5636 2464 5673 2493
rect 5637 2462 5673 2464
rect 5048 2456 5084 2457
rect 4896 2426 4905 2446
rect 4925 2426 4933 2446
rect 4896 2416 4933 2426
rect 4992 2446 5140 2456
rect 5240 2453 5336 2455
rect 4992 2426 5001 2446
rect 5021 2426 5111 2446
rect 5131 2426 5140 2446
rect 4992 2417 5140 2426
rect 5198 2446 5336 2453
rect 5198 2426 5207 2446
rect 5227 2426 5336 2446
rect 5637 2440 5828 2462
rect 5854 2461 5891 2493
rect 6167 2489 6231 2501
rect 5854 2460 6129 2461
rect 6271 2460 6298 2641
rect 5854 2435 6298 2460
rect 6434 2466 6473 4281
rect 6775 4268 6808 4601
rect 6872 4633 7040 4634
rect 7166 4633 7206 4857
rect 7669 4861 7837 4862
rect 8078 4861 8113 4878
rect 8470 4868 8517 4879
rect 7669 4835 8113 4861
rect 7669 4833 7837 4835
rect 8033 4834 8113 4835
rect 8268 4834 8335 4860
rect 8474 4834 8517 4868
rect 7669 4655 7696 4833
rect 7736 4795 7800 4807
rect 8076 4803 8113 4834
rect 8294 4803 8331 4834
rect 8476 4809 8517 4834
rect 8921 4892 8962 4917
rect 9107 4892 9144 4923
rect 9325 4892 9362 4923
rect 9638 4919 9702 4931
rect 9742 4893 9769 5071
rect 8921 4858 8964 4892
rect 9103 4866 9170 4892
rect 9325 4891 9405 4892
rect 9601 4891 9769 4893
rect 9325 4865 9769 4891
rect 8921 4847 8968 4858
rect 9325 4848 9360 4865
rect 9601 4864 9769 4865
rect 10232 4869 10272 5093
rect 10398 5092 10566 5093
rect 10630 5125 10663 5458
rect 10965 5445 11004 7260
rect 11140 7266 11584 7291
rect 11140 7085 11167 7266
rect 11309 7265 11584 7266
rect 11207 7225 11271 7237
rect 11547 7233 11584 7265
rect 11610 7264 11801 7286
rect 12102 7280 12211 7300
rect 12231 7280 12240 7300
rect 12102 7273 12240 7280
rect 12298 7300 12446 7309
rect 12298 7280 12307 7300
rect 12327 7280 12417 7300
rect 12437 7280 12446 7300
rect 12102 7271 12198 7273
rect 12298 7270 12446 7280
rect 12505 7300 12542 7310
rect 12505 7280 12513 7300
rect 12533 7280 12542 7300
rect 12354 7269 12390 7270
rect 11765 7262 11801 7264
rect 11765 7233 11802 7262
rect 11207 7224 11242 7225
rect 11184 7219 11242 7224
rect 11184 7199 11187 7219
rect 11207 7205 11242 7219
rect 11262 7205 11271 7225
rect 11207 7197 11271 7205
rect 11233 7196 11271 7197
rect 11234 7195 11271 7196
rect 11337 7229 11373 7230
rect 11445 7229 11481 7230
rect 11337 7221 11481 7229
rect 11337 7201 11345 7221
rect 11365 7219 11453 7221
rect 11365 7201 11398 7219
rect 11337 7197 11398 7201
rect 11421 7201 11453 7219
rect 11473 7201 11481 7221
rect 11421 7197 11481 7201
rect 11337 7195 11481 7197
rect 11547 7225 11585 7233
rect 11663 7229 11699 7230
rect 11547 7205 11556 7225
rect 11576 7205 11585 7225
rect 11547 7196 11585 7205
rect 11614 7221 11699 7229
rect 11614 7201 11671 7221
rect 11691 7201 11699 7221
rect 11547 7195 11584 7196
rect 11614 7195 11699 7201
rect 11765 7225 11803 7233
rect 11765 7205 11774 7225
rect 11794 7205 11803 7225
rect 12505 7213 12542 7280
rect 12577 7309 12608 7360
rect 12890 7348 12908 7366
rect 12926 7348 12942 7366
rect 12627 7309 12664 7310
rect 12577 7300 12664 7309
rect 12577 7280 12635 7300
rect 12655 7280 12664 7300
rect 12577 7270 12664 7280
rect 12723 7300 12760 7310
rect 12723 7280 12731 7300
rect 12751 7280 12760 7300
rect 12577 7269 12608 7270
rect 12202 7210 12239 7211
rect 12505 7210 12544 7213
rect 12201 7209 12544 7210
rect 12723 7209 12760 7280
rect 11765 7196 11803 7205
rect 12126 7204 12544 7209
rect 11765 7195 11802 7196
rect 11226 7167 11316 7173
rect 11226 7147 11242 7167
rect 11262 7165 11316 7167
rect 11262 7147 11287 7165
rect 11226 7145 11287 7147
rect 11307 7145 11316 7165
rect 11226 7139 11316 7145
rect 11239 7085 11276 7086
rect 11335 7085 11372 7086
rect 11391 7085 11427 7195
rect 11614 7174 11645 7195
rect 12126 7184 12129 7204
rect 12149 7184 12544 7204
rect 12573 7185 12760 7209
rect 11610 7173 11645 7174
rect 11488 7163 11645 7173
rect 11488 7143 11505 7163
rect 11525 7143 11645 7163
rect 11488 7136 11645 7143
rect 11712 7166 11861 7174
rect 11712 7146 11723 7166
rect 11743 7146 11782 7166
rect 11802 7146 11861 7166
rect 11712 7139 11861 7146
rect 12505 7159 12544 7184
rect 12890 7159 12942 7348
rect 13334 7376 13344 7394
rect 13362 7376 13374 7394
rect 13506 7392 13515 7412
rect 13535 7392 13544 7412
rect 13506 7384 13544 7392
rect 13610 7416 13695 7422
rect 13725 7421 13762 7422
rect 13610 7396 13618 7416
rect 13638 7396 13695 7416
rect 13610 7388 13695 7396
rect 13724 7412 13762 7421
rect 13724 7392 13733 7412
rect 13753 7392 13762 7412
rect 13610 7387 13646 7388
rect 13724 7384 13762 7392
rect 13828 7416 13972 7422
rect 13828 7396 13836 7416
rect 13856 7396 13889 7416
rect 13909 7396 13944 7416
rect 13964 7396 13972 7416
rect 13828 7388 13972 7396
rect 13828 7387 13864 7388
rect 13936 7387 13972 7388
rect 14038 7421 14075 7422
rect 14038 7420 14076 7421
rect 14038 7412 14102 7420
rect 14038 7392 14047 7412
rect 14067 7398 14102 7412
rect 14122 7398 14125 7418
rect 14067 7393 14125 7398
rect 14067 7392 14102 7393
rect 13334 7320 13374 7376
rect 13507 7355 13544 7384
rect 13508 7353 13544 7355
rect 13508 7331 13699 7353
rect 13725 7352 13762 7384
rect 14038 7380 14102 7392
rect 14142 7354 14169 7532
rect 15027 7507 15069 7552
rect 14001 7352 14169 7354
rect 13725 7342 14169 7352
rect 14310 7448 14497 7472
rect 14528 7453 14921 7473
rect 14941 7453 14944 7473
rect 14528 7448 14944 7453
rect 14310 7377 14347 7448
rect 14528 7447 14869 7448
rect 14462 7387 14493 7388
rect 14310 7357 14319 7377
rect 14339 7357 14347 7377
rect 14310 7347 14347 7357
rect 14406 7377 14493 7387
rect 14406 7357 14415 7377
rect 14435 7357 14493 7377
rect 14406 7348 14493 7357
rect 14406 7347 14443 7348
rect 13331 7315 13374 7320
rect 13722 7326 14169 7342
rect 13722 7320 13750 7326
rect 14001 7325 14169 7326
rect 13331 7312 13481 7315
rect 13722 7312 13749 7320
rect 13331 7310 13749 7312
rect 13331 7292 13340 7310
rect 13358 7292 13749 7310
rect 14462 7297 14493 7348
rect 14528 7377 14565 7447
rect 14831 7446 14868 7447
rect 14680 7387 14716 7388
rect 14528 7357 14537 7377
rect 14557 7357 14565 7377
rect 14528 7347 14565 7357
rect 14624 7377 14772 7387
rect 14872 7384 14968 7386
rect 14624 7357 14633 7377
rect 14653 7357 14743 7377
rect 14763 7357 14772 7377
rect 14624 7348 14772 7357
rect 14830 7377 14968 7384
rect 14830 7357 14839 7377
rect 14859 7357 14968 7377
rect 14830 7348 14968 7357
rect 14624 7347 14661 7348
rect 14354 7294 14395 7295
rect 13331 7289 13749 7292
rect 13331 7283 13374 7289
rect 13334 7280 13374 7283
rect 14249 7287 14395 7294
rect 13731 7271 13771 7272
rect 13442 7254 13771 7271
rect 14249 7267 14305 7287
rect 14325 7267 14364 7287
rect 14384 7267 14395 7287
rect 14249 7259 14395 7267
rect 14462 7290 14619 7297
rect 14462 7270 14582 7290
rect 14602 7270 14619 7290
rect 14462 7260 14619 7270
rect 14462 7259 14497 7260
rect 13326 7211 13369 7222
rect 13326 7193 13338 7211
rect 13356 7193 13369 7211
rect 13326 7167 13369 7193
rect 13442 7167 13469 7254
rect 13731 7245 13771 7254
rect 12505 7141 12944 7159
rect 11712 7138 11753 7139
rect 11446 7085 11483 7086
rect 11139 7076 11277 7085
rect 11139 7056 11248 7076
rect 11268 7056 11277 7076
rect 11139 7049 11277 7056
rect 11335 7076 11483 7085
rect 11335 7056 11344 7076
rect 11364 7056 11454 7076
rect 11474 7056 11483 7076
rect 11139 7047 11235 7049
rect 11335 7046 11483 7056
rect 11542 7076 11579 7086
rect 11542 7056 11550 7076
rect 11570 7056 11579 7076
rect 11391 7045 11427 7046
rect 11239 6986 11276 6987
rect 11542 6986 11579 7056
rect 11614 7085 11645 7136
rect 12505 7123 12905 7141
rect 12923 7123 12944 7141
rect 12505 7117 12944 7123
rect 12511 7113 12944 7117
rect 13326 7146 13469 7167
rect 13513 7219 13547 7235
rect 13731 7225 14124 7245
rect 14144 7225 14147 7245
rect 14462 7238 14493 7259
rect 14680 7238 14716 7348
rect 14735 7347 14772 7348
rect 14831 7347 14868 7348
rect 14791 7288 14881 7294
rect 14791 7268 14800 7288
rect 14820 7286 14881 7288
rect 14820 7268 14845 7286
rect 14791 7266 14845 7268
rect 14865 7266 14881 7286
rect 14791 7260 14881 7266
rect 14305 7237 14342 7238
rect 13731 7220 14147 7225
rect 14304 7228 14342 7237
rect 13731 7219 14072 7220
rect 13513 7149 13550 7219
rect 13665 7159 13696 7160
rect 13326 7144 13463 7146
rect 12890 7111 12942 7113
rect 13326 7102 13369 7144
rect 13513 7129 13522 7149
rect 13542 7129 13550 7149
rect 13513 7119 13550 7129
rect 13609 7149 13696 7159
rect 13609 7129 13618 7149
rect 13638 7129 13696 7149
rect 13609 7120 13696 7129
rect 13609 7119 13646 7120
rect 13324 7092 13369 7102
rect 11664 7085 11701 7086
rect 11614 7076 11701 7085
rect 11614 7056 11672 7076
rect 11692 7056 11701 7076
rect 11614 7046 11701 7056
rect 11760 7076 11797 7086
rect 11760 7056 11768 7076
rect 11788 7056 11797 7076
rect 13324 7074 13333 7092
rect 13351 7074 13369 7092
rect 13324 7068 13369 7074
rect 13665 7069 13696 7120
rect 13731 7149 13768 7219
rect 14034 7218 14071 7219
rect 14304 7208 14313 7228
rect 14333 7208 14342 7228
rect 14304 7200 14342 7208
rect 14408 7232 14493 7238
rect 14523 7237 14560 7238
rect 14408 7212 14416 7232
rect 14436 7212 14493 7232
rect 14408 7204 14493 7212
rect 14522 7228 14560 7237
rect 14522 7208 14531 7228
rect 14551 7208 14560 7228
rect 14408 7203 14444 7204
rect 14522 7200 14560 7208
rect 14626 7232 14770 7238
rect 14626 7212 14634 7232
rect 14654 7229 14742 7232
rect 14654 7212 14689 7229
rect 14626 7211 14689 7212
rect 14708 7212 14742 7229
rect 14762 7212 14770 7232
rect 14708 7211 14770 7212
rect 14626 7204 14770 7211
rect 14626 7203 14662 7204
rect 14734 7203 14770 7204
rect 14836 7237 14873 7238
rect 14836 7236 14874 7237
rect 14896 7236 14923 7240
rect 14836 7234 14923 7236
rect 14836 7228 14900 7234
rect 14836 7208 14845 7228
rect 14865 7214 14900 7228
rect 14920 7214 14923 7234
rect 14865 7209 14923 7214
rect 14865 7208 14900 7209
rect 14305 7171 14342 7200
rect 14306 7169 14342 7171
rect 13883 7159 13919 7160
rect 13731 7129 13740 7149
rect 13760 7129 13768 7149
rect 13731 7119 13768 7129
rect 13827 7149 13975 7159
rect 14075 7156 14171 7158
rect 13827 7129 13836 7149
rect 13856 7129 13946 7149
rect 13966 7129 13975 7149
rect 13827 7120 13975 7129
rect 14033 7149 14171 7156
rect 14033 7129 14042 7149
rect 14062 7129 14171 7149
rect 14306 7147 14497 7169
rect 14523 7168 14560 7200
rect 14836 7196 14900 7208
rect 14940 7170 14967 7348
rect 14799 7168 14967 7170
rect 14523 7142 14967 7168
rect 14033 7120 14171 7129
rect 13827 7119 13864 7120
rect 13324 7065 13361 7068
rect 13557 7066 13598 7067
rect 11614 7045 11645 7046
rect 11238 6985 11579 6986
rect 11760 6985 11797 7056
rect 13449 7059 13598 7066
rect 12893 7046 12930 7051
rect 11163 6980 11579 6985
rect 11163 6960 11166 6980
rect 11186 6960 11579 6980
rect 11610 6961 11797 6985
rect 12884 7042 12931 7046
rect 12884 7024 12903 7042
rect 12921 7024 12931 7042
rect 13449 7039 13508 7059
rect 13528 7039 13567 7059
rect 13587 7039 13598 7059
rect 13449 7031 13598 7039
rect 13665 7062 13822 7069
rect 13665 7042 13785 7062
rect 13805 7042 13822 7062
rect 13665 7032 13822 7042
rect 13665 7031 13700 7032
rect 12884 6976 12931 7024
rect 13665 7010 13696 7031
rect 13883 7010 13919 7120
rect 13938 7119 13975 7120
rect 14034 7119 14071 7120
rect 13994 7060 14084 7066
rect 13994 7040 14003 7060
rect 14023 7058 14084 7060
rect 14023 7040 14048 7058
rect 13994 7038 14048 7040
rect 14068 7038 14084 7058
rect 13994 7032 14084 7038
rect 13508 7009 13545 7010
rect 12508 6973 12931 6976
rect 11383 6959 11448 6960
rect 12486 6943 12931 6973
rect 13320 7001 13358 7003
rect 13320 6993 13363 7001
rect 13320 6975 13331 6993
rect 13349 6975 13363 6993
rect 13320 6948 13363 6975
rect 13507 7000 13545 7009
rect 13507 6980 13516 7000
rect 13536 6980 13545 7000
rect 13507 6972 13545 6980
rect 13611 7004 13696 7010
rect 13726 7009 13763 7010
rect 13611 6984 13619 7004
rect 13639 6984 13696 7004
rect 13611 6976 13696 6984
rect 13725 7000 13763 7009
rect 13725 6980 13734 7000
rect 13754 6980 13763 7000
rect 13611 6975 13647 6976
rect 13725 6972 13763 6980
rect 13829 7008 13973 7010
rect 13829 7004 13881 7008
rect 13829 6984 13837 7004
rect 13857 6988 13881 7004
rect 13901 7004 13973 7008
rect 13901 6988 13945 7004
rect 13857 6984 13945 6988
rect 13965 6984 13973 7004
rect 13829 6976 13973 6984
rect 13829 6975 13865 6976
rect 13937 6975 13973 6976
rect 14039 7009 14076 7010
rect 14039 7008 14077 7009
rect 14039 7000 14103 7008
rect 14039 6980 14048 7000
rect 14068 6986 14103 7000
rect 14123 6986 14126 7006
rect 14068 6981 14126 6986
rect 14068 6980 14103 6981
rect 11579 6927 11619 6935
rect 11579 6905 11587 6927
rect 11611 6905 11619 6927
rect 11184 6676 11221 6682
rect 11184 6657 11192 6676
rect 11213 6657 11221 6676
rect 11184 6649 11221 6657
rect 11188 6316 11221 6649
rect 11285 6681 11453 6682
rect 11579 6681 11619 6905
rect 12082 6909 12250 6910
rect 12486 6909 12527 6943
rect 12884 6922 12931 6943
rect 12082 6899 12527 6909
rect 12599 6907 12742 6908
rect 12082 6883 12526 6899
rect 12082 6881 12250 6883
rect 12446 6882 12526 6883
rect 12599 6882 12744 6907
rect 12886 6882 12931 6922
rect 12082 6703 12109 6881
rect 12149 6843 12213 6855
rect 12489 6851 12526 6882
rect 12707 6851 12744 6882
rect 12889 6875 12931 6882
rect 13321 6941 13363 6948
rect 13508 6941 13545 6972
rect 13726 6941 13763 6972
rect 14039 6968 14103 6980
rect 14143 6942 14170 7120
rect 13321 6901 13366 6941
rect 13508 6916 13653 6941
rect 13726 6940 13806 6941
rect 14002 6940 14170 6942
rect 13726 6924 14170 6940
rect 13510 6915 13653 6916
rect 13725 6914 14170 6924
rect 13321 6880 13368 6901
rect 13725 6880 13766 6914
rect 14002 6913 14170 6914
rect 14633 6918 14673 7142
rect 14799 7141 14967 7142
rect 15031 7174 15064 7507
rect 15669 7506 15696 7684
rect 15736 7646 15800 7658
rect 16076 7654 16113 7686
rect 16139 7685 16330 7707
rect 16465 7705 16574 7725
rect 16594 7705 16603 7725
rect 16465 7698 16603 7705
rect 16661 7725 16809 7734
rect 16661 7705 16670 7725
rect 16690 7705 16780 7725
rect 16800 7705 16809 7725
rect 16465 7696 16561 7698
rect 16661 7695 16809 7705
rect 16868 7725 16905 7735
rect 16868 7705 16876 7725
rect 16896 7705 16905 7725
rect 16717 7694 16753 7695
rect 16294 7683 16330 7685
rect 16294 7654 16331 7683
rect 15736 7645 15771 7646
rect 15713 7640 15771 7645
rect 15713 7620 15716 7640
rect 15736 7626 15771 7640
rect 15791 7626 15800 7646
rect 15736 7618 15800 7626
rect 15762 7617 15800 7618
rect 15763 7616 15800 7617
rect 15866 7650 15902 7651
rect 15974 7650 16010 7651
rect 15866 7642 16010 7650
rect 15866 7622 15874 7642
rect 15894 7641 15982 7642
rect 15894 7622 15929 7641
rect 15950 7622 15982 7641
rect 16002 7622 16010 7642
rect 15866 7616 16010 7622
rect 16076 7646 16114 7654
rect 16192 7650 16228 7651
rect 16076 7626 16085 7646
rect 16105 7626 16114 7646
rect 16076 7617 16114 7626
rect 16143 7642 16228 7650
rect 16143 7622 16200 7642
rect 16220 7622 16228 7642
rect 16076 7616 16113 7617
rect 16143 7616 16228 7622
rect 16294 7646 16332 7654
rect 16294 7626 16303 7646
rect 16323 7626 16332 7646
rect 16565 7635 16602 7636
rect 16868 7635 16905 7705
rect 16940 7734 16971 7785
rect 17267 7780 17312 7786
rect 17267 7762 17285 7780
rect 17303 7762 17312 7780
rect 17607 7773 17617 7791
rect 17635 7773 17654 7791
rect 17607 7769 17654 7773
rect 17608 7764 17645 7769
rect 17267 7752 17312 7762
rect 18675 7761 18712 7832
rect 18893 7831 19234 7832
rect 18827 7771 18858 7772
rect 16990 7734 17027 7735
rect 16940 7725 17027 7734
rect 16940 7705 16998 7725
rect 17018 7705 17027 7725
rect 16940 7695 17027 7705
rect 17086 7725 17123 7735
rect 17086 7705 17094 7725
rect 17114 7705 17123 7725
rect 17267 7710 17310 7752
rect 18675 7741 18684 7761
rect 18704 7741 18712 7761
rect 18675 7731 18712 7741
rect 18771 7761 18858 7771
rect 18771 7741 18780 7761
rect 18800 7741 18858 7761
rect 18771 7732 18858 7741
rect 18771 7731 18808 7732
rect 17173 7708 17310 7710
rect 16940 7694 16971 7695
rect 17086 7635 17123 7705
rect 16564 7634 16905 7635
rect 16294 7617 16332 7626
rect 16489 7629 16905 7634
rect 16294 7616 16331 7617
rect 15755 7588 15845 7594
rect 15755 7568 15771 7588
rect 15791 7586 15845 7588
rect 15791 7568 15816 7586
rect 15755 7566 15816 7568
rect 15836 7566 15845 7586
rect 15755 7560 15845 7566
rect 15768 7506 15805 7507
rect 15864 7506 15901 7507
rect 15920 7506 15956 7616
rect 16143 7595 16174 7616
rect 16489 7609 16492 7629
rect 16512 7609 16905 7629
rect 17089 7619 17123 7635
rect 17167 7687 17310 7708
rect 17596 7702 17648 7704
rect 16865 7600 16905 7609
rect 17167 7600 17194 7687
rect 17267 7661 17310 7687
rect 17267 7643 17280 7661
rect 17298 7643 17310 7661
rect 17594 7698 18027 7702
rect 17594 7692 18033 7698
rect 17594 7674 17615 7692
rect 17633 7674 18033 7692
rect 18827 7681 18858 7732
rect 18893 7761 18930 7831
rect 19196 7830 19233 7831
rect 19045 7771 19081 7772
rect 18893 7741 18902 7761
rect 18922 7741 18930 7761
rect 18893 7731 18930 7741
rect 18989 7761 19137 7771
rect 19237 7768 19333 7770
rect 18989 7741 18998 7761
rect 19018 7741 19108 7761
rect 19128 7741 19137 7761
rect 18989 7732 19137 7741
rect 19195 7761 19333 7768
rect 19195 7741 19204 7761
rect 19224 7741 19333 7761
rect 19195 7732 19333 7741
rect 18989 7731 19026 7732
rect 18719 7678 18760 7679
rect 17594 7656 18033 7674
rect 17267 7632 17310 7643
rect 16139 7594 16174 7595
rect 16017 7584 16174 7594
rect 16017 7564 16034 7584
rect 16054 7564 16174 7584
rect 16017 7557 16174 7564
rect 16241 7587 16390 7595
rect 16241 7567 16252 7587
rect 16272 7567 16311 7587
rect 16331 7567 16390 7587
rect 16865 7583 17194 7600
rect 16865 7582 16905 7583
rect 16241 7560 16390 7567
rect 17262 7571 17302 7574
rect 17262 7565 17305 7571
rect 16887 7562 17305 7565
rect 16241 7559 16282 7560
rect 15975 7506 16012 7507
rect 15668 7497 15806 7506
rect 15531 7487 15567 7493
rect 15531 7469 15536 7487
rect 15558 7469 15567 7487
rect 15531 7465 15567 7469
rect 15668 7477 15777 7497
rect 15797 7477 15806 7497
rect 15668 7470 15806 7477
rect 15864 7497 16012 7506
rect 15864 7477 15873 7497
rect 15893 7477 15983 7497
rect 16003 7477 16012 7497
rect 15668 7468 15764 7470
rect 15864 7467 16012 7477
rect 16071 7497 16108 7507
rect 16071 7477 16079 7497
rect 16099 7477 16108 7497
rect 15920 7466 15956 7467
rect 15534 7306 15567 7465
rect 15768 7407 15805 7408
rect 16071 7407 16108 7477
rect 16143 7506 16174 7557
rect 16887 7544 17278 7562
rect 17296 7544 17305 7562
rect 16887 7542 17305 7544
rect 16887 7534 16914 7542
rect 17155 7539 17305 7542
rect 16467 7528 16635 7529
rect 16886 7528 16914 7534
rect 16467 7512 16914 7528
rect 17262 7534 17305 7539
rect 16193 7506 16230 7507
rect 16143 7497 16230 7506
rect 16143 7477 16201 7497
rect 16221 7477 16230 7497
rect 16143 7467 16230 7477
rect 16289 7497 16326 7507
rect 16289 7477 16297 7497
rect 16317 7477 16326 7497
rect 16143 7466 16174 7467
rect 15767 7406 16108 7407
rect 16289 7406 16326 7477
rect 15692 7401 16108 7406
rect 15692 7381 15695 7401
rect 15715 7381 16108 7401
rect 16139 7382 16326 7406
rect 16467 7502 16911 7512
rect 16467 7500 16635 7502
rect 16467 7322 16494 7500
rect 16534 7462 16598 7474
rect 16874 7470 16911 7502
rect 16937 7501 17128 7523
rect 17092 7499 17128 7501
rect 17092 7470 17129 7499
rect 17262 7478 17302 7534
rect 16534 7461 16569 7462
rect 16511 7456 16569 7461
rect 16511 7436 16514 7456
rect 16534 7442 16569 7456
rect 16589 7442 16598 7462
rect 16534 7434 16598 7442
rect 16560 7433 16598 7434
rect 16561 7432 16598 7433
rect 16664 7466 16700 7467
rect 16772 7466 16808 7467
rect 16664 7458 16808 7466
rect 16664 7438 16672 7458
rect 16692 7438 16727 7458
rect 16747 7438 16780 7458
rect 16800 7438 16808 7458
rect 16664 7432 16808 7438
rect 16874 7462 16912 7470
rect 16990 7466 17026 7467
rect 16874 7442 16883 7462
rect 16903 7442 16912 7462
rect 16874 7433 16912 7442
rect 16941 7458 17026 7466
rect 16941 7438 16998 7458
rect 17018 7438 17026 7458
rect 16874 7432 16911 7433
rect 16941 7432 17026 7438
rect 17092 7462 17130 7470
rect 17092 7442 17101 7462
rect 17121 7442 17130 7462
rect 17262 7460 17274 7478
rect 17292 7460 17302 7478
rect 17262 7450 17302 7460
rect 17596 7467 17648 7656
rect 17994 7631 18033 7656
rect 18611 7671 18760 7678
rect 18611 7651 18670 7671
rect 18690 7651 18729 7671
rect 18749 7651 18760 7671
rect 18611 7643 18760 7651
rect 18827 7674 18984 7681
rect 18827 7654 18947 7674
rect 18967 7654 18984 7674
rect 18827 7644 18984 7654
rect 18827 7643 18862 7644
rect 17778 7606 17965 7630
rect 17994 7611 18389 7631
rect 18409 7611 18412 7631
rect 18827 7622 18858 7643
rect 19045 7622 19081 7732
rect 19100 7731 19137 7732
rect 19196 7731 19233 7732
rect 19156 7672 19246 7678
rect 19156 7652 19165 7672
rect 19185 7670 19246 7672
rect 19185 7652 19210 7670
rect 19156 7650 19210 7652
rect 19230 7650 19246 7670
rect 19156 7644 19246 7650
rect 18670 7621 18707 7622
rect 17994 7606 18412 7611
rect 18669 7612 18707 7621
rect 17778 7535 17815 7606
rect 17994 7605 18337 7606
rect 17994 7602 18033 7605
rect 18299 7604 18336 7605
rect 17930 7545 17961 7546
rect 17778 7515 17787 7535
rect 17807 7515 17815 7535
rect 17778 7505 17815 7515
rect 17874 7535 17961 7545
rect 17874 7515 17883 7535
rect 17903 7515 17961 7535
rect 17874 7506 17961 7515
rect 17874 7505 17911 7506
rect 17092 7433 17130 7442
rect 17596 7449 17612 7467
rect 17630 7449 17648 7467
rect 17930 7455 17961 7506
rect 17996 7535 18033 7602
rect 18669 7592 18678 7612
rect 18698 7592 18707 7612
rect 18669 7584 18707 7592
rect 18773 7616 18858 7622
rect 18888 7621 18925 7622
rect 18773 7596 18781 7616
rect 18801 7596 18858 7616
rect 18773 7588 18858 7596
rect 18887 7612 18925 7621
rect 18887 7592 18896 7612
rect 18916 7592 18925 7612
rect 18773 7587 18809 7588
rect 18887 7584 18925 7592
rect 18991 7617 19135 7622
rect 18991 7616 19053 7617
rect 18991 7596 18999 7616
rect 19019 7598 19053 7616
rect 19074 7616 19135 7617
rect 19074 7598 19107 7616
rect 19019 7596 19107 7598
rect 19127 7596 19135 7616
rect 18991 7588 19135 7596
rect 18991 7587 19027 7588
rect 19099 7587 19135 7588
rect 19201 7621 19238 7622
rect 19201 7620 19239 7621
rect 19201 7612 19265 7620
rect 19201 7592 19210 7612
rect 19230 7598 19265 7612
rect 19285 7598 19288 7618
rect 19230 7593 19288 7598
rect 19230 7592 19265 7593
rect 18670 7555 18707 7584
rect 18671 7553 18707 7555
rect 18148 7545 18184 7546
rect 17996 7515 18005 7535
rect 18025 7515 18033 7535
rect 17996 7505 18033 7515
rect 18092 7535 18240 7545
rect 18340 7542 18436 7544
rect 18092 7515 18101 7535
rect 18121 7515 18211 7535
rect 18231 7515 18240 7535
rect 18092 7506 18240 7515
rect 18298 7535 18436 7542
rect 18298 7515 18307 7535
rect 18327 7515 18436 7535
rect 18671 7531 18862 7553
rect 18888 7552 18925 7584
rect 19201 7580 19265 7592
rect 19305 7554 19332 7732
rect 19164 7552 19332 7554
rect 18888 7538 19332 7552
rect 19935 7686 20103 7687
rect 20229 7686 20269 7910
rect 20732 7914 20900 7915
rect 21135 7914 21175 7947
rect 21531 7914 21578 7947
rect 21969 7946 22010 7971
rect 22155 7946 22192 7977
rect 22373 7946 22410 7977
rect 22686 7973 22750 7985
rect 22790 7947 22817 8125
rect 21969 7919 22018 7946
rect 22154 7920 22203 7946
rect 22372 7945 22453 7946
rect 22649 7945 22817 7947
rect 22372 7920 22817 7945
rect 22373 7919 22817 7920
rect 20732 7913 21176 7914
rect 20732 7888 21177 7913
rect 20732 7886 20900 7888
rect 21096 7887 21177 7888
rect 21346 7887 21395 7913
rect 21531 7887 21580 7914
rect 20732 7708 20759 7886
rect 20799 7848 20863 7860
rect 21139 7856 21176 7887
rect 21357 7856 21394 7887
rect 21539 7862 21580 7887
rect 21971 7886 22018 7919
rect 22374 7886 22414 7919
rect 22649 7918 22817 7919
rect 23280 7923 23320 8147
rect 23446 8146 23614 8147
rect 24217 8281 24661 8295
rect 24217 8279 24385 8281
rect 24217 8101 24244 8279
rect 24284 8241 24348 8253
rect 24624 8249 24661 8281
rect 24687 8280 24878 8302
rect 25113 8298 25222 8318
rect 25242 8298 25251 8318
rect 25113 8291 25251 8298
rect 25309 8318 25457 8327
rect 25309 8298 25318 8318
rect 25338 8298 25428 8318
rect 25448 8298 25457 8318
rect 25113 8289 25209 8291
rect 25309 8288 25457 8298
rect 25516 8318 25553 8328
rect 25516 8298 25524 8318
rect 25544 8298 25553 8318
rect 25365 8287 25401 8288
rect 24842 8278 24878 8280
rect 24842 8249 24879 8278
rect 24284 8240 24319 8241
rect 24261 8235 24319 8240
rect 24261 8215 24264 8235
rect 24284 8221 24319 8235
rect 24339 8221 24348 8241
rect 24284 8213 24348 8221
rect 24310 8212 24348 8213
rect 24311 8211 24348 8212
rect 24414 8245 24450 8246
rect 24522 8245 24558 8246
rect 24414 8239 24558 8245
rect 24414 8237 24475 8239
rect 24414 8217 24422 8237
rect 24442 8222 24475 8237
rect 24494 8237 24558 8239
rect 24494 8222 24530 8237
rect 24442 8217 24530 8222
rect 24550 8217 24558 8237
rect 24414 8211 24558 8217
rect 24624 8241 24662 8249
rect 24740 8245 24776 8246
rect 24624 8221 24633 8241
rect 24653 8221 24662 8241
rect 24624 8212 24662 8221
rect 24691 8237 24776 8245
rect 24691 8217 24748 8237
rect 24768 8217 24776 8237
rect 24624 8211 24661 8212
rect 24691 8211 24776 8217
rect 24842 8241 24880 8249
rect 24842 8221 24851 8241
rect 24871 8221 24880 8241
rect 25516 8231 25553 8298
rect 25588 8327 25619 8378
rect 25901 8366 25919 8384
rect 25937 8366 25953 8384
rect 25638 8327 25675 8328
rect 25588 8318 25675 8327
rect 25588 8298 25646 8318
rect 25666 8298 25675 8318
rect 25588 8288 25675 8298
rect 25734 8318 25771 8328
rect 25734 8298 25742 8318
rect 25762 8298 25771 8318
rect 25588 8287 25619 8288
rect 25213 8228 25250 8229
rect 25516 8228 25555 8231
rect 25212 8227 25555 8228
rect 25734 8227 25771 8298
rect 24842 8212 24880 8221
rect 25137 8222 25555 8227
rect 24842 8211 24879 8212
rect 24303 8183 24393 8189
rect 24303 8163 24319 8183
rect 24339 8181 24393 8183
rect 24339 8163 24364 8181
rect 24303 8161 24364 8163
rect 24384 8161 24393 8181
rect 24303 8155 24393 8161
rect 24316 8101 24353 8102
rect 24412 8101 24449 8102
rect 24468 8101 24504 8211
rect 24691 8190 24722 8211
rect 25137 8202 25140 8222
rect 25160 8202 25555 8222
rect 25584 8203 25771 8227
rect 24687 8189 24722 8190
rect 24565 8179 24722 8189
rect 24565 8159 24582 8179
rect 24602 8159 24722 8179
rect 24565 8152 24722 8159
rect 24789 8182 24938 8190
rect 24789 8162 24800 8182
rect 24820 8162 24859 8182
rect 24879 8162 24938 8182
rect 24789 8155 24938 8162
rect 25516 8177 25555 8202
rect 25901 8177 25953 8366
rect 26358 8393 26368 8411
rect 26386 8393 26398 8411
rect 26530 8409 26539 8429
rect 26559 8409 26568 8429
rect 26530 8401 26568 8409
rect 26634 8433 26719 8439
rect 26749 8438 26786 8439
rect 26634 8413 26642 8433
rect 26662 8413 26719 8433
rect 26634 8405 26719 8413
rect 26748 8429 26786 8438
rect 26748 8409 26757 8429
rect 26777 8409 26786 8429
rect 26634 8404 26670 8405
rect 26748 8401 26786 8409
rect 26852 8433 26996 8439
rect 26852 8413 26860 8433
rect 26880 8413 26913 8433
rect 26933 8413 26968 8433
rect 26988 8413 26996 8433
rect 26852 8405 26996 8413
rect 26852 8404 26888 8405
rect 26960 8404 26996 8405
rect 27062 8438 27099 8439
rect 27062 8437 27100 8438
rect 27062 8429 27126 8437
rect 27062 8409 27071 8429
rect 27091 8415 27126 8429
rect 27146 8415 27149 8435
rect 27091 8410 27149 8415
rect 27091 8409 27126 8410
rect 26358 8337 26398 8393
rect 26531 8372 26568 8401
rect 26532 8370 26568 8372
rect 26532 8348 26723 8370
rect 26749 8369 26786 8401
rect 27062 8397 27126 8409
rect 27166 8371 27193 8549
rect 27025 8369 27193 8371
rect 26749 8359 27193 8369
rect 27334 8465 27521 8489
rect 27552 8470 27945 8490
rect 27965 8470 27968 8490
rect 27552 8465 27968 8470
rect 27334 8394 27371 8465
rect 27552 8464 27893 8465
rect 27486 8404 27517 8405
rect 27334 8374 27343 8394
rect 27363 8374 27371 8394
rect 27334 8364 27371 8374
rect 27430 8394 27517 8404
rect 27430 8374 27439 8394
rect 27459 8374 27517 8394
rect 27430 8365 27517 8374
rect 27430 8364 27467 8365
rect 26355 8332 26398 8337
rect 26746 8343 27193 8359
rect 26746 8337 26774 8343
rect 27025 8342 27193 8343
rect 26355 8329 26505 8332
rect 26746 8329 26773 8337
rect 26355 8327 26773 8329
rect 26355 8309 26364 8327
rect 26382 8309 26773 8327
rect 27486 8314 27517 8365
rect 27552 8394 27589 8464
rect 27855 8463 27892 8464
rect 27704 8404 27740 8405
rect 27552 8374 27561 8394
rect 27581 8374 27589 8394
rect 27552 8364 27589 8374
rect 27648 8394 27796 8404
rect 27896 8401 27992 8403
rect 27648 8374 27657 8394
rect 27677 8374 27767 8394
rect 27787 8374 27796 8394
rect 27648 8365 27796 8374
rect 27854 8394 27992 8401
rect 27854 8374 27863 8394
rect 27883 8374 27992 8394
rect 27854 8365 27992 8374
rect 27648 8364 27685 8365
rect 27378 8311 27419 8312
rect 26355 8306 26773 8309
rect 26355 8300 26398 8306
rect 26358 8297 26398 8300
rect 27270 8304 27419 8311
rect 26755 8288 26795 8289
rect 26466 8271 26795 8288
rect 27270 8284 27329 8304
rect 27349 8284 27388 8304
rect 27408 8284 27419 8304
rect 27270 8276 27419 8284
rect 27486 8307 27643 8314
rect 27486 8287 27606 8307
rect 27626 8287 27643 8307
rect 27486 8277 27643 8287
rect 27486 8276 27521 8277
rect 26350 8228 26393 8239
rect 26350 8210 26362 8228
rect 26380 8210 26393 8228
rect 26350 8184 26393 8210
rect 26466 8184 26493 8271
rect 26755 8262 26795 8271
rect 25516 8159 25955 8177
rect 24789 8154 24830 8155
rect 24523 8101 24560 8102
rect 24216 8092 24354 8101
rect 24216 8072 24325 8092
rect 24345 8072 24354 8092
rect 24216 8065 24354 8072
rect 24412 8092 24560 8101
rect 24412 8072 24421 8092
rect 24441 8072 24531 8092
rect 24551 8072 24560 8092
rect 24216 8063 24312 8065
rect 24412 8062 24560 8072
rect 24619 8092 24656 8102
rect 24619 8072 24627 8092
rect 24647 8072 24656 8092
rect 24468 8061 24504 8062
rect 24316 8002 24353 8003
rect 24619 8002 24656 8072
rect 24691 8101 24722 8152
rect 25516 8141 25916 8159
rect 25934 8141 25955 8159
rect 25516 8135 25955 8141
rect 25522 8131 25955 8135
rect 26350 8163 26493 8184
rect 26537 8236 26571 8252
rect 26755 8242 27148 8262
rect 27168 8242 27171 8262
rect 27486 8255 27517 8276
rect 27704 8255 27740 8365
rect 27759 8364 27796 8365
rect 27855 8364 27892 8365
rect 27815 8305 27905 8311
rect 27815 8285 27824 8305
rect 27844 8303 27905 8305
rect 27844 8285 27869 8303
rect 27815 8283 27869 8285
rect 27889 8283 27905 8303
rect 27815 8277 27905 8283
rect 27329 8254 27366 8255
rect 26755 8237 27171 8242
rect 27328 8245 27366 8254
rect 26755 8236 27096 8237
rect 26537 8166 26574 8236
rect 26689 8176 26720 8177
rect 26350 8161 26487 8163
rect 25901 8129 25953 8131
rect 26350 8119 26393 8161
rect 26537 8146 26546 8166
rect 26566 8146 26574 8166
rect 26537 8136 26574 8146
rect 26633 8166 26720 8176
rect 26633 8146 26642 8166
rect 26662 8146 26720 8166
rect 26633 8137 26720 8146
rect 26633 8136 26670 8137
rect 26348 8109 26393 8119
rect 24741 8101 24778 8102
rect 24691 8092 24778 8101
rect 24691 8072 24749 8092
rect 24769 8072 24778 8092
rect 24691 8062 24778 8072
rect 24837 8092 24874 8102
rect 24837 8072 24845 8092
rect 24865 8072 24874 8092
rect 26348 8091 26357 8109
rect 26375 8091 26393 8109
rect 26348 8085 26393 8091
rect 26689 8086 26720 8137
rect 26755 8166 26792 8236
rect 27058 8235 27095 8236
rect 27328 8225 27337 8245
rect 27357 8225 27366 8245
rect 27328 8217 27366 8225
rect 27432 8249 27517 8255
rect 27547 8254 27584 8255
rect 27432 8229 27440 8249
rect 27460 8229 27517 8249
rect 27432 8221 27517 8229
rect 27546 8245 27584 8254
rect 27546 8225 27555 8245
rect 27575 8225 27584 8245
rect 27432 8220 27468 8221
rect 27546 8217 27584 8225
rect 27650 8249 27794 8255
rect 27650 8229 27658 8249
rect 27678 8230 27710 8249
rect 27731 8230 27766 8249
rect 27678 8229 27766 8230
rect 27786 8229 27794 8249
rect 27650 8221 27794 8229
rect 27650 8220 27686 8221
rect 27758 8220 27794 8221
rect 27860 8254 27897 8255
rect 27860 8253 27898 8254
rect 27860 8245 27924 8253
rect 27860 8225 27869 8245
rect 27889 8231 27924 8245
rect 27944 8231 27947 8251
rect 27889 8226 27947 8231
rect 27889 8225 27924 8226
rect 27329 8188 27366 8217
rect 27330 8186 27366 8188
rect 26907 8176 26943 8177
rect 26755 8146 26764 8166
rect 26784 8146 26792 8166
rect 26755 8136 26792 8146
rect 26851 8166 26999 8176
rect 27099 8173 27195 8175
rect 26851 8146 26860 8166
rect 26880 8146 26970 8166
rect 26990 8146 26999 8166
rect 26851 8137 26999 8146
rect 27057 8166 27195 8173
rect 27057 8146 27066 8166
rect 27086 8146 27195 8166
rect 27330 8164 27521 8186
rect 27547 8185 27584 8217
rect 27860 8213 27924 8225
rect 27964 8187 27991 8365
rect 28596 8364 28629 8697
rect 28693 8729 28861 8730
rect 28987 8729 29027 8953
rect 29490 8957 29658 8958
rect 29891 8957 29936 8978
rect 29490 8931 29936 8957
rect 29490 8929 29658 8931
rect 29854 8930 29936 8931
rect 30071 8930 30152 8956
rect 30296 8943 30777 8978
rect 33351 8966 33359 8988
rect 33383 8966 33391 8988
rect 29490 8751 29517 8929
rect 29557 8891 29621 8903
rect 29897 8899 29934 8930
rect 30115 8899 30152 8930
rect 30299 8924 30338 8943
rect 30297 8905 30338 8924
rect 29557 8890 29592 8891
rect 29534 8885 29592 8890
rect 29534 8865 29537 8885
rect 29557 8871 29592 8885
rect 29612 8871 29621 8891
rect 29557 8863 29621 8871
rect 29583 8862 29621 8863
rect 29584 8861 29621 8862
rect 29687 8895 29723 8896
rect 29795 8895 29831 8896
rect 29687 8887 29831 8895
rect 29687 8867 29695 8887
rect 29715 8883 29803 8887
rect 29715 8867 29759 8883
rect 29687 8863 29759 8867
rect 29779 8867 29803 8883
rect 29823 8867 29831 8887
rect 29779 8863 29831 8867
rect 29687 8861 29831 8863
rect 29897 8891 29935 8899
rect 30013 8895 30049 8896
rect 29897 8871 29906 8891
rect 29926 8871 29935 8891
rect 29897 8862 29935 8871
rect 29964 8887 30049 8895
rect 29964 8867 30021 8887
rect 30041 8867 30049 8887
rect 29897 8861 29934 8862
rect 29964 8861 30049 8867
rect 30115 8891 30153 8899
rect 30115 8871 30124 8891
rect 30144 8871 30153 8891
rect 30115 8862 30153 8871
rect 30297 8896 30339 8905
rect 30297 8878 30311 8896
rect 30329 8878 30339 8896
rect 30297 8870 30339 8878
rect 30302 8868 30339 8870
rect 30115 8861 30152 8862
rect 29576 8833 29666 8839
rect 29576 8813 29592 8833
rect 29612 8831 29666 8833
rect 29612 8813 29637 8831
rect 29576 8811 29637 8813
rect 29657 8811 29666 8831
rect 29576 8805 29666 8811
rect 29589 8751 29626 8752
rect 29685 8751 29722 8752
rect 29741 8751 29777 8861
rect 29964 8840 29995 8861
rect 30729 8847 30776 8943
rect 29960 8839 29995 8840
rect 29838 8829 29995 8839
rect 29838 8809 29855 8829
rect 29875 8809 29995 8829
rect 29838 8802 29995 8809
rect 30062 8832 30211 8840
rect 30062 8812 30073 8832
rect 30093 8812 30132 8832
rect 30152 8812 30211 8832
rect 30729 8829 30739 8847
rect 30757 8829 30776 8847
rect 30729 8825 30776 8829
rect 30730 8820 30767 8825
rect 30062 8805 30211 8812
rect 30062 8804 30103 8805
rect 30299 8803 30336 8806
rect 29796 8751 29833 8752
rect 29489 8742 29627 8751
rect 28693 8703 29137 8729
rect 28693 8701 28861 8703
rect 28693 8523 28720 8701
rect 28760 8663 28824 8675
rect 29100 8671 29137 8703
rect 29163 8702 29354 8724
rect 29489 8722 29598 8742
rect 29618 8722 29627 8742
rect 29489 8715 29627 8722
rect 29685 8742 29833 8751
rect 29685 8722 29694 8742
rect 29714 8722 29804 8742
rect 29824 8722 29833 8742
rect 29489 8713 29585 8715
rect 29685 8712 29833 8722
rect 29892 8742 29929 8752
rect 29892 8722 29900 8742
rect 29920 8722 29929 8742
rect 29741 8711 29777 8712
rect 29318 8700 29354 8702
rect 29318 8671 29355 8700
rect 28760 8662 28795 8663
rect 28737 8657 28795 8662
rect 28737 8637 28740 8657
rect 28760 8643 28795 8657
rect 28815 8643 28824 8663
rect 28760 8637 28824 8643
rect 28737 8635 28824 8637
rect 28737 8631 28764 8635
rect 28786 8634 28824 8635
rect 28787 8633 28824 8634
rect 28890 8667 28926 8668
rect 28998 8667 29034 8668
rect 28890 8660 29034 8667
rect 28890 8659 28952 8660
rect 28890 8639 28898 8659
rect 28918 8642 28952 8659
rect 28971 8659 29034 8660
rect 28971 8642 29006 8659
rect 28918 8639 29006 8642
rect 29026 8639 29034 8659
rect 28890 8633 29034 8639
rect 29100 8663 29138 8671
rect 29216 8667 29252 8668
rect 29100 8643 29109 8663
rect 29129 8643 29138 8663
rect 29100 8634 29138 8643
rect 29167 8659 29252 8667
rect 29167 8639 29224 8659
rect 29244 8639 29252 8659
rect 29100 8633 29137 8634
rect 29167 8633 29252 8639
rect 29318 8663 29356 8671
rect 29318 8643 29327 8663
rect 29347 8643 29356 8663
rect 29589 8652 29626 8653
rect 29892 8652 29929 8722
rect 29964 8751 29995 8802
rect 30291 8797 30336 8803
rect 30291 8779 30309 8797
rect 30327 8779 30336 8797
rect 30291 8769 30336 8779
rect 30014 8751 30051 8752
rect 29964 8742 30051 8751
rect 29964 8722 30022 8742
rect 30042 8722 30051 8742
rect 29964 8712 30051 8722
rect 30110 8742 30147 8752
rect 30110 8722 30118 8742
rect 30138 8722 30147 8742
rect 30291 8727 30334 8769
rect 30718 8758 30770 8760
rect 30197 8725 30334 8727
rect 29964 8711 29995 8712
rect 30110 8652 30147 8722
rect 29588 8651 29929 8652
rect 29318 8634 29356 8643
rect 29513 8646 29929 8651
rect 29318 8633 29355 8634
rect 28779 8605 28869 8611
rect 28779 8585 28795 8605
rect 28815 8603 28869 8605
rect 28815 8585 28840 8603
rect 28779 8583 28840 8585
rect 28860 8583 28869 8603
rect 28779 8577 28869 8583
rect 28792 8523 28829 8524
rect 28888 8523 28925 8524
rect 28944 8523 28980 8633
rect 29167 8612 29198 8633
rect 29513 8626 29516 8646
rect 29536 8626 29929 8646
rect 30113 8636 30147 8652
rect 30191 8704 30334 8725
rect 30716 8754 31149 8758
rect 30716 8748 31155 8754
rect 30716 8730 30737 8748
rect 30755 8730 31155 8748
rect 30716 8712 31155 8730
rect 29889 8617 29929 8626
rect 30191 8617 30218 8704
rect 30291 8678 30334 8704
rect 30291 8660 30304 8678
rect 30322 8660 30334 8678
rect 30291 8649 30334 8660
rect 29163 8611 29198 8612
rect 29041 8601 29198 8611
rect 29041 8581 29058 8601
rect 29078 8581 29198 8601
rect 29041 8574 29198 8581
rect 29265 8604 29411 8612
rect 29265 8584 29276 8604
rect 29296 8584 29335 8604
rect 29355 8584 29411 8604
rect 29889 8600 30218 8617
rect 29889 8599 29929 8600
rect 29265 8577 29411 8584
rect 30286 8588 30326 8591
rect 30286 8582 30329 8588
rect 29911 8579 30329 8582
rect 29265 8576 29306 8577
rect 28999 8523 29036 8524
rect 28692 8514 28830 8523
rect 28692 8494 28801 8514
rect 28821 8494 28830 8514
rect 28692 8487 28830 8494
rect 28888 8514 29036 8523
rect 28888 8494 28897 8514
rect 28917 8494 29007 8514
rect 29027 8494 29036 8514
rect 28692 8485 28788 8487
rect 28888 8484 29036 8494
rect 29095 8514 29132 8524
rect 29095 8494 29103 8514
rect 29123 8494 29132 8514
rect 28944 8483 28980 8484
rect 28792 8424 28829 8425
rect 29095 8424 29132 8494
rect 29167 8523 29198 8574
rect 29911 8561 30302 8579
rect 30320 8561 30329 8579
rect 29911 8559 30329 8561
rect 29911 8551 29938 8559
rect 30179 8556 30329 8559
rect 29491 8545 29659 8546
rect 29910 8545 29938 8551
rect 29491 8529 29938 8545
rect 30286 8551 30329 8556
rect 29217 8523 29254 8524
rect 29167 8514 29254 8523
rect 29167 8494 29225 8514
rect 29245 8494 29254 8514
rect 29167 8484 29254 8494
rect 29313 8514 29350 8524
rect 29313 8494 29321 8514
rect 29341 8494 29350 8514
rect 29167 8483 29198 8484
rect 28791 8423 29132 8424
rect 29313 8423 29350 8494
rect 28716 8418 29132 8423
rect 28716 8398 28719 8418
rect 28739 8398 29132 8418
rect 29163 8399 29350 8423
rect 29491 8519 29935 8529
rect 29491 8517 29659 8519
rect 28591 8319 28633 8364
rect 29491 8339 29518 8517
rect 29558 8479 29622 8491
rect 29898 8487 29935 8519
rect 29961 8518 30152 8540
rect 30116 8516 30152 8518
rect 30116 8487 30153 8516
rect 30286 8495 30326 8551
rect 29558 8478 29593 8479
rect 29535 8473 29593 8478
rect 29535 8453 29538 8473
rect 29558 8459 29593 8473
rect 29613 8459 29622 8479
rect 29558 8451 29622 8459
rect 29584 8450 29622 8451
rect 29585 8449 29622 8450
rect 29688 8483 29724 8484
rect 29796 8483 29832 8484
rect 29688 8475 29832 8483
rect 29688 8455 29696 8475
rect 29716 8455 29751 8475
rect 29771 8455 29804 8475
rect 29824 8455 29832 8475
rect 29688 8449 29832 8455
rect 29898 8479 29936 8487
rect 30014 8483 30050 8484
rect 29898 8459 29907 8479
rect 29927 8459 29936 8479
rect 29898 8450 29936 8459
rect 29965 8475 30050 8483
rect 29965 8455 30022 8475
rect 30042 8455 30050 8475
rect 29898 8449 29935 8450
rect 29965 8449 30050 8455
rect 30116 8479 30154 8487
rect 30116 8459 30125 8479
rect 30145 8459 30154 8479
rect 30286 8477 30298 8495
rect 30316 8477 30326 8495
rect 30718 8523 30770 8712
rect 31116 8687 31155 8712
rect 32956 8737 32993 8743
rect 32956 8718 32964 8737
rect 32985 8718 32993 8737
rect 32956 8710 32993 8718
rect 30900 8662 31087 8686
rect 31116 8667 31511 8687
rect 31531 8667 31534 8687
rect 31116 8662 31534 8667
rect 30900 8591 30937 8662
rect 31116 8661 31459 8662
rect 31116 8658 31155 8661
rect 31421 8660 31458 8661
rect 31052 8601 31083 8602
rect 30900 8571 30909 8591
rect 30929 8571 30937 8591
rect 30900 8561 30937 8571
rect 30996 8591 31083 8601
rect 30996 8571 31005 8591
rect 31025 8571 31083 8591
rect 30996 8562 31083 8571
rect 30996 8561 31033 8562
rect 30718 8505 30734 8523
rect 30752 8505 30770 8523
rect 31052 8511 31083 8562
rect 31118 8591 31155 8658
rect 31270 8601 31306 8602
rect 31118 8571 31127 8591
rect 31147 8571 31155 8591
rect 31118 8561 31155 8571
rect 31214 8591 31362 8601
rect 31462 8598 31558 8600
rect 31214 8571 31223 8591
rect 31243 8571 31333 8591
rect 31353 8571 31362 8591
rect 31214 8562 31362 8571
rect 31420 8591 31558 8598
rect 31420 8571 31429 8591
rect 31449 8571 31558 8591
rect 31420 8562 31558 8571
rect 31214 8561 31251 8562
rect 30944 8508 30985 8509
rect 30718 8487 30770 8505
rect 30836 8501 30985 8508
rect 30286 8467 30326 8477
rect 30836 8481 30895 8501
rect 30915 8481 30954 8501
rect 30974 8481 30985 8501
rect 30836 8473 30985 8481
rect 31052 8504 31209 8511
rect 31052 8484 31172 8504
rect 31192 8484 31209 8504
rect 31052 8474 31209 8484
rect 31052 8473 31087 8474
rect 30116 8450 30154 8459
rect 31052 8452 31083 8473
rect 31270 8452 31306 8562
rect 31325 8561 31362 8562
rect 31421 8561 31458 8562
rect 31381 8502 31471 8508
rect 31381 8482 31390 8502
rect 31410 8500 31471 8502
rect 31410 8482 31435 8500
rect 31381 8480 31435 8482
rect 31455 8480 31471 8500
rect 31381 8474 31471 8480
rect 30895 8451 30932 8452
rect 30116 8449 30153 8450
rect 29577 8421 29667 8427
rect 29577 8401 29593 8421
rect 29613 8419 29667 8421
rect 29613 8401 29638 8419
rect 29577 8399 29638 8401
rect 29658 8399 29667 8419
rect 29577 8393 29667 8399
rect 29590 8339 29627 8340
rect 29686 8339 29723 8340
rect 29742 8339 29778 8449
rect 29965 8428 29996 8449
rect 30894 8442 30932 8451
rect 29961 8427 29996 8428
rect 29839 8417 29996 8427
rect 29839 8397 29856 8417
rect 29876 8397 29996 8417
rect 29839 8390 29996 8397
rect 30063 8420 30212 8428
rect 30063 8400 30074 8420
rect 30094 8400 30133 8420
rect 30153 8400 30212 8420
rect 30722 8424 30762 8434
rect 30063 8393 30212 8400
rect 30278 8396 30330 8414
rect 30063 8392 30104 8393
rect 29797 8339 29834 8340
rect 29490 8330 29628 8339
rect 28962 8319 28995 8321
rect 28591 8307 29038 8319
rect 27823 8185 27991 8187
rect 27547 8159 27991 8185
rect 27057 8137 27195 8146
rect 26851 8136 26888 8137
rect 26348 8082 26385 8085
rect 26581 8083 26622 8084
rect 24691 8061 24722 8062
rect 24315 8001 24656 8002
rect 24837 8001 24874 8072
rect 26473 8076 26622 8083
rect 25904 8064 25941 8069
rect 25895 8060 25942 8064
rect 25895 8042 25914 8060
rect 25932 8042 25942 8060
rect 26473 8056 26532 8076
rect 26552 8056 26591 8076
rect 26611 8056 26622 8076
rect 26473 8048 26622 8056
rect 26689 8079 26846 8086
rect 26689 8059 26809 8079
rect 26829 8059 26846 8079
rect 26689 8049 26846 8059
rect 26689 8048 26724 8049
rect 24240 7996 24656 8001
rect 24240 7976 24243 7996
rect 24263 7976 24656 7996
rect 24687 7977 24874 8001
rect 25499 7999 25539 8004
rect 25895 7999 25942 8042
rect 26689 8027 26720 8048
rect 26907 8027 26943 8137
rect 26962 8136 26999 8137
rect 27058 8136 27095 8137
rect 27018 8077 27108 8083
rect 27018 8057 27027 8077
rect 27047 8075 27108 8077
rect 27047 8057 27072 8075
rect 27018 8055 27072 8057
rect 27092 8055 27108 8075
rect 27018 8049 27108 8055
rect 26532 8026 26569 8027
rect 25499 7960 25942 7999
rect 26345 8018 26382 8020
rect 26345 8010 26387 8018
rect 26345 7992 26355 8010
rect 26373 7992 26387 8010
rect 26345 7983 26387 7992
rect 26531 8017 26569 8026
rect 26531 7997 26540 8017
rect 26560 7997 26569 8017
rect 26531 7989 26569 7997
rect 26635 8021 26720 8027
rect 26750 8026 26787 8027
rect 26635 8001 26643 8021
rect 26663 8001 26720 8021
rect 26635 7993 26720 8001
rect 26749 8017 26787 8026
rect 26749 7997 26758 8017
rect 26778 7997 26787 8017
rect 26635 7992 26671 7993
rect 26749 7989 26787 7997
rect 26853 8025 26997 8027
rect 26853 8021 26905 8025
rect 26853 8001 26861 8021
rect 26881 8005 26905 8021
rect 26925 8021 26997 8025
rect 26925 8005 26969 8021
rect 26881 8001 26969 8005
rect 26989 8001 26997 8021
rect 26853 7993 26997 8001
rect 26853 7992 26889 7993
rect 26961 7992 26997 7993
rect 27063 8026 27100 8027
rect 27063 8025 27101 8026
rect 27063 8017 27127 8025
rect 27063 7997 27072 8017
rect 27092 8003 27127 8017
rect 27147 8003 27150 8023
rect 27092 7998 27150 8003
rect 27092 7997 27127 7998
rect 23280 7901 23288 7923
rect 23312 7901 23320 7923
rect 23280 7893 23320 7901
rect 24593 7945 24633 7953
rect 24593 7923 24601 7945
rect 24625 7923 24633 7945
rect 20799 7847 20834 7848
rect 20776 7842 20834 7847
rect 20776 7822 20779 7842
rect 20799 7828 20834 7842
rect 20854 7828 20863 7848
rect 20799 7820 20863 7828
rect 20825 7819 20863 7820
rect 20826 7818 20863 7819
rect 20929 7852 20965 7853
rect 21037 7852 21073 7853
rect 20929 7844 21073 7852
rect 20929 7824 20937 7844
rect 20957 7840 21045 7844
rect 20957 7824 21001 7840
rect 20929 7820 21001 7824
rect 21021 7824 21045 7840
rect 21065 7824 21073 7844
rect 21021 7820 21073 7824
rect 20929 7818 21073 7820
rect 21139 7848 21177 7856
rect 21255 7852 21291 7853
rect 21139 7828 21148 7848
rect 21168 7828 21177 7848
rect 21139 7819 21177 7828
rect 21206 7844 21291 7852
rect 21206 7824 21263 7844
rect 21283 7824 21291 7844
rect 21139 7818 21176 7819
rect 21206 7818 21291 7824
rect 21357 7848 21395 7856
rect 21357 7828 21366 7848
rect 21386 7828 21395 7848
rect 21357 7819 21395 7828
rect 21539 7853 21581 7862
rect 21539 7835 21553 7853
rect 21571 7835 21581 7853
rect 21539 7827 21581 7835
rect 21544 7825 21581 7827
rect 21971 7847 22414 7886
rect 21357 7818 21394 7819
rect 20818 7790 20908 7796
rect 20818 7770 20834 7790
rect 20854 7788 20908 7790
rect 20854 7770 20879 7788
rect 20818 7768 20879 7770
rect 20899 7768 20908 7788
rect 20818 7762 20908 7768
rect 20831 7708 20868 7709
rect 20927 7708 20964 7709
rect 20983 7708 21019 7818
rect 21206 7797 21237 7818
rect 21971 7804 22018 7847
rect 22374 7842 22414 7847
rect 23039 7845 23226 7869
rect 23257 7850 23650 7870
rect 23670 7850 23673 7870
rect 23257 7845 23673 7850
rect 21202 7796 21237 7797
rect 21080 7786 21237 7796
rect 21080 7766 21097 7786
rect 21117 7766 21237 7786
rect 21080 7759 21237 7766
rect 21304 7789 21453 7797
rect 21304 7769 21315 7789
rect 21335 7769 21374 7789
rect 21394 7769 21453 7789
rect 21971 7786 21981 7804
rect 21999 7786 22018 7804
rect 21971 7782 22018 7786
rect 21972 7777 22009 7782
rect 21304 7762 21453 7769
rect 23039 7774 23076 7845
rect 23257 7844 23598 7845
rect 23191 7784 23222 7785
rect 21304 7761 21345 7762
rect 21541 7760 21578 7763
rect 21038 7708 21075 7709
rect 20731 7699 20869 7708
rect 19935 7660 20379 7686
rect 19935 7658 20103 7660
rect 18888 7526 19335 7538
rect 18931 7524 18964 7526
rect 18298 7506 18436 7515
rect 18092 7505 18129 7506
rect 17822 7452 17863 7453
rect 17092 7432 17129 7433
rect 16553 7404 16643 7410
rect 16553 7384 16569 7404
rect 16589 7402 16643 7404
rect 16589 7384 16614 7402
rect 16553 7382 16614 7384
rect 16634 7382 16643 7402
rect 16553 7376 16643 7382
rect 16566 7322 16603 7323
rect 16662 7322 16699 7323
rect 16718 7322 16754 7432
rect 16941 7411 16972 7432
rect 17596 7431 17648 7449
rect 17714 7445 17863 7452
rect 17714 7425 17773 7445
rect 17793 7425 17832 7445
rect 17852 7425 17863 7445
rect 17714 7417 17863 7425
rect 17930 7448 18087 7455
rect 17930 7428 18050 7448
rect 18070 7428 18087 7448
rect 17930 7418 18087 7428
rect 17930 7417 17965 7418
rect 16937 7410 16972 7411
rect 16815 7400 16972 7410
rect 16815 7380 16832 7400
rect 16852 7380 16972 7400
rect 16815 7373 16972 7380
rect 17039 7403 17188 7411
rect 17039 7383 17050 7403
rect 17070 7383 17109 7403
rect 17129 7383 17188 7403
rect 17039 7376 17188 7383
rect 17254 7379 17306 7397
rect 17930 7396 17961 7417
rect 18148 7396 18184 7506
rect 18203 7505 18240 7506
rect 18299 7505 18336 7506
rect 18259 7446 18349 7452
rect 18259 7426 18268 7446
rect 18288 7444 18349 7446
rect 18288 7426 18313 7444
rect 18259 7424 18313 7426
rect 18333 7424 18349 7444
rect 18259 7418 18349 7424
rect 17773 7395 17810 7396
rect 17039 7375 17080 7376
rect 16773 7322 16810 7323
rect 16466 7313 16604 7322
rect 15533 7305 15570 7306
rect 15504 7304 15672 7305
rect 15798 7304 15838 7306
rect 15329 7295 15368 7301
rect 15329 7273 15337 7295
rect 15361 7273 15368 7295
rect 15031 7166 15068 7174
rect 15031 7147 15039 7166
rect 15060 7147 15068 7166
rect 15031 7141 15068 7147
rect 14633 6896 14641 6918
rect 14665 6896 14673 6918
rect 14633 6888 14673 6896
rect 12149 6842 12184 6843
rect 12126 6837 12184 6842
rect 12126 6817 12129 6837
rect 12149 6823 12184 6837
rect 12204 6823 12213 6843
rect 12149 6815 12213 6823
rect 12175 6814 12213 6815
rect 12176 6813 12213 6814
rect 12279 6847 12315 6848
rect 12387 6847 12423 6848
rect 12279 6839 12423 6847
rect 12279 6819 12287 6839
rect 12307 6835 12395 6839
rect 12307 6819 12351 6835
rect 12279 6815 12351 6819
rect 12371 6819 12395 6835
rect 12415 6819 12423 6839
rect 12371 6815 12423 6819
rect 12279 6813 12423 6815
rect 12489 6843 12527 6851
rect 12605 6847 12641 6848
rect 12489 6823 12498 6843
rect 12518 6823 12527 6843
rect 12489 6814 12527 6823
rect 12556 6839 12641 6847
rect 12556 6819 12613 6839
rect 12633 6819 12641 6839
rect 12489 6813 12526 6814
rect 12556 6813 12641 6819
rect 12707 6843 12745 6851
rect 12707 6823 12716 6843
rect 12736 6823 12745 6843
rect 12707 6814 12745 6823
rect 12889 6848 12932 6875
rect 12889 6830 12903 6848
rect 12921 6830 12932 6848
rect 12889 6822 12932 6830
rect 12894 6820 12932 6822
rect 13321 6850 13766 6880
rect 14804 6863 14869 6864
rect 13321 6847 13744 6850
rect 12707 6813 12744 6814
rect 12168 6785 12258 6791
rect 12168 6765 12184 6785
rect 12204 6783 12258 6785
rect 12204 6765 12229 6783
rect 12168 6763 12229 6765
rect 12249 6763 12258 6783
rect 12168 6757 12258 6763
rect 12181 6703 12218 6704
rect 12277 6703 12314 6704
rect 12333 6703 12369 6813
rect 12556 6792 12587 6813
rect 13321 6799 13368 6847
rect 12552 6791 12587 6792
rect 12430 6781 12587 6791
rect 12430 6761 12447 6781
rect 12467 6761 12587 6781
rect 12430 6754 12587 6761
rect 12654 6784 12803 6792
rect 12654 6764 12665 6784
rect 12685 6764 12724 6784
rect 12744 6764 12803 6784
rect 13321 6781 13331 6799
rect 13349 6781 13368 6799
rect 13321 6777 13368 6781
rect 14455 6838 14642 6862
rect 14673 6843 15066 6863
rect 15086 6843 15089 6863
rect 14673 6838 15089 6843
rect 13322 6772 13359 6777
rect 12654 6757 12803 6764
rect 14455 6767 14492 6838
rect 14673 6837 15014 6838
rect 14607 6777 14638 6778
rect 12654 6756 12695 6757
rect 12891 6755 12928 6758
rect 12388 6703 12425 6704
rect 12081 6694 12219 6703
rect 11285 6655 11729 6681
rect 11285 6653 11453 6655
rect 11285 6475 11312 6653
rect 11352 6615 11416 6627
rect 11692 6623 11729 6655
rect 11755 6654 11946 6676
rect 12081 6674 12190 6694
rect 12210 6674 12219 6694
rect 12081 6667 12219 6674
rect 12277 6694 12425 6703
rect 12277 6674 12286 6694
rect 12306 6674 12396 6694
rect 12416 6674 12425 6694
rect 12081 6665 12177 6667
rect 12277 6664 12425 6674
rect 12484 6694 12521 6704
rect 12484 6674 12492 6694
rect 12512 6674 12521 6694
rect 12333 6663 12369 6664
rect 11910 6652 11946 6654
rect 11910 6623 11947 6652
rect 11352 6614 11387 6615
rect 11329 6609 11387 6614
rect 11329 6589 11332 6609
rect 11352 6595 11387 6609
rect 11407 6595 11416 6615
rect 11352 6589 11416 6595
rect 11329 6587 11416 6589
rect 11329 6583 11356 6587
rect 11378 6586 11416 6587
rect 11379 6585 11416 6586
rect 11482 6619 11518 6620
rect 11590 6619 11626 6620
rect 11482 6612 11626 6619
rect 11482 6611 11544 6612
rect 11482 6591 11490 6611
rect 11510 6594 11544 6611
rect 11563 6611 11626 6612
rect 11563 6594 11598 6611
rect 11510 6591 11598 6594
rect 11618 6591 11626 6611
rect 11482 6585 11626 6591
rect 11692 6615 11730 6623
rect 11808 6619 11844 6620
rect 11692 6595 11701 6615
rect 11721 6595 11730 6615
rect 11692 6586 11730 6595
rect 11759 6611 11844 6619
rect 11759 6591 11816 6611
rect 11836 6591 11844 6611
rect 11692 6585 11729 6586
rect 11759 6585 11844 6591
rect 11910 6615 11948 6623
rect 11910 6595 11919 6615
rect 11939 6595 11948 6615
rect 12181 6604 12218 6605
rect 12484 6604 12521 6674
rect 12556 6703 12587 6754
rect 12883 6749 12928 6755
rect 12883 6731 12901 6749
rect 12919 6731 12928 6749
rect 14455 6747 14464 6767
rect 14484 6747 14492 6767
rect 14455 6737 14492 6747
rect 14551 6767 14638 6777
rect 14551 6747 14560 6767
rect 14580 6747 14638 6767
rect 14551 6738 14638 6747
rect 14551 6737 14588 6738
rect 12883 6721 12928 6731
rect 12606 6703 12643 6704
rect 12556 6694 12643 6703
rect 12556 6674 12614 6694
rect 12634 6674 12643 6694
rect 12556 6664 12643 6674
rect 12702 6694 12739 6704
rect 12702 6674 12710 6694
rect 12730 6674 12739 6694
rect 12883 6679 12926 6721
rect 13310 6710 13362 6712
rect 12789 6677 12926 6679
rect 12556 6663 12587 6664
rect 12702 6604 12739 6674
rect 12180 6603 12521 6604
rect 11910 6586 11948 6595
rect 12105 6598 12521 6603
rect 11910 6585 11947 6586
rect 11371 6557 11461 6563
rect 11371 6537 11387 6557
rect 11407 6555 11461 6557
rect 11407 6537 11432 6555
rect 11371 6535 11432 6537
rect 11452 6535 11461 6555
rect 11371 6529 11461 6535
rect 11384 6475 11421 6476
rect 11480 6475 11517 6476
rect 11536 6475 11572 6585
rect 11759 6564 11790 6585
rect 12105 6578 12108 6598
rect 12128 6578 12521 6598
rect 12705 6588 12739 6604
rect 12783 6656 12926 6677
rect 13308 6706 13741 6710
rect 13308 6700 13747 6706
rect 13308 6682 13329 6700
rect 13347 6682 13747 6700
rect 14607 6687 14638 6738
rect 14673 6767 14710 6837
rect 14976 6836 15013 6837
rect 14825 6777 14861 6778
rect 14673 6747 14682 6767
rect 14702 6747 14710 6767
rect 14673 6737 14710 6747
rect 14769 6767 14917 6777
rect 15017 6774 15113 6776
rect 14769 6747 14778 6767
rect 14798 6747 14888 6767
rect 14908 6747 14917 6767
rect 14769 6738 14917 6747
rect 14975 6767 15113 6774
rect 14975 6747 14984 6767
rect 15004 6747 15113 6767
rect 14975 6738 15113 6747
rect 14769 6737 14806 6738
rect 14499 6684 14540 6685
rect 13308 6664 13747 6682
rect 12481 6569 12521 6578
rect 12783 6569 12810 6656
rect 12883 6630 12926 6656
rect 12883 6612 12896 6630
rect 12914 6612 12926 6630
rect 12883 6601 12926 6612
rect 11755 6563 11790 6564
rect 11633 6553 11790 6563
rect 11633 6533 11650 6553
rect 11670 6533 11790 6553
rect 11633 6526 11790 6533
rect 11857 6556 12003 6564
rect 11857 6536 11868 6556
rect 11888 6536 11927 6556
rect 11947 6536 12003 6556
rect 12481 6552 12810 6569
rect 12481 6551 12521 6552
rect 11857 6529 12003 6536
rect 12878 6540 12918 6543
rect 12878 6534 12921 6540
rect 12503 6531 12921 6534
rect 11857 6528 11898 6529
rect 11591 6475 11628 6476
rect 11284 6466 11422 6475
rect 11284 6446 11393 6466
rect 11413 6446 11422 6466
rect 11284 6439 11422 6446
rect 11480 6466 11628 6475
rect 11480 6446 11489 6466
rect 11509 6446 11599 6466
rect 11619 6446 11628 6466
rect 11284 6437 11380 6439
rect 11480 6436 11628 6446
rect 11687 6466 11724 6476
rect 11687 6446 11695 6466
rect 11715 6446 11724 6466
rect 11536 6435 11572 6436
rect 11384 6376 11421 6377
rect 11687 6376 11724 6446
rect 11759 6475 11790 6526
rect 12503 6513 12894 6531
rect 12912 6513 12921 6531
rect 12503 6511 12921 6513
rect 12503 6503 12530 6511
rect 12771 6508 12921 6511
rect 12083 6497 12251 6498
rect 12502 6497 12530 6503
rect 12083 6481 12530 6497
rect 12878 6503 12921 6508
rect 11809 6475 11846 6476
rect 11759 6466 11846 6475
rect 11759 6446 11817 6466
rect 11837 6446 11846 6466
rect 11759 6436 11846 6446
rect 11905 6466 11942 6476
rect 11905 6446 11913 6466
rect 11933 6446 11942 6466
rect 11759 6435 11790 6436
rect 11383 6375 11724 6376
rect 11905 6375 11942 6446
rect 11308 6370 11724 6375
rect 11308 6350 11311 6370
rect 11331 6350 11724 6370
rect 11755 6351 11942 6375
rect 12083 6471 12527 6481
rect 12083 6469 12251 6471
rect 11183 6271 11225 6316
rect 12083 6291 12110 6469
rect 12150 6431 12214 6443
rect 12490 6439 12527 6471
rect 12553 6470 12744 6492
rect 12708 6468 12744 6470
rect 12708 6439 12745 6468
rect 12878 6447 12918 6503
rect 12150 6430 12185 6431
rect 12127 6425 12185 6430
rect 12127 6405 12130 6425
rect 12150 6411 12185 6425
rect 12205 6411 12214 6431
rect 12150 6403 12214 6411
rect 12176 6402 12214 6403
rect 12177 6401 12214 6402
rect 12280 6435 12316 6436
rect 12388 6435 12424 6436
rect 12280 6427 12424 6435
rect 12280 6407 12288 6427
rect 12308 6407 12343 6427
rect 12363 6407 12396 6427
rect 12416 6407 12424 6427
rect 12280 6401 12424 6407
rect 12490 6431 12528 6439
rect 12606 6435 12642 6436
rect 12490 6411 12499 6431
rect 12519 6411 12528 6431
rect 12490 6402 12528 6411
rect 12557 6427 12642 6435
rect 12557 6407 12614 6427
rect 12634 6407 12642 6427
rect 12490 6401 12527 6402
rect 12557 6401 12642 6407
rect 12708 6431 12746 6439
rect 12708 6411 12717 6431
rect 12737 6411 12746 6431
rect 12878 6429 12890 6447
rect 12908 6429 12918 6447
rect 13310 6475 13362 6664
rect 13708 6639 13747 6664
rect 14391 6677 14540 6684
rect 14391 6657 14450 6677
rect 14470 6657 14509 6677
rect 14529 6657 14540 6677
rect 14391 6649 14540 6657
rect 14607 6680 14764 6687
rect 14607 6660 14727 6680
rect 14747 6660 14764 6680
rect 14607 6650 14764 6660
rect 14607 6649 14642 6650
rect 13492 6614 13679 6638
rect 13708 6619 14103 6639
rect 14123 6619 14126 6639
rect 14607 6628 14638 6649
rect 14825 6628 14861 6738
rect 14880 6737 14917 6738
rect 14976 6737 15013 6738
rect 14936 6678 15026 6684
rect 14936 6658 14945 6678
rect 14965 6676 15026 6678
rect 14965 6658 14990 6676
rect 14936 6656 14990 6658
rect 15010 6656 15026 6676
rect 14936 6650 15026 6656
rect 14450 6627 14487 6628
rect 13708 6614 14126 6619
rect 14449 6618 14487 6627
rect 13492 6543 13529 6614
rect 13708 6613 14051 6614
rect 13708 6610 13747 6613
rect 14013 6612 14050 6613
rect 13644 6553 13675 6554
rect 13492 6523 13501 6543
rect 13521 6523 13529 6543
rect 13492 6513 13529 6523
rect 13588 6543 13675 6553
rect 13588 6523 13597 6543
rect 13617 6523 13675 6543
rect 13588 6514 13675 6523
rect 13588 6513 13625 6514
rect 13310 6457 13326 6475
rect 13344 6457 13362 6475
rect 13644 6463 13675 6514
rect 13710 6543 13747 6610
rect 14449 6598 14458 6618
rect 14478 6598 14487 6618
rect 14449 6590 14487 6598
rect 14553 6622 14638 6628
rect 14668 6627 14705 6628
rect 14553 6602 14561 6622
rect 14581 6602 14638 6622
rect 14553 6594 14638 6602
rect 14667 6618 14705 6627
rect 14667 6598 14676 6618
rect 14696 6598 14705 6618
rect 14553 6593 14589 6594
rect 14667 6590 14705 6598
rect 14771 6622 14915 6628
rect 14771 6602 14779 6622
rect 14799 6621 14887 6622
rect 14799 6603 14834 6621
rect 14852 6603 14887 6621
rect 14799 6602 14887 6603
rect 14907 6602 14915 6622
rect 14771 6594 14915 6602
rect 14771 6593 14807 6594
rect 14879 6593 14915 6594
rect 14981 6627 15018 6628
rect 14981 6626 15019 6627
rect 14981 6618 15045 6626
rect 14981 6598 14990 6618
rect 15010 6604 15045 6618
rect 15065 6604 15068 6624
rect 15010 6599 15068 6604
rect 15010 6598 15045 6599
rect 14450 6561 14487 6590
rect 14451 6559 14487 6561
rect 13862 6553 13898 6554
rect 13710 6523 13719 6543
rect 13739 6523 13747 6543
rect 13710 6513 13747 6523
rect 13806 6543 13954 6553
rect 14054 6550 14150 6552
rect 13806 6523 13815 6543
rect 13835 6523 13925 6543
rect 13945 6523 13954 6543
rect 13806 6514 13954 6523
rect 14012 6543 14150 6550
rect 14012 6523 14021 6543
rect 14041 6523 14150 6543
rect 14451 6537 14642 6559
rect 14668 6558 14705 6590
rect 14981 6586 15045 6598
rect 15085 6562 15112 6738
rect 15031 6560 15112 6562
rect 14944 6558 15112 6560
rect 14668 6532 15112 6558
rect 14778 6530 14818 6532
rect 14944 6531 15112 6532
rect 14012 6514 14150 6523
rect 15053 6529 15112 6531
rect 13806 6513 13843 6514
rect 13536 6460 13577 6461
rect 13310 6439 13362 6457
rect 13428 6453 13577 6460
rect 12878 6419 12918 6429
rect 13428 6433 13487 6453
rect 13507 6433 13546 6453
rect 13566 6433 13577 6453
rect 13428 6425 13577 6433
rect 13644 6456 13801 6463
rect 13644 6436 13764 6456
rect 13784 6436 13801 6456
rect 13644 6426 13801 6436
rect 13644 6425 13679 6426
rect 12708 6402 12746 6411
rect 13644 6404 13675 6425
rect 13862 6404 13898 6514
rect 13917 6513 13954 6514
rect 14013 6513 14050 6514
rect 13973 6454 14063 6460
rect 13973 6434 13982 6454
rect 14002 6452 14063 6454
rect 14002 6434 14027 6452
rect 13973 6432 14027 6434
rect 14047 6432 14063 6452
rect 13973 6426 14063 6432
rect 13487 6403 13524 6404
rect 12708 6401 12745 6402
rect 12169 6373 12259 6379
rect 12169 6353 12185 6373
rect 12205 6371 12259 6373
rect 12205 6353 12230 6371
rect 12169 6351 12230 6353
rect 12250 6351 12259 6371
rect 12169 6345 12259 6351
rect 12182 6291 12219 6292
rect 12278 6291 12315 6292
rect 12334 6291 12370 6401
rect 12557 6380 12588 6401
rect 13486 6394 13524 6403
rect 12553 6379 12588 6380
rect 12431 6369 12588 6379
rect 12431 6349 12448 6369
rect 12468 6349 12588 6369
rect 12431 6342 12588 6349
rect 12655 6372 12804 6380
rect 12655 6352 12666 6372
rect 12686 6352 12725 6372
rect 12745 6352 12804 6372
rect 13314 6376 13354 6386
rect 12655 6345 12804 6352
rect 12870 6348 12922 6366
rect 12655 6344 12696 6345
rect 12389 6291 12426 6292
rect 12082 6282 12220 6291
rect 11554 6271 11587 6273
rect 11183 6259 11630 6271
rect 11186 6245 11630 6259
rect 11186 6243 11354 6245
rect 11186 6065 11213 6243
rect 11253 6205 11317 6217
rect 11593 6213 11630 6245
rect 11656 6244 11847 6266
rect 12082 6262 12191 6282
rect 12211 6262 12220 6282
rect 12082 6255 12220 6262
rect 12278 6282 12426 6291
rect 12278 6262 12287 6282
rect 12307 6262 12397 6282
rect 12417 6262 12426 6282
rect 12082 6253 12178 6255
rect 12278 6252 12426 6262
rect 12485 6282 12522 6292
rect 12485 6262 12493 6282
rect 12513 6262 12522 6282
rect 12334 6251 12370 6252
rect 11811 6242 11847 6244
rect 11811 6213 11848 6242
rect 11253 6204 11288 6205
rect 11230 6199 11288 6204
rect 11230 6179 11233 6199
rect 11253 6185 11288 6199
rect 11308 6185 11317 6205
rect 11253 6177 11317 6185
rect 11279 6176 11317 6177
rect 11280 6175 11317 6176
rect 11383 6209 11419 6210
rect 11491 6209 11527 6210
rect 11383 6201 11527 6209
rect 11383 6181 11391 6201
rect 11411 6199 11499 6201
rect 11411 6181 11444 6199
rect 11383 6180 11444 6181
rect 11465 6181 11499 6199
rect 11519 6181 11527 6201
rect 11465 6180 11527 6181
rect 11383 6175 11527 6180
rect 11593 6205 11631 6213
rect 11709 6209 11745 6210
rect 11593 6185 11602 6205
rect 11622 6185 11631 6205
rect 11593 6176 11631 6185
rect 11660 6201 11745 6209
rect 11660 6181 11717 6201
rect 11737 6181 11745 6201
rect 11593 6175 11630 6176
rect 11660 6175 11745 6181
rect 11811 6205 11849 6213
rect 11811 6185 11820 6205
rect 11840 6185 11849 6205
rect 12485 6195 12522 6262
rect 12557 6291 12588 6342
rect 12870 6330 12888 6348
rect 12906 6330 12922 6348
rect 12607 6291 12644 6292
rect 12557 6282 12644 6291
rect 12557 6262 12615 6282
rect 12635 6262 12644 6282
rect 12557 6252 12644 6262
rect 12703 6282 12740 6292
rect 12703 6262 12711 6282
rect 12731 6262 12740 6282
rect 12557 6251 12588 6252
rect 12182 6192 12219 6193
rect 12485 6192 12524 6195
rect 12181 6191 12524 6192
rect 12703 6191 12740 6262
rect 11811 6176 11849 6185
rect 12106 6186 12524 6191
rect 11811 6175 11848 6176
rect 11272 6147 11362 6153
rect 11272 6127 11288 6147
rect 11308 6145 11362 6147
rect 11308 6127 11333 6145
rect 11272 6125 11333 6127
rect 11353 6125 11362 6145
rect 11272 6119 11362 6125
rect 11285 6065 11322 6066
rect 11381 6065 11418 6066
rect 11437 6065 11473 6175
rect 11660 6154 11691 6175
rect 12106 6166 12109 6186
rect 12129 6166 12524 6186
rect 12553 6167 12740 6191
rect 11656 6153 11691 6154
rect 11534 6143 11691 6153
rect 11534 6123 11551 6143
rect 11571 6123 11691 6143
rect 11534 6116 11691 6123
rect 11758 6146 11907 6154
rect 11758 6126 11769 6146
rect 11789 6126 11828 6146
rect 11848 6126 11907 6146
rect 11758 6119 11907 6126
rect 12485 6141 12524 6166
rect 12870 6141 12922 6330
rect 13314 6358 13324 6376
rect 13342 6358 13354 6376
rect 13486 6374 13495 6394
rect 13515 6374 13524 6394
rect 13486 6366 13524 6374
rect 13590 6398 13675 6404
rect 13705 6403 13742 6404
rect 13590 6378 13598 6398
rect 13618 6378 13675 6398
rect 13590 6370 13675 6378
rect 13704 6394 13742 6403
rect 13704 6374 13713 6394
rect 13733 6374 13742 6394
rect 13590 6369 13626 6370
rect 13704 6366 13742 6374
rect 13808 6398 13952 6404
rect 13808 6378 13816 6398
rect 13836 6378 13869 6398
rect 13889 6378 13924 6398
rect 13944 6378 13952 6398
rect 13808 6370 13952 6378
rect 13808 6369 13844 6370
rect 13916 6369 13952 6370
rect 14018 6403 14055 6404
rect 14018 6402 14056 6403
rect 14018 6394 14082 6402
rect 14018 6374 14027 6394
rect 14047 6380 14082 6394
rect 14102 6380 14105 6400
rect 14047 6375 14105 6380
rect 14047 6374 14082 6375
rect 13314 6302 13354 6358
rect 13487 6337 13524 6366
rect 13488 6335 13524 6337
rect 13488 6313 13679 6335
rect 13705 6334 13742 6366
rect 14018 6362 14082 6374
rect 14122 6336 14149 6514
rect 15053 6511 15082 6529
rect 13981 6334 14149 6336
rect 13705 6324 14149 6334
rect 14290 6430 14477 6454
rect 14508 6435 14901 6455
rect 14921 6435 14924 6455
rect 14508 6430 14924 6435
rect 14290 6359 14327 6430
rect 14508 6429 14849 6430
rect 14442 6369 14473 6370
rect 14290 6339 14299 6359
rect 14319 6339 14327 6359
rect 14290 6329 14327 6339
rect 14386 6359 14473 6369
rect 14386 6339 14395 6359
rect 14415 6339 14473 6359
rect 14386 6330 14473 6339
rect 14386 6329 14423 6330
rect 13311 6297 13354 6302
rect 13702 6308 14149 6324
rect 13702 6302 13730 6308
rect 13981 6307 14149 6308
rect 13311 6294 13461 6297
rect 13702 6294 13729 6302
rect 13311 6292 13729 6294
rect 13311 6274 13320 6292
rect 13338 6274 13729 6292
rect 14442 6279 14473 6330
rect 14508 6359 14545 6429
rect 14811 6428 14848 6429
rect 14660 6369 14696 6370
rect 14508 6339 14517 6359
rect 14537 6339 14545 6359
rect 14508 6329 14545 6339
rect 14604 6359 14752 6369
rect 14852 6366 14948 6368
rect 14604 6339 14613 6359
rect 14633 6339 14723 6359
rect 14743 6339 14752 6359
rect 14604 6330 14752 6339
rect 14810 6359 14948 6366
rect 14810 6339 14819 6359
rect 14839 6339 14948 6359
rect 14810 6330 14948 6339
rect 14604 6329 14641 6330
rect 14334 6276 14375 6277
rect 13311 6271 13729 6274
rect 13311 6265 13354 6271
rect 13314 6262 13354 6265
rect 14226 6269 14375 6276
rect 13711 6253 13751 6254
rect 13422 6236 13751 6253
rect 14226 6249 14285 6269
rect 14305 6249 14344 6269
rect 14364 6249 14375 6269
rect 14226 6241 14375 6249
rect 14442 6272 14599 6279
rect 14442 6252 14562 6272
rect 14582 6252 14599 6272
rect 14442 6242 14599 6252
rect 14442 6241 14477 6242
rect 13306 6193 13349 6204
rect 13306 6175 13318 6193
rect 13336 6175 13349 6193
rect 13306 6149 13349 6175
rect 13422 6149 13449 6236
rect 13711 6227 13751 6236
rect 12485 6123 12924 6141
rect 11758 6118 11799 6119
rect 11492 6065 11529 6066
rect 11185 6056 11323 6065
rect 11185 6036 11294 6056
rect 11314 6036 11323 6056
rect 11185 6029 11323 6036
rect 11381 6056 11529 6065
rect 11381 6036 11390 6056
rect 11410 6036 11500 6056
rect 11520 6036 11529 6056
rect 11185 6027 11281 6029
rect 11381 6026 11529 6036
rect 11588 6056 11625 6066
rect 11588 6036 11596 6056
rect 11616 6036 11625 6056
rect 11437 6025 11473 6026
rect 11285 5966 11322 5967
rect 11588 5966 11625 6036
rect 11660 6065 11691 6116
rect 12485 6105 12885 6123
rect 12903 6105 12924 6123
rect 12485 6099 12924 6105
rect 12491 6095 12924 6099
rect 13306 6128 13449 6149
rect 13493 6201 13527 6217
rect 13711 6207 14104 6227
rect 14124 6207 14127 6227
rect 14442 6220 14473 6241
rect 14660 6220 14696 6330
rect 14715 6329 14752 6330
rect 14811 6329 14848 6330
rect 14771 6270 14861 6276
rect 14771 6250 14780 6270
rect 14800 6268 14861 6270
rect 14800 6250 14825 6268
rect 14771 6248 14825 6250
rect 14845 6248 14861 6268
rect 14771 6242 14861 6248
rect 14285 6219 14322 6220
rect 13711 6202 14127 6207
rect 14284 6210 14322 6219
rect 13711 6201 14052 6202
rect 13493 6131 13530 6201
rect 13645 6141 13676 6142
rect 13306 6126 13443 6128
rect 12870 6093 12922 6095
rect 13306 6084 13349 6126
rect 13493 6111 13502 6131
rect 13522 6111 13530 6131
rect 13493 6101 13530 6111
rect 13589 6131 13676 6141
rect 13589 6111 13598 6131
rect 13618 6111 13676 6131
rect 13589 6102 13676 6111
rect 13589 6101 13626 6102
rect 13304 6074 13349 6084
rect 11710 6065 11747 6066
rect 11660 6056 11747 6065
rect 11660 6036 11718 6056
rect 11738 6036 11747 6056
rect 11660 6026 11747 6036
rect 11806 6056 11843 6066
rect 11806 6036 11814 6056
rect 11834 6036 11843 6056
rect 13304 6056 13313 6074
rect 13331 6056 13349 6074
rect 13304 6050 13349 6056
rect 13645 6051 13676 6102
rect 13711 6131 13748 6201
rect 14014 6200 14051 6201
rect 14284 6190 14293 6210
rect 14313 6190 14322 6210
rect 14284 6182 14322 6190
rect 14388 6214 14473 6220
rect 14503 6219 14540 6220
rect 14388 6194 14396 6214
rect 14416 6194 14473 6214
rect 14388 6186 14473 6194
rect 14502 6210 14540 6219
rect 14502 6190 14511 6210
rect 14531 6190 14540 6210
rect 14388 6185 14424 6186
rect 14502 6182 14540 6190
rect 14606 6214 14750 6220
rect 14606 6194 14614 6214
rect 14634 6195 14666 6214
rect 14687 6195 14722 6214
rect 14634 6194 14722 6195
rect 14742 6194 14750 6214
rect 14606 6186 14750 6194
rect 14606 6185 14642 6186
rect 14714 6185 14750 6186
rect 14816 6219 14853 6220
rect 14816 6218 14854 6219
rect 14816 6210 14880 6218
rect 14816 6190 14825 6210
rect 14845 6196 14880 6210
rect 14900 6196 14903 6216
rect 14845 6191 14903 6196
rect 14845 6190 14880 6191
rect 14285 6153 14322 6182
rect 14286 6151 14322 6153
rect 13863 6141 13899 6142
rect 13711 6111 13720 6131
rect 13740 6111 13748 6131
rect 13711 6101 13748 6111
rect 13807 6131 13955 6141
rect 14055 6138 14151 6140
rect 13807 6111 13816 6131
rect 13836 6111 13926 6131
rect 13946 6111 13955 6131
rect 13807 6102 13955 6111
rect 14013 6131 14151 6138
rect 14013 6111 14022 6131
rect 14042 6111 14151 6131
rect 14286 6129 14477 6151
rect 14503 6150 14540 6182
rect 14816 6178 14880 6190
rect 14920 6152 14947 6330
rect 14779 6150 14947 6152
rect 14503 6124 14947 6150
rect 14013 6102 14151 6111
rect 13807 6101 13844 6102
rect 13304 6047 13341 6050
rect 13537 6048 13578 6049
rect 11660 6025 11691 6026
rect 11284 5965 11625 5966
rect 11806 5965 11843 6036
rect 13429 6041 13578 6048
rect 12873 6028 12910 6033
rect 12864 6024 12911 6028
rect 12864 6006 12883 6024
rect 12901 6006 12911 6024
rect 13429 6021 13488 6041
rect 13508 6021 13547 6041
rect 13567 6021 13578 6041
rect 13429 6013 13578 6021
rect 13645 6044 13802 6051
rect 13645 6024 13765 6044
rect 13785 6024 13802 6044
rect 13645 6014 13802 6024
rect 13645 6013 13680 6014
rect 11209 5960 11625 5965
rect 11209 5940 11212 5960
rect 11232 5940 11625 5960
rect 11656 5941 11843 5965
rect 12468 5963 12508 5968
rect 12864 5963 12911 6006
rect 13645 5992 13676 6013
rect 13863 5992 13899 6102
rect 13918 6101 13955 6102
rect 14014 6101 14051 6102
rect 13974 6042 14064 6048
rect 13974 6022 13983 6042
rect 14003 6040 14064 6042
rect 14003 6022 14028 6040
rect 13974 6020 14028 6022
rect 14048 6020 14064 6040
rect 13974 6014 14064 6020
rect 13488 5991 13525 5992
rect 12468 5924 12911 5963
rect 13301 5983 13338 5985
rect 13301 5975 13343 5983
rect 13301 5957 13311 5975
rect 13329 5957 13343 5975
rect 13301 5948 13343 5957
rect 13487 5982 13525 5991
rect 13487 5962 13496 5982
rect 13516 5962 13525 5982
rect 13487 5954 13525 5962
rect 13591 5986 13676 5992
rect 13706 5991 13743 5992
rect 13591 5966 13599 5986
rect 13619 5966 13676 5986
rect 13591 5958 13676 5966
rect 13705 5982 13743 5991
rect 13705 5962 13714 5982
rect 13734 5962 13743 5982
rect 13591 5957 13627 5958
rect 13705 5954 13743 5962
rect 13809 5990 13953 5992
rect 13809 5986 13861 5990
rect 13809 5966 13817 5986
rect 13837 5970 13861 5986
rect 13881 5986 13953 5990
rect 13881 5970 13925 5986
rect 13837 5966 13925 5970
rect 13945 5966 13953 5986
rect 13809 5958 13953 5966
rect 13809 5957 13845 5958
rect 13917 5957 13953 5958
rect 14019 5991 14056 5992
rect 14019 5990 14057 5991
rect 14019 5982 14083 5990
rect 14019 5962 14028 5982
rect 14048 5968 14083 5982
rect 14103 5968 14106 5988
rect 14048 5963 14106 5968
rect 14048 5962 14083 5963
rect 11562 5909 11602 5917
rect 11562 5887 11570 5909
rect 11594 5887 11602 5909
rect 11268 5663 11436 5664
rect 11562 5663 11602 5887
rect 12065 5891 12233 5892
rect 12468 5891 12508 5924
rect 12864 5891 12911 5924
rect 13302 5923 13343 5948
rect 13488 5923 13525 5954
rect 13706 5923 13743 5954
rect 14019 5950 14083 5962
rect 14123 5924 14150 6102
rect 13302 5896 13351 5923
rect 13487 5897 13536 5923
rect 13705 5922 13786 5923
rect 13982 5922 14150 5924
rect 13705 5897 14150 5922
rect 13706 5896 14150 5897
rect 12065 5890 12509 5891
rect 12065 5865 12510 5890
rect 12065 5863 12233 5865
rect 12429 5864 12510 5865
rect 12679 5864 12728 5890
rect 12864 5864 12913 5891
rect 12065 5685 12092 5863
rect 12132 5825 12196 5837
rect 12472 5833 12509 5864
rect 12690 5833 12727 5864
rect 12872 5839 12913 5864
rect 13304 5863 13351 5896
rect 13707 5863 13747 5896
rect 13982 5895 14150 5896
rect 14613 5900 14653 6124
rect 14779 6123 14947 6124
rect 14613 5878 14621 5900
rect 14645 5878 14653 5900
rect 14613 5870 14653 5878
rect 12132 5824 12167 5825
rect 12109 5819 12167 5824
rect 12109 5799 12112 5819
rect 12132 5805 12167 5819
rect 12187 5805 12196 5825
rect 12132 5797 12196 5805
rect 12158 5796 12196 5797
rect 12159 5795 12196 5796
rect 12262 5829 12298 5830
rect 12370 5829 12406 5830
rect 12262 5821 12406 5829
rect 12262 5801 12270 5821
rect 12290 5817 12378 5821
rect 12290 5801 12334 5817
rect 12262 5797 12334 5801
rect 12354 5801 12378 5817
rect 12398 5801 12406 5821
rect 12354 5797 12406 5801
rect 12262 5795 12406 5797
rect 12472 5825 12510 5833
rect 12588 5829 12624 5830
rect 12472 5805 12481 5825
rect 12501 5805 12510 5825
rect 12472 5796 12510 5805
rect 12539 5821 12624 5829
rect 12539 5801 12596 5821
rect 12616 5801 12624 5821
rect 12472 5795 12509 5796
rect 12539 5795 12624 5801
rect 12690 5825 12728 5833
rect 12690 5805 12699 5825
rect 12719 5805 12728 5825
rect 12690 5796 12728 5805
rect 12872 5830 12914 5839
rect 12872 5812 12886 5830
rect 12904 5812 12914 5830
rect 12872 5804 12914 5812
rect 12877 5802 12914 5804
rect 13304 5824 13747 5863
rect 12690 5795 12727 5796
rect 12151 5767 12241 5773
rect 12151 5747 12167 5767
rect 12187 5765 12241 5767
rect 12187 5747 12212 5765
rect 12151 5745 12212 5747
rect 12232 5745 12241 5765
rect 12151 5739 12241 5745
rect 12164 5685 12201 5686
rect 12260 5685 12297 5686
rect 12316 5685 12352 5795
rect 12539 5774 12570 5795
rect 13304 5781 13351 5824
rect 13707 5819 13747 5824
rect 14372 5822 14559 5846
rect 14590 5827 14983 5847
rect 15003 5827 15006 5847
rect 14590 5822 15006 5827
rect 12535 5773 12570 5774
rect 12413 5763 12570 5773
rect 12413 5743 12430 5763
rect 12450 5743 12570 5763
rect 12413 5736 12570 5743
rect 12637 5766 12786 5774
rect 12637 5746 12648 5766
rect 12668 5746 12707 5766
rect 12727 5746 12786 5766
rect 13304 5763 13314 5781
rect 13332 5763 13351 5781
rect 13304 5759 13351 5763
rect 13305 5754 13342 5759
rect 12637 5739 12786 5746
rect 14372 5751 14409 5822
rect 14590 5821 14931 5822
rect 14524 5761 14555 5762
rect 12637 5738 12678 5739
rect 12874 5737 12911 5740
rect 12371 5685 12408 5686
rect 12064 5676 12202 5685
rect 11268 5637 11712 5663
rect 11268 5635 11436 5637
rect 11268 5457 11295 5635
rect 11335 5597 11399 5609
rect 11675 5605 11712 5637
rect 11738 5636 11929 5658
rect 12064 5656 12173 5676
rect 12193 5656 12202 5676
rect 12064 5649 12202 5656
rect 12260 5676 12408 5685
rect 12260 5656 12269 5676
rect 12289 5656 12379 5676
rect 12399 5656 12408 5676
rect 12064 5647 12160 5649
rect 12260 5646 12408 5656
rect 12467 5676 12504 5686
rect 12467 5656 12475 5676
rect 12495 5656 12504 5676
rect 12316 5645 12352 5646
rect 11893 5634 11929 5636
rect 11893 5605 11930 5634
rect 11335 5596 11370 5597
rect 11312 5591 11370 5596
rect 11312 5571 11315 5591
rect 11335 5577 11370 5591
rect 11390 5577 11399 5597
rect 11335 5569 11399 5577
rect 11361 5568 11399 5569
rect 11362 5567 11399 5568
rect 11465 5601 11501 5602
rect 11573 5601 11609 5602
rect 11465 5593 11609 5601
rect 11465 5573 11473 5593
rect 11493 5592 11581 5593
rect 11493 5573 11528 5592
rect 11549 5573 11581 5592
rect 11601 5573 11609 5593
rect 11465 5567 11609 5573
rect 11675 5597 11713 5605
rect 11791 5601 11827 5602
rect 11675 5577 11684 5597
rect 11704 5577 11713 5597
rect 11675 5568 11713 5577
rect 11742 5593 11827 5601
rect 11742 5573 11799 5593
rect 11819 5573 11827 5593
rect 11675 5567 11712 5568
rect 11742 5567 11827 5573
rect 11893 5597 11931 5605
rect 11893 5577 11902 5597
rect 11922 5577 11931 5597
rect 12164 5586 12201 5587
rect 12467 5586 12504 5656
rect 12539 5685 12570 5736
rect 12866 5731 12911 5737
rect 12866 5713 12884 5731
rect 12902 5713 12911 5731
rect 14372 5731 14381 5751
rect 14401 5731 14409 5751
rect 14372 5721 14409 5731
rect 14468 5751 14555 5761
rect 14468 5731 14477 5751
rect 14497 5731 14555 5751
rect 14468 5722 14555 5731
rect 14468 5721 14505 5722
rect 12866 5703 12911 5713
rect 12589 5685 12626 5686
rect 12539 5676 12626 5685
rect 12539 5656 12597 5676
rect 12617 5656 12626 5676
rect 12539 5646 12626 5656
rect 12685 5676 12722 5686
rect 12685 5656 12693 5676
rect 12713 5656 12722 5676
rect 12866 5661 12909 5703
rect 13293 5692 13345 5694
rect 12772 5659 12909 5661
rect 12539 5645 12570 5646
rect 12685 5586 12722 5656
rect 12163 5585 12504 5586
rect 11893 5568 11931 5577
rect 12088 5580 12504 5585
rect 11893 5567 11930 5568
rect 11354 5539 11444 5545
rect 11354 5519 11370 5539
rect 11390 5537 11444 5539
rect 11390 5519 11415 5537
rect 11354 5517 11415 5519
rect 11435 5517 11444 5537
rect 11354 5511 11444 5517
rect 11367 5457 11404 5458
rect 11463 5457 11500 5458
rect 11519 5457 11555 5567
rect 11742 5546 11773 5567
rect 12088 5560 12091 5580
rect 12111 5560 12504 5580
rect 12688 5570 12722 5586
rect 12766 5638 12909 5659
rect 13291 5688 13724 5692
rect 13291 5682 13730 5688
rect 13291 5664 13312 5682
rect 13330 5664 13730 5682
rect 14524 5671 14555 5722
rect 14590 5751 14627 5821
rect 14893 5820 14930 5821
rect 14742 5761 14778 5762
rect 14590 5731 14599 5751
rect 14619 5731 14627 5751
rect 14590 5721 14627 5731
rect 14686 5751 14834 5761
rect 14934 5758 15030 5760
rect 14686 5731 14695 5751
rect 14715 5731 14805 5751
rect 14825 5731 14834 5751
rect 14686 5722 14834 5731
rect 14892 5751 15030 5758
rect 14892 5731 14901 5751
rect 14921 5731 15030 5751
rect 14892 5722 15030 5731
rect 14686 5721 14723 5722
rect 14416 5668 14457 5669
rect 13291 5646 13730 5664
rect 12464 5551 12504 5560
rect 12766 5551 12793 5638
rect 12866 5612 12909 5638
rect 12866 5594 12879 5612
rect 12897 5594 12909 5612
rect 12866 5583 12909 5594
rect 11738 5545 11773 5546
rect 11616 5535 11773 5545
rect 11616 5515 11633 5535
rect 11653 5515 11773 5535
rect 11616 5508 11773 5515
rect 11840 5538 11989 5546
rect 11840 5518 11851 5538
rect 11871 5518 11910 5538
rect 11930 5518 11989 5538
rect 12464 5534 12793 5551
rect 12464 5533 12504 5534
rect 11840 5511 11989 5518
rect 12861 5522 12901 5525
rect 12861 5516 12904 5522
rect 12486 5513 12904 5516
rect 11840 5510 11881 5511
rect 11574 5457 11611 5458
rect 11267 5448 11405 5457
rect 10965 5273 11005 5445
rect 11267 5428 11376 5448
rect 11396 5428 11405 5448
rect 11267 5421 11405 5428
rect 11463 5448 11611 5457
rect 11463 5428 11472 5448
rect 11492 5428 11582 5448
rect 11602 5428 11611 5448
rect 11267 5419 11363 5421
rect 11463 5418 11611 5428
rect 11670 5448 11707 5458
rect 11670 5428 11678 5448
rect 11698 5428 11707 5448
rect 11519 5417 11555 5418
rect 11367 5358 11404 5359
rect 11670 5358 11707 5428
rect 11742 5457 11773 5508
rect 12486 5495 12877 5513
rect 12895 5495 12904 5513
rect 12486 5493 12904 5495
rect 12486 5485 12513 5493
rect 12754 5490 12904 5493
rect 12066 5479 12234 5480
rect 12485 5479 12513 5485
rect 12066 5463 12513 5479
rect 12861 5485 12904 5490
rect 11792 5457 11829 5458
rect 11742 5448 11829 5457
rect 11742 5428 11800 5448
rect 11820 5428 11829 5448
rect 11742 5418 11829 5428
rect 11888 5448 11925 5458
rect 11888 5428 11896 5448
rect 11916 5428 11925 5448
rect 11742 5417 11773 5418
rect 11366 5357 11707 5358
rect 11888 5357 11925 5428
rect 11291 5352 11707 5357
rect 11291 5332 11294 5352
rect 11314 5332 11707 5352
rect 11738 5333 11925 5357
rect 12066 5453 12510 5463
rect 12066 5451 12234 5453
rect 12066 5273 12093 5451
rect 12133 5413 12197 5425
rect 12473 5421 12510 5453
rect 12536 5452 12727 5474
rect 12691 5450 12727 5452
rect 12691 5421 12728 5450
rect 12861 5429 12901 5485
rect 12133 5412 12168 5413
rect 12110 5407 12168 5412
rect 12110 5387 12113 5407
rect 12133 5393 12168 5407
rect 12188 5393 12197 5413
rect 12133 5385 12197 5393
rect 12159 5384 12197 5385
rect 12160 5383 12197 5384
rect 12263 5417 12299 5418
rect 12371 5417 12407 5418
rect 12263 5409 12407 5417
rect 12263 5389 12271 5409
rect 12291 5389 12326 5409
rect 12346 5389 12379 5409
rect 12399 5389 12407 5409
rect 12263 5383 12407 5389
rect 12473 5413 12511 5421
rect 12589 5417 12625 5418
rect 12473 5393 12482 5413
rect 12502 5393 12511 5413
rect 12473 5384 12511 5393
rect 12540 5409 12625 5417
rect 12540 5389 12597 5409
rect 12617 5389 12625 5409
rect 12473 5383 12510 5384
rect 12540 5383 12625 5389
rect 12691 5413 12729 5421
rect 12691 5393 12700 5413
rect 12720 5393 12729 5413
rect 12861 5411 12873 5429
rect 12891 5411 12901 5429
rect 13293 5457 13345 5646
rect 13691 5621 13730 5646
rect 14308 5661 14457 5668
rect 14308 5641 14367 5661
rect 14387 5641 14426 5661
rect 14446 5641 14457 5661
rect 14308 5633 14457 5641
rect 14524 5664 14681 5671
rect 14524 5644 14644 5664
rect 14664 5644 14681 5664
rect 14524 5634 14681 5644
rect 14524 5633 14559 5634
rect 13475 5596 13662 5620
rect 13691 5601 14086 5621
rect 14106 5601 14109 5621
rect 14524 5612 14555 5633
rect 14742 5612 14778 5722
rect 14797 5721 14834 5722
rect 14893 5721 14930 5722
rect 14853 5662 14943 5668
rect 14853 5642 14862 5662
rect 14882 5660 14943 5662
rect 14882 5642 14907 5660
rect 14853 5640 14907 5642
rect 14927 5640 14943 5660
rect 14853 5634 14943 5640
rect 14367 5611 14404 5612
rect 13691 5596 14109 5601
rect 14366 5602 14404 5611
rect 13475 5525 13512 5596
rect 13691 5595 14034 5596
rect 13691 5592 13730 5595
rect 13996 5594 14033 5595
rect 13627 5535 13658 5536
rect 13475 5505 13484 5525
rect 13504 5505 13512 5525
rect 13475 5495 13512 5505
rect 13571 5525 13658 5535
rect 13571 5505 13580 5525
rect 13600 5505 13658 5525
rect 13571 5496 13658 5505
rect 13571 5495 13608 5496
rect 13293 5439 13309 5457
rect 13327 5439 13345 5457
rect 13627 5445 13658 5496
rect 13693 5525 13730 5592
rect 14366 5582 14375 5602
rect 14395 5582 14404 5602
rect 14366 5574 14404 5582
rect 14470 5606 14555 5612
rect 14585 5611 14622 5612
rect 14470 5586 14478 5606
rect 14498 5586 14555 5606
rect 14470 5578 14555 5586
rect 14584 5602 14622 5611
rect 14584 5582 14593 5602
rect 14613 5582 14622 5602
rect 14470 5577 14506 5578
rect 14584 5574 14622 5582
rect 14688 5606 14832 5612
rect 14688 5586 14696 5606
rect 14716 5601 14804 5606
rect 14716 5586 14752 5601
rect 14688 5584 14752 5586
rect 14771 5586 14804 5601
rect 14824 5586 14832 5606
rect 14771 5584 14832 5586
rect 14688 5578 14832 5584
rect 14688 5577 14724 5578
rect 14796 5577 14832 5578
rect 14898 5611 14935 5612
rect 14898 5610 14936 5611
rect 14898 5602 14962 5610
rect 14898 5582 14907 5602
rect 14927 5588 14962 5602
rect 14982 5588 14985 5608
rect 14927 5583 14985 5588
rect 14927 5582 14962 5583
rect 14367 5545 14404 5574
rect 14368 5543 14404 5545
rect 13845 5535 13881 5536
rect 13693 5505 13702 5525
rect 13722 5505 13730 5525
rect 13693 5495 13730 5505
rect 13789 5525 13937 5535
rect 14037 5532 14133 5534
rect 13789 5505 13798 5525
rect 13818 5505 13908 5525
rect 13928 5505 13937 5525
rect 13789 5496 13937 5505
rect 13995 5525 14133 5532
rect 13995 5505 14004 5525
rect 14024 5505 14133 5525
rect 14368 5521 14559 5543
rect 14585 5542 14622 5574
rect 14898 5570 14962 5582
rect 15002 5544 15029 5722
rect 14861 5542 15029 5544
rect 14585 5528 15029 5542
rect 15053 5565 15081 6511
rect 15053 5535 15098 5565
rect 14585 5516 15032 5528
rect 14628 5514 14661 5516
rect 13995 5496 14133 5505
rect 13789 5495 13826 5496
rect 13519 5442 13560 5443
rect 13293 5421 13345 5439
rect 13411 5435 13560 5442
rect 12861 5401 12901 5411
rect 13411 5415 13470 5435
rect 13490 5415 13529 5435
rect 13549 5415 13560 5435
rect 13411 5407 13560 5415
rect 13627 5438 13784 5445
rect 13627 5418 13747 5438
rect 13767 5418 13784 5438
rect 13627 5408 13784 5418
rect 13627 5407 13662 5408
rect 12691 5384 12729 5393
rect 13627 5386 13658 5407
rect 13845 5386 13881 5496
rect 13900 5495 13937 5496
rect 13996 5495 14033 5496
rect 13956 5436 14046 5442
rect 13956 5416 13965 5436
rect 13985 5434 14046 5436
rect 13985 5416 14010 5434
rect 13956 5414 14010 5416
rect 14030 5414 14046 5434
rect 13956 5408 14046 5414
rect 13470 5385 13507 5386
rect 12691 5383 12728 5384
rect 12152 5355 12242 5361
rect 12152 5335 12168 5355
rect 12188 5353 12242 5355
rect 12188 5335 12213 5353
rect 12152 5333 12213 5335
rect 12233 5333 12242 5353
rect 12152 5327 12242 5333
rect 12165 5273 12202 5274
rect 12261 5273 12298 5274
rect 12317 5273 12353 5383
rect 12540 5362 12571 5383
rect 13469 5376 13507 5385
rect 12536 5361 12571 5362
rect 12414 5351 12571 5361
rect 12414 5331 12431 5351
rect 12451 5331 12571 5351
rect 12414 5324 12571 5331
rect 12638 5354 12787 5362
rect 12638 5334 12649 5354
rect 12669 5334 12708 5354
rect 12728 5334 12787 5354
rect 13297 5358 13337 5368
rect 12638 5327 12787 5334
rect 12853 5330 12905 5348
rect 12638 5326 12679 5327
rect 12372 5273 12409 5274
rect 10966 5258 11005 5273
rect 12065 5264 12203 5273
rect 10966 5257 11132 5258
rect 11258 5257 11298 5259
rect 10966 5231 11408 5257
rect 10966 5229 11132 5231
rect 10630 5117 10667 5125
rect 10630 5098 10638 5117
rect 10659 5098 10667 5117
rect 10630 5092 10667 5098
rect 10966 5051 10991 5229
rect 11031 5191 11095 5203
rect 11371 5199 11408 5231
rect 11434 5230 11625 5252
rect 12065 5244 12174 5264
rect 12194 5244 12203 5264
rect 12065 5237 12203 5244
rect 12261 5264 12409 5273
rect 12261 5244 12270 5264
rect 12290 5244 12380 5264
rect 12400 5244 12409 5264
rect 12065 5235 12161 5237
rect 12261 5234 12409 5244
rect 12468 5264 12505 5274
rect 12468 5244 12476 5264
rect 12496 5244 12505 5264
rect 12317 5233 12353 5234
rect 11589 5228 11625 5230
rect 11589 5199 11626 5228
rect 11031 5190 11066 5191
rect 11008 5185 11066 5190
rect 11008 5165 11011 5185
rect 11031 5171 11066 5185
rect 11086 5171 11095 5191
rect 11031 5163 11095 5171
rect 11057 5162 11095 5163
rect 11058 5161 11095 5162
rect 11161 5195 11197 5196
rect 11269 5195 11305 5196
rect 11161 5190 11305 5195
rect 11161 5187 11223 5190
rect 11161 5167 11169 5187
rect 11189 5167 11223 5187
rect 11161 5164 11223 5167
rect 11249 5187 11305 5190
rect 11249 5167 11277 5187
rect 11297 5167 11305 5187
rect 11249 5164 11305 5167
rect 11161 5161 11305 5164
rect 11371 5191 11409 5199
rect 11487 5195 11523 5196
rect 11371 5171 11380 5191
rect 11400 5171 11409 5191
rect 11371 5162 11409 5171
rect 11438 5187 11523 5195
rect 11438 5167 11495 5187
rect 11515 5167 11523 5187
rect 11371 5161 11408 5162
rect 11438 5161 11523 5167
rect 11589 5191 11627 5199
rect 11589 5171 11598 5191
rect 11618 5171 11627 5191
rect 12468 5177 12505 5244
rect 12540 5273 12571 5324
rect 12853 5312 12871 5330
rect 12889 5312 12905 5330
rect 12590 5273 12627 5274
rect 12540 5264 12627 5273
rect 12540 5244 12598 5264
rect 12618 5244 12627 5264
rect 12540 5234 12627 5244
rect 12686 5264 12723 5274
rect 12686 5244 12694 5264
rect 12714 5244 12723 5264
rect 12540 5233 12571 5234
rect 12165 5174 12202 5175
rect 12468 5174 12507 5177
rect 12164 5173 12507 5174
rect 12686 5173 12723 5244
rect 11589 5162 11627 5171
rect 12089 5168 12507 5173
rect 11589 5161 11626 5162
rect 11050 5133 11140 5139
rect 11050 5113 11066 5133
rect 11086 5131 11140 5133
rect 11086 5113 11111 5131
rect 11050 5111 11111 5113
rect 11131 5111 11140 5131
rect 11050 5105 11140 5111
rect 11063 5051 11100 5052
rect 11159 5051 11196 5052
rect 11215 5051 11251 5161
rect 11438 5140 11469 5161
rect 12089 5148 12092 5168
rect 12112 5148 12507 5168
rect 12536 5149 12723 5173
rect 11434 5139 11469 5140
rect 11312 5129 11469 5139
rect 11312 5109 11329 5129
rect 11349 5109 11469 5129
rect 11312 5102 11469 5109
rect 11536 5132 11685 5140
rect 11536 5112 11547 5132
rect 11567 5112 11606 5132
rect 11626 5112 11685 5132
rect 11536 5105 11685 5112
rect 12468 5123 12507 5148
rect 12853 5123 12905 5312
rect 13297 5340 13307 5358
rect 13325 5340 13337 5358
rect 13469 5356 13478 5376
rect 13498 5356 13507 5376
rect 13469 5348 13507 5356
rect 13573 5380 13658 5386
rect 13688 5385 13725 5386
rect 13573 5360 13581 5380
rect 13601 5360 13658 5380
rect 13573 5352 13658 5360
rect 13687 5376 13725 5385
rect 13687 5356 13696 5376
rect 13716 5356 13725 5376
rect 13573 5351 13609 5352
rect 13687 5348 13725 5356
rect 13791 5380 13935 5386
rect 13791 5360 13799 5380
rect 13819 5360 13852 5380
rect 13872 5360 13907 5380
rect 13927 5360 13935 5380
rect 13791 5352 13935 5360
rect 13791 5351 13827 5352
rect 13899 5351 13935 5352
rect 14001 5385 14038 5386
rect 14001 5384 14039 5385
rect 14001 5376 14065 5384
rect 14001 5356 14010 5376
rect 14030 5362 14065 5376
rect 14085 5362 14088 5382
rect 14030 5357 14088 5362
rect 14030 5356 14065 5357
rect 13297 5284 13337 5340
rect 13470 5319 13507 5348
rect 13471 5317 13507 5319
rect 13471 5295 13662 5317
rect 13688 5316 13725 5348
rect 14001 5344 14065 5356
rect 14105 5318 14132 5496
rect 14990 5471 15032 5516
rect 15053 5517 15064 5535
rect 15086 5517 15098 5535
rect 15053 5511 15098 5517
rect 15054 5510 15098 5511
rect 13964 5316 14132 5318
rect 13688 5306 14132 5316
rect 14273 5412 14460 5436
rect 14491 5417 14884 5437
rect 14904 5417 14907 5437
rect 14491 5412 14907 5417
rect 14273 5341 14310 5412
rect 14491 5411 14832 5412
rect 14425 5351 14456 5352
rect 14273 5321 14282 5341
rect 14302 5321 14310 5341
rect 14273 5311 14310 5321
rect 14369 5341 14456 5351
rect 14369 5321 14378 5341
rect 14398 5321 14456 5341
rect 14369 5312 14456 5321
rect 14369 5311 14406 5312
rect 13294 5279 13337 5284
rect 13685 5290 14132 5306
rect 13685 5284 13713 5290
rect 13964 5289 14132 5290
rect 13294 5276 13444 5279
rect 13685 5276 13712 5284
rect 13294 5274 13712 5276
rect 13294 5256 13303 5274
rect 13321 5256 13712 5274
rect 14425 5261 14456 5312
rect 14491 5341 14528 5411
rect 14794 5410 14831 5411
rect 14643 5351 14679 5352
rect 14491 5321 14500 5341
rect 14520 5321 14528 5341
rect 14491 5311 14528 5321
rect 14587 5341 14735 5351
rect 14835 5348 14931 5350
rect 14587 5321 14596 5341
rect 14616 5321 14706 5341
rect 14726 5321 14735 5341
rect 14587 5312 14735 5321
rect 14793 5341 14931 5348
rect 14793 5321 14802 5341
rect 14822 5321 14931 5341
rect 14793 5312 14931 5321
rect 14587 5311 14624 5312
rect 14317 5258 14358 5259
rect 13294 5253 13712 5256
rect 13294 5247 13337 5253
rect 13297 5244 13337 5247
rect 14212 5251 14358 5258
rect 13694 5235 13734 5236
rect 13405 5218 13734 5235
rect 14212 5231 14268 5251
rect 14288 5231 14327 5251
rect 14347 5231 14358 5251
rect 14212 5223 14358 5231
rect 14425 5254 14582 5261
rect 14425 5234 14545 5254
rect 14565 5234 14582 5254
rect 14425 5224 14582 5234
rect 14425 5223 14460 5224
rect 13289 5175 13332 5186
rect 13289 5157 13301 5175
rect 13319 5157 13332 5175
rect 13289 5131 13332 5157
rect 13405 5131 13432 5218
rect 13694 5209 13734 5218
rect 12468 5105 12907 5123
rect 11536 5104 11577 5105
rect 11270 5051 11307 5052
rect 10966 5042 11101 5051
rect 10966 5022 11072 5042
rect 11092 5022 11101 5042
rect 10966 5015 11101 5022
rect 11159 5042 11307 5051
rect 11159 5022 11168 5042
rect 11188 5022 11278 5042
rect 11298 5022 11307 5042
rect 10966 5013 11059 5015
rect 11159 5012 11307 5022
rect 11366 5042 11403 5052
rect 11366 5022 11374 5042
rect 11394 5022 11403 5042
rect 11215 5011 11251 5012
rect 11063 4952 11100 4953
rect 11366 4952 11403 5022
rect 11438 5051 11469 5102
rect 12468 5087 12868 5105
rect 12886 5087 12907 5105
rect 12468 5081 12907 5087
rect 12474 5077 12907 5081
rect 13289 5110 13432 5131
rect 13476 5183 13510 5199
rect 13694 5189 14087 5209
rect 14107 5189 14110 5209
rect 14425 5202 14456 5223
rect 14643 5202 14679 5312
rect 14698 5311 14735 5312
rect 14794 5311 14831 5312
rect 14754 5252 14844 5258
rect 14754 5232 14763 5252
rect 14783 5250 14844 5252
rect 14783 5232 14808 5250
rect 14754 5230 14808 5232
rect 14828 5230 14844 5250
rect 14754 5224 14844 5230
rect 14268 5201 14305 5202
rect 13694 5184 14110 5189
rect 14267 5192 14305 5201
rect 13694 5183 14035 5184
rect 13476 5113 13513 5183
rect 13628 5123 13659 5124
rect 13289 5108 13426 5110
rect 12853 5075 12905 5077
rect 13289 5066 13332 5108
rect 13476 5093 13485 5113
rect 13505 5093 13513 5113
rect 13476 5083 13513 5093
rect 13572 5113 13659 5123
rect 13572 5093 13581 5113
rect 13601 5093 13659 5113
rect 13572 5084 13659 5093
rect 13572 5083 13609 5084
rect 13287 5056 13332 5066
rect 11488 5051 11525 5052
rect 11438 5042 11525 5051
rect 11438 5022 11496 5042
rect 11516 5022 11525 5042
rect 11438 5012 11525 5022
rect 11584 5042 11621 5052
rect 11584 5022 11592 5042
rect 11612 5022 11621 5042
rect 13287 5038 13296 5056
rect 13314 5038 13332 5056
rect 13287 5032 13332 5038
rect 13628 5033 13659 5084
rect 13694 5113 13731 5183
rect 13997 5182 14034 5183
rect 14267 5172 14276 5192
rect 14296 5172 14305 5192
rect 14267 5164 14305 5172
rect 14371 5196 14456 5202
rect 14486 5201 14523 5202
rect 14371 5176 14379 5196
rect 14399 5176 14456 5196
rect 14371 5168 14456 5176
rect 14485 5192 14523 5201
rect 14485 5172 14494 5192
rect 14514 5172 14523 5192
rect 14371 5167 14407 5168
rect 14485 5164 14523 5172
rect 14589 5196 14733 5202
rect 14589 5176 14597 5196
rect 14617 5193 14705 5196
rect 14617 5176 14652 5193
rect 14589 5175 14652 5176
rect 14671 5176 14705 5193
rect 14725 5176 14733 5196
rect 14671 5175 14733 5176
rect 14589 5168 14733 5175
rect 14589 5167 14625 5168
rect 14697 5167 14733 5168
rect 14799 5201 14836 5202
rect 14799 5200 14837 5201
rect 14859 5200 14886 5204
rect 14799 5198 14886 5200
rect 14799 5192 14863 5198
rect 14799 5172 14808 5192
rect 14828 5178 14863 5192
rect 14883 5178 14886 5198
rect 14828 5173 14886 5178
rect 14828 5172 14863 5173
rect 14268 5135 14305 5164
rect 14269 5133 14305 5135
rect 13846 5123 13882 5124
rect 13694 5093 13703 5113
rect 13723 5093 13731 5113
rect 13694 5083 13731 5093
rect 13790 5113 13938 5123
rect 14038 5120 14134 5122
rect 13790 5093 13799 5113
rect 13819 5093 13909 5113
rect 13929 5093 13938 5113
rect 13790 5084 13938 5093
rect 13996 5113 14134 5120
rect 13996 5093 14005 5113
rect 14025 5093 14134 5113
rect 14269 5111 14460 5133
rect 14486 5132 14523 5164
rect 14799 5160 14863 5172
rect 14903 5134 14930 5312
rect 14762 5132 14930 5134
rect 14486 5106 14930 5132
rect 13996 5084 14134 5093
rect 13790 5083 13827 5084
rect 13287 5029 13324 5032
rect 13520 5030 13561 5031
rect 11438 5011 11469 5012
rect 11062 4951 11403 4952
rect 11584 4951 11621 5022
rect 13412 5023 13561 5030
rect 12856 5010 12893 5015
rect 10987 4946 11403 4951
rect 10987 4926 10990 4946
rect 11010 4926 11403 4946
rect 11434 4927 11621 4951
rect 12847 5006 12894 5010
rect 12847 4988 12866 5006
rect 12884 4988 12894 5006
rect 13412 5003 13471 5023
rect 13491 5003 13530 5023
rect 13550 5003 13561 5023
rect 13412 4995 13561 5003
rect 13628 5026 13785 5033
rect 13628 5006 13748 5026
rect 13768 5006 13785 5026
rect 13628 4996 13785 5006
rect 13628 4995 13663 4996
rect 12455 4929 12493 4930
rect 12847 4929 12894 4988
rect 13628 4974 13659 4995
rect 13846 4974 13882 5084
rect 13901 5083 13938 5084
rect 13997 5083 14034 5084
rect 13957 5024 14047 5030
rect 13957 5004 13966 5024
rect 13986 5022 14047 5024
rect 13986 5004 14011 5022
rect 13957 5002 14011 5004
rect 14031 5002 14047 5022
rect 13957 4996 14047 5002
rect 13471 4973 13508 4974
rect 13284 4965 13321 4967
rect 13284 4957 13326 4965
rect 13284 4939 13294 4957
rect 13312 4939 13326 4957
rect 13284 4930 13326 4939
rect 13470 4964 13508 4973
rect 13470 4944 13479 4964
rect 13499 4944 13508 4964
rect 13470 4936 13508 4944
rect 13574 4968 13659 4974
rect 13689 4973 13726 4974
rect 13574 4948 13582 4968
rect 13602 4948 13659 4968
rect 13574 4940 13659 4948
rect 13688 4964 13726 4973
rect 13688 4944 13697 4964
rect 13717 4944 13726 4964
rect 13574 4939 13610 4940
rect 13688 4936 13726 4944
rect 13792 4972 13936 4974
rect 13792 4968 13844 4972
rect 13792 4948 13800 4968
rect 13820 4952 13844 4968
rect 13864 4968 13936 4972
rect 13864 4952 13908 4968
rect 13820 4948 13908 4952
rect 13928 4948 13936 4968
rect 13792 4940 13936 4948
rect 13792 4939 13828 4940
rect 13900 4939 13936 4940
rect 14002 4973 14039 4974
rect 14002 4972 14040 4973
rect 14002 4964 14066 4972
rect 14002 4944 14011 4964
rect 14031 4950 14066 4964
rect 14086 4950 14089 4970
rect 14031 4945 14089 4950
rect 14031 4944 14066 4945
rect 11207 4925 11272 4926
rect 9322 4847 9360 4848
rect 8921 4809 9360 4847
rect 10232 4847 10240 4869
rect 10264 4847 10272 4869
rect 10232 4839 10272 4847
rect 11543 4891 11583 4899
rect 11543 4869 11551 4891
rect 11575 4869 11583 4891
rect 12455 4891 12894 4929
rect 12455 4890 12493 4891
rect 10543 4812 10608 4813
rect 7736 4794 7771 4795
rect 7713 4789 7771 4794
rect 7713 4769 7716 4789
rect 7736 4775 7771 4789
rect 7791 4775 7800 4795
rect 7736 4767 7800 4775
rect 7762 4766 7800 4767
rect 7763 4765 7800 4766
rect 7866 4799 7902 4800
rect 7974 4799 8010 4800
rect 7866 4791 8010 4799
rect 7866 4771 7874 4791
rect 7894 4787 7982 4791
rect 7894 4771 7938 4787
rect 7866 4767 7938 4771
rect 7958 4771 7982 4787
rect 8002 4771 8010 4791
rect 7958 4767 8010 4771
rect 7866 4765 8010 4767
rect 8076 4795 8114 4803
rect 8192 4799 8228 4800
rect 8076 4775 8085 4795
rect 8105 4775 8114 4795
rect 8076 4766 8114 4775
rect 8143 4791 8228 4799
rect 8143 4771 8200 4791
rect 8220 4771 8228 4791
rect 8076 4765 8113 4766
rect 8143 4765 8228 4771
rect 8294 4795 8332 4803
rect 8294 4775 8303 4795
rect 8323 4775 8332 4795
rect 8294 4766 8332 4775
rect 8476 4800 8518 4809
rect 8476 4782 8490 4800
rect 8508 4782 8518 4800
rect 8476 4774 8518 4782
rect 8481 4772 8518 4774
rect 8294 4765 8331 4766
rect 7755 4737 7845 4743
rect 7755 4717 7771 4737
rect 7791 4735 7845 4737
rect 7791 4717 7816 4735
rect 7755 4715 7816 4717
rect 7836 4715 7845 4735
rect 7755 4709 7845 4715
rect 7768 4655 7805 4656
rect 7864 4655 7901 4656
rect 7920 4655 7956 4765
rect 8143 4744 8174 4765
rect 8921 4750 8968 4809
rect 9322 4808 9360 4809
rect 8139 4743 8174 4744
rect 8017 4733 8174 4743
rect 8017 4713 8034 4733
rect 8054 4713 8174 4733
rect 8017 4706 8174 4713
rect 8241 4736 8390 4744
rect 8241 4716 8252 4736
rect 8272 4716 8311 4736
rect 8331 4716 8390 4736
rect 8921 4732 8931 4750
rect 8949 4732 8968 4750
rect 8921 4728 8968 4732
rect 10194 4787 10381 4811
rect 10412 4792 10805 4812
rect 10825 4792 10828 4812
rect 10412 4787 10828 4792
rect 8922 4723 8959 4728
rect 8241 4709 8390 4716
rect 10194 4716 10231 4787
rect 10412 4786 10753 4787
rect 10346 4726 10377 4727
rect 8241 4708 8282 4709
rect 8478 4707 8515 4710
rect 7975 4655 8012 4656
rect 7668 4646 7806 4655
rect 6872 4607 7316 4633
rect 6872 4605 7040 4607
rect 6872 4427 6899 4605
rect 6939 4567 7003 4579
rect 7279 4575 7316 4607
rect 7342 4606 7533 4628
rect 7668 4626 7777 4646
rect 7797 4626 7806 4646
rect 7668 4619 7806 4626
rect 7864 4646 8012 4655
rect 7864 4626 7873 4646
rect 7893 4626 7983 4646
rect 8003 4626 8012 4646
rect 7668 4617 7764 4619
rect 7864 4616 8012 4626
rect 8071 4646 8108 4656
rect 8071 4626 8079 4646
rect 8099 4626 8108 4646
rect 7920 4615 7956 4616
rect 7497 4604 7533 4606
rect 7497 4575 7534 4604
rect 6939 4566 6974 4567
rect 6916 4561 6974 4566
rect 6916 4541 6919 4561
rect 6939 4547 6974 4561
rect 6994 4547 7003 4567
rect 6939 4541 7003 4547
rect 6916 4539 7003 4541
rect 6916 4535 6943 4539
rect 6965 4538 7003 4539
rect 6966 4537 7003 4538
rect 7069 4571 7105 4572
rect 7177 4571 7213 4572
rect 7069 4564 7213 4571
rect 7069 4563 7131 4564
rect 7069 4543 7077 4563
rect 7097 4546 7131 4563
rect 7150 4563 7213 4564
rect 7150 4546 7185 4563
rect 7097 4543 7185 4546
rect 7205 4543 7213 4563
rect 7069 4537 7213 4543
rect 7279 4567 7317 4575
rect 7395 4571 7431 4572
rect 7279 4547 7288 4567
rect 7308 4547 7317 4567
rect 7279 4538 7317 4547
rect 7346 4563 7431 4571
rect 7346 4543 7403 4563
rect 7423 4543 7431 4563
rect 7279 4537 7316 4538
rect 7346 4537 7431 4543
rect 7497 4567 7535 4575
rect 7497 4547 7506 4567
rect 7526 4547 7535 4567
rect 7768 4556 7805 4557
rect 8071 4556 8108 4626
rect 8143 4655 8174 4706
rect 8470 4701 8515 4707
rect 8470 4683 8488 4701
rect 8506 4683 8515 4701
rect 10194 4696 10203 4716
rect 10223 4696 10231 4716
rect 10194 4686 10231 4696
rect 10290 4716 10377 4726
rect 10290 4696 10299 4716
rect 10319 4696 10377 4716
rect 10290 4687 10377 4696
rect 10290 4686 10327 4687
rect 8470 4673 8515 4683
rect 8193 4655 8230 4656
rect 8143 4646 8230 4655
rect 8143 4626 8201 4646
rect 8221 4626 8230 4646
rect 8143 4616 8230 4626
rect 8289 4646 8326 4656
rect 8289 4626 8297 4646
rect 8317 4626 8326 4646
rect 8470 4631 8513 4673
rect 8910 4661 8962 4663
rect 8376 4629 8513 4631
rect 8143 4615 8174 4616
rect 8289 4556 8326 4626
rect 7767 4555 8108 4556
rect 7497 4538 7535 4547
rect 7692 4550 8108 4555
rect 7497 4537 7534 4538
rect 6958 4509 7048 4515
rect 6958 4489 6974 4509
rect 6994 4507 7048 4509
rect 6994 4489 7019 4507
rect 6958 4487 7019 4489
rect 7039 4487 7048 4507
rect 6958 4481 7048 4487
rect 6971 4427 7008 4428
rect 7067 4427 7104 4428
rect 7123 4427 7159 4537
rect 7346 4516 7377 4537
rect 7692 4530 7695 4550
rect 7715 4530 8108 4550
rect 8292 4540 8326 4556
rect 8370 4608 8513 4629
rect 8908 4657 9341 4661
rect 8908 4651 9347 4657
rect 8908 4633 8929 4651
rect 8947 4633 9347 4651
rect 10346 4636 10377 4687
rect 10412 4716 10449 4786
rect 10715 4785 10752 4786
rect 10564 4726 10600 4727
rect 10412 4696 10421 4716
rect 10441 4696 10449 4716
rect 10412 4686 10449 4696
rect 10508 4716 10656 4726
rect 10756 4723 10852 4725
rect 10508 4696 10517 4716
rect 10537 4696 10627 4716
rect 10647 4696 10656 4716
rect 10508 4687 10656 4696
rect 10714 4716 10852 4723
rect 10714 4696 10723 4716
rect 10743 4696 10852 4716
rect 10714 4687 10852 4696
rect 10508 4686 10545 4687
rect 10238 4633 10279 4634
rect 8908 4615 9347 4633
rect 8068 4521 8108 4530
rect 8370 4521 8397 4608
rect 8470 4582 8513 4608
rect 8470 4564 8483 4582
rect 8501 4564 8513 4582
rect 8470 4553 8513 4564
rect 7342 4515 7377 4516
rect 7220 4505 7377 4515
rect 7220 4485 7237 4505
rect 7257 4485 7377 4505
rect 7220 4478 7377 4485
rect 7444 4508 7590 4516
rect 7444 4488 7455 4508
rect 7475 4488 7514 4508
rect 7534 4488 7590 4508
rect 8068 4504 8397 4521
rect 8068 4503 8108 4504
rect 7444 4481 7590 4488
rect 8465 4492 8505 4495
rect 8465 4486 8508 4492
rect 8090 4483 8508 4486
rect 7444 4480 7485 4481
rect 7178 4427 7215 4428
rect 6871 4418 7009 4427
rect 6871 4398 6980 4418
rect 7000 4398 7009 4418
rect 6871 4391 7009 4398
rect 7067 4418 7215 4427
rect 7067 4398 7076 4418
rect 7096 4398 7186 4418
rect 7206 4398 7215 4418
rect 6871 4389 6967 4391
rect 7067 4388 7215 4398
rect 7274 4418 7311 4428
rect 7274 4398 7282 4418
rect 7302 4398 7311 4418
rect 7123 4387 7159 4388
rect 6971 4328 7008 4329
rect 7274 4328 7311 4398
rect 7346 4427 7377 4478
rect 8090 4465 8481 4483
rect 8499 4465 8508 4483
rect 8090 4463 8508 4465
rect 8090 4455 8117 4463
rect 8358 4460 8508 4463
rect 7670 4449 7838 4450
rect 8089 4449 8117 4455
rect 7670 4433 8117 4449
rect 8465 4455 8508 4460
rect 7396 4427 7433 4428
rect 7346 4418 7433 4427
rect 7346 4398 7404 4418
rect 7424 4398 7433 4418
rect 7346 4388 7433 4398
rect 7492 4418 7529 4428
rect 7492 4398 7500 4418
rect 7520 4398 7529 4418
rect 7346 4387 7377 4388
rect 6970 4327 7311 4328
rect 7492 4327 7529 4398
rect 6895 4322 7311 4327
rect 6895 4302 6898 4322
rect 6918 4302 7311 4322
rect 7342 4303 7529 4327
rect 7670 4423 8114 4433
rect 7670 4421 7838 4423
rect 6704 4228 6748 4229
rect 6704 4222 6749 4228
rect 6704 4204 6716 4222
rect 6738 4204 6749 4222
rect 6770 4223 6812 4268
rect 7670 4243 7697 4421
rect 7737 4383 7801 4395
rect 8077 4391 8114 4423
rect 8140 4422 8331 4444
rect 8295 4420 8331 4422
rect 8295 4391 8332 4420
rect 8465 4399 8505 4455
rect 7737 4382 7772 4383
rect 7714 4377 7772 4382
rect 7714 4357 7717 4377
rect 7737 4363 7772 4377
rect 7792 4363 7801 4383
rect 7737 4355 7801 4363
rect 7763 4354 7801 4355
rect 7764 4353 7801 4354
rect 7867 4387 7903 4388
rect 7975 4387 8011 4388
rect 7867 4379 8011 4387
rect 7867 4359 7875 4379
rect 7895 4359 7930 4379
rect 7950 4359 7983 4379
rect 8003 4359 8011 4379
rect 7867 4353 8011 4359
rect 8077 4383 8115 4391
rect 8193 4387 8229 4388
rect 8077 4363 8086 4383
rect 8106 4363 8115 4383
rect 8077 4354 8115 4363
rect 8144 4379 8229 4387
rect 8144 4359 8201 4379
rect 8221 4359 8229 4379
rect 8077 4353 8114 4354
rect 8144 4353 8229 4359
rect 8295 4383 8333 4391
rect 8295 4363 8304 4383
rect 8324 4363 8333 4383
rect 8465 4381 8477 4399
rect 8495 4381 8505 4399
rect 8910 4426 8962 4615
rect 9308 4590 9347 4615
rect 10130 4626 10279 4633
rect 10130 4606 10189 4626
rect 10209 4606 10248 4626
rect 10268 4606 10279 4626
rect 10130 4598 10279 4606
rect 10346 4629 10503 4636
rect 10346 4609 10466 4629
rect 10486 4609 10503 4629
rect 10346 4599 10503 4609
rect 10346 4598 10381 4599
rect 9092 4565 9279 4589
rect 9308 4570 9703 4590
rect 9723 4570 9726 4590
rect 10346 4577 10377 4598
rect 10564 4577 10600 4687
rect 10619 4686 10656 4687
rect 10715 4686 10752 4687
rect 10675 4627 10765 4633
rect 10675 4607 10684 4627
rect 10704 4625 10765 4627
rect 10704 4607 10729 4625
rect 10675 4605 10729 4607
rect 10749 4605 10765 4625
rect 10675 4599 10765 4605
rect 10189 4576 10226 4577
rect 9308 4565 9726 4570
rect 10188 4567 10226 4576
rect 9092 4494 9129 4565
rect 9308 4564 9651 4565
rect 9308 4561 9347 4564
rect 9613 4563 9650 4564
rect 9244 4504 9275 4505
rect 9092 4474 9101 4494
rect 9121 4474 9129 4494
rect 9092 4464 9129 4474
rect 9188 4494 9275 4504
rect 9188 4474 9197 4494
rect 9217 4474 9275 4494
rect 9188 4465 9275 4474
rect 9188 4464 9225 4465
rect 8910 4408 8926 4426
rect 8944 4408 8962 4426
rect 9244 4414 9275 4465
rect 9310 4494 9347 4561
rect 10188 4547 10197 4567
rect 10217 4547 10226 4567
rect 10188 4539 10226 4547
rect 10292 4571 10377 4577
rect 10407 4576 10444 4577
rect 10292 4551 10300 4571
rect 10320 4551 10377 4571
rect 10292 4543 10377 4551
rect 10406 4567 10444 4576
rect 10406 4547 10415 4567
rect 10435 4547 10444 4567
rect 10292 4542 10328 4543
rect 10406 4539 10444 4547
rect 10510 4571 10654 4577
rect 10510 4551 10518 4571
rect 10538 4565 10626 4571
rect 10538 4551 10567 4565
rect 10510 4543 10567 4551
rect 10510 4542 10546 4543
rect 10590 4551 10626 4565
rect 10646 4551 10654 4571
rect 10590 4543 10654 4551
rect 10618 4542 10654 4543
rect 10720 4576 10757 4577
rect 10720 4575 10758 4576
rect 10720 4567 10784 4575
rect 10720 4547 10729 4567
rect 10749 4553 10784 4567
rect 10804 4553 10807 4573
rect 10749 4548 10807 4553
rect 10749 4547 10784 4548
rect 10189 4510 10226 4539
rect 10190 4508 10226 4510
rect 9462 4504 9498 4505
rect 9310 4474 9319 4494
rect 9339 4474 9347 4494
rect 9310 4464 9347 4474
rect 9406 4494 9554 4504
rect 9654 4501 9750 4503
rect 9406 4474 9415 4494
rect 9435 4474 9525 4494
rect 9545 4474 9554 4494
rect 9406 4465 9554 4474
rect 9612 4494 9750 4501
rect 9612 4474 9621 4494
rect 9641 4474 9750 4494
rect 10190 4486 10381 4508
rect 10407 4507 10444 4539
rect 10720 4535 10784 4547
rect 10824 4509 10851 4687
rect 11148 4640 11185 4646
rect 11148 4621 11156 4640
rect 11177 4621 11185 4640
rect 11148 4613 11185 4621
rect 10683 4507 10851 4509
rect 10407 4481 10851 4507
rect 10517 4479 10557 4481
rect 10683 4480 10851 4481
rect 9612 4465 9750 4474
rect 10810 4475 10851 4480
rect 9406 4464 9443 4465
rect 9136 4411 9177 4412
rect 8910 4390 8962 4408
rect 9028 4404 9177 4411
rect 8465 4371 8505 4381
rect 9028 4384 9087 4404
rect 9107 4384 9146 4404
rect 9166 4384 9177 4404
rect 9028 4376 9177 4384
rect 9244 4407 9401 4414
rect 9244 4387 9364 4407
rect 9384 4387 9401 4407
rect 9244 4377 9401 4387
rect 9244 4376 9279 4377
rect 8295 4354 8333 4363
rect 9244 4355 9275 4376
rect 9462 4355 9498 4465
rect 9517 4464 9554 4465
rect 9613 4464 9650 4465
rect 9573 4405 9663 4411
rect 9573 4385 9582 4405
rect 9602 4403 9663 4405
rect 9602 4385 9627 4403
rect 9573 4383 9627 4385
rect 9647 4383 9663 4403
rect 9573 4377 9663 4383
rect 9087 4354 9124 4355
rect 8295 4353 8332 4354
rect 7756 4325 7846 4331
rect 7756 4305 7772 4325
rect 7792 4323 7846 4325
rect 7792 4305 7817 4323
rect 7756 4303 7817 4305
rect 7837 4303 7846 4323
rect 7756 4297 7846 4303
rect 7769 4243 7806 4244
rect 7865 4243 7902 4244
rect 7921 4243 7957 4353
rect 8144 4332 8175 4353
rect 9086 4345 9124 4354
rect 8140 4331 8175 4332
rect 8018 4321 8175 4331
rect 8018 4301 8035 4321
rect 8055 4301 8175 4321
rect 8018 4294 8175 4301
rect 8242 4324 8391 4332
rect 8242 4304 8253 4324
rect 8273 4304 8312 4324
rect 8332 4304 8391 4324
rect 8914 4327 8954 4337
rect 8242 4297 8391 4304
rect 8457 4300 8509 4318
rect 8242 4296 8283 4297
rect 7976 4243 8013 4244
rect 7669 4234 7807 4243
rect 7141 4223 7174 4225
rect 6770 4211 7217 4223
rect 6704 4174 6749 4204
rect 6721 3228 6749 4174
rect 6773 4197 7217 4211
rect 6773 4195 6941 4197
rect 6773 4017 6800 4195
rect 6840 4157 6904 4169
rect 7180 4165 7217 4197
rect 7243 4196 7434 4218
rect 7669 4214 7778 4234
rect 7798 4214 7807 4234
rect 7669 4207 7807 4214
rect 7865 4234 8013 4243
rect 7865 4214 7874 4234
rect 7894 4214 7984 4234
rect 8004 4214 8013 4234
rect 7669 4205 7765 4207
rect 7865 4204 8013 4214
rect 8072 4234 8109 4244
rect 8072 4214 8080 4234
rect 8100 4214 8109 4234
rect 7921 4203 7957 4204
rect 7398 4194 7434 4196
rect 7398 4165 7435 4194
rect 6840 4156 6875 4157
rect 6817 4151 6875 4156
rect 6817 4131 6820 4151
rect 6840 4137 6875 4151
rect 6895 4137 6904 4157
rect 6840 4129 6904 4137
rect 6866 4128 6904 4129
rect 6867 4127 6904 4128
rect 6970 4161 7006 4162
rect 7078 4161 7114 4162
rect 6970 4155 7114 4161
rect 6970 4153 7031 4155
rect 6970 4133 6978 4153
rect 6998 4138 7031 4153
rect 7050 4153 7114 4155
rect 7050 4138 7086 4153
rect 6998 4133 7086 4138
rect 7106 4133 7114 4153
rect 6970 4127 7114 4133
rect 7180 4157 7218 4165
rect 7296 4161 7332 4162
rect 7180 4137 7189 4157
rect 7209 4137 7218 4157
rect 7180 4128 7218 4137
rect 7247 4153 7332 4161
rect 7247 4133 7304 4153
rect 7324 4133 7332 4153
rect 7180 4127 7217 4128
rect 7247 4127 7332 4133
rect 7398 4157 7436 4165
rect 7398 4137 7407 4157
rect 7427 4137 7436 4157
rect 8072 4147 8109 4214
rect 8144 4243 8175 4294
rect 8457 4282 8475 4300
rect 8493 4282 8509 4300
rect 8194 4243 8231 4244
rect 8144 4234 8231 4243
rect 8144 4214 8202 4234
rect 8222 4214 8231 4234
rect 8144 4204 8231 4214
rect 8290 4234 8327 4244
rect 8290 4214 8298 4234
rect 8318 4214 8327 4234
rect 8144 4203 8175 4204
rect 7769 4144 7806 4145
rect 8072 4144 8111 4147
rect 7768 4143 8111 4144
rect 8290 4143 8327 4214
rect 7398 4128 7436 4137
rect 7693 4138 8111 4143
rect 7398 4127 7435 4128
rect 6859 4099 6949 4105
rect 6859 4079 6875 4099
rect 6895 4097 6949 4099
rect 6895 4079 6920 4097
rect 6859 4077 6920 4079
rect 6940 4077 6949 4097
rect 6859 4071 6949 4077
rect 6872 4017 6909 4018
rect 6968 4017 7005 4018
rect 7024 4017 7060 4127
rect 7247 4106 7278 4127
rect 7693 4118 7696 4138
rect 7716 4118 8111 4138
rect 8140 4119 8327 4143
rect 7243 4105 7278 4106
rect 7121 4095 7278 4105
rect 7121 4075 7138 4095
rect 7158 4075 7278 4095
rect 7121 4068 7278 4075
rect 7345 4098 7494 4106
rect 7345 4078 7356 4098
rect 7376 4078 7415 4098
rect 7435 4078 7494 4098
rect 7345 4071 7494 4078
rect 8072 4093 8111 4118
rect 8457 4093 8509 4282
rect 8914 4309 8924 4327
rect 8942 4309 8954 4327
rect 9086 4325 9095 4345
rect 9115 4325 9124 4345
rect 9086 4317 9124 4325
rect 9190 4349 9275 4355
rect 9305 4354 9342 4355
rect 9190 4329 9198 4349
rect 9218 4329 9275 4349
rect 9190 4321 9275 4329
rect 9304 4345 9342 4354
rect 9304 4325 9313 4345
rect 9333 4325 9342 4345
rect 9190 4320 9226 4321
rect 9304 4317 9342 4325
rect 9408 4349 9552 4355
rect 9408 4329 9416 4349
rect 9436 4329 9469 4349
rect 9489 4329 9524 4349
rect 9544 4329 9552 4349
rect 9408 4321 9552 4329
rect 9408 4320 9444 4321
rect 9516 4320 9552 4321
rect 9618 4354 9655 4355
rect 9618 4353 9656 4354
rect 9618 4345 9682 4353
rect 9618 4325 9627 4345
rect 9647 4331 9682 4345
rect 9702 4331 9705 4351
rect 9647 4326 9705 4331
rect 9647 4325 9682 4326
rect 8914 4253 8954 4309
rect 9087 4288 9124 4317
rect 9088 4286 9124 4288
rect 9088 4264 9279 4286
rect 9305 4285 9342 4317
rect 9618 4313 9682 4325
rect 9722 4287 9749 4465
rect 9581 4285 9749 4287
rect 9305 4275 9749 4285
rect 9890 4381 10077 4405
rect 10108 4386 10501 4406
rect 10521 4386 10524 4406
rect 10108 4381 10524 4386
rect 9890 4310 9927 4381
rect 10108 4380 10449 4381
rect 10042 4320 10073 4321
rect 9890 4290 9899 4310
rect 9919 4290 9927 4310
rect 9890 4280 9927 4290
rect 9986 4310 10073 4320
rect 9986 4290 9995 4310
rect 10015 4290 10073 4310
rect 9986 4281 10073 4290
rect 9986 4280 10023 4281
rect 8911 4248 8954 4253
rect 9302 4259 9749 4275
rect 9302 4253 9330 4259
rect 9581 4258 9749 4259
rect 8911 4245 9061 4248
rect 9302 4245 9329 4253
rect 8911 4243 9329 4245
rect 8911 4225 8920 4243
rect 8938 4225 9329 4243
rect 10042 4230 10073 4281
rect 10108 4310 10145 4380
rect 10411 4379 10448 4380
rect 10260 4320 10296 4321
rect 10108 4290 10117 4310
rect 10137 4290 10145 4310
rect 10108 4280 10145 4290
rect 10204 4310 10352 4320
rect 10452 4317 10548 4319
rect 10204 4290 10213 4310
rect 10233 4290 10323 4310
rect 10343 4290 10352 4310
rect 10204 4281 10352 4290
rect 10410 4310 10548 4317
rect 10410 4290 10419 4310
rect 10439 4290 10548 4310
rect 10810 4293 10850 4475
rect 10410 4281 10548 4290
rect 10204 4280 10241 4281
rect 9934 4227 9975 4228
rect 8911 4222 9329 4225
rect 8911 4216 8954 4222
rect 8914 4213 8954 4216
rect 9826 4220 9975 4227
rect 9311 4204 9351 4205
rect 9022 4187 9351 4204
rect 9826 4200 9885 4220
rect 9905 4200 9944 4220
rect 9964 4200 9975 4220
rect 9826 4192 9975 4200
rect 10042 4223 10199 4230
rect 10042 4203 10162 4223
rect 10182 4203 10199 4223
rect 10042 4193 10199 4203
rect 10042 4192 10077 4193
rect 8906 4144 8949 4155
rect 8906 4126 8918 4144
rect 8936 4126 8949 4144
rect 8906 4100 8949 4126
rect 9022 4100 9049 4187
rect 9311 4178 9351 4187
rect 8072 4075 8511 4093
rect 7345 4070 7386 4071
rect 7079 4017 7116 4018
rect 6772 4008 6910 4017
rect 6772 3988 6881 4008
rect 6901 3988 6910 4008
rect 6772 3981 6910 3988
rect 6968 4008 7116 4017
rect 6968 3988 6977 4008
rect 6997 3988 7087 4008
rect 7107 3988 7116 4008
rect 6772 3979 6868 3981
rect 6968 3978 7116 3988
rect 7175 4008 7212 4018
rect 7175 3988 7183 4008
rect 7203 3988 7212 4008
rect 7024 3977 7060 3978
rect 6872 3918 6909 3919
rect 7175 3918 7212 3988
rect 7247 4017 7278 4068
rect 8072 4057 8472 4075
rect 8490 4057 8511 4075
rect 8072 4051 8511 4057
rect 8078 4047 8511 4051
rect 8906 4079 9049 4100
rect 9093 4152 9127 4168
rect 9311 4158 9704 4178
rect 9724 4158 9727 4178
rect 10042 4171 10073 4192
rect 10260 4171 10296 4281
rect 10315 4280 10352 4281
rect 10411 4280 10448 4281
rect 10371 4221 10461 4227
rect 10371 4201 10380 4221
rect 10400 4219 10461 4221
rect 10400 4201 10425 4219
rect 10371 4199 10425 4201
rect 10445 4199 10461 4219
rect 10371 4193 10461 4199
rect 9885 4170 9922 4171
rect 9311 4153 9727 4158
rect 9884 4161 9922 4170
rect 9311 4152 9652 4153
rect 9093 4082 9130 4152
rect 9245 4092 9276 4093
rect 8906 4077 9043 4079
rect 8457 4045 8509 4047
rect 8906 4035 8949 4077
rect 9093 4062 9102 4082
rect 9122 4062 9130 4082
rect 9093 4052 9130 4062
rect 9189 4082 9276 4092
rect 9189 4062 9198 4082
rect 9218 4062 9276 4082
rect 9189 4053 9276 4062
rect 9189 4052 9226 4053
rect 8904 4025 8949 4035
rect 7297 4017 7334 4018
rect 7247 4008 7334 4017
rect 7247 3988 7305 4008
rect 7325 3988 7334 4008
rect 7247 3978 7334 3988
rect 7393 4008 7430 4018
rect 7393 3988 7401 4008
rect 7421 3988 7430 4008
rect 8904 4007 8913 4025
rect 8931 4007 8949 4025
rect 8904 4001 8949 4007
rect 9245 4002 9276 4053
rect 9311 4082 9348 4152
rect 9614 4151 9651 4152
rect 9884 4141 9893 4161
rect 9913 4141 9922 4161
rect 9884 4133 9922 4141
rect 9988 4165 10073 4171
rect 10103 4170 10140 4171
rect 9988 4145 9996 4165
rect 10016 4145 10073 4165
rect 9988 4137 10073 4145
rect 10102 4161 10140 4170
rect 10102 4141 10111 4161
rect 10131 4141 10140 4161
rect 9988 4136 10024 4137
rect 10102 4133 10140 4141
rect 10206 4165 10350 4171
rect 10206 4145 10214 4165
rect 10234 4146 10266 4165
rect 10287 4146 10322 4165
rect 10234 4145 10322 4146
rect 10342 4145 10350 4165
rect 10206 4137 10350 4145
rect 10206 4136 10242 4137
rect 10314 4136 10350 4137
rect 10416 4170 10453 4171
rect 10416 4169 10454 4170
rect 10416 4161 10480 4169
rect 10416 4141 10425 4161
rect 10445 4147 10480 4161
rect 10500 4147 10503 4167
rect 10445 4142 10503 4147
rect 10445 4141 10480 4142
rect 9885 4104 9922 4133
rect 9886 4102 9922 4104
rect 9463 4092 9499 4093
rect 9311 4062 9320 4082
rect 9340 4062 9348 4082
rect 9311 4052 9348 4062
rect 9407 4082 9555 4092
rect 9655 4089 9751 4091
rect 9407 4062 9416 4082
rect 9436 4062 9526 4082
rect 9546 4062 9555 4082
rect 9407 4053 9555 4062
rect 9613 4082 9751 4089
rect 9613 4062 9622 4082
rect 9642 4062 9751 4082
rect 9886 4080 10077 4102
rect 10103 4101 10140 4133
rect 10416 4129 10480 4141
rect 10520 4103 10547 4281
rect 10379 4101 10547 4103
rect 10103 4075 10547 4101
rect 9613 4053 9751 4062
rect 9407 4052 9444 4053
rect 8904 3998 8941 4001
rect 9137 3999 9178 4000
rect 7247 3977 7278 3978
rect 6871 3917 7212 3918
rect 7393 3917 7430 3988
rect 9029 3992 9178 3999
rect 8460 3980 8497 3985
rect 8451 3976 8498 3980
rect 8451 3958 8470 3976
rect 8488 3958 8498 3976
rect 9029 3972 9088 3992
rect 9108 3972 9147 3992
rect 9167 3972 9178 3992
rect 9029 3964 9178 3972
rect 9245 3995 9402 4002
rect 9245 3975 9365 3995
rect 9385 3975 9402 3995
rect 9245 3965 9402 3975
rect 9245 3964 9280 3965
rect 6796 3912 7212 3917
rect 6796 3892 6799 3912
rect 6819 3892 7212 3912
rect 7243 3893 7430 3917
rect 8055 3915 8095 3920
rect 8451 3915 8498 3958
rect 9245 3943 9276 3964
rect 9463 3943 9499 4053
rect 9518 4052 9555 4053
rect 9614 4052 9651 4053
rect 9574 3993 9664 3999
rect 9574 3973 9583 3993
rect 9603 3991 9664 3993
rect 9603 3973 9628 3991
rect 9574 3971 9628 3973
rect 9648 3971 9664 3991
rect 9574 3965 9664 3971
rect 9088 3942 9125 3943
rect 8055 3876 8498 3915
rect 8901 3934 8938 3936
rect 8901 3926 8943 3934
rect 8901 3908 8911 3926
rect 8929 3908 8943 3926
rect 8901 3899 8943 3908
rect 9087 3933 9125 3942
rect 9087 3913 9096 3933
rect 9116 3913 9125 3933
rect 9087 3905 9125 3913
rect 9191 3937 9276 3943
rect 9306 3942 9343 3943
rect 9191 3917 9199 3937
rect 9219 3917 9276 3937
rect 9191 3909 9276 3917
rect 9305 3933 9343 3942
rect 9305 3913 9314 3933
rect 9334 3913 9343 3933
rect 9191 3908 9227 3909
rect 9305 3905 9343 3913
rect 9409 3941 9553 3943
rect 9409 3937 9461 3941
rect 9409 3917 9417 3937
rect 9437 3921 9461 3937
rect 9481 3937 9553 3941
rect 9481 3921 9525 3937
rect 9437 3917 9525 3921
rect 9545 3917 9553 3937
rect 9409 3909 9553 3917
rect 9409 3908 9445 3909
rect 9517 3908 9553 3909
rect 9619 3942 9656 3943
rect 9619 3941 9657 3942
rect 9619 3933 9683 3941
rect 9619 3913 9628 3933
rect 9648 3919 9683 3933
rect 9703 3919 9706 3939
rect 9648 3914 9706 3919
rect 9648 3913 9683 3914
rect 7149 3861 7189 3869
rect 7149 3839 7157 3861
rect 7181 3839 7189 3861
rect 6855 3615 7023 3616
rect 7149 3615 7189 3839
rect 7652 3843 7820 3844
rect 8055 3843 8095 3876
rect 8451 3843 8498 3876
rect 8902 3874 8943 3899
rect 9088 3874 9125 3905
rect 9306 3874 9343 3905
rect 9619 3901 9683 3913
rect 9723 3875 9750 4053
rect 8902 3847 8951 3874
rect 9087 3848 9136 3874
rect 9305 3873 9386 3874
rect 9582 3873 9750 3875
rect 9305 3848 9750 3873
rect 9306 3847 9750 3848
rect 7652 3842 8096 3843
rect 7652 3817 8097 3842
rect 7652 3815 7820 3817
rect 8016 3816 8097 3817
rect 8266 3816 8315 3842
rect 8451 3816 8500 3843
rect 7652 3637 7679 3815
rect 7719 3777 7783 3789
rect 8059 3785 8096 3816
rect 8277 3785 8314 3816
rect 8459 3791 8500 3816
rect 8904 3814 8951 3847
rect 9307 3814 9347 3847
rect 9582 3846 9750 3847
rect 10213 3851 10253 4075
rect 10379 4074 10547 4075
rect 10213 3829 10221 3851
rect 10245 3829 10253 3851
rect 10213 3821 10253 3829
rect 7719 3776 7754 3777
rect 7696 3771 7754 3776
rect 7696 3751 7699 3771
rect 7719 3757 7754 3771
rect 7774 3757 7783 3777
rect 7719 3749 7783 3757
rect 7745 3748 7783 3749
rect 7746 3747 7783 3748
rect 7849 3781 7885 3782
rect 7957 3781 7993 3782
rect 7849 3773 7993 3781
rect 7849 3753 7857 3773
rect 7877 3769 7965 3773
rect 7877 3753 7921 3769
rect 7849 3749 7921 3753
rect 7941 3753 7965 3769
rect 7985 3753 7993 3773
rect 7941 3749 7993 3753
rect 7849 3747 7993 3749
rect 8059 3777 8097 3785
rect 8175 3781 8211 3782
rect 8059 3757 8068 3777
rect 8088 3757 8097 3777
rect 8059 3748 8097 3757
rect 8126 3773 8211 3781
rect 8126 3753 8183 3773
rect 8203 3753 8211 3773
rect 8059 3747 8096 3748
rect 8126 3747 8211 3753
rect 8277 3777 8315 3785
rect 8277 3757 8286 3777
rect 8306 3757 8315 3777
rect 8277 3748 8315 3757
rect 8459 3782 8501 3791
rect 8459 3764 8473 3782
rect 8491 3764 8501 3782
rect 8459 3756 8501 3764
rect 8464 3754 8501 3756
rect 8904 3775 9347 3814
rect 8277 3747 8314 3748
rect 7738 3719 7828 3725
rect 7738 3699 7754 3719
rect 7774 3717 7828 3719
rect 7774 3699 7799 3717
rect 7738 3697 7799 3699
rect 7819 3697 7828 3717
rect 7738 3691 7828 3697
rect 7751 3637 7788 3638
rect 7847 3637 7884 3638
rect 7903 3637 7939 3747
rect 8126 3726 8157 3747
rect 8904 3732 8951 3775
rect 9307 3770 9347 3775
rect 9972 3773 10159 3797
rect 10190 3778 10583 3798
rect 10603 3778 10606 3798
rect 10190 3773 10606 3778
rect 8122 3725 8157 3726
rect 8000 3715 8157 3725
rect 8000 3695 8017 3715
rect 8037 3695 8157 3715
rect 8000 3688 8157 3695
rect 8224 3718 8373 3726
rect 8224 3698 8235 3718
rect 8255 3698 8294 3718
rect 8314 3698 8373 3718
rect 8904 3714 8914 3732
rect 8932 3714 8951 3732
rect 8904 3710 8951 3714
rect 8905 3705 8942 3710
rect 8224 3691 8373 3698
rect 9972 3702 10009 3773
rect 10190 3772 10531 3773
rect 10124 3712 10155 3713
rect 8224 3690 8265 3691
rect 8461 3689 8498 3692
rect 7958 3637 7995 3638
rect 7651 3628 7789 3637
rect 6855 3589 7299 3615
rect 6855 3587 7023 3589
rect 6855 3409 6882 3587
rect 6922 3549 6986 3561
rect 7262 3557 7299 3589
rect 7325 3588 7516 3610
rect 7651 3608 7760 3628
rect 7780 3608 7789 3628
rect 7651 3601 7789 3608
rect 7847 3628 7995 3637
rect 7847 3608 7856 3628
rect 7876 3608 7966 3628
rect 7986 3608 7995 3628
rect 7651 3599 7747 3601
rect 7847 3598 7995 3608
rect 8054 3628 8091 3638
rect 8054 3608 8062 3628
rect 8082 3608 8091 3628
rect 7903 3597 7939 3598
rect 7480 3586 7516 3588
rect 7480 3557 7517 3586
rect 6922 3548 6957 3549
rect 6899 3543 6957 3548
rect 6899 3523 6902 3543
rect 6922 3529 6957 3543
rect 6977 3529 6986 3549
rect 6922 3521 6986 3529
rect 6948 3520 6986 3521
rect 6949 3519 6986 3520
rect 7052 3553 7088 3554
rect 7160 3553 7196 3554
rect 7052 3545 7196 3553
rect 7052 3525 7060 3545
rect 7080 3544 7168 3545
rect 7080 3525 7115 3544
rect 7136 3525 7168 3544
rect 7188 3525 7196 3545
rect 7052 3519 7196 3525
rect 7262 3549 7300 3557
rect 7378 3553 7414 3554
rect 7262 3529 7271 3549
rect 7291 3529 7300 3549
rect 7262 3520 7300 3529
rect 7329 3545 7414 3553
rect 7329 3525 7386 3545
rect 7406 3525 7414 3545
rect 7262 3519 7299 3520
rect 7329 3519 7414 3525
rect 7480 3549 7518 3557
rect 7480 3529 7489 3549
rect 7509 3529 7518 3549
rect 7751 3538 7788 3539
rect 8054 3538 8091 3608
rect 8126 3637 8157 3688
rect 8453 3683 8498 3689
rect 8453 3665 8471 3683
rect 8489 3665 8498 3683
rect 9972 3682 9981 3702
rect 10001 3682 10009 3702
rect 9972 3672 10009 3682
rect 10068 3702 10155 3712
rect 10068 3682 10077 3702
rect 10097 3682 10155 3702
rect 10068 3673 10155 3682
rect 10068 3672 10105 3673
rect 8453 3655 8498 3665
rect 8176 3637 8213 3638
rect 8126 3628 8213 3637
rect 8126 3608 8184 3628
rect 8204 3608 8213 3628
rect 8126 3598 8213 3608
rect 8272 3628 8309 3638
rect 8272 3608 8280 3628
rect 8300 3608 8309 3628
rect 8453 3613 8496 3655
rect 8893 3643 8945 3645
rect 8359 3611 8496 3613
rect 8126 3597 8157 3598
rect 8272 3538 8309 3608
rect 7750 3537 8091 3538
rect 7480 3520 7518 3529
rect 7675 3532 8091 3537
rect 7480 3519 7517 3520
rect 6941 3491 7031 3497
rect 6941 3471 6957 3491
rect 6977 3489 7031 3491
rect 6977 3471 7002 3489
rect 6941 3469 7002 3471
rect 7022 3469 7031 3489
rect 6941 3463 7031 3469
rect 6954 3409 6991 3410
rect 7050 3409 7087 3410
rect 7106 3409 7142 3519
rect 7329 3498 7360 3519
rect 7675 3512 7678 3532
rect 7698 3512 8091 3532
rect 8275 3522 8309 3538
rect 8353 3590 8496 3611
rect 8891 3639 9324 3643
rect 8891 3633 9330 3639
rect 8891 3615 8912 3633
rect 8930 3615 9330 3633
rect 10124 3622 10155 3673
rect 10190 3702 10227 3772
rect 10493 3771 10530 3772
rect 10342 3712 10378 3713
rect 10190 3682 10199 3702
rect 10219 3682 10227 3702
rect 10190 3672 10227 3682
rect 10286 3702 10434 3712
rect 10534 3709 10630 3711
rect 10286 3682 10295 3702
rect 10315 3682 10405 3702
rect 10425 3682 10434 3702
rect 10286 3673 10434 3682
rect 10492 3702 10630 3709
rect 10492 3682 10501 3702
rect 10521 3682 10630 3702
rect 10492 3673 10630 3682
rect 10286 3672 10323 3673
rect 10016 3619 10057 3620
rect 8891 3597 9330 3615
rect 8051 3503 8091 3512
rect 8353 3503 8380 3590
rect 8453 3564 8496 3590
rect 8453 3546 8466 3564
rect 8484 3546 8496 3564
rect 8453 3535 8496 3546
rect 7325 3497 7360 3498
rect 7203 3487 7360 3497
rect 7203 3467 7220 3487
rect 7240 3467 7360 3487
rect 7203 3460 7360 3467
rect 7427 3490 7576 3498
rect 7427 3470 7438 3490
rect 7458 3470 7497 3490
rect 7517 3470 7576 3490
rect 8051 3486 8380 3503
rect 8051 3485 8091 3486
rect 7427 3463 7576 3470
rect 8448 3474 8488 3477
rect 8448 3468 8491 3474
rect 8073 3465 8491 3468
rect 7427 3462 7468 3463
rect 7161 3409 7198 3410
rect 6854 3400 6992 3409
rect 6854 3380 6963 3400
rect 6983 3380 6992 3400
rect 6854 3373 6992 3380
rect 7050 3400 7198 3409
rect 7050 3380 7059 3400
rect 7079 3380 7169 3400
rect 7189 3380 7198 3400
rect 6854 3371 6950 3373
rect 7050 3370 7198 3380
rect 7257 3400 7294 3410
rect 7257 3380 7265 3400
rect 7285 3380 7294 3400
rect 7106 3369 7142 3370
rect 6954 3310 6991 3311
rect 7257 3310 7294 3380
rect 7329 3409 7360 3460
rect 8073 3447 8464 3465
rect 8482 3447 8491 3465
rect 8073 3445 8491 3447
rect 8073 3437 8100 3445
rect 8341 3442 8491 3445
rect 7653 3431 7821 3432
rect 8072 3431 8100 3437
rect 7653 3415 8100 3431
rect 8448 3437 8491 3442
rect 7379 3409 7416 3410
rect 7329 3400 7416 3409
rect 7329 3380 7387 3400
rect 7407 3380 7416 3400
rect 7329 3370 7416 3380
rect 7475 3400 7512 3410
rect 7475 3380 7483 3400
rect 7503 3380 7512 3400
rect 7329 3369 7360 3370
rect 6953 3309 7294 3310
rect 7475 3309 7512 3380
rect 6878 3304 7294 3309
rect 6878 3284 6881 3304
rect 6901 3284 7294 3304
rect 7325 3285 7512 3309
rect 7653 3405 8097 3415
rect 7653 3403 7821 3405
rect 6720 3210 6749 3228
rect 7653 3225 7680 3403
rect 7720 3365 7784 3377
rect 8060 3373 8097 3405
rect 8123 3404 8314 3426
rect 8278 3402 8314 3404
rect 8278 3373 8315 3402
rect 8448 3381 8488 3437
rect 7720 3364 7755 3365
rect 7697 3359 7755 3364
rect 7697 3339 7700 3359
rect 7720 3345 7755 3359
rect 7775 3345 7784 3365
rect 7720 3337 7784 3345
rect 7746 3336 7784 3337
rect 7747 3335 7784 3336
rect 7850 3369 7886 3370
rect 7958 3369 7994 3370
rect 7850 3361 7994 3369
rect 7850 3341 7858 3361
rect 7878 3341 7913 3361
rect 7933 3341 7966 3361
rect 7986 3341 7994 3361
rect 7850 3335 7994 3341
rect 8060 3365 8098 3373
rect 8176 3369 8212 3370
rect 8060 3345 8069 3365
rect 8089 3345 8098 3365
rect 8060 3336 8098 3345
rect 8127 3361 8212 3369
rect 8127 3341 8184 3361
rect 8204 3341 8212 3361
rect 8060 3335 8097 3336
rect 8127 3335 8212 3341
rect 8278 3365 8316 3373
rect 8278 3345 8287 3365
rect 8307 3345 8316 3365
rect 8448 3363 8460 3381
rect 8478 3363 8488 3381
rect 8893 3408 8945 3597
rect 9291 3572 9330 3597
rect 9908 3612 10057 3619
rect 9908 3592 9967 3612
rect 9987 3592 10026 3612
rect 10046 3592 10057 3612
rect 9908 3584 10057 3592
rect 10124 3615 10281 3622
rect 10124 3595 10244 3615
rect 10264 3595 10281 3615
rect 10124 3585 10281 3595
rect 10124 3584 10159 3585
rect 9075 3547 9262 3571
rect 9291 3552 9686 3572
rect 9706 3552 9709 3572
rect 10124 3563 10155 3584
rect 10342 3563 10378 3673
rect 10397 3672 10434 3673
rect 10493 3672 10530 3673
rect 10453 3613 10543 3619
rect 10453 3593 10462 3613
rect 10482 3611 10543 3613
rect 10482 3593 10507 3611
rect 10453 3591 10507 3593
rect 10527 3591 10543 3611
rect 10453 3585 10543 3591
rect 9967 3562 10004 3563
rect 9291 3547 9709 3552
rect 9966 3553 10004 3562
rect 9075 3476 9112 3547
rect 9291 3546 9634 3547
rect 9291 3543 9330 3546
rect 9596 3545 9633 3546
rect 9227 3486 9258 3487
rect 9075 3456 9084 3476
rect 9104 3456 9112 3476
rect 9075 3446 9112 3456
rect 9171 3476 9258 3486
rect 9171 3456 9180 3476
rect 9200 3456 9258 3476
rect 9171 3447 9258 3456
rect 9171 3446 9208 3447
rect 8893 3390 8909 3408
rect 8927 3390 8945 3408
rect 9227 3396 9258 3447
rect 9293 3476 9330 3543
rect 9966 3533 9975 3553
rect 9995 3533 10004 3553
rect 9966 3525 10004 3533
rect 10070 3557 10155 3563
rect 10185 3562 10222 3563
rect 10070 3537 10078 3557
rect 10098 3537 10155 3557
rect 10070 3529 10155 3537
rect 10184 3553 10222 3562
rect 10184 3533 10193 3553
rect 10213 3533 10222 3553
rect 10070 3528 10106 3529
rect 10184 3525 10222 3533
rect 10288 3558 10432 3563
rect 10288 3557 10350 3558
rect 10288 3537 10296 3557
rect 10316 3539 10350 3557
rect 10371 3557 10432 3558
rect 10371 3539 10404 3557
rect 10316 3537 10404 3539
rect 10424 3537 10432 3557
rect 10288 3529 10432 3537
rect 10288 3528 10324 3529
rect 10396 3528 10432 3529
rect 10498 3562 10535 3563
rect 10498 3561 10536 3562
rect 10498 3553 10562 3561
rect 10498 3533 10507 3553
rect 10527 3539 10562 3553
rect 10582 3539 10585 3559
rect 10527 3534 10585 3539
rect 10527 3533 10562 3534
rect 9967 3496 10004 3525
rect 9968 3494 10004 3496
rect 9445 3486 9481 3487
rect 9293 3456 9302 3476
rect 9322 3456 9330 3476
rect 9293 3446 9330 3456
rect 9389 3476 9537 3486
rect 9637 3483 9733 3485
rect 9389 3456 9398 3476
rect 9418 3456 9508 3476
rect 9528 3456 9537 3476
rect 9389 3447 9537 3456
rect 9595 3476 9733 3483
rect 9595 3456 9604 3476
rect 9624 3456 9733 3476
rect 9968 3472 10159 3494
rect 10185 3493 10222 3525
rect 10498 3521 10562 3533
rect 10602 3495 10629 3673
rect 10461 3493 10629 3495
rect 10185 3479 10629 3493
rect 10185 3467 10632 3479
rect 10228 3465 10261 3467
rect 9595 3447 9733 3456
rect 9389 3446 9426 3447
rect 9119 3393 9160 3394
rect 8893 3372 8945 3390
rect 9011 3386 9160 3393
rect 8448 3353 8488 3363
rect 9011 3366 9070 3386
rect 9090 3366 9129 3386
rect 9149 3366 9160 3386
rect 9011 3358 9160 3366
rect 9227 3389 9384 3396
rect 9227 3369 9347 3389
rect 9367 3369 9384 3389
rect 9227 3359 9384 3369
rect 9227 3358 9262 3359
rect 8278 3336 8316 3345
rect 9227 3337 9258 3358
rect 9445 3337 9481 3447
rect 9500 3446 9537 3447
rect 9596 3446 9633 3447
rect 9556 3387 9646 3393
rect 9556 3367 9565 3387
rect 9585 3385 9646 3387
rect 9585 3367 9610 3385
rect 9556 3365 9610 3367
rect 9630 3365 9646 3385
rect 9556 3359 9646 3365
rect 9070 3336 9107 3337
rect 8278 3335 8315 3336
rect 7739 3307 7829 3313
rect 7739 3287 7755 3307
rect 7775 3305 7829 3307
rect 7775 3287 7800 3305
rect 7739 3285 7800 3287
rect 7820 3285 7829 3305
rect 7739 3279 7829 3285
rect 7752 3225 7789 3226
rect 7848 3225 7885 3226
rect 7904 3225 7940 3335
rect 8127 3314 8158 3335
rect 9069 3327 9107 3336
rect 8123 3313 8158 3314
rect 8001 3303 8158 3313
rect 8001 3283 8018 3303
rect 8038 3283 8158 3303
rect 8001 3276 8158 3283
rect 8225 3306 8374 3314
rect 8225 3286 8236 3306
rect 8256 3286 8295 3306
rect 8315 3286 8374 3306
rect 8897 3309 8937 3319
rect 8225 3279 8374 3286
rect 8440 3282 8492 3300
rect 8225 3278 8266 3279
rect 7959 3225 7996 3226
rect 6690 3208 6749 3210
rect 7652 3216 7790 3225
rect 6690 3207 6858 3208
rect 6984 3207 7024 3209
rect 6690 3181 7134 3207
rect 6690 3179 6858 3181
rect 6690 3177 6771 3179
rect 6690 3001 6717 3177
rect 6757 3141 6821 3153
rect 7097 3149 7134 3181
rect 7160 3180 7351 3202
rect 7652 3196 7761 3216
rect 7781 3196 7790 3216
rect 7652 3189 7790 3196
rect 7848 3216 7996 3225
rect 7848 3196 7857 3216
rect 7877 3196 7967 3216
rect 7987 3196 7996 3216
rect 7652 3187 7748 3189
rect 7848 3186 7996 3196
rect 8055 3216 8092 3226
rect 8055 3196 8063 3216
rect 8083 3196 8092 3216
rect 7904 3185 7940 3186
rect 7315 3178 7351 3180
rect 7315 3149 7352 3178
rect 6757 3140 6792 3141
rect 6734 3135 6792 3140
rect 6734 3115 6737 3135
rect 6757 3121 6792 3135
rect 6812 3121 6821 3141
rect 6757 3113 6821 3121
rect 6783 3112 6821 3113
rect 6784 3111 6821 3112
rect 6887 3145 6923 3146
rect 6995 3145 7031 3146
rect 6887 3137 7031 3145
rect 6887 3117 6895 3137
rect 6915 3136 7003 3137
rect 6915 3118 6950 3136
rect 6968 3118 7003 3136
rect 6915 3117 7003 3118
rect 7023 3117 7031 3137
rect 6887 3111 7031 3117
rect 7097 3141 7135 3149
rect 7213 3145 7249 3146
rect 7097 3121 7106 3141
rect 7126 3121 7135 3141
rect 7097 3112 7135 3121
rect 7164 3137 7249 3145
rect 7164 3117 7221 3137
rect 7241 3117 7249 3137
rect 7097 3111 7134 3112
rect 7164 3111 7249 3117
rect 7315 3141 7353 3149
rect 7315 3121 7324 3141
rect 7344 3121 7353 3141
rect 8055 3129 8092 3196
rect 8127 3225 8158 3276
rect 8440 3264 8458 3282
rect 8476 3264 8492 3282
rect 8177 3225 8214 3226
rect 8127 3216 8214 3225
rect 8127 3196 8185 3216
rect 8205 3196 8214 3216
rect 8127 3186 8214 3196
rect 8273 3216 8310 3226
rect 8273 3196 8281 3216
rect 8301 3196 8310 3216
rect 8127 3185 8158 3186
rect 7752 3126 7789 3127
rect 8055 3126 8094 3129
rect 7751 3125 8094 3126
rect 8273 3125 8310 3196
rect 7315 3112 7353 3121
rect 7676 3120 8094 3125
rect 7315 3111 7352 3112
rect 6776 3083 6866 3089
rect 6776 3063 6792 3083
rect 6812 3081 6866 3083
rect 6812 3063 6837 3081
rect 6776 3061 6837 3063
rect 6857 3061 6866 3081
rect 6776 3055 6866 3061
rect 6789 3001 6826 3002
rect 6885 3001 6922 3002
rect 6941 3001 6977 3111
rect 7164 3090 7195 3111
rect 7676 3100 7679 3120
rect 7699 3100 8094 3120
rect 8123 3101 8310 3125
rect 7160 3089 7195 3090
rect 7038 3079 7195 3089
rect 7038 3059 7055 3079
rect 7075 3059 7195 3079
rect 7038 3052 7195 3059
rect 7262 3082 7411 3090
rect 7262 3062 7273 3082
rect 7293 3062 7332 3082
rect 7352 3062 7411 3082
rect 7262 3055 7411 3062
rect 8055 3075 8094 3100
rect 8440 3075 8492 3264
rect 8897 3291 8907 3309
rect 8925 3291 8937 3309
rect 9069 3307 9078 3327
rect 9098 3307 9107 3327
rect 9069 3299 9107 3307
rect 9173 3331 9258 3337
rect 9288 3336 9325 3337
rect 9173 3311 9181 3331
rect 9201 3311 9258 3331
rect 9173 3303 9258 3311
rect 9287 3327 9325 3336
rect 9287 3307 9296 3327
rect 9316 3307 9325 3327
rect 9173 3302 9209 3303
rect 9287 3299 9325 3307
rect 9391 3331 9535 3337
rect 9391 3311 9399 3331
rect 9419 3311 9452 3331
rect 9472 3311 9507 3331
rect 9527 3311 9535 3331
rect 9391 3303 9535 3311
rect 9391 3302 9427 3303
rect 9499 3302 9535 3303
rect 9601 3336 9638 3337
rect 9601 3335 9639 3336
rect 9601 3327 9665 3335
rect 9601 3307 9610 3327
rect 9630 3313 9665 3327
rect 9685 3313 9688 3333
rect 9630 3308 9688 3313
rect 9630 3307 9665 3308
rect 8897 3235 8937 3291
rect 9070 3270 9107 3299
rect 9071 3268 9107 3270
rect 9071 3246 9262 3268
rect 9288 3267 9325 3299
rect 9601 3295 9665 3307
rect 9705 3269 9732 3447
rect 10590 3422 10632 3467
rect 9564 3267 9732 3269
rect 9288 3257 9732 3267
rect 9873 3363 10060 3387
rect 10091 3368 10484 3388
rect 10504 3368 10507 3388
rect 10091 3363 10507 3368
rect 9873 3292 9910 3363
rect 10091 3362 10432 3363
rect 10025 3302 10056 3303
rect 9873 3272 9882 3292
rect 9902 3272 9910 3292
rect 9873 3262 9910 3272
rect 9969 3292 10056 3302
rect 9969 3272 9978 3292
rect 9998 3272 10056 3292
rect 9969 3263 10056 3272
rect 9969 3262 10006 3263
rect 8894 3230 8937 3235
rect 9285 3241 9732 3257
rect 9285 3235 9313 3241
rect 9564 3240 9732 3241
rect 8894 3227 9044 3230
rect 9285 3227 9312 3235
rect 8894 3225 9312 3227
rect 8894 3207 8903 3225
rect 8921 3207 9312 3225
rect 10025 3212 10056 3263
rect 10091 3292 10128 3362
rect 10394 3361 10431 3362
rect 10243 3302 10279 3303
rect 10091 3272 10100 3292
rect 10120 3272 10128 3292
rect 10091 3262 10128 3272
rect 10187 3292 10335 3302
rect 10435 3299 10531 3301
rect 10187 3272 10196 3292
rect 10216 3272 10306 3292
rect 10326 3272 10335 3292
rect 10187 3263 10335 3272
rect 10393 3292 10531 3299
rect 10393 3272 10402 3292
rect 10422 3272 10531 3292
rect 10393 3263 10531 3272
rect 10187 3262 10224 3263
rect 9917 3209 9958 3210
rect 8894 3204 9312 3207
rect 8894 3198 8937 3204
rect 8897 3195 8937 3198
rect 9812 3202 9958 3209
rect 9294 3186 9334 3187
rect 9005 3169 9334 3186
rect 9812 3182 9868 3202
rect 9888 3182 9927 3202
rect 9947 3182 9958 3202
rect 9812 3174 9958 3182
rect 10025 3205 10182 3212
rect 10025 3185 10145 3205
rect 10165 3185 10182 3205
rect 10025 3175 10182 3185
rect 10025 3174 10060 3175
rect 8889 3126 8932 3137
rect 8889 3108 8901 3126
rect 8919 3108 8932 3126
rect 8889 3082 8932 3108
rect 9005 3082 9032 3169
rect 9294 3160 9334 3169
rect 8055 3057 8494 3075
rect 7262 3054 7303 3055
rect 6996 3001 7033 3002
rect 6689 2992 6827 3001
rect 6689 2972 6798 2992
rect 6818 2972 6827 2992
rect 6689 2965 6827 2972
rect 6885 2992 7033 3001
rect 6885 2972 6894 2992
rect 6914 2972 7004 2992
rect 7024 2972 7033 2992
rect 6689 2963 6785 2965
rect 6885 2962 7033 2972
rect 7092 2992 7129 3002
rect 7092 2972 7100 2992
rect 7120 2972 7129 2992
rect 6941 2961 6977 2962
rect 6789 2902 6826 2903
rect 7092 2902 7129 2972
rect 7164 3001 7195 3052
rect 8055 3039 8455 3057
rect 8473 3039 8494 3057
rect 8055 3033 8494 3039
rect 8061 3029 8494 3033
rect 8889 3061 9032 3082
rect 9076 3134 9110 3150
rect 9294 3140 9687 3160
rect 9707 3140 9710 3160
rect 10025 3153 10056 3174
rect 10243 3153 10279 3263
rect 10298 3262 10335 3263
rect 10394 3262 10431 3263
rect 10354 3203 10444 3209
rect 10354 3183 10363 3203
rect 10383 3201 10444 3203
rect 10383 3183 10408 3201
rect 10354 3181 10408 3183
rect 10428 3181 10444 3201
rect 10354 3175 10444 3181
rect 9868 3152 9905 3153
rect 9294 3135 9710 3140
rect 9867 3143 9905 3152
rect 9294 3134 9635 3135
rect 9076 3064 9113 3134
rect 9228 3074 9259 3075
rect 8889 3059 9026 3061
rect 8440 3027 8492 3029
rect 8889 3017 8932 3059
rect 9076 3044 9085 3064
rect 9105 3044 9113 3064
rect 9076 3034 9113 3044
rect 9172 3064 9259 3074
rect 9172 3044 9181 3064
rect 9201 3044 9259 3064
rect 9172 3035 9259 3044
rect 9172 3034 9209 3035
rect 8887 3007 8932 3017
rect 7214 3001 7251 3002
rect 7164 2992 7251 3001
rect 7164 2972 7222 2992
rect 7242 2972 7251 2992
rect 7164 2962 7251 2972
rect 7310 2992 7347 3002
rect 7310 2972 7318 2992
rect 7338 2972 7347 2992
rect 8887 2989 8896 3007
rect 8914 2989 8932 3007
rect 8887 2983 8932 2989
rect 9228 2984 9259 3035
rect 9294 3064 9331 3134
rect 9597 3133 9634 3134
rect 9867 3123 9876 3143
rect 9896 3123 9905 3143
rect 9867 3115 9905 3123
rect 9971 3147 10056 3153
rect 10086 3152 10123 3153
rect 9971 3127 9979 3147
rect 9999 3127 10056 3147
rect 9971 3119 10056 3127
rect 10085 3143 10123 3152
rect 10085 3123 10094 3143
rect 10114 3123 10123 3143
rect 9971 3118 10007 3119
rect 10085 3115 10123 3123
rect 10189 3147 10333 3153
rect 10189 3127 10197 3147
rect 10217 3144 10305 3147
rect 10217 3127 10252 3144
rect 10189 3126 10252 3127
rect 10271 3127 10305 3144
rect 10325 3127 10333 3147
rect 10271 3126 10333 3127
rect 10189 3119 10333 3126
rect 10189 3118 10225 3119
rect 10297 3118 10333 3119
rect 10399 3152 10436 3153
rect 10399 3151 10437 3152
rect 10459 3151 10486 3155
rect 10399 3149 10486 3151
rect 10399 3143 10463 3149
rect 10399 3123 10408 3143
rect 10428 3129 10463 3143
rect 10483 3129 10486 3149
rect 10428 3124 10486 3129
rect 10428 3123 10463 3124
rect 9868 3086 9905 3115
rect 9869 3084 9905 3086
rect 9446 3074 9482 3075
rect 9294 3044 9303 3064
rect 9323 3044 9331 3064
rect 9294 3034 9331 3044
rect 9390 3064 9538 3074
rect 9638 3071 9734 3073
rect 9390 3044 9399 3064
rect 9419 3044 9509 3064
rect 9529 3044 9538 3064
rect 9390 3035 9538 3044
rect 9596 3064 9734 3071
rect 9596 3044 9605 3064
rect 9625 3044 9734 3064
rect 9869 3062 10060 3084
rect 10086 3083 10123 3115
rect 10399 3111 10463 3123
rect 10503 3085 10530 3263
rect 10362 3083 10530 3085
rect 10086 3057 10530 3083
rect 9596 3035 9734 3044
rect 9390 3034 9427 3035
rect 8887 2980 8924 2983
rect 9120 2981 9161 2982
rect 7164 2961 7195 2962
rect 6788 2901 7129 2902
rect 7310 2901 7347 2972
rect 9012 2974 9161 2981
rect 8443 2962 8480 2967
rect 6713 2896 7129 2901
rect 6713 2876 6716 2896
rect 6736 2876 7129 2896
rect 7160 2877 7347 2901
rect 8434 2958 8481 2962
rect 8434 2940 8453 2958
rect 8471 2940 8481 2958
rect 9012 2954 9071 2974
rect 9091 2954 9130 2974
rect 9150 2954 9161 2974
rect 9012 2946 9161 2954
rect 9228 2977 9385 2984
rect 9228 2957 9348 2977
rect 9368 2957 9385 2977
rect 9228 2947 9385 2957
rect 9228 2946 9263 2947
rect 8434 2892 8481 2940
rect 9228 2925 9259 2946
rect 9446 2925 9482 3035
rect 9501 3034 9538 3035
rect 9597 3034 9634 3035
rect 9557 2975 9647 2981
rect 9557 2955 9566 2975
rect 9586 2973 9647 2975
rect 9586 2955 9611 2973
rect 9557 2953 9611 2955
rect 9631 2953 9647 2973
rect 9557 2947 9647 2953
rect 9071 2924 9108 2925
rect 8058 2889 8481 2892
rect 6933 2875 6998 2876
rect 8036 2859 8481 2889
rect 8883 2916 8921 2918
rect 8883 2908 8926 2916
rect 8883 2890 8894 2908
rect 8912 2890 8926 2908
rect 8883 2863 8926 2890
rect 9070 2915 9108 2924
rect 9070 2895 9079 2915
rect 9099 2895 9108 2915
rect 9070 2887 9108 2895
rect 9174 2919 9259 2925
rect 9289 2924 9326 2925
rect 9174 2899 9182 2919
rect 9202 2899 9259 2919
rect 9174 2891 9259 2899
rect 9288 2915 9326 2924
rect 9288 2895 9297 2915
rect 9317 2895 9326 2915
rect 9174 2890 9210 2891
rect 9288 2887 9326 2895
rect 9392 2923 9536 2925
rect 9392 2919 9444 2923
rect 9392 2899 9400 2919
rect 9420 2903 9444 2919
rect 9464 2919 9536 2923
rect 9464 2903 9508 2919
rect 9420 2899 9508 2903
rect 9528 2899 9536 2919
rect 9392 2891 9536 2899
rect 9392 2890 9428 2891
rect 9500 2890 9536 2891
rect 9602 2924 9639 2925
rect 9602 2923 9640 2924
rect 9602 2915 9666 2923
rect 9602 2895 9611 2915
rect 9631 2901 9666 2915
rect 9686 2901 9689 2921
rect 9631 2896 9689 2901
rect 9631 2895 9666 2896
rect 7129 2843 7169 2851
rect 7129 2821 7137 2843
rect 7161 2821 7169 2843
rect 6734 2592 6771 2598
rect 6734 2573 6742 2592
rect 6763 2573 6771 2592
rect 6734 2565 6771 2573
rect 6434 2444 6441 2466
rect 6465 2444 6473 2466
rect 6434 2438 6473 2444
rect 5964 2433 6004 2435
rect 6130 2434 6298 2435
rect 6232 2433 6269 2434
rect 5198 2417 5336 2426
rect 4992 2416 5029 2417
rect 4722 2363 4763 2364
rect 4496 2342 4548 2360
rect 4614 2356 4763 2363
rect 4064 2322 4104 2332
rect 4614 2336 4673 2356
rect 4693 2336 4732 2356
rect 4752 2336 4763 2356
rect 4614 2328 4763 2336
rect 4830 2359 4987 2366
rect 4830 2339 4950 2359
rect 4970 2339 4987 2359
rect 4830 2329 4987 2339
rect 4830 2328 4865 2329
rect 3894 2305 3932 2314
rect 4830 2307 4861 2328
rect 5048 2307 5084 2417
rect 5103 2416 5140 2417
rect 5199 2416 5236 2417
rect 5159 2357 5249 2363
rect 5159 2337 5168 2357
rect 5188 2355 5249 2357
rect 5188 2337 5213 2355
rect 5159 2335 5213 2337
rect 5233 2335 5249 2355
rect 5159 2329 5249 2335
rect 4673 2306 4710 2307
rect 3894 2304 3931 2305
rect 3355 2276 3445 2282
rect 3355 2256 3371 2276
rect 3391 2274 3445 2276
rect 3391 2256 3416 2274
rect 3355 2254 3416 2256
rect 3436 2254 3445 2274
rect 3355 2248 3445 2254
rect 3368 2194 3405 2195
rect 3464 2194 3501 2195
rect 3520 2194 3556 2304
rect 3743 2283 3774 2304
rect 4672 2297 4710 2306
rect 3739 2282 3774 2283
rect 3617 2272 3774 2282
rect 3617 2252 3634 2272
rect 3654 2252 3774 2272
rect 3617 2245 3774 2252
rect 3841 2275 3990 2283
rect 3841 2255 3852 2275
rect 3872 2255 3911 2275
rect 3931 2255 3990 2275
rect 4500 2279 4540 2289
rect 3841 2248 3990 2255
rect 4056 2251 4108 2269
rect 3841 2247 3882 2248
rect 3575 2194 3612 2195
rect 3268 2185 3406 2194
rect 2740 2174 2773 2176
rect 2369 2162 2816 2174
rect 1601 2040 1769 2042
rect 1325 2014 1769 2040
rect 835 1992 973 2001
rect 629 1991 666 1992
rect 126 1937 163 1940
rect 359 1938 400 1939
rect 251 1931 400 1938
rect 251 1911 310 1931
rect 330 1911 369 1931
rect 389 1911 400 1931
rect 251 1903 400 1911
rect 467 1934 624 1941
rect 467 1914 587 1934
rect 607 1914 624 1934
rect 467 1904 624 1914
rect 467 1903 502 1904
rect 467 1882 498 1903
rect 685 1882 721 1992
rect 740 1991 777 1992
rect 836 1991 873 1992
rect 796 1932 886 1938
rect 796 1912 805 1932
rect 825 1930 886 1932
rect 825 1912 850 1930
rect 796 1910 850 1912
rect 870 1910 886 1930
rect 796 1904 886 1910
rect 310 1881 347 1882
rect 123 1873 160 1875
rect 123 1865 165 1873
rect 123 1847 133 1865
rect 151 1847 165 1865
rect 123 1838 165 1847
rect 309 1872 347 1881
rect 309 1852 318 1872
rect 338 1852 347 1872
rect 309 1844 347 1852
rect 413 1876 498 1882
rect 528 1881 565 1882
rect 413 1856 421 1876
rect 441 1856 498 1876
rect 413 1848 498 1856
rect 527 1872 565 1881
rect 527 1852 536 1872
rect 556 1852 565 1872
rect 413 1847 449 1848
rect 527 1844 565 1852
rect 631 1880 775 1882
rect 631 1876 683 1880
rect 631 1856 639 1876
rect 659 1860 683 1876
rect 703 1876 775 1880
rect 703 1860 747 1876
rect 659 1856 747 1860
rect 767 1856 775 1876
rect 631 1848 775 1856
rect 631 1847 667 1848
rect 739 1847 775 1848
rect 841 1881 878 1882
rect 841 1880 879 1881
rect 841 1872 905 1880
rect 841 1852 850 1872
rect 870 1858 905 1872
rect 925 1858 928 1878
rect 870 1853 928 1858
rect 870 1852 905 1853
rect 124 1813 165 1838
rect 310 1813 347 1844
rect 528 1813 565 1844
rect 841 1840 905 1852
rect 945 1814 972 1992
rect 124 1786 173 1813
rect 309 1787 358 1813
rect 527 1812 608 1813
rect 804 1812 972 1814
rect 527 1787 972 1812
rect 528 1786 972 1787
rect 126 1753 173 1786
rect 529 1753 569 1786
rect 804 1785 972 1786
rect 1435 1790 1475 2014
rect 1601 2013 1769 2014
rect 2372 2148 2816 2162
rect 2372 2146 2540 2148
rect 2372 1968 2399 2146
rect 2439 2108 2503 2120
rect 2779 2116 2816 2148
rect 2842 2147 3033 2169
rect 3268 2165 3377 2185
rect 3397 2165 3406 2185
rect 3268 2158 3406 2165
rect 3464 2185 3612 2194
rect 3464 2165 3473 2185
rect 3493 2165 3583 2185
rect 3603 2165 3612 2185
rect 3268 2156 3364 2158
rect 3464 2155 3612 2165
rect 3671 2185 3708 2195
rect 3671 2165 3679 2185
rect 3699 2165 3708 2185
rect 3520 2154 3556 2155
rect 2997 2145 3033 2147
rect 2997 2116 3034 2145
rect 2439 2107 2474 2108
rect 2416 2102 2474 2107
rect 2416 2082 2419 2102
rect 2439 2088 2474 2102
rect 2494 2088 2503 2108
rect 2439 2080 2503 2088
rect 2465 2079 2503 2080
rect 2466 2078 2503 2079
rect 2569 2112 2605 2113
rect 2677 2112 2713 2113
rect 2569 2104 2713 2112
rect 2569 2084 2577 2104
rect 2597 2102 2685 2104
rect 2597 2084 2630 2102
rect 2569 2083 2630 2084
rect 2651 2084 2685 2102
rect 2705 2084 2713 2104
rect 2651 2083 2713 2084
rect 2569 2078 2713 2083
rect 2779 2108 2817 2116
rect 2895 2112 2931 2113
rect 2779 2088 2788 2108
rect 2808 2088 2817 2108
rect 2779 2079 2817 2088
rect 2846 2104 2931 2112
rect 2846 2084 2903 2104
rect 2923 2084 2931 2104
rect 2779 2078 2816 2079
rect 2846 2078 2931 2084
rect 2997 2108 3035 2116
rect 2997 2088 3006 2108
rect 3026 2088 3035 2108
rect 3671 2098 3708 2165
rect 3743 2194 3774 2245
rect 4056 2233 4074 2251
rect 4092 2233 4108 2251
rect 3793 2194 3830 2195
rect 3743 2185 3830 2194
rect 3743 2165 3801 2185
rect 3821 2165 3830 2185
rect 3743 2155 3830 2165
rect 3889 2185 3926 2195
rect 3889 2165 3897 2185
rect 3917 2165 3926 2185
rect 3743 2154 3774 2155
rect 3368 2095 3405 2096
rect 3671 2095 3710 2098
rect 3367 2094 3710 2095
rect 3889 2094 3926 2165
rect 2997 2079 3035 2088
rect 3292 2089 3710 2094
rect 2997 2078 3034 2079
rect 2458 2050 2548 2056
rect 2458 2030 2474 2050
rect 2494 2048 2548 2050
rect 2494 2030 2519 2048
rect 2458 2028 2519 2030
rect 2539 2028 2548 2048
rect 2458 2022 2548 2028
rect 2471 1968 2508 1969
rect 2567 1968 2604 1969
rect 2623 1968 2659 2078
rect 2846 2057 2877 2078
rect 3292 2069 3295 2089
rect 3315 2069 3710 2089
rect 3739 2070 3926 2094
rect 2842 2056 2877 2057
rect 2720 2046 2877 2056
rect 2720 2026 2737 2046
rect 2757 2026 2877 2046
rect 2720 2019 2877 2026
rect 2944 2049 3093 2057
rect 2944 2029 2955 2049
rect 2975 2029 3014 2049
rect 3034 2029 3093 2049
rect 2944 2022 3093 2029
rect 3671 2044 3710 2069
rect 4056 2044 4108 2233
rect 4500 2261 4510 2279
rect 4528 2261 4540 2279
rect 4672 2277 4681 2297
rect 4701 2277 4710 2297
rect 4672 2269 4710 2277
rect 4776 2301 4861 2307
rect 4891 2306 4928 2307
rect 4776 2281 4784 2301
rect 4804 2281 4861 2301
rect 4776 2273 4861 2281
rect 4890 2297 4928 2306
rect 4890 2277 4899 2297
rect 4919 2277 4928 2297
rect 4776 2272 4812 2273
rect 4890 2269 4928 2277
rect 4994 2301 5138 2307
rect 4994 2281 5002 2301
rect 5022 2281 5055 2301
rect 5075 2281 5110 2301
rect 5130 2281 5138 2301
rect 4994 2273 5138 2281
rect 4994 2272 5030 2273
rect 5102 2272 5138 2273
rect 5204 2306 5241 2307
rect 5204 2305 5242 2306
rect 5204 2297 5268 2305
rect 5204 2277 5213 2297
rect 5233 2283 5268 2297
rect 5288 2283 5291 2303
rect 5233 2278 5291 2283
rect 5233 2277 5268 2278
rect 4500 2205 4540 2261
rect 4673 2240 4710 2269
rect 4674 2238 4710 2240
rect 4674 2216 4865 2238
rect 4891 2237 4928 2269
rect 5204 2265 5268 2277
rect 5308 2239 5335 2417
rect 5167 2237 5335 2239
rect 4891 2227 5335 2237
rect 5476 2333 5663 2357
rect 5694 2338 6087 2358
rect 6107 2338 6110 2358
rect 5694 2333 6110 2338
rect 5476 2262 5513 2333
rect 5694 2332 6035 2333
rect 5628 2272 5659 2273
rect 5476 2242 5485 2262
rect 5505 2242 5513 2262
rect 5476 2232 5513 2242
rect 5572 2262 5659 2272
rect 5572 2242 5581 2262
rect 5601 2242 5659 2262
rect 5572 2233 5659 2242
rect 5572 2232 5609 2233
rect 4497 2200 4540 2205
rect 4888 2211 5335 2227
rect 4888 2205 4916 2211
rect 5167 2210 5335 2211
rect 4497 2197 4647 2200
rect 4888 2197 4915 2205
rect 4497 2195 4915 2197
rect 4497 2177 4506 2195
rect 4524 2177 4915 2195
rect 5628 2182 5659 2233
rect 5694 2262 5731 2332
rect 5997 2331 6034 2332
rect 6235 2274 6268 2433
rect 5846 2272 5882 2273
rect 5694 2242 5703 2262
rect 5723 2242 5731 2262
rect 5694 2232 5731 2242
rect 5790 2262 5938 2272
rect 6038 2269 6134 2271
rect 5790 2242 5799 2262
rect 5819 2242 5909 2262
rect 5929 2242 5938 2262
rect 5790 2233 5938 2242
rect 5996 2262 6134 2269
rect 5996 2242 6005 2262
rect 6025 2242 6134 2262
rect 6235 2270 6271 2274
rect 6235 2252 6244 2270
rect 6266 2252 6271 2270
rect 6235 2246 6271 2252
rect 5996 2233 6134 2242
rect 5790 2232 5827 2233
rect 5520 2179 5561 2180
rect 4497 2174 4915 2177
rect 4497 2168 4540 2174
rect 4500 2165 4540 2168
rect 5412 2172 5561 2179
rect 4897 2156 4937 2157
rect 4608 2139 4937 2156
rect 5412 2152 5471 2172
rect 5491 2152 5530 2172
rect 5550 2152 5561 2172
rect 5412 2144 5561 2152
rect 5628 2175 5785 2182
rect 5628 2155 5748 2175
rect 5768 2155 5785 2175
rect 5628 2145 5785 2155
rect 5628 2144 5663 2145
rect 4492 2096 4535 2107
rect 4492 2078 4504 2096
rect 4522 2078 4535 2096
rect 4492 2052 4535 2078
rect 4608 2052 4635 2139
rect 4897 2130 4937 2139
rect 3671 2026 4110 2044
rect 2944 2021 2985 2022
rect 2678 1968 2715 1969
rect 2371 1959 2509 1968
rect 2371 1939 2480 1959
rect 2500 1939 2509 1959
rect 2371 1932 2509 1939
rect 2567 1959 2715 1968
rect 2567 1939 2576 1959
rect 2596 1939 2686 1959
rect 2706 1939 2715 1959
rect 2371 1930 2467 1932
rect 2567 1929 2715 1939
rect 2774 1959 2811 1969
rect 2774 1939 2782 1959
rect 2802 1939 2811 1959
rect 2623 1928 2659 1929
rect 2471 1869 2508 1870
rect 2774 1869 2811 1939
rect 2846 1968 2877 2019
rect 3671 2008 4071 2026
rect 4089 2008 4110 2026
rect 3671 2002 4110 2008
rect 3677 1998 4110 2002
rect 4492 2031 4635 2052
rect 4679 2104 4713 2120
rect 4897 2110 5290 2130
rect 5310 2110 5313 2130
rect 5628 2123 5659 2144
rect 5846 2123 5882 2233
rect 5901 2232 5938 2233
rect 5997 2232 6034 2233
rect 5957 2173 6047 2179
rect 5957 2153 5966 2173
rect 5986 2171 6047 2173
rect 5986 2153 6011 2171
rect 5957 2151 6011 2153
rect 6031 2151 6047 2171
rect 5957 2145 6047 2151
rect 5471 2122 5508 2123
rect 4897 2105 5313 2110
rect 5470 2113 5508 2122
rect 4897 2104 5238 2105
rect 4679 2034 4716 2104
rect 4831 2044 4862 2045
rect 4492 2029 4629 2031
rect 4056 1996 4108 1998
rect 4492 1987 4535 2029
rect 4679 2014 4688 2034
rect 4708 2014 4716 2034
rect 4679 2004 4716 2014
rect 4775 2034 4862 2044
rect 4775 2014 4784 2034
rect 4804 2014 4862 2034
rect 4775 2005 4862 2014
rect 4775 2004 4812 2005
rect 4490 1977 4535 1987
rect 2896 1968 2933 1969
rect 2846 1959 2933 1968
rect 2846 1939 2904 1959
rect 2924 1939 2933 1959
rect 2846 1929 2933 1939
rect 2992 1959 3029 1969
rect 2992 1939 3000 1959
rect 3020 1939 3029 1959
rect 4490 1959 4499 1977
rect 4517 1959 4535 1977
rect 4490 1953 4535 1959
rect 4831 1954 4862 2005
rect 4897 2034 4934 2104
rect 5200 2103 5237 2104
rect 5470 2093 5479 2113
rect 5499 2093 5508 2113
rect 5470 2085 5508 2093
rect 5574 2117 5659 2123
rect 5689 2122 5726 2123
rect 5574 2097 5582 2117
rect 5602 2097 5659 2117
rect 5574 2089 5659 2097
rect 5688 2113 5726 2122
rect 5688 2093 5697 2113
rect 5717 2093 5726 2113
rect 5574 2088 5610 2089
rect 5688 2085 5726 2093
rect 5792 2117 5936 2123
rect 5792 2097 5800 2117
rect 5820 2098 5852 2117
rect 5873 2098 5908 2117
rect 5820 2097 5908 2098
rect 5928 2097 5936 2117
rect 5792 2089 5936 2097
rect 5792 2088 5828 2089
rect 5900 2088 5936 2089
rect 6002 2122 6039 2123
rect 6002 2121 6040 2122
rect 6002 2113 6066 2121
rect 6002 2093 6011 2113
rect 6031 2099 6066 2113
rect 6086 2099 6089 2119
rect 6031 2094 6089 2099
rect 6031 2093 6066 2094
rect 5471 2056 5508 2085
rect 5472 2054 5508 2056
rect 5049 2044 5085 2045
rect 4897 2014 4906 2034
rect 4926 2014 4934 2034
rect 4897 2004 4934 2014
rect 4993 2034 5141 2044
rect 5241 2041 5337 2043
rect 4993 2014 5002 2034
rect 5022 2014 5112 2034
rect 5132 2014 5141 2034
rect 4993 2005 5141 2014
rect 5199 2034 5337 2041
rect 5199 2014 5208 2034
rect 5228 2014 5337 2034
rect 5472 2032 5663 2054
rect 5689 2053 5726 2085
rect 6002 2081 6066 2093
rect 6106 2055 6133 2233
rect 6738 2232 6771 2565
rect 6835 2597 7003 2598
rect 7129 2597 7169 2821
rect 7632 2825 7800 2826
rect 8036 2825 8077 2859
rect 8434 2838 8481 2859
rect 7632 2815 8077 2825
rect 8149 2823 8292 2824
rect 7632 2799 8076 2815
rect 7632 2797 7800 2799
rect 7996 2798 8076 2799
rect 8149 2798 8294 2823
rect 8436 2798 8481 2838
rect 7632 2619 7659 2797
rect 7699 2759 7763 2771
rect 8039 2767 8076 2798
rect 8257 2767 8294 2798
rect 8439 2791 8481 2798
rect 8884 2856 8926 2863
rect 9071 2856 9108 2887
rect 9289 2856 9326 2887
rect 9602 2883 9666 2895
rect 9706 2857 9733 3035
rect 8884 2816 8929 2856
rect 9071 2831 9216 2856
rect 9289 2855 9369 2856
rect 9565 2855 9733 2857
rect 9289 2839 9733 2855
rect 9073 2830 9216 2831
rect 9288 2829 9733 2839
rect 8884 2795 8931 2816
rect 9288 2795 9329 2829
rect 9565 2828 9733 2829
rect 10196 2833 10236 3057
rect 10362 3056 10530 3057
rect 10594 3089 10627 3422
rect 10594 3081 10631 3089
rect 10594 3062 10602 3081
rect 10623 3062 10631 3081
rect 10594 3056 10631 3062
rect 10196 2811 10204 2833
rect 10228 2811 10236 2833
rect 10196 2803 10236 2811
rect 7699 2758 7734 2759
rect 7676 2753 7734 2758
rect 7676 2733 7679 2753
rect 7699 2739 7734 2753
rect 7754 2739 7763 2759
rect 7699 2731 7763 2739
rect 7725 2730 7763 2731
rect 7726 2729 7763 2730
rect 7829 2763 7865 2764
rect 7937 2763 7973 2764
rect 7829 2755 7973 2763
rect 7829 2735 7837 2755
rect 7857 2751 7945 2755
rect 7857 2735 7901 2751
rect 7829 2731 7901 2735
rect 7921 2735 7945 2751
rect 7965 2735 7973 2755
rect 7921 2731 7973 2735
rect 7829 2729 7973 2731
rect 8039 2759 8077 2767
rect 8155 2763 8191 2764
rect 8039 2739 8048 2759
rect 8068 2739 8077 2759
rect 8039 2730 8077 2739
rect 8106 2755 8191 2763
rect 8106 2735 8163 2755
rect 8183 2735 8191 2755
rect 8039 2729 8076 2730
rect 8106 2729 8191 2735
rect 8257 2759 8295 2767
rect 8257 2739 8266 2759
rect 8286 2739 8295 2759
rect 8257 2730 8295 2739
rect 8439 2764 8482 2791
rect 8439 2746 8453 2764
rect 8471 2746 8482 2764
rect 8439 2738 8482 2746
rect 8444 2736 8482 2738
rect 8884 2765 9329 2795
rect 10367 2778 10432 2779
rect 8884 2762 9307 2765
rect 8257 2729 8294 2730
rect 7718 2701 7808 2707
rect 7718 2681 7734 2701
rect 7754 2699 7808 2701
rect 7754 2681 7779 2699
rect 7718 2679 7779 2681
rect 7799 2679 7808 2699
rect 7718 2673 7808 2679
rect 7731 2619 7768 2620
rect 7827 2619 7864 2620
rect 7883 2619 7919 2729
rect 8106 2708 8137 2729
rect 8884 2714 8931 2762
rect 8102 2707 8137 2708
rect 7980 2697 8137 2707
rect 7980 2677 7997 2697
rect 8017 2677 8137 2697
rect 7980 2670 8137 2677
rect 8204 2700 8353 2708
rect 8204 2680 8215 2700
rect 8235 2680 8274 2700
rect 8294 2680 8353 2700
rect 8884 2696 8894 2714
rect 8912 2696 8931 2714
rect 8884 2692 8931 2696
rect 10018 2753 10205 2777
rect 10236 2758 10629 2778
rect 10649 2758 10652 2778
rect 10236 2753 10652 2758
rect 8885 2687 8922 2692
rect 8204 2673 8353 2680
rect 10018 2682 10055 2753
rect 10236 2752 10577 2753
rect 10170 2692 10201 2693
rect 8204 2672 8245 2673
rect 8441 2671 8478 2674
rect 7938 2619 7975 2620
rect 7631 2610 7769 2619
rect 6835 2571 7279 2597
rect 6835 2569 7003 2571
rect 6835 2391 6862 2569
rect 6902 2531 6966 2543
rect 7242 2539 7279 2571
rect 7305 2570 7496 2592
rect 7631 2590 7740 2610
rect 7760 2590 7769 2610
rect 7631 2583 7769 2590
rect 7827 2610 7975 2619
rect 7827 2590 7836 2610
rect 7856 2590 7946 2610
rect 7966 2590 7975 2610
rect 7631 2581 7727 2583
rect 7827 2580 7975 2590
rect 8034 2610 8071 2620
rect 8034 2590 8042 2610
rect 8062 2590 8071 2610
rect 7883 2579 7919 2580
rect 7460 2568 7496 2570
rect 7460 2539 7497 2568
rect 6902 2530 6937 2531
rect 6879 2525 6937 2530
rect 6879 2505 6882 2525
rect 6902 2511 6937 2525
rect 6957 2511 6966 2531
rect 6902 2505 6966 2511
rect 6879 2503 6966 2505
rect 6879 2499 6906 2503
rect 6928 2502 6966 2503
rect 6929 2501 6966 2502
rect 7032 2535 7068 2536
rect 7140 2535 7176 2536
rect 7032 2528 7176 2535
rect 7032 2527 7094 2528
rect 7032 2507 7040 2527
rect 7060 2510 7094 2527
rect 7113 2527 7176 2528
rect 7113 2510 7148 2527
rect 7060 2507 7148 2510
rect 7168 2507 7176 2527
rect 7032 2501 7176 2507
rect 7242 2531 7280 2539
rect 7358 2535 7394 2536
rect 7242 2511 7251 2531
rect 7271 2511 7280 2531
rect 7242 2502 7280 2511
rect 7309 2527 7394 2535
rect 7309 2507 7366 2527
rect 7386 2507 7394 2527
rect 7242 2501 7279 2502
rect 7309 2501 7394 2507
rect 7460 2531 7498 2539
rect 7460 2511 7469 2531
rect 7489 2511 7498 2531
rect 7731 2520 7768 2521
rect 8034 2520 8071 2590
rect 8106 2619 8137 2670
rect 8433 2665 8478 2671
rect 8433 2647 8451 2665
rect 8469 2647 8478 2665
rect 10018 2662 10027 2682
rect 10047 2662 10055 2682
rect 10018 2652 10055 2662
rect 10114 2682 10201 2692
rect 10114 2662 10123 2682
rect 10143 2662 10201 2682
rect 10114 2653 10201 2662
rect 10114 2652 10151 2653
rect 8433 2637 8478 2647
rect 8156 2619 8193 2620
rect 8106 2610 8193 2619
rect 8106 2590 8164 2610
rect 8184 2590 8193 2610
rect 8106 2580 8193 2590
rect 8252 2610 8289 2620
rect 8252 2590 8260 2610
rect 8280 2590 8289 2610
rect 8433 2595 8476 2637
rect 8873 2625 8925 2627
rect 8339 2593 8476 2595
rect 8106 2579 8137 2580
rect 8252 2520 8289 2590
rect 7730 2519 8071 2520
rect 7460 2502 7498 2511
rect 7655 2514 8071 2519
rect 7460 2501 7497 2502
rect 6921 2473 7011 2479
rect 6921 2453 6937 2473
rect 6957 2471 7011 2473
rect 6957 2453 6982 2471
rect 6921 2451 6982 2453
rect 7002 2451 7011 2471
rect 6921 2445 7011 2451
rect 6934 2391 6971 2392
rect 7030 2391 7067 2392
rect 7086 2391 7122 2501
rect 7309 2480 7340 2501
rect 7655 2494 7658 2514
rect 7678 2494 8071 2514
rect 8255 2504 8289 2520
rect 8333 2572 8476 2593
rect 8871 2621 9304 2625
rect 8871 2615 9310 2621
rect 8871 2597 8892 2615
rect 8910 2597 9310 2615
rect 10170 2602 10201 2653
rect 10236 2682 10273 2752
rect 10539 2751 10576 2752
rect 10388 2692 10424 2693
rect 10236 2662 10245 2682
rect 10265 2662 10273 2682
rect 10236 2652 10273 2662
rect 10332 2682 10480 2692
rect 10580 2689 10676 2691
rect 10332 2662 10341 2682
rect 10361 2662 10451 2682
rect 10471 2662 10480 2682
rect 10332 2653 10480 2662
rect 10538 2682 10676 2689
rect 10538 2662 10547 2682
rect 10567 2662 10676 2682
rect 10538 2653 10676 2662
rect 10332 2652 10369 2653
rect 10062 2599 10103 2600
rect 8871 2579 9310 2597
rect 8031 2485 8071 2494
rect 8333 2485 8360 2572
rect 8433 2546 8476 2572
rect 8433 2528 8446 2546
rect 8464 2528 8476 2546
rect 8433 2517 8476 2528
rect 7305 2479 7340 2480
rect 7183 2469 7340 2479
rect 7183 2449 7200 2469
rect 7220 2449 7340 2469
rect 7183 2442 7340 2449
rect 7407 2472 7553 2480
rect 7407 2452 7418 2472
rect 7438 2452 7477 2472
rect 7497 2452 7553 2472
rect 8031 2468 8360 2485
rect 8031 2467 8071 2468
rect 7407 2445 7553 2452
rect 8428 2456 8468 2459
rect 8428 2450 8471 2456
rect 8053 2447 8471 2450
rect 7407 2444 7448 2445
rect 7141 2391 7178 2392
rect 6834 2382 6972 2391
rect 6834 2362 6943 2382
rect 6963 2362 6972 2382
rect 6834 2355 6972 2362
rect 7030 2382 7178 2391
rect 7030 2362 7039 2382
rect 7059 2362 7149 2382
rect 7169 2362 7178 2382
rect 6834 2353 6930 2355
rect 7030 2352 7178 2362
rect 7237 2382 7274 2392
rect 7237 2362 7245 2382
rect 7265 2362 7274 2382
rect 7086 2351 7122 2352
rect 6934 2292 6971 2293
rect 7237 2292 7274 2362
rect 7309 2391 7340 2442
rect 8053 2429 8444 2447
rect 8462 2429 8471 2447
rect 8053 2427 8471 2429
rect 8053 2419 8080 2427
rect 8321 2424 8471 2427
rect 7633 2413 7801 2414
rect 8052 2413 8080 2419
rect 7633 2397 8080 2413
rect 8428 2419 8471 2424
rect 7359 2391 7396 2392
rect 7309 2382 7396 2391
rect 7309 2362 7367 2382
rect 7387 2362 7396 2382
rect 7309 2352 7396 2362
rect 7455 2382 7492 2392
rect 7455 2362 7463 2382
rect 7483 2362 7492 2382
rect 7309 2351 7340 2352
rect 6933 2291 7274 2292
rect 7455 2291 7492 2362
rect 6858 2286 7274 2291
rect 6858 2266 6861 2286
rect 6881 2266 7274 2286
rect 7305 2267 7492 2291
rect 7633 2387 8077 2397
rect 7633 2385 7801 2387
rect 6733 2187 6775 2232
rect 7633 2207 7660 2385
rect 7700 2347 7764 2359
rect 8040 2355 8077 2387
rect 8103 2386 8294 2408
rect 8258 2384 8294 2386
rect 8258 2355 8295 2384
rect 8428 2363 8468 2419
rect 7700 2346 7735 2347
rect 7677 2341 7735 2346
rect 7677 2321 7680 2341
rect 7700 2327 7735 2341
rect 7755 2327 7764 2347
rect 7700 2319 7764 2327
rect 7726 2318 7764 2319
rect 7727 2317 7764 2318
rect 7830 2351 7866 2352
rect 7938 2351 7974 2352
rect 7830 2343 7974 2351
rect 7830 2323 7838 2343
rect 7858 2323 7893 2343
rect 7913 2323 7946 2343
rect 7966 2323 7974 2343
rect 7830 2317 7974 2323
rect 8040 2347 8078 2355
rect 8156 2351 8192 2352
rect 8040 2327 8049 2347
rect 8069 2327 8078 2347
rect 8040 2318 8078 2327
rect 8107 2343 8192 2351
rect 8107 2323 8164 2343
rect 8184 2323 8192 2343
rect 8040 2317 8077 2318
rect 8107 2317 8192 2323
rect 8258 2347 8296 2355
rect 8258 2327 8267 2347
rect 8287 2327 8296 2347
rect 8428 2345 8440 2363
rect 8458 2345 8468 2363
rect 8873 2390 8925 2579
rect 9271 2554 9310 2579
rect 9954 2592 10103 2599
rect 9954 2572 10013 2592
rect 10033 2572 10072 2592
rect 10092 2572 10103 2592
rect 9954 2564 10103 2572
rect 10170 2595 10327 2602
rect 10170 2575 10290 2595
rect 10310 2575 10327 2595
rect 10170 2565 10327 2575
rect 10170 2564 10205 2565
rect 9055 2529 9242 2553
rect 9271 2534 9666 2554
rect 9686 2534 9689 2554
rect 10170 2543 10201 2564
rect 10388 2543 10424 2653
rect 10443 2652 10480 2653
rect 10539 2652 10576 2653
rect 10499 2593 10589 2599
rect 10499 2573 10508 2593
rect 10528 2591 10589 2593
rect 10528 2573 10553 2591
rect 10499 2571 10553 2573
rect 10573 2571 10589 2591
rect 10499 2565 10589 2571
rect 10013 2542 10050 2543
rect 9271 2529 9689 2534
rect 10012 2533 10050 2542
rect 9055 2458 9092 2529
rect 9271 2528 9614 2529
rect 9271 2525 9310 2528
rect 9576 2527 9613 2528
rect 9207 2468 9238 2469
rect 9055 2438 9064 2458
rect 9084 2438 9092 2458
rect 9055 2428 9092 2438
rect 9151 2458 9238 2468
rect 9151 2438 9160 2458
rect 9180 2438 9238 2458
rect 9151 2429 9238 2438
rect 9151 2428 9188 2429
rect 8873 2372 8889 2390
rect 8907 2372 8925 2390
rect 9207 2378 9238 2429
rect 9273 2458 9310 2525
rect 10012 2513 10021 2533
rect 10041 2513 10050 2533
rect 10012 2505 10050 2513
rect 10116 2537 10201 2543
rect 10231 2542 10268 2543
rect 10116 2517 10124 2537
rect 10144 2517 10201 2537
rect 10116 2509 10201 2517
rect 10230 2533 10268 2542
rect 10230 2513 10239 2533
rect 10259 2513 10268 2533
rect 10116 2508 10152 2509
rect 10230 2505 10268 2513
rect 10334 2541 10478 2543
rect 10334 2537 10394 2541
rect 10334 2517 10342 2537
rect 10362 2519 10394 2537
rect 10417 2537 10478 2541
rect 10417 2519 10450 2537
rect 10362 2517 10450 2519
rect 10470 2517 10478 2537
rect 10334 2509 10478 2517
rect 10334 2508 10370 2509
rect 10442 2508 10478 2509
rect 10544 2542 10581 2543
rect 10544 2541 10582 2542
rect 10544 2533 10608 2541
rect 10544 2513 10553 2533
rect 10573 2519 10608 2533
rect 10628 2519 10631 2539
rect 10573 2514 10631 2519
rect 10573 2513 10608 2514
rect 10013 2476 10050 2505
rect 10014 2474 10050 2476
rect 9425 2468 9461 2469
rect 9273 2438 9282 2458
rect 9302 2438 9310 2458
rect 9273 2428 9310 2438
rect 9369 2458 9517 2468
rect 9617 2465 9713 2467
rect 9369 2438 9378 2458
rect 9398 2438 9488 2458
rect 9508 2438 9517 2458
rect 9369 2429 9517 2438
rect 9575 2458 9713 2465
rect 9575 2438 9584 2458
rect 9604 2438 9713 2458
rect 10014 2452 10205 2474
rect 10231 2473 10268 2505
rect 10544 2501 10608 2513
rect 10231 2472 10506 2473
rect 10648 2472 10675 2653
rect 10231 2447 10675 2472
rect 10811 2478 10850 4293
rect 11152 4280 11185 4613
rect 11249 4645 11417 4646
rect 11543 4645 11583 4869
rect 12046 4873 12214 4874
rect 12455 4873 12490 4890
rect 12847 4880 12894 4891
rect 12046 4847 12490 4873
rect 12046 4845 12214 4847
rect 12410 4846 12490 4847
rect 12645 4846 12712 4872
rect 12851 4846 12894 4880
rect 12046 4667 12073 4845
rect 12113 4807 12177 4819
rect 12453 4815 12490 4846
rect 12671 4815 12708 4846
rect 12853 4821 12894 4846
rect 13285 4905 13326 4930
rect 13471 4905 13508 4936
rect 13689 4905 13726 4936
rect 14002 4932 14066 4944
rect 14106 4906 14133 5084
rect 13285 4871 13328 4905
rect 13467 4879 13534 4905
rect 13689 4904 13769 4905
rect 13965 4904 14133 4906
rect 13689 4878 14133 4904
rect 13285 4860 13332 4871
rect 13689 4861 13724 4878
rect 13965 4877 14133 4878
rect 14596 4882 14636 5106
rect 14762 5105 14930 5106
rect 14994 5138 15027 5471
rect 15329 5458 15368 7273
rect 15504 7279 15948 7304
rect 15504 7098 15531 7279
rect 15673 7278 15948 7279
rect 15571 7238 15635 7250
rect 15911 7246 15948 7278
rect 15974 7277 16165 7299
rect 16466 7293 16575 7313
rect 16595 7293 16604 7313
rect 16466 7286 16604 7293
rect 16662 7313 16810 7322
rect 16662 7293 16671 7313
rect 16691 7293 16781 7313
rect 16801 7293 16810 7313
rect 16466 7284 16562 7286
rect 16662 7283 16810 7293
rect 16869 7313 16906 7323
rect 16869 7293 16877 7313
rect 16897 7293 16906 7313
rect 16718 7282 16754 7283
rect 16129 7275 16165 7277
rect 16129 7246 16166 7275
rect 15571 7237 15606 7238
rect 15548 7232 15606 7237
rect 15548 7212 15551 7232
rect 15571 7218 15606 7232
rect 15626 7218 15635 7238
rect 15571 7210 15635 7218
rect 15597 7209 15635 7210
rect 15598 7208 15635 7209
rect 15701 7242 15737 7243
rect 15809 7242 15845 7243
rect 15701 7234 15845 7242
rect 15701 7214 15709 7234
rect 15729 7232 15817 7234
rect 15729 7214 15762 7232
rect 15701 7210 15762 7214
rect 15785 7214 15817 7232
rect 15837 7214 15845 7234
rect 15785 7210 15845 7214
rect 15701 7208 15845 7210
rect 15911 7238 15949 7246
rect 16027 7242 16063 7243
rect 15911 7218 15920 7238
rect 15940 7218 15949 7238
rect 15911 7209 15949 7218
rect 15978 7234 16063 7242
rect 15978 7214 16035 7234
rect 16055 7214 16063 7234
rect 15911 7208 15948 7209
rect 15978 7208 16063 7214
rect 16129 7238 16167 7246
rect 16129 7218 16138 7238
rect 16158 7218 16167 7238
rect 16869 7226 16906 7293
rect 16941 7322 16972 7373
rect 17254 7361 17272 7379
rect 17290 7361 17306 7379
rect 17772 7386 17810 7395
rect 16991 7322 17028 7323
rect 16941 7313 17028 7322
rect 16941 7293 16999 7313
rect 17019 7293 17028 7313
rect 16941 7283 17028 7293
rect 17087 7313 17124 7323
rect 17087 7293 17095 7313
rect 17115 7293 17124 7313
rect 16941 7282 16972 7283
rect 16566 7223 16603 7224
rect 16869 7223 16908 7226
rect 16565 7222 16908 7223
rect 17087 7222 17124 7293
rect 16129 7209 16167 7218
rect 16490 7217 16908 7222
rect 16129 7208 16166 7209
rect 15590 7180 15680 7186
rect 15590 7160 15606 7180
rect 15626 7178 15680 7180
rect 15626 7160 15651 7178
rect 15590 7158 15651 7160
rect 15671 7158 15680 7178
rect 15590 7152 15680 7158
rect 15603 7098 15640 7099
rect 15699 7098 15736 7099
rect 15755 7098 15791 7208
rect 15978 7187 16009 7208
rect 16490 7197 16493 7217
rect 16513 7197 16908 7217
rect 16937 7198 17124 7222
rect 15974 7186 16009 7187
rect 15852 7176 16009 7186
rect 15852 7156 15869 7176
rect 15889 7156 16009 7176
rect 15852 7149 16009 7156
rect 16076 7179 16225 7187
rect 16076 7159 16087 7179
rect 16107 7159 16146 7179
rect 16166 7159 16225 7179
rect 16076 7152 16225 7159
rect 16869 7172 16908 7197
rect 17254 7172 17306 7361
rect 17600 7368 17640 7378
rect 17600 7350 17610 7368
rect 17628 7350 17640 7368
rect 17772 7366 17781 7386
rect 17801 7366 17810 7386
rect 17772 7358 17810 7366
rect 17876 7390 17961 7396
rect 17991 7395 18028 7396
rect 17876 7370 17884 7390
rect 17904 7370 17961 7390
rect 17876 7362 17961 7370
rect 17990 7386 18028 7395
rect 17990 7366 17999 7386
rect 18019 7366 18028 7386
rect 17876 7361 17912 7362
rect 17990 7358 18028 7366
rect 18094 7390 18238 7396
rect 18094 7370 18102 7390
rect 18122 7370 18155 7390
rect 18175 7370 18210 7390
rect 18230 7370 18238 7390
rect 18094 7362 18238 7370
rect 18094 7361 18130 7362
rect 18202 7361 18238 7362
rect 18304 7395 18341 7396
rect 18304 7394 18342 7395
rect 18304 7386 18368 7394
rect 18304 7366 18313 7386
rect 18333 7372 18368 7386
rect 18388 7372 18391 7392
rect 18333 7367 18391 7372
rect 18333 7366 18368 7367
rect 17600 7294 17640 7350
rect 17773 7329 17810 7358
rect 17774 7327 17810 7329
rect 17774 7305 17965 7327
rect 17991 7326 18028 7358
rect 18304 7354 18368 7366
rect 18408 7328 18435 7506
rect 19293 7481 19335 7526
rect 18267 7326 18435 7328
rect 17991 7316 18435 7326
rect 18576 7422 18763 7446
rect 18794 7427 19187 7447
rect 19207 7427 19210 7447
rect 18794 7422 19210 7427
rect 18576 7351 18613 7422
rect 18794 7421 19135 7422
rect 18728 7361 18759 7362
rect 18576 7331 18585 7351
rect 18605 7331 18613 7351
rect 18576 7321 18613 7331
rect 18672 7351 18759 7361
rect 18672 7331 18681 7351
rect 18701 7331 18759 7351
rect 18672 7322 18759 7331
rect 18672 7321 18709 7322
rect 17597 7289 17640 7294
rect 17988 7300 18435 7316
rect 17988 7294 18016 7300
rect 18267 7299 18435 7300
rect 17597 7286 17747 7289
rect 17988 7286 18015 7294
rect 17597 7284 18015 7286
rect 17597 7266 17606 7284
rect 17624 7266 18015 7284
rect 18728 7271 18759 7322
rect 18794 7351 18831 7421
rect 19097 7420 19134 7421
rect 18946 7361 18982 7362
rect 18794 7331 18803 7351
rect 18823 7331 18831 7351
rect 18794 7321 18831 7331
rect 18890 7351 19038 7361
rect 19138 7358 19234 7360
rect 18890 7331 18899 7351
rect 18919 7331 19009 7351
rect 19029 7331 19038 7351
rect 18890 7322 19038 7331
rect 19096 7351 19234 7358
rect 19096 7331 19105 7351
rect 19125 7331 19234 7351
rect 19096 7322 19234 7331
rect 18890 7321 18927 7322
rect 18620 7268 18661 7269
rect 17597 7263 18015 7266
rect 17597 7257 17640 7263
rect 17600 7254 17640 7257
rect 18515 7261 18661 7268
rect 17997 7245 18037 7246
rect 17708 7228 18037 7245
rect 18515 7241 18571 7261
rect 18591 7241 18630 7261
rect 18650 7241 18661 7261
rect 18515 7233 18661 7241
rect 18728 7264 18885 7271
rect 18728 7244 18848 7264
rect 18868 7244 18885 7264
rect 18728 7234 18885 7244
rect 18728 7233 18763 7234
rect 17592 7185 17635 7196
rect 16869 7154 17308 7172
rect 16076 7151 16117 7152
rect 15810 7098 15847 7099
rect 15503 7089 15641 7098
rect 15503 7069 15612 7089
rect 15632 7069 15641 7089
rect 15503 7062 15641 7069
rect 15699 7089 15847 7098
rect 15699 7069 15708 7089
rect 15728 7069 15818 7089
rect 15838 7069 15847 7089
rect 15503 7060 15599 7062
rect 15699 7059 15847 7069
rect 15906 7089 15943 7099
rect 15906 7069 15914 7089
rect 15934 7069 15943 7089
rect 15755 7058 15791 7059
rect 15603 6999 15640 7000
rect 15906 6999 15943 7069
rect 15978 7098 16009 7149
rect 16869 7136 17269 7154
rect 17287 7136 17308 7154
rect 16869 7130 17308 7136
rect 16875 7126 17308 7130
rect 17592 7167 17604 7185
rect 17622 7167 17635 7185
rect 17592 7141 17635 7167
rect 17708 7141 17735 7228
rect 17997 7219 18037 7228
rect 17254 7124 17306 7126
rect 17592 7120 17735 7141
rect 17779 7193 17813 7209
rect 17997 7199 18390 7219
rect 18410 7199 18413 7219
rect 18728 7212 18759 7233
rect 18946 7212 18982 7322
rect 19001 7321 19038 7322
rect 19097 7321 19134 7322
rect 19057 7262 19147 7268
rect 19057 7242 19066 7262
rect 19086 7260 19147 7262
rect 19086 7242 19111 7260
rect 19057 7240 19111 7242
rect 19131 7240 19147 7260
rect 19057 7234 19147 7240
rect 18571 7211 18608 7212
rect 17997 7194 18413 7199
rect 18570 7202 18608 7211
rect 17997 7193 18338 7194
rect 17779 7123 17816 7193
rect 17931 7133 17962 7134
rect 17592 7118 17729 7120
rect 16028 7098 16065 7099
rect 15978 7089 16065 7098
rect 15978 7069 16036 7089
rect 16056 7069 16065 7089
rect 15978 7059 16065 7069
rect 16124 7089 16161 7099
rect 16124 7069 16132 7089
rect 16152 7069 16161 7089
rect 17592 7076 17635 7118
rect 17779 7103 17788 7123
rect 17808 7103 17816 7123
rect 17779 7093 17816 7103
rect 17875 7123 17962 7133
rect 17875 7103 17884 7123
rect 17904 7103 17962 7123
rect 17875 7094 17962 7103
rect 17875 7093 17912 7094
rect 15978 7058 16009 7059
rect 15602 6998 15943 6999
rect 16124 6998 16161 7069
rect 17590 7066 17635 7076
rect 17257 7059 17294 7064
rect 15527 6993 15943 6998
rect 15527 6973 15530 6993
rect 15550 6973 15943 6993
rect 15974 6974 16161 6998
rect 17248 7055 17295 7059
rect 17248 7037 17267 7055
rect 17285 7037 17295 7055
rect 17590 7048 17599 7066
rect 17617 7048 17635 7066
rect 17590 7042 17635 7048
rect 17931 7043 17962 7094
rect 17997 7123 18034 7193
rect 18300 7192 18337 7193
rect 18570 7182 18579 7202
rect 18599 7182 18608 7202
rect 18570 7174 18608 7182
rect 18674 7206 18759 7212
rect 18789 7211 18826 7212
rect 18674 7186 18682 7206
rect 18702 7186 18759 7206
rect 18674 7178 18759 7186
rect 18788 7202 18826 7211
rect 18788 7182 18797 7202
rect 18817 7182 18826 7202
rect 18674 7177 18710 7178
rect 18788 7174 18826 7182
rect 18892 7206 19036 7212
rect 18892 7186 18900 7206
rect 18920 7203 19008 7206
rect 18920 7186 18955 7203
rect 18892 7185 18955 7186
rect 18974 7186 19008 7203
rect 19028 7186 19036 7206
rect 18974 7185 19036 7186
rect 18892 7178 19036 7185
rect 18892 7177 18928 7178
rect 19000 7177 19036 7178
rect 19102 7211 19139 7212
rect 19102 7210 19140 7211
rect 19162 7210 19189 7214
rect 19102 7208 19189 7210
rect 19102 7202 19166 7208
rect 19102 7182 19111 7202
rect 19131 7188 19166 7202
rect 19186 7188 19189 7208
rect 19131 7183 19189 7188
rect 19131 7182 19166 7183
rect 18571 7145 18608 7174
rect 18572 7143 18608 7145
rect 18149 7133 18185 7134
rect 17997 7103 18006 7123
rect 18026 7103 18034 7123
rect 17997 7093 18034 7103
rect 18093 7123 18241 7133
rect 18341 7130 18437 7132
rect 18093 7103 18102 7123
rect 18122 7103 18212 7123
rect 18232 7103 18241 7123
rect 18093 7094 18241 7103
rect 18299 7123 18437 7130
rect 18299 7103 18308 7123
rect 18328 7103 18437 7123
rect 18572 7121 18763 7143
rect 18789 7142 18826 7174
rect 19102 7170 19166 7182
rect 19206 7144 19233 7322
rect 19065 7142 19233 7144
rect 18789 7116 19233 7142
rect 18299 7094 18437 7103
rect 18093 7093 18130 7094
rect 17590 7039 17627 7042
rect 17823 7040 17864 7041
rect 17248 6989 17295 7037
rect 17715 7033 17864 7040
rect 17715 7013 17774 7033
rect 17794 7013 17833 7033
rect 17853 7013 17864 7033
rect 17715 7005 17864 7013
rect 17931 7036 18088 7043
rect 17931 7016 18051 7036
rect 18071 7016 18088 7036
rect 17931 7006 18088 7016
rect 17931 7005 17966 7006
rect 16872 6986 17295 6989
rect 15747 6972 15812 6973
rect 16850 6956 17295 6986
rect 17931 6984 17962 7005
rect 18149 6984 18185 7094
rect 18204 7093 18241 7094
rect 18300 7093 18337 7094
rect 18260 7034 18350 7040
rect 18260 7014 18269 7034
rect 18289 7032 18350 7034
rect 18289 7014 18314 7032
rect 18260 7012 18314 7014
rect 18334 7012 18350 7032
rect 18260 7006 18350 7012
rect 17774 6983 17811 6984
rect 15943 6940 15983 6948
rect 15943 6918 15951 6940
rect 15975 6918 15983 6940
rect 15548 6689 15585 6695
rect 15548 6670 15556 6689
rect 15577 6670 15585 6689
rect 15548 6662 15585 6670
rect 15552 6329 15585 6662
rect 15649 6694 15817 6695
rect 15943 6694 15983 6918
rect 16446 6922 16614 6923
rect 16850 6922 16891 6956
rect 17248 6935 17295 6956
rect 16446 6912 16891 6922
rect 16963 6920 17106 6921
rect 16446 6896 16890 6912
rect 16446 6894 16614 6896
rect 16810 6895 16890 6896
rect 16963 6895 17108 6920
rect 17250 6895 17295 6935
rect 17586 6975 17624 6977
rect 17586 6967 17629 6975
rect 17586 6949 17597 6967
rect 17615 6949 17629 6967
rect 17586 6922 17629 6949
rect 17773 6974 17811 6983
rect 17773 6954 17782 6974
rect 17802 6954 17811 6974
rect 17773 6946 17811 6954
rect 17877 6978 17962 6984
rect 17992 6983 18029 6984
rect 17877 6958 17885 6978
rect 17905 6958 17962 6978
rect 17877 6950 17962 6958
rect 17991 6974 18029 6983
rect 17991 6954 18000 6974
rect 18020 6954 18029 6974
rect 17877 6949 17913 6950
rect 17991 6946 18029 6954
rect 18095 6982 18239 6984
rect 18095 6978 18147 6982
rect 18095 6958 18103 6978
rect 18123 6962 18147 6978
rect 18167 6978 18239 6982
rect 18167 6962 18211 6978
rect 18123 6958 18211 6962
rect 18231 6958 18239 6978
rect 18095 6950 18239 6958
rect 18095 6949 18131 6950
rect 18203 6949 18239 6950
rect 18305 6983 18342 6984
rect 18305 6982 18343 6983
rect 18305 6974 18369 6982
rect 18305 6954 18314 6974
rect 18334 6960 18369 6974
rect 18389 6960 18392 6980
rect 18334 6955 18392 6960
rect 18334 6954 18369 6955
rect 16446 6716 16473 6894
rect 16513 6856 16577 6868
rect 16853 6864 16890 6895
rect 17071 6864 17108 6895
rect 17253 6888 17295 6895
rect 17587 6915 17629 6922
rect 17774 6915 17811 6946
rect 17992 6915 18029 6946
rect 18305 6942 18369 6954
rect 18409 6916 18436 7094
rect 16513 6855 16548 6856
rect 16490 6850 16548 6855
rect 16490 6830 16493 6850
rect 16513 6836 16548 6850
rect 16568 6836 16577 6856
rect 16513 6828 16577 6836
rect 16539 6827 16577 6828
rect 16540 6826 16577 6827
rect 16643 6860 16679 6861
rect 16751 6860 16787 6861
rect 16643 6852 16787 6860
rect 16643 6832 16651 6852
rect 16671 6848 16759 6852
rect 16671 6832 16715 6848
rect 16643 6828 16715 6832
rect 16735 6832 16759 6848
rect 16779 6832 16787 6852
rect 16735 6828 16787 6832
rect 16643 6826 16787 6828
rect 16853 6856 16891 6864
rect 16969 6860 17005 6861
rect 16853 6836 16862 6856
rect 16882 6836 16891 6856
rect 16853 6827 16891 6836
rect 16920 6852 17005 6860
rect 16920 6832 16977 6852
rect 16997 6832 17005 6852
rect 16853 6826 16890 6827
rect 16920 6826 17005 6832
rect 17071 6856 17109 6864
rect 17071 6836 17080 6856
rect 17100 6836 17109 6856
rect 17071 6827 17109 6836
rect 17253 6861 17296 6888
rect 17253 6843 17267 6861
rect 17285 6843 17296 6861
rect 17253 6835 17296 6843
rect 17258 6833 17296 6835
rect 17587 6875 17632 6915
rect 17774 6890 17919 6915
rect 17992 6914 18072 6915
rect 18268 6914 18436 6916
rect 17992 6898 18436 6914
rect 17776 6889 17919 6890
rect 17991 6888 18436 6898
rect 17587 6854 17634 6875
rect 17991 6854 18032 6888
rect 18268 6887 18436 6888
rect 18899 6892 18939 7116
rect 19065 7115 19233 7116
rect 19297 7148 19330 7481
rect 19935 7480 19962 7658
rect 20002 7620 20066 7632
rect 20342 7628 20379 7660
rect 20405 7659 20596 7681
rect 20731 7679 20840 7699
rect 20860 7679 20869 7699
rect 20731 7672 20869 7679
rect 20927 7699 21075 7708
rect 20927 7679 20936 7699
rect 20956 7679 21046 7699
rect 21066 7679 21075 7699
rect 20731 7670 20827 7672
rect 20927 7669 21075 7679
rect 21134 7699 21171 7709
rect 21134 7679 21142 7699
rect 21162 7679 21171 7699
rect 20983 7668 21019 7669
rect 20560 7657 20596 7659
rect 20560 7628 20597 7657
rect 20002 7619 20037 7620
rect 19979 7614 20037 7619
rect 19979 7594 19982 7614
rect 20002 7600 20037 7614
rect 20057 7600 20066 7620
rect 20002 7592 20066 7600
rect 20028 7591 20066 7592
rect 20029 7590 20066 7591
rect 20132 7624 20168 7625
rect 20240 7624 20276 7625
rect 20132 7616 20276 7624
rect 20132 7596 20140 7616
rect 20160 7615 20248 7616
rect 20160 7596 20195 7615
rect 20216 7596 20248 7615
rect 20268 7596 20276 7616
rect 20132 7590 20276 7596
rect 20342 7620 20380 7628
rect 20458 7624 20494 7625
rect 20342 7600 20351 7620
rect 20371 7600 20380 7620
rect 20342 7591 20380 7600
rect 20409 7616 20494 7624
rect 20409 7596 20466 7616
rect 20486 7596 20494 7616
rect 20342 7590 20379 7591
rect 20409 7590 20494 7596
rect 20560 7620 20598 7628
rect 20560 7600 20569 7620
rect 20589 7600 20598 7620
rect 20831 7609 20868 7610
rect 21134 7609 21171 7679
rect 21206 7708 21237 7759
rect 21533 7754 21578 7760
rect 21533 7736 21551 7754
rect 21569 7736 21578 7754
rect 23039 7754 23048 7774
rect 23068 7754 23076 7774
rect 23039 7744 23076 7754
rect 23135 7774 23222 7784
rect 23135 7754 23144 7774
rect 23164 7754 23222 7774
rect 23135 7745 23222 7754
rect 23135 7744 23172 7745
rect 21533 7726 21578 7736
rect 21256 7708 21293 7709
rect 21206 7699 21293 7708
rect 21206 7679 21264 7699
rect 21284 7679 21293 7699
rect 21206 7669 21293 7679
rect 21352 7699 21389 7709
rect 21352 7679 21360 7699
rect 21380 7679 21389 7699
rect 21533 7684 21576 7726
rect 21960 7715 22012 7717
rect 21439 7682 21576 7684
rect 21206 7668 21237 7669
rect 21352 7609 21389 7679
rect 20830 7608 21171 7609
rect 20560 7591 20598 7600
rect 20755 7603 21171 7608
rect 20560 7590 20597 7591
rect 20021 7562 20111 7568
rect 20021 7542 20037 7562
rect 20057 7560 20111 7562
rect 20057 7542 20082 7560
rect 20021 7540 20082 7542
rect 20102 7540 20111 7560
rect 20021 7534 20111 7540
rect 20034 7480 20071 7481
rect 20130 7480 20167 7481
rect 20186 7480 20222 7590
rect 20409 7569 20440 7590
rect 20755 7583 20758 7603
rect 20778 7583 21171 7603
rect 21355 7593 21389 7609
rect 21433 7661 21576 7682
rect 21958 7711 22391 7715
rect 21958 7705 22397 7711
rect 21958 7687 21979 7705
rect 21997 7687 22397 7705
rect 23191 7694 23222 7745
rect 23257 7774 23294 7844
rect 23560 7843 23597 7844
rect 23409 7784 23445 7785
rect 23257 7754 23266 7774
rect 23286 7754 23294 7774
rect 23257 7744 23294 7754
rect 23353 7774 23501 7784
rect 23601 7781 23697 7783
rect 23353 7754 23362 7774
rect 23382 7754 23472 7774
rect 23492 7754 23501 7774
rect 23353 7745 23501 7754
rect 23559 7774 23697 7781
rect 23559 7754 23568 7774
rect 23588 7754 23697 7774
rect 23559 7745 23697 7754
rect 23353 7744 23390 7745
rect 23083 7691 23124 7692
rect 21958 7669 22397 7687
rect 21131 7574 21171 7583
rect 21433 7574 21460 7661
rect 21533 7635 21576 7661
rect 21533 7617 21546 7635
rect 21564 7617 21576 7635
rect 21533 7606 21576 7617
rect 20405 7568 20440 7569
rect 20283 7558 20440 7568
rect 20283 7538 20300 7558
rect 20320 7538 20440 7558
rect 20283 7531 20440 7538
rect 20507 7561 20656 7569
rect 20507 7541 20518 7561
rect 20538 7541 20577 7561
rect 20597 7541 20656 7561
rect 21131 7557 21460 7574
rect 21131 7556 21171 7557
rect 20507 7534 20656 7541
rect 21528 7545 21568 7548
rect 21528 7539 21571 7545
rect 21153 7536 21571 7539
rect 20507 7533 20548 7534
rect 20241 7480 20278 7481
rect 19934 7471 20072 7480
rect 19797 7461 19833 7467
rect 19797 7443 19802 7461
rect 19824 7443 19833 7461
rect 19797 7439 19833 7443
rect 19934 7451 20043 7471
rect 20063 7451 20072 7471
rect 19934 7444 20072 7451
rect 20130 7471 20278 7480
rect 20130 7451 20139 7471
rect 20159 7451 20249 7471
rect 20269 7451 20278 7471
rect 19934 7442 20030 7444
rect 20130 7441 20278 7451
rect 20337 7471 20374 7481
rect 20337 7451 20345 7471
rect 20365 7451 20374 7471
rect 20186 7440 20222 7441
rect 19800 7280 19833 7439
rect 20034 7381 20071 7382
rect 20337 7381 20374 7451
rect 20409 7480 20440 7531
rect 21153 7518 21544 7536
rect 21562 7518 21571 7536
rect 21153 7516 21571 7518
rect 21153 7508 21180 7516
rect 21421 7513 21571 7516
rect 20733 7502 20901 7503
rect 21152 7502 21180 7508
rect 20733 7486 21180 7502
rect 21528 7508 21571 7513
rect 20459 7480 20496 7481
rect 20409 7471 20496 7480
rect 20409 7451 20467 7471
rect 20487 7451 20496 7471
rect 20409 7441 20496 7451
rect 20555 7471 20592 7481
rect 20555 7451 20563 7471
rect 20583 7451 20592 7471
rect 20409 7440 20440 7441
rect 20033 7380 20374 7381
rect 20555 7380 20592 7451
rect 19958 7375 20374 7380
rect 19958 7355 19961 7375
rect 19981 7355 20374 7375
rect 20405 7356 20592 7380
rect 20733 7476 21177 7486
rect 20733 7474 20901 7476
rect 20733 7296 20760 7474
rect 20800 7436 20864 7448
rect 21140 7444 21177 7476
rect 21203 7475 21394 7497
rect 21358 7473 21394 7475
rect 21358 7444 21395 7473
rect 21528 7452 21568 7508
rect 20800 7435 20835 7436
rect 20777 7430 20835 7435
rect 20777 7410 20780 7430
rect 20800 7416 20835 7430
rect 20855 7416 20864 7436
rect 20800 7408 20864 7416
rect 20826 7407 20864 7408
rect 20827 7406 20864 7407
rect 20930 7440 20966 7441
rect 21038 7440 21074 7441
rect 20930 7432 21074 7440
rect 20930 7412 20938 7432
rect 20958 7412 20993 7432
rect 21013 7412 21046 7432
rect 21066 7412 21074 7432
rect 20930 7406 21074 7412
rect 21140 7436 21178 7444
rect 21256 7440 21292 7441
rect 21140 7416 21149 7436
rect 21169 7416 21178 7436
rect 21140 7407 21178 7416
rect 21207 7432 21292 7440
rect 21207 7412 21264 7432
rect 21284 7412 21292 7432
rect 21140 7406 21177 7407
rect 21207 7406 21292 7412
rect 21358 7436 21396 7444
rect 21358 7416 21367 7436
rect 21387 7416 21396 7436
rect 21528 7434 21540 7452
rect 21558 7434 21568 7452
rect 21960 7480 22012 7669
rect 22358 7644 22397 7669
rect 22975 7684 23124 7691
rect 22975 7664 23034 7684
rect 23054 7664 23093 7684
rect 23113 7664 23124 7684
rect 22975 7656 23124 7664
rect 23191 7687 23348 7694
rect 23191 7667 23311 7687
rect 23331 7667 23348 7687
rect 23191 7657 23348 7667
rect 23191 7656 23226 7657
rect 22142 7619 22329 7643
rect 22358 7624 22753 7644
rect 22773 7624 22776 7644
rect 23191 7635 23222 7656
rect 23409 7635 23445 7745
rect 23464 7744 23501 7745
rect 23560 7744 23597 7745
rect 23520 7685 23610 7691
rect 23520 7665 23529 7685
rect 23549 7683 23610 7685
rect 23549 7665 23574 7683
rect 23520 7663 23574 7665
rect 23594 7663 23610 7683
rect 23520 7657 23610 7663
rect 23034 7634 23071 7635
rect 22358 7619 22776 7624
rect 23033 7625 23071 7634
rect 22142 7548 22179 7619
rect 22358 7618 22701 7619
rect 22358 7615 22397 7618
rect 22663 7617 22700 7618
rect 22294 7558 22325 7559
rect 22142 7528 22151 7548
rect 22171 7528 22179 7548
rect 22142 7518 22179 7528
rect 22238 7548 22325 7558
rect 22238 7528 22247 7548
rect 22267 7528 22325 7548
rect 22238 7519 22325 7528
rect 22238 7518 22275 7519
rect 21960 7462 21976 7480
rect 21994 7462 22012 7480
rect 22294 7468 22325 7519
rect 22360 7548 22397 7615
rect 23033 7605 23042 7625
rect 23062 7605 23071 7625
rect 23033 7597 23071 7605
rect 23137 7629 23222 7635
rect 23252 7634 23289 7635
rect 23137 7609 23145 7629
rect 23165 7609 23222 7629
rect 23137 7601 23222 7609
rect 23251 7625 23289 7634
rect 23251 7605 23260 7625
rect 23280 7605 23289 7625
rect 23137 7600 23173 7601
rect 23251 7597 23289 7605
rect 23355 7630 23499 7635
rect 23355 7629 23417 7630
rect 23355 7609 23363 7629
rect 23383 7611 23417 7629
rect 23438 7629 23499 7630
rect 23438 7611 23471 7629
rect 23383 7609 23471 7611
rect 23491 7609 23499 7629
rect 23355 7601 23499 7609
rect 23355 7600 23391 7601
rect 23463 7600 23499 7601
rect 23565 7634 23602 7635
rect 23565 7633 23603 7634
rect 23565 7625 23629 7633
rect 23565 7605 23574 7625
rect 23594 7611 23629 7625
rect 23649 7611 23652 7631
rect 23594 7606 23652 7611
rect 23594 7605 23629 7606
rect 23034 7568 23071 7597
rect 23035 7566 23071 7568
rect 22512 7558 22548 7559
rect 22360 7528 22369 7548
rect 22389 7528 22397 7548
rect 22360 7518 22397 7528
rect 22456 7548 22604 7558
rect 22704 7555 22800 7557
rect 22456 7528 22465 7548
rect 22485 7528 22575 7548
rect 22595 7528 22604 7548
rect 22456 7519 22604 7528
rect 22662 7548 22800 7555
rect 22662 7528 22671 7548
rect 22691 7528 22800 7548
rect 23035 7544 23226 7566
rect 23252 7565 23289 7597
rect 23565 7593 23629 7605
rect 23669 7567 23696 7745
rect 23528 7565 23696 7567
rect 23252 7551 23696 7565
rect 24299 7699 24467 7700
rect 24593 7699 24633 7923
rect 25096 7927 25264 7928
rect 25499 7927 25539 7960
rect 25895 7927 25942 7960
rect 26346 7958 26387 7983
rect 26532 7958 26569 7989
rect 26750 7958 26787 7989
rect 27063 7985 27127 7997
rect 27167 7959 27194 8137
rect 26346 7931 26395 7958
rect 26531 7932 26580 7958
rect 26749 7957 26830 7958
rect 27026 7957 27194 7959
rect 26749 7932 27194 7957
rect 26750 7931 27194 7932
rect 25096 7926 25540 7927
rect 25096 7901 25541 7926
rect 25096 7899 25264 7901
rect 25460 7900 25541 7901
rect 25710 7900 25759 7926
rect 25895 7900 25944 7927
rect 25096 7721 25123 7899
rect 25163 7861 25227 7873
rect 25503 7869 25540 7900
rect 25721 7869 25758 7900
rect 25903 7875 25944 7900
rect 26348 7898 26395 7931
rect 26751 7898 26791 7931
rect 27026 7930 27194 7931
rect 27657 7935 27697 8159
rect 27823 8158 27991 8159
rect 28594 8293 29038 8307
rect 28594 8291 28762 8293
rect 28594 8113 28621 8291
rect 28661 8253 28725 8265
rect 29001 8261 29038 8293
rect 29064 8292 29255 8314
rect 29490 8310 29599 8330
rect 29619 8310 29628 8330
rect 29490 8303 29628 8310
rect 29686 8330 29834 8339
rect 29686 8310 29695 8330
rect 29715 8310 29805 8330
rect 29825 8310 29834 8330
rect 29490 8301 29586 8303
rect 29686 8300 29834 8310
rect 29893 8330 29930 8340
rect 29893 8310 29901 8330
rect 29921 8310 29930 8330
rect 29742 8299 29778 8300
rect 29219 8290 29255 8292
rect 29219 8261 29256 8290
rect 28661 8252 28696 8253
rect 28638 8247 28696 8252
rect 28638 8227 28641 8247
rect 28661 8233 28696 8247
rect 28716 8233 28725 8253
rect 28661 8225 28725 8233
rect 28687 8224 28725 8225
rect 28688 8223 28725 8224
rect 28791 8257 28827 8258
rect 28899 8257 28935 8258
rect 28791 8251 28935 8257
rect 28791 8249 28852 8251
rect 28791 8229 28799 8249
rect 28819 8234 28852 8249
rect 28871 8249 28935 8251
rect 28871 8234 28907 8249
rect 28819 8229 28907 8234
rect 28927 8229 28935 8249
rect 28791 8223 28935 8229
rect 29001 8253 29039 8261
rect 29117 8257 29153 8258
rect 29001 8233 29010 8253
rect 29030 8233 29039 8253
rect 29001 8224 29039 8233
rect 29068 8249 29153 8257
rect 29068 8229 29125 8249
rect 29145 8229 29153 8249
rect 29001 8223 29038 8224
rect 29068 8223 29153 8229
rect 29219 8253 29257 8261
rect 29219 8233 29228 8253
rect 29248 8233 29257 8253
rect 29893 8243 29930 8310
rect 29965 8339 29996 8390
rect 30278 8378 30296 8396
rect 30314 8378 30330 8396
rect 30015 8339 30052 8340
rect 29965 8330 30052 8339
rect 29965 8310 30023 8330
rect 30043 8310 30052 8330
rect 29965 8300 30052 8310
rect 30111 8330 30148 8340
rect 30111 8310 30119 8330
rect 30139 8310 30148 8330
rect 29965 8299 29996 8300
rect 29590 8240 29627 8241
rect 29893 8240 29932 8243
rect 29589 8239 29932 8240
rect 30111 8239 30148 8310
rect 29219 8224 29257 8233
rect 29514 8234 29932 8239
rect 29219 8223 29256 8224
rect 28680 8195 28770 8201
rect 28680 8175 28696 8195
rect 28716 8193 28770 8195
rect 28716 8175 28741 8193
rect 28680 8173 28741 8175
rect 28761 8173 28770 8193
rect 28680 8167 28770 8173
rect 28693 8113 28730 8114
rect 28789 8113 28826 8114
rect 28845 8113 28881 8223
rect 29068 8202 29099 8223
rect 29514 8214 29517 8234
rect 29537 8214 29932 8234
rect 29961 8215 30148 8239
rect 29064 8201 29099 8202
rect 28942 8191 29099 8201
rect 28942 8171 28959 8191
rect 28979 8171 29099 8191
rect 28942 8164 29099 8171
rect 29166 8194 29315 8202
rect 29166 8174 29177 8194
rect 29197 8174 29236 8194
rect 29256 8174 29315 8194
rect 29166 8167 29315 8174
rect 29893 8189 29932 8214
rect 30278 8189 30330 8378
rect 30722 8406 30732 8424
rect 30750 8406 30762 8424
rect 30894 8422 30903 8442
rect 30923 8422 30932 8442
rect 30894 8414 30932 8422
rect 30998 8446 31083 8452
rect 31113 8451 31150 8452
rect 30998 8426 31006 8446
rect 31026 8426 31083 8446
rect 30998 8418 31083 8426
rect 31112 8442 31150 8451
rect 31112 8422 31121 8442
rect 31141 8422 31150 8442
rect 30998 8417 31034 8418
rect 31112 8414 31150 8422
rect 31216 8446 31360 8452
rect 31216 8426 31224 8446
rect 31244 8426 31277 8446
rect 31297 8426 31332 8446
rect 31352 8426 31360 8446
rect 31216 8418 31360 8426
rect 31216 8417 31252 8418
rect 31324 8417 31360 8418
rect 31426 8451 31463 8452
rect 31426 8450 31464 8451
rect 31426 8442 31490 8450
rect 31426 8422 31435 8442
rect 31455 8428 31490 8442
rect 31510 8428 31513 8448
rect 31455 8423 31513 8428
rect 31455 8422 31490 8423
rect 30722 8350 30762 8406
rect 30895 8385 30932 8414
rect 30896 8383 30932 8385
rect 30896 8361 31087 8383
rect 31113 8382 31150 8414
rect 31426 8410 31490 8422
rect 31530 8384 31557 8562
rect 31389 8382 31557 8384
rect 31113 8372 31557 8382
rect 31698 8478 31885 8502
rect 31916 8483 32309 8503
rect 32329 8483 32332 8503
rect 31916 8478 32332 8483
rect 31698 8407 31735 8478
rect 31916 8477 32257 8478
rect 31850 8417 31881 8418
rect 31698 8387 31707 8407
rect 31727 8387 31735 8407
rect 31698 8377 31735 8387
rect 31794 8407 31881 8417
rect 31794 8387 31803 8407
rect 31823 8387 31881 8407
rect 31794 8378 31881 8387
rect 31794 8377 31831 8378
rect 30719 8345 30762 8350
rect 31110 8356 31557 8372
rect 31110 8350 31138 8356
rect 31389 8355 31557 8356
rect 30719 8342 30869 8345
rect 31110 8342 31137 8350
rect 30719 8340 31137 8342
rect 30719 8322 30728 8340
rect 30746 8322 31137 8340
rect 31850 8327 31881 8378
rect 31916 8407 31953 8477
rect 32219 8476 32256 8477
rect 32068 8417 32104 8418
rect 31916 8387 31925 8407
rect 31945 8387 31953 8407
rect 31916 8377 31953 8387
rect 32012 8407 32160 8417
rect 32260 8414 32356 8416
rect 32012 8387 32021 8407
rect 32041 8387 32131 8407
rect 32151 8387 32160 8407
rect 32012 8378 32160 8387
rect 32218 8407 32356 8414
rect 32218 8387 32227 8407
rect 32247 8387 32356 8407
rect 32218 8378 32356 8387
rect 32012 8377 32049 8378
rect 31742 8324 31783 8325
rect 30719 8319 31137 8322
rect 30719 8313 30762 8319
rect 30722 8310 30762 8313
rect 31634 8317 31783 8324
rect 31119 8301 31159 8302
rect 30830 8284 31159 8301
rect 31634 8297 31693 8317
rect 31713 8297 31752 8317
rect 31772 8297 31783 8317
rect 31634 8289 31783 8297
rect 31850 8320 32007 8327
rect 31850 8300 31970 8320
rect 31990 8300 32007 8320
rect 31850 8290 32007 8300
rect 31850 8289 31885 8290
rect 30714 8241 30757 8252
rect 30714 8223 30726 8241
rect 30744 8223 30757 8241
rect 30714 8197 30757 8223
rect 30830 8197 30857 8284
rect 31119 8275 31159 8284
rect 29893 8171 30332 8189
rect 29166 8166 29207 8167
rect 28900 8113 28937 8114
rect 28593 8104 28731 8113
rect 28593 8084 28702 8104
rect 28722 8084 28731 8104
rect 28593 8077 28731 8084
rect 28789 8104 28937 8113
rect 28789 8084 28798 8104
rect 28818 8084 28908 8104
rect 28928 8084 28937 8104
rect 28593 8075 28689 8077
rect 28789 8074 28937 8084
rect 28996 8104 29033 8114
rect 28996 8084 29004 8104
rect 29024 8084 29033 8104
rect 28845 8073 28881 8074
rect 28693 8014 28730 8015
rect 28996 8014 29033 8084
rect 29068 8113 29099 8164
rect 29893 8153 30293 8171
rect 30311 8153 30332 8171
rect 29893 8147 30332 8153
rect 29899 8143 30332 8147
rect 30714 8176 30857 8197
rect 30901 8249 30935 8265
rect 31119 8255 31512 8275
rect 31532 8255 31535 8275
rect 31850 8268 31881 8289
rect 32068 8268 32104 8378
rect 32123 8377 32160 8378
rect 32219 8377 32256 8378
rect 32179 8318 32269 8324
rect 32179 8298 32188 8318
rect 32208 8316 32269 8318
rect 32208 8298 32233 8316
rect 32179 8296 32233 8298
rect 32253 8296 32269 8316
rect 32179 8290 32269 8296
rect 31693 8267 31730 8268
rect 31119 8250 31535 8255
rect 31692 8258 31730 8267
rect 31119 8249 31460 8250
rect 30901 8179 30938 8249
rect 31053 8189 31084 8190
rect 30714 8174 30851 8176
rect 30278 8141 30330 8143
rect 30714 8132 30757 8174
rect 30901 8159 30910 8179
rect 30930 8159 30938 8179
rect 30901 8149 30938 8159
rect 30997 8179 31084 8189
rect 30997 8159 31006 8179
rect 31026 8159 31084 8179
rect 30997 8150 31084 8159
rect 30997 8149 31034 8150
rect 30712 8122 30757 8132
rect 29118 8113 29155 8114
rect 29068 8104 29155 8113
rect 29068 8084 29126 8104
rect 29146 8084 29155 8104
rect 29068 8074 29155 8084
rect 29214 8104 29251 8114
rect 29214 8084 29222 8104
rect 29242 8084 29251 8104
rect 30712 8104 30721 8122
rect 30739 8104 30757 8122
rect 30712 8098 30757 8104
rect 31053 8099 31084 8150
rect 31119 8179 31156 8249
rect 31422 8248 31459 8249
rect 31692 8238 31701 8258
rect 31721 8238 31730 8258
rect 31692 8230 31730 8238
rect 31796 8262 31881 8268
rect 31911 8267 31948 8268
rect 31796 8242 31804 8262
rect 31824 8242 31881 8262
rect 31796 8234 31881 8242
rect 31910 8258 31948 8267
rect 31910 8238 31919 8258
rect 31939 8238 31948 8258
rect 31796 8233 31832 8234
rect 31910 8230 31948 8238
rect 32014 8262 32158 8268
rect 32014 8242 32022 8262
rect 32042 8243 32074 8262
rect 32095 8243 32130 8262
rect 32042 8242 32130 8243
rect 32150 8242 32158 8262
rect 32014 8234 32158 8242
rect 32014 8233 32050 8234
rect 32122 8233 32158 8234
rect 32224 8267 32261 8268
rect 32224 8266 32262 8267
rect 32224 8258 32288 8266
rect 32224 8238 32233 8258
rect 32253 8244 32288 8258
rect 32308 8244 32311 8264
rect 32253 8239 32311 8244
rect 32253 8238 32288 8239
rect 31693 8201 31730 8230
rect 31694 8199 31730 8201
rect 31271 8189 31307 8190
rect 31119 8159 31128 8179
rect 31148 8159 31156 8179
rect 31119 8149 31156 8159
rect 31215 8179 31363 8189
rect 31463 8186 31559 8188
rect 31215 8159 31224 8179
rect 31244 8159 31334 8179
rect 31354 8159 31363 8179
rect 31215 8150 31363 8159
rect 31421 8179 31559 8186
rect 31421 8159 31430 8179
rect 31450 8159 31559 8179
rect 31694 8177 31885 8199
rect 31911 8198 31948 8230
rect 32224 8226 32288 8238
rect 32328 8200 32355 8378
rect 32960 8377 32993 8710
rect 33057 8742 33225 8743
rect 33351 8742 33391 8966
rect 33854 8970 34022 8971
rect 33854 8969 34298 8970
rect 34661 8969 34702 8970
rect 33854 8944 34702 8969
rect 33854 8942 34022 8944
rect 34218 8943 34702 8944
rect 33854 8764 33881 8942
rect 33921 8904 33985 8916
rect 34261 8912 34298 8943
rect 34479 8912 34516 8943
rect 34661 8918 34702 8943
rect 33921 8903 33956 8904
rect 33898 8898 33956 8903
rect 33898 8878 33901 8898
rect 33921 8884 33956 8898
rect 33976 8884 33985 8904
rect 33921 8876 33985 8884
rect 33947 8875 33985 8876
rect 33948 8874 33985 8875
rect 34051 8908 34087 8909
rect 34159 8908 34195 8909
rect 34051 8900 34195 8908
rect 34051 8880 34059 8900
rect 34079 8896 34167 8900
rect 34079 8880 34123 8896
rect 34051 8876 34123 8880
rect 34143 8880 34167 8896
rect 34187 8880 34195 8900
rect 34143 8876 34195 8880
rect 34051 8874 34195 8876
rect 34261 8904 34299 8912
rect 34377 8908 34413 8909
rect 34261 8884 34270 8904
rect 34290 8884 34299 8904
rect 34261 8875 34299 8884
rect 34328 8900 34413 8908
rect 34328 8880 34385 8900
rect 34405 8880 34413 8900
rect 34261 8874 34298 8875
rect 34328 8874 34413 8880
rect 34479 8904 34517 8912
rect 34479 8884 34488 8904
rect 34508 8884 34517 8904
rect 34479 8875 34517 8884
rect 34661 8909 34703 8918
rect 34661 8891 34675 8909
rect 34693 8891 34703 8909
rect 34661 8883 34703 8891
rect 34666 8881 34703 8883
rect 34479 8874 34516 8875
rect 33940 8846 34030 8852
rect 33940 8826 33956 8846
rect 33976 8844 34030 8846
rect 33976 8826 34001 8844
rect 33940 8824 34001 8826
rect 34021 8824 34030 8844
rect 33940 8818 34030 8824
rect 33953 8764 33990 8765
rect 34049 8764 34086 8765
rect 34105 8764 34141 8874
rect 34328 8853 34359 8874
rect 34324 8852 34359 8853
rect 34202 8842 34359 8852
rect 34202 8822 34219 8842
rect 34239 8822 34359 8842
rect 34202 8815 34359 8822
rect 34426 8845 34575 8853
rect 34426 8825 34437 8845
rect 34457 8825 34496 8845
rect 34516 8825 34575 8845
rect 34426 8818 34575 8825
rect 34426 8817 34467 8818
rect 34663 8816 34700 8819
rect 34160 8764 34197 8765
rect 33853 8755 33991 8764
rect 33057 8716 33501 8742
rect 33057 8714 33225 8716
rect 33057 8536 33084 8714
rect 33124 8676 33188 8688
rect 33464 8684 33501 8716
rect 33527 8715 33718 8737
rect 33853 8735 33962 8755
rect 33982 8735 33991 8755
rect 33853 8728 33991 8735
rect 34049 8755 34197 8764
rect 34049 8735 34058 8755
rect 34078 8735 34168 8755
rect 34188 8735 34197 8755
rect 33853 8726 33949 8728
rect 34049 8725 34197 8735
rect 34256 8755 34293 8765
rect 34256 8735 34264 8755
rect 34284 8735 34293 8755
rect 34105 8724 34141 8725
rect 33682 8713 33718 8715
rect 33682 8684 33719 8713
rect 33124 8675 33159 8676
rect 33101 8670 33159 8675
rect 33101 8650 33104 8670
rect 33124 8656 33159 8670
rect 33179 8656 33188 8676
rect 33124 8650 33188 8656
rect 33101 8648 33188 8650
rect 33101 8644 33128 8648
rect 33150 8647 33188 8648
rect 33151 8646 33188 8647
rect 33254 8680 33290 8681
rect 33362 8680 33398 8681
rect 33254 8673 33398 8680
rect 33254 8672 33316 8673
rect 33254 8652 33262 8672
rect 33282 8655 33316 8672
rect 33335 8672 33398 8673
rect 33335 8655 33370 8672
rect 33282 8652 33370 8655
rect 33390 8652 33398 8672
rect 33254 8646 33398 8652
rect 33464 8676 33502 8684
rect 33580 8680 33616 8681
rect 33464 8656 33473 8676
rect 33493 8656 33502 8676
rect 33464 8647 33502 8656
rect 33531 8672 33616 8680
rect 33531 8652 33588 8672
rect 33608 8652 33616 8672
rect 33464 8646 33501 8647
rect 33531 8646 33616 8652
rect 33682 8676 33720 8684
rect 33682 8656 33691 8676
rect 33711 8656 33720 8676
rect 33953 8665 33990 8666
rect 34256 8665 34293 8735
rect 34328 8764 34359 8815
rect 34655 8810 34700 8816
rect 34655 8792 34673 8810
rect 34691 8792 34700 8810
rect 34655 8782 34700 8792
rect 34378 8764 34415 8765
rect 34328 8755 34415 8764
rect 34328 8735 34386 8755
rect 34406 8735 34415 8755
rect 34328 8725 34415 8735
rect 34474 8755 34511 8765
rect 34474 8735 34482 8755
rect 34502 8735 34511 8755
rect 34655 8740 34698 8782
rect 34561 8738 34698 8740
rect 34328 8724 34359 8725
rect 34474 8665 34511 8735
rect 33952 8664 34293 8665
rect 33682 8647 33720 8656
rect 33877 8659 34293 8664
rect 33682 8646 33719 8647
rect 33143 8618 33233 8624
rect 33143 8598 33159 8618
rect 33179 8616 33233 8618
rect 33179 8598 33204 8616
rect 33143 8596 33204 8598
rect 33224 8596 33233 8616
rect 33143 8590 33233 8596
rect 33156 8536 33193 8537
rect 33252 8536 33289 8537
rect 33308 8536 33344 8646
rect 33531 8625 33562 8646
rect 33877 8639 33880 8659
rect 33900 8639 34293 8659
rect 34477 8649 34511 8665
rect 34555 8717 34698 8738
rect 34253 8630 34293 8639
rect 34555 8630 34582 8717
rect 34655 8691 34698 8717
rect 34655 8673 34668 8691
rect 34686 8673 34698 8691
rect 34655 8662 34698 8673
rect 33527 8624 33562 8625
rect 33405 8614 33562 8624
rect 33405 8594 33422 8614
rect 33442 8594 33562 8614
rect 33405 8587 33562 8594
rect 33629 8617 33775 8625
rect 33629 8597 33640 8617
rect 33660 8597 33699 8617
rect 33719 8597 33775 8617
rect 34253 8613 34582 8630
rect 34253 8612 34293 8613
rect 33629 8590 33775 8597
rect 34650 8601 34690 8604
rect 34650 8595 34693 8601
rect 34275 8592 34693 8595
rect 33629 8589 33670 8590
rect 33363 8536 33400 8537
rect 33056 8527 33194 8536
rect 33056 8507 33165 8527
rect 33185 8507 33194 8527
rect 33056 8500 33194 8507
rect 33252 8527 33400 8536
rect 33252 8507 33261 8527
rect 33281 8507 33371 8527
rect 33391 8507 33400 8527
rect 33056 8498 33152 8500
rect 33252 8497 33400 8507
rect 33459 8527 33496 8537
rect 33459 8507 33467 8527
rect 33487 8507 33496 8527
rect 33308 8496 33344 8497
rect 33156 8437 33193 8438
rect 33459 8437 33496 8507
rect 33531 8536 33562 8587
rect 34275 8574 34666 8592
rect 34684 8574 34693 8592
rect 34275 8572 34693 8574
rect 34275 8564 34302 8572
rect 34543 8569 34693 8572
rect 33855 8558 34023 8559
rect 34274 8558 34302 8564
rect 33855 8542 34302 8558
rect 34650 8564 34693 8569
rect 33581 8536 33618 8537
rect 33531 8527 33618 8536
rect 33531 8507 33589 8527
rect 33609 8507 33618 8527
rect 33531 8497 33618 8507
rect 33677 8527 33714 8537
rect 33677 8507 33685 8527
rect 33705 8507 33714 8527
rect 33531 8496 33562 8497
rect 33155 8436 33496 8437
rect 33677 8436 33714 8507
rect 33080 8431 33496 8436
rect 33080 8411 33083 8431
rect 33103 8411 33496 8431
rect 33527 8412 33714 8436
rect 33855 8532 34299 8542
rect 33855 8530 34023 8532
rect 32955 8332 32997 8377
rect 33855 8352 33882 8530
rect 33922 8492 33986 8504
rect 34262 8500 34299 8532
rect 34325 8531 34516 8553
rect 34480 8529 34516 8531
rect 34480 8500 34517 8529
rect 34650 8508 34690 8564
rect 33922 8491 33957 8492
rect 33899 8486 33957 8491
rect 33899 8466 33902 8486
rect 33922 8472 33957 8486
rect 33977 8472 33986 8492
rect 33922 8464 33986 8472
rect 33948 8463 33986 8464
rect 33949 8462 33986 8463
rect 34052 8496 34088 8497
rect 34160 8496 34196 8497
rect 34052 8488 34196 8496
rect 34052 8468 34060 8488
rect 34080 8468 34115 8488
rect 34135 8468 34168 8488
rect 34188 8468 34196 8488
rect 34052 8462 34196 8468
rect 34262 8492 34300 8500
rect 34378 8496 34414 8497
rect 34262 8472 34271 8492
rect 34291 8472 34300 8492
rect 34262 8463 34300 8472
rect 34329 8488 34414 8496
rect 34329 8468 34386 8488
rect 34406 8468 34414 8488
rect 34262 8462 34299 8463
rect 34329 8462 34414 8468
rect 34480 8492 34518 8500
rect 34480 8472 34489 8492
rect 34509 8472 34518 8492
rect 34650 8490 34662 8508
rect 34680 8490 34690 8508
rect 34650 8480 34690 8490
rect 34480 8463 34518 8472
rect 34480 8462 34517 8463
rect 33941 8434 34031 8440
rect 33941 8414 33957 8434
rect 33977 8432 34031 8434
rect 33977 8414 34002 8432
rect 33941 8412 34002 8414
rect 34022 8412 34031 8432
rect 33941 8406 34031 8412
rect 33954 8352 33991 8353
rect 34050 8352 34087 8353
rect 34106 8352 34142 8462
rect 34329 8441 34360 8462
rect 34325 8440 34360 8441
rect 34203 8430 34360 8440
rect 34203 8410 34220 8430
rect 34240 8410 34360 8430
rect 34203 8403 34360 8410
rect 34427 8433 34576 8441
rect 34427 8413 34438 8433
rect 34458 8413 34497 8433
rect 34517 8413 34576 8433
rect 34427 8406 34576 8413
rect 34642 8409 34694 8427
rect 34427 8405 34468 8406
rect 34161 8352 34198 8353
rect 33854 8343 33992 8352
rect 33326 8332 33359 8334
rect 32955 8320 33402 8332
rect 32187 8198 32355 8200
rect 31911 8172 32355 8198
rect 31421 8150 31559 8159
rect 31215 8149 31252 8150
rect 30712 8095 30749 8098
rect 30945 8096 30986 8097
rect 29068 8073 29099 8074
rect 28692 8013 29033 8014
rect 29214 8013 29251 8084
rect 30837 8089 30986 8096
rect 30281 8076 30318 8081
rect 30272 8072 30319 8076
rect 30272 8054 30291 8072
rect 30309 8054 30319 8072
rect 30837 8069 30896 8089
rect 30916 8069 30955 8089
rect 30975 8069 30986 8089
rect 30837 8061 30986 8069
rect 31053 8092 31210 8099
rect 31053 8072 31173 8092
rect 31193 8072 31210 8092
rect 31053 8062 31210 8072
rect 31053 8061 31088 8062
rect 28617 8008 29033 8013
rect 28617 7988 28620 8008
rect 28640 7988 29033 8008
rect 29064 7989 29251 8013
rect 29876 8011 29916 8016
rect 30272 8011 30319 8054
rect 31053 8040 31084 8061
rect 31271 8040 31307 8150
rect 31326 8149 31363 8150
rect 31422 8149 31459 8150
rect 31382 8090 31472 8096
rect 31382 8070 31391 8090
rect 31411 8088 31472 8090
rect 31411 8070 31436 8088
rect 31382 8068 31436 8070
rect 31456 8068 31472 8088
rect 31382 8062 31472 8068
rect 30896 8039 30933 8040
rect 29876 7972 30319 8011
rect 30709 8031 30746 8033
rect 30709 8023 30751 8031
rect 30709 8005 30719 8023
rect 30737 8005 30751 8023
rect 30709 7996 30751 8005
rect 30895 8030 30933 8039
rect 30895 8010 30904 8030
rect 30924 8010 30933 8030
rect 30895 8002 30933 8010
rect 30999 8034 31084 8040
rect 31114 8039 31151 8040
rect 30999 8014 31007 8034
rect 31027 8014 31084 8034
rect 30999 8006 31084 8014
rect 31113 8030 31151 8039
rect 31113 8010 31122 8030
rect 31142 8010 31151 8030
rect 30999 8005 31035 8006
rect 31113 8002 31151 8010
rect 31217 8038 31361 8040
rect 31217 8034 31269 8038
rect 31217 8014 31225 8034
rect 31245 8018 31269 8034
rect 31289 8034 31361 8038
rect 31289 8018 31333 8034
rect 31245 8014 31333 8018
rect 31353 8014 31361 8034
rect 31217 8006 31361 8014
rect 31217 8005 31253 8006
rect 31325 8005 31361 8006
rect 31427 8039 31464 8040
rect 31427 8038 31465 8039
rect 31427 8030 31491 8038
rect 31427 8010 31436 8030
rect 31456 8016 31491 8030
rect 31511 8016 31514 8036
rect 31456 8011 31514 8016
rect 31456 8010 31491 8011
rect 27657 7913 27665 7935
rect 27689 7913 27697 7935
rect 27657 7905 27697 7913
rect 28970 7957 29010 7965
rect 28970 7935 28978 7957
rect 29002 7935 29010 7957
rect 25163 7860 25198 7861
rect 25140 7855 25198 7860
rect 25140 7835 25143 7855
rect 25163 7841 25198 7855
rect 25218 7841 25227 7861
rect 25163 7833 25227 7841
rect 25189 7832 25227 7833
rect 25190 7831 25227 7832
rect 25293 7865 25329 7866
rect 25401 7865 25437 7866
rect 25293 7857 25437 7865
rect 25293 7837 25301 7857
rect 25321 7853 25409 7857
rect 25321 7837 25365 7853
rect 25293 7833 25365 7837
rect 25385 7837 25409 7853
rect 25429 7837 25437 7857
rect 25385 7833 25437 7837
rect 25293 7831 25437 7833
rect 25503 7861 25541 7869
rect 25619 7865 25655 7866
rect 25503 7841 25512 7861
rect 25532 7841 25541 7861
rect 25503 7832 25541 7841
rect 25570 7857 25655 7865
rect 25570 7837 25627 7857
rect 25647 7837 25655 7857
rect 25503 7831 25540 7832
rect 25570 7831 25655 7837
rect 25721 7861 25759 7869
rect 25721 7841 25730 7861
rect 25750 7841 25759 7861
rect 25721 7832 25759 7841
rect 25903 7866 25945 7875
rect 25903 7848 25917 7866
rect 25935 7848 25945 7866
rect 25903 7840 25945 7848
rect 25908 7838 25945 7840
rect 26348 7859 26791 7898
rect 25721 7831 25758 7832
rect 25182 7803 25272 7809
rect 25182 7783 25198 7803
rect 25218 7801 25272 7803
rect 25218 7783 25243 7801
rect 25182 7781 25243 7783
rect 25263 7781 25272 7801
rect 25182 7775 25272 7781
rect 25195 7721 25232 7722
rect 25291 7721 25328 7722
rect 25347 7721 25383 7831
rect 25570 7810 25601 7831
rect 26348 7816 26395 7859
rect 26751 7854 26791 7859
rect 27416 7857 27603 7881
rect 27634 7862 28027 7882
rect 28047 7862 28050 7882
rect 27634 7857 28050 7862
rect 25566 7809 25601 7810
rect 25444 7799 25601 7809
rect 25444 7779 25461 7799
rect 25481 7779 25601 7799
rect 25444 7772 25601 7779
rect 25668 7802 25817 7810
rect 25668 7782 25679 7802
rect 25699 7782 25738 7802
rect 25758 7782 25817 7802
rect 26348 7798 26358 7816
rect 26376 7798 26395 7816
rect 26348 7794 26395 7798
rect 26349 7789 26386 7794
rect 25668 7775 25817 7782
rect 27416 7786 27453 7857
rect 27634 7856 27975 7857
rect 27568 7796 27599 7797
rect 25668 7774 25709 7775
rect 25905 7773 25942 7776
rect 25402 7721 25439 7722
rect 25095 7712 25233 7721
rect 24299 7673 24743 7699
rect 24299 7671 24467 7673
rect 23252 7539 23699 7551
rect 23295 7537 23328 7539
rect 22662 7519 22800 7528
rect 22456 7518 22493 7519
rect 22186 7465 22227 7466
rect 21960 7444 22012 7462
rect 22078 7458 22227 7465
rect 21528 7424 21568 7434
rect 22078 7438 22137 7458
rect 22157 7438 22196 7458
rect 22216 7438 22227 7458
rect 22078 7430 22227 7438
rect 22294 7461 22451 7468
rect 22294 7441 22414 7461
rect 22434 7441 22451 7461
rect 22294 7431 22451 7441
rect 22294 7430 22329 7431
rect 21358 7407 21396 7416
rect 22294 7409 22325 7430
rect 22512 7409 22548 7519
rect 22567 7518 22604 7519
rect 22663 7518 22700 7519
rect 22623 7459 22713 7465
rect 22623 7439 22632 7459
rect 22652 7457 22713 7459
rect 22652 7439 22677 7457
rect 22623 7437 22677 7439
rect 22697 7437 22713 7457
rect 22623 7431 22713 7437
rect 22137 7408 22174 7409
rect 21358 7406 21395 7407
rect 20819 7378 20909 7384
rect 20819 7358 20835 7378
rect 20855 7376 20909 7378
rect 20855 7358 20880 7376
rect 20819 7356 20880 7358
rect 20900 7356 20909 7376
rect 20819 7350 20909 7356
rect 20832 7296 20869 7297
rect 20928 7296 20965 7297
rect 20984 7296 21020 7406
rect 21207 7385 21238 7406
rect 22136 7399 22174 7408
rect 21203 7384 21238 7385
rect 21081 7374 21238 7384
rect 21081 7354 21098 7374
rect 21118 7354 21238 7374
rect 21081 7347 21238 7354
rect 21305 7377 21454 7385
rect 21305 7357 21316 7377
rect 21336 7357 21375 7377
rect 21395 7357 21454 7377
rect 21964 7381 22004 7391
rect 21305 7350 21454 7357
rect 21520 7353 21572 7371
rect 21305 7349 21346 7350
rect 21039 7296 21076 7297
rect 20732 7287 20870 7296
rect 19799 7279 19836 7280
rect 19770 7278 19938 7279
rect 20064 7278 20104 7280
rect 19595 7269 19634 7275
rect 19595 7247 19603 7269
rect 19627 7247 19634 7269
rect 19297 7140 19334 7148
rect 19297 7121 19305 7140
rect 19326 7121 19334 7140
rect 19297 7115 19334 7121
rect 18899 6870 18907 6892
rect 18931 6870 18939 6892
rect 18899 6862 18939 6870
rect 17071 6826 17108 6827
rect 16532 6798 16622 6804
rect 16532 6778 16548 6798
rect 16568 6796 16622 6798
rect 16568 6778 16593 6796
rect 16532 6776 16593 6778
rect 16613 6776 16622 6796
rect 16532 6770 16622 6776
rect 16545 6716 16582 6717
rect 16641 6716 16678 6717
rect 16697 6716 16733 6826
rect 16920 6805 16951 6826
rect 17587 6824 18032 6854
rect 19070 6837 19135 6838
rect 17587 6821 18010 6824
rect 16916 6804 16951 6805
rect 16794 6794 16951 6804
rect 16794 6774 16811 6794
rect 16831 6774 16951 6794
rect 16794 6767 16951 6774
rect 17018 6797 17167 6805
rect 17018 6777 17029 6797
rect 17049 6777 17088 6797
rect 17108 6777 17167 6797
rect 17018 6770 17167 6777
rect 17587 6773 17634 6821
rect 17018 6769 17059 6770
rect 17255 6768 17292 6771
rect 16752 6716 16789 6717
rect 16445 6707 16583 6716
rect 15649 6668 16093 6694
rect 15649 6666 15817 6668
rect 15649 6488 15676 6666
rect 15716 6628 15780 6640
rect 16056 6636 16093 6668
rect 16119 6667 16310 6689
rect 16445 6687 16554 6707
rect 16574 6687 16583 6707
rect 16445 6680 16583 6687
rect 16641 6707 16789 6716
rect 16641 6687 16650 6707
rect 16670 6687 16760 6707
rect 16780 6687 16789 6707
rect 16445 6678 16541 6680
rect 16641 6677 16789 6687
rect 16848 6707 16885 6717
rect 16848 6687 16856 6707
rect 16876 6687 16885 6707
rect 16697 6676 16733 6677
rect 16274 6665 16310 6667
rect 16274 6636 16311 6665
rect 15716 6627 15751 6628
rect 15693 6622 15751 6627
rect 15693 6602 15696 6622
rect 15716 6608 15751 6622
rect 15771 6608 15780 6628
rect 15716 6602 15780 6608
rect 15693 6600 15780 6602
rect 15693 6596 15720 6600
rect 15742 6599 15780 6600
rect 15743 6598 15780 6599
rect 15846 6632 15882 6633
rect 15954 6632 15990 6633
rect 15846 6625 15990 6632
rect 15846 6624 15908 6625
rect 15846 6604 15854 6624
rect 15874 6607 15908 6624
rect 15927 6624 15990 6625
rect 15927 6607 15962 6624
rect 15874 6604 15962 6607
rect 15982 6604 15990 6624
rect 15846 6598 15990 6604
rect 16056 6628 16094 6636
rect 16172 6632 16208 6633
rect 16056 6608 16065 6628
rect 16085 6608 16094 6628
rect 16056 6599 16094 6608
rect 16123 6624 16208 6632
rect 16123 6604 16180 6624
rect 16200 6604 16208 6624
rect 16056 6598 16093 6599
rect 16123 6598 16208 6604
rect 16274 6628 16312 6636
rect 16274 6608 16283 6628
rect 16303 6608 16312 6628
rect 16545 6617 16582 6618
rect 16848 6617 16885 6687
rect 16920 6716 16951 6767
rect 17247 6762 17292 6768
rect 17247 6744 17265 6762
rect 17283 6744 17292 6762
rect 17587 6755 17597 6773
rect 17615 6755 17634 6773
rect 17587 6751 17634 6755
rect 18721 6812 18908 6836
rect 18939 6817 19332 6837
rect 19352 6817 19355 6837
rect 18939 6812 19355 6817
rect 17588 6746 17625 6751
rect 17247 6734 17292 6744
rect 18721 6741 18758 6812
rect 18939 6811 19280 6812
rect 18873 6751 18904 6752
rect 16970 6716 17007 6717
rect 16920 6707 17007 6716
rect 16920 6687 16978 6707
rect 16998 6687 17007 6707
rect 16920 6677 17007 6687
rect 17066 6707 17103 6717
rect 17066 6687 17074 6707
rect 17094 6687 17103 6707
rect 17247 6692 17290 6734
rect 18721 6721 18730 6741
rect 18750 6721 18758 6741
rect 18721 6711 18758 6721
rect 18817 6741 18904 6751
rect 18817 6721 18826 6741
rect 18846 6721 18904 6741
rect 18817 6712 18904 6721
rect 18817 6711 18854 6712
rect 17153 6690 17290 6692
rect 16920 6676 16951 6677
rect 17066 6617 17103 6687
rect 16544 6616 16885 6617
rect 16274 6599 16312 6608
rect 16469 6611 16885 6616
rect 16274 6598 16311 6599
rect 15735 6570 15825 6576
rect 15735 6550 15751 6570
rect 15771 6568 15825 6570
rect 15771 6550 15796 6568
rect 15735 6548 15796 6550
rect 15816 6548 15825 6568
rect 15735 6542 15825 6548
rect 15748 6488 15785 6489
rect 15844 6488 15881 6489
rect 15900 6488 15936 6598
rect 16123 6577 16154 6598
rect 16469 6591 16472 6611
rect 16492 6591 16885 6611
rect 17069 6601 17103 6617
rect 17147 6669 17290 6690
rect 17576 6684 17628 6686
rect 16845 6582 16885 6591
rect 17147 6582 17174 6669
rect 17247 6643 17290 6669
rect 17247 6625 17260 6643
rect 17278 6625 17290 6643
rect 17574 6680 18007 6684
rect 17574 6674 18013 6680
rect 17574 6656 17595 6674
rect 17613 6656 18013 6674
rect 18873 6661 18904 6712
rect 18939 6741 18976 6811
rect 19242 6810 19279 6811
rect 19091 6751 19127 6752
rect 18939 6721 18948 6741
rect 18968 6721 18976 6741
rect 18939 6711 18976 6721
rect 19035 6741 19183 6751
rect 19283 6748 19379 6750
rect 19035 6721 19044 6741
rect 19064 6721 19154 6741
rect 19174 6721 19183 6741
rect 19035 6712 19183 6721
rect 19241 6741 19379 6748
rect 19241 6721 19250 6741
rect 19270 6721 19379 6741
rect 19241 6712 19379 6721
rect 19035 6711 19072 6712
rect 18765 6658 18806 6659
rect 17574 6638 18013 6656
rect 17247 6614 17290 6625
rect 16119 6576 16154 6577
rect 15997 6566 16154 6576
rect 15997 6546 16014 6566
rect 16034 6546 16154 6566
rect 15997 6539 16154 6546
rect 16221 6569 16367 6577
rect 16221 6549 16232 6569
rect 16252 6549 16291 6569
rect 16311 6549 16367 6569
rect 16845 6565 17174 6582
rect 16845 6564 16885 6565
rect 16221 6542 16367 6549
rect 17242 6553 17282 6556
rect 17242 6547 17285 6553
rect 16867 6544 17285 6547
rect 16221 6541 16262 6542
rect 15955 6488 15992 6489
rect 15648 6479 15786 6488
rect 15648 6459 15757 6479
rect 15777 6459 15786 6479
rect 15648 6452 15786 6459
rect 15844 6479 15992 6488
rect 15844 6459 15853 6479
rect 15873 6459 15963 6479
rect 15983 6459 15992 6479
rect 15648 6450 15744 6452
rect 15844 6449 15992 6459
rect 16051 6479 16088 6489
rect 16051 6459 16059 6479
rect 16079 6459 16088 6479
rect 15900 6448 15936 6449
rect 15748 6389 15785 6390
rect 16051 6389 16088 6459
rect 16123 6488 16154 6539
rect 16867 6526 17258 6544
rect 17276 6526 17285 6544
rect 16867 6524 17285 6526
rect 16867 6516 16894 6524
rect 17135 6521 17285 6524
rect 16447 6510 16615 6511
rect 16866 6510 16894 6516
rect 16447 6494 16894 6510
rect 17242 6516 17285 6521
rect 16173 6488 16210 6489
rect 16123 6479 16210 6488
rect 16123 6459 16181 6479
rect 16201 6459 16210 6479
rect 16123 6449 16210 6459
rect 16269 6479 16306 6489
rect 16269 6459 16277 6479
rect 16297 6459 16306 6479
rect 16123 6448 16154 6449
rect 15747 6388 16088 6389
rect 16269 6388 16306 6459
rect 15672 6383 16088 6388
rect 15672 6363 15675 6383
rect 15695 6363 16088 6383
rect 16119 6364 16306 6388
rect 16447 6484 16891 6494
rect 16447 6482 16615 6484
rect 15547 6284 15589 6329
rect 16447 6304 16474 6482
rect 16514 6444 16578 6456
rect 16854 6452 16891 6484
rect 16917 6483 17108 6505
rect 17072 6481 17108 6483
rect 17072 6452 17109 6481
rect 17242 6460 17282 6516
rect 16514 6443 16549 6444
rect 16491 6438 16549 6443
rect 16491 6418 16494 6438
rect 16514 6424 16549 6438
rect 16569 6424 16578 6444
rect 16514 6416 16578 6424
rect 16540 6415 16578 6416
rect 16541 6414 16578 6415
rect 16644 6448 16680 6449
rect 16752 6448 16788 6449
rect 16644 6440 16788 6448
rect 16644 6420 16652 6440
rect 16672 6420 16707 6440
rect 16727 6420 16760 6440
rect 16780 6420 16788 6440
rect 16644 6414 16788 6420
rect 16854 6444 16892 6452
rect 16970 6448 17006 6449
rect 16854 6424 16863 6444
rect 16883 6424 16892 6444
rect 16854 6415 16892 6424
rect 16921 6440 17006 6448
rect 16921 6420 16978 6440
rect 16998 6420 17006 6440
rect 16854 6414 16891 6415
rect 16921 6414 17006 6420
rect 17072 6444 17110 6452
rect 17072 6424 17081 6444
rect 17101 6424 17110 6444
rect 17242 6442 17254 6460
rect 17272 6442 17282 6460
rect 17242 6432 17282 6442
rect 17576 6449 17628 6638
rect 17974 6613 18013 6638
rect 18657 6651 18806 6658
rect 18657 6631 18716 6651
rect 18736 6631 18775 6651
rect 18795 6631 18806 6651
rect 18657 6623 18806 6631
rect 18873 6654 19030 6661
rect 18873 6634 18993 6654
rect 19013 6634 19030 6654
rect 18873 6624 19030 6634
rect 18873 6623 18908 6624
rect 17758 6588 17945 6612
rect 17974 6593 18369 6613
rect 18389 6593 18392 6613
rect 18873 6602 18904 6623
rect 19091 6602 19127 6712
rect 19146 6711 19183 6712
rect 19242 6711 19279 6712
rect 19202 6652 19292 6658
rect 19202 6632 19211 6652
rect 19231 6650 19292 6652
rect 19231 6632 19256 6650
rect 19202 6630 19256 6632
rect 19276 6630 19292 6650
rect 19202 6624 19292 6630
rect 18716 6601 18753 6602
rect 17974 6588 18392 6593
rect 18715 6592 18753 6601
rect 17758 6517 17795 6588
rect 17974 6587 18317 6588
rect 17974 6584 18013 6587
rect 18279 6586 18316 6587
rect 17910 6527 17941 6528
rect 17758 6497 17767 6517
rect 17787 6497 17795 6517
rect 17758 6487 17795 6497
rect 17854 6517 17941 6527
rect 17854 6497 17863 6517
rect 17883 6497 17941 6517
rect 17854 6488 17941 6497
rect 17854 6487 17891 6488
rect 17072 6415 17110 6424
rect 17576 6431 17592 6449
rect 17610 6431 17628 6449
rect 17910 6437 17941 6488
rect 17976 6517 18013 6584
rect 18715 6572 18724 6592
rect 18744 6572 18753 6592
rect 18715 6564 18753 6572
rect 18819 6596 18904 6602
rect 18934 6601 18971 6602
rect 18819 6576 18827 6596
rect 18847 6576 18904 6596
rect 18819 6568 18904 6576
rect 18933 6592 18971 6601
rect 18933 6572 18942 6592
rect 18962 6572 18971 6592
rect 18819 6567 18855 6568
rect 18933 6564 18971 6572
rect 19037 6596 19181 6602
rect 19037 6576 19045 6596
rect 19065 6595 19153 6596
rect 19065 6577 19100 6595
rect 19118 6577 19153 6595
rect 19065 6576 19153 6577
rect 19173 6576 19181 6596
rect 19037 6568 19181 6576
rect 19037 6567 19073 6568
rect 19145 6567 19181 6568
rect 19247 6601 19284 6602
rect 19247 6600 19285 6601
rect 19247 6592 19311 6600
rect 19247 6572 19256 6592
rect 19276 6578 19311 6592
rect 19331 6578 19334 6598
rect 19276 6573 19334 6578
rect 19276 6572 19311 6573
rect 18716 6535 18753 6564
rect 18717 6533 18753 6535
rect 18128 6527 18164 6528
rect 17976 6497 17985 6517
rect 18005 6497 18013 6517
rect 17976 6487 18013 6497
rect 18072 6517 18220 6527
rect 18320 6524 18416 6526
rect 18072 6497 18081 6517
rect 18101 6497 18191 6517
rect 18211 6497 18220 6517
rect 18072 6488 18220 6497
rect 18278 6517 18416 6524
rect 18278 6497 18287 6517
rect 18307 6497 18416 6517
rect 18717 6511 18908 6533
rect 18934 6532 18971 6564
rect 19247 6560 19311 6572
rect 19351 6536 19378 6712
rect 19297 6534 19378 6536
rect 19210 6532 19378 6534
rect 18934 6506 19378 6532
rect 19044 6504 19084 6506
rect 19210 6505 19378 6506
rect 18278 6488 18416 6497
rect 19319 6503 19378 6505
rect 18072 6487 18109 6488
rect 17802 6434 17843 6435
rect 17072 6414 17109 6415
rect 16533 6386 16623 6392
rect 16533 6366 16549 6386
rect 16569 6384 16623 6386
rect 16569 6366 16594 6384
rect 16533 6364 16594 6366
rect 16614 6364 16623 6384
rect 16533 6358 16623 6364
rect 16546 6304 16583 6305
rect 16642 6304 16679 6305
rect 16698 6304 16734 6414
rect 16921 6393 16952 6414
rect 17576 6413 17628 6431
rect 17694 6427 17843 6434
rect 17694 6407 17753 6427
rect 17773 6407 17812 6427
rect 17832 6407 17843 6427
rect 17694 6399 17843 6407
rect 17910 6430 18067 6437
rect 17910 6410 18030 6430
rect 18050 6410 18067 6430
rect 17910 6400 18067 6410
rect 17910 6399 17945 6400
rect 16917 6392 16952 6393
rect 16795 6382 16952 6392
rect 16795 6362 16812 6382
rect 16832 6362 16952 6382
rect 16795 6355 16952 6362
rect 17019 6385 17168 6393
rect 17019 6365 17030 6385
rect 17050 6365 17089 6385
rect 17109 6365 17168 6385
rect 17019 6358 17168 6365
rect 17234 6361 17286 6379
rect 17910 6378 17941 6399
rect 18128 6378 18164 6488
rect 18183 6487 18220 6488
rect 18279 6487 18316 6488
rect 18239 6428 18329 6434
rect 18239 6408 18248 6428
rect 18268 6426 18329 6428
rect 18268 6408 18293 6426
rect 18239 6406 18293 6408
rect 18313 6406 18329 6426
rect 18239 6400 18329 6406
rect 17753 6377 17790 6378
rect 17019 6357 17060 6358
rect 16753 6304 16790 6305
rect 16446 6295 16584 6304
rect 15918 6284 15951 6286
rect 15547 6272 15994 6284
rect 15550 6258 15994 6272
rect 15550 6256 15718 6258
rect 15550 6078 15577 6256
rect 15617 6218 15681 6230
rect 15957 6226 15994 6258
rect 16020 6257 16211 6279
rect 16446 6275 16555 6295
rect 16575 6275 16584 6295
rect 16446 6268 16584 6275
rect 16642 6295 16790 6304
rect 16642 6275 16651 6295
rect 16671 6275 16761 6295
rect 16781 6275 16790 6295
rect 16446 6266 16542 6268
rect 16642 6265 16790 6275
rect 16849 6295 16886 6305
rect 16849 6275 16857 6295
rect 16877 6275 16886 6295
rect 16698 6264 16734 6265
rect 16175 6255 16211 6257
rect 16175 6226 16212 6255
rect 15617 6217 15652 6218
rect 15594 6212 15652 6217
rect 15594 6192 15597 6212
rect 15617 6198 15652 6212
rect 15672 6198 15681 6218
rect 15617 6190 15681 6198
rect 15643 6189 15681 6190
rect 15644 6188 15681 6189
rect 15747 6222 15783 6223
rect 15855 6222 15891 6223
rect 15747 6214 15891 6222
rect 15747 6194 15755 6214
rect 15775 6212 15863 6214
rect 15775 6194 15808 6212
rect 15747 6193 15808 6194
rect 15829 6194 15863 6212
rect 15883 6194 15891 6214
rect 15829 6193 15891 6194
rect 15747 6188 15891 6193
rect 15957 6218 15995 6226
rect 16073 6222 16109 6223
rect 15957 6198 15966 6218
rect 15986 6198 15995 6218
rect 15957 6189 15995 6198
rect 16024 6214 16109 6222
rect 16024 6194 16081 6214
rect 16101 6194 16109 6214
rect 15957 6188 15994 6189
rect 16024 6188 16109 6194
rect 16175 6218 16213 6226
rect 16175 6198 16184 6218
rect 16204 6198 16213 6218
rect 16849 6208 16886 6275
rect 16921 6304 16952 6355
rect 17234 6343 17252 6361
rect 17270 6343 17286 6361
rect 17752 6368 17790 6377
rect 16971 6304 17008 6305
rect 16921 6295 17008 6304
rect 16921 6275 16979 6295
rect 16999 6275 17008 6295
rect 16921 6265 17008 6275
rect 17067 6295 17104 6305
rect 17067 6275 17075 6295
rect 17095 6275 17104 6295
rect 16921 6264 16952 6265
rect 16546 6205 16583 6206
rect 16849 6205 16888 6208
rect 16545 6204 16888 6205
rect 17067 6204 17104 6275
rect 16175 6189 16213 6198
rect 16470 6199 16888 6204
rect 16175 6188 16212 6189
rect 15636 6160 15726 6166
rect 15636 6140 15652 6160
rect 15672 6158 15726 6160
rect 15672 6140 15697 6158
rect 15636 6138 15697 6140
rect 15717 6138 15726 6158
rect 15636 6132 15726 6138
rect 15649 6078 15686 6079
rect 15745 6078 15782 6079
rect 15801 6078 15837 6188
rect 16024 6167 16055 6188
rect 16470 6179 16473 6199
rect 16493 6179 16888 6199
rect 16917 6180 17104 6204
rect 16020 6166 16055 6167
rect 15898 6156 16055 6166
rect 15898 6136 15915 6156
rect 15935 6136 16055 6156
rect 15898 6129 16055 6136
rect 16122 6159 16271 6167
rect 16122 6139 16133 6159
rect 16153 6139 16192 6159
rect 16212 6139 16271 6159
rect 16122 6132 16271 6139
rect 16849 6154 16888 6179
rect 17234 6154 17286 6343
rect 17580 6350 17620 6360
rect 17580 6332 17590 6350
rect 17608 6332 17620 6350
rect 17752 6348 17761 6368
rect 17781 6348 17790 6368
rect 17752 6340 17790 6348
rect 17856 6372 17941 6378
rect 17971 6377 18008 6378
rect 17856 6352 17864 6372
rect 17884 6352 17941 6372
rect 17856 6344 17941 6352
rect 17970 6368 18008 6377
rect 17970 6348 17979 6368
rect 17999 6348 18008 6368
rect 17856 6343 17892 6344
rect 17970 6340 18008 6348
rect 18074 6372 18218 6378
rect 18074 6352 18082 6372
rect 18102 6352 18135 6372
rect 18155 6352 18190 6372
rect 18210 6352 18218 6372
rect 18074 6344 18218 6352
rect 18074 6343 18110 6344
rect 18182 6343 18218 6344
rect 18284 6377 18321 6378
rect 18284 6376 18322 6377
rect 18284 6368 18348 6376
rect 18284 6348 18293 6368
rect 18313 6354 18348 6368
rect 18368 6354 18371 6374
rect 18313 6349 18371 6354
rect 18313 6348 18348 6349
rect 17580 6276 17620 6332
rect 17753 6311 17790 6340
rect 17754 6309 17790 6311
rect 17754 6287 17945 6309
rect 17971 6308 18008 6340
rect 18284 6336 18348 6348
rect 18388 6310 18415 6488
rect 19319 6485 19348 6503
rect 18247 6308 18415 6310
rect 17971 6298 18415 6308
rect 18556 6404 18743 6428
rect 18774 6409 19167 6429
rect 19187 6409 19190 6429
rect 18774 6404 19190 6409
rect 18556 6333 18593 6404
rect 18774 6403 19115 6404
rect 18708 6343 18739 6344
rect 18556 6313 18565 6333
rect 18585 6313 18593 6333
rect 18556 6303 18593 6313
rect 18652 6333 18739 6343
rect 18652 6313 18661 6333
rect 18681 6313 18739 6333
rect 18652 6304 18739 6313
rect 18652 6303 18689 6304
rect 17577 6271 17620 6276
rect 17968 6282 18415 6298
rect 17968 6276 17996 6282
rect 18247 6281 18415 6282
rect 17577 6268 17727 6271
rect 17968 6268 17995 6276
rect 17577 6266 17995 6268
rect 17577 6248 17586 6266
rect 17604 6248 17995 6266
rect 18708 6253 18739 6304
rect 18774 6333 18811 6403
rect 19077 6402 19114 6403
rect 18926 6343 18962 6344
rect 18774 6313 18783 6333
rect 18803 6313 18811 6333
rect 18774 6303 18811 6313
rect 18870 6333 19018 6343
rect 19118 6340 19214 6342
rect 18870 6313 18879 6333
rect 18899 6313 18989 6333
rect 19009 6313 19018 6333
rect 18870 6304 19018 6313
rect 19076 6333 19214 6340
rect 19076 6313 19085 6333
rect 19105 6313 19214 6333
rect 19076 6304 19214 6313
rect 18870 6303 18907 6304
rect 18600 6250 18641 6251
rect 17577 6245 17995 6248
rect 17577 6239 17620 6245
rect 17580 6236 17620 6239
rect 18492 6243 18641 6250
rect 17977 6227 18017 6228
rect 17688 6210 18017 6227
rect 18492 6223 18551 6243
rect 18571 6223 18610 6243
rect 18630 6223 18641 6243
rect 18492 6215 18641 6223
rect 18708 6246 18865 6253
rect 18708 6226 18828 6246
rect 18848 6226 18865 6246
rect 18708 6216 18865 6226
rect 18708 6215 18743 6216
rect 17572 6167 17615 6178
rect 16849 6136 17288 6154
rect 16122 6131 16163 6132
rect 15856 6078 15893 6079
rect 15549 6069 15687 6078
rect 15549 6049 15658 6069
rect 15678 6049 15687 6069
rect 15549 6042 15687 6049
rect 15745 6069 15893 6078
rect 15745 6049 15754 6069
rect 15774 6049 15864 6069
rect 15884 6049 15893 6069
rect 15549 6040 15645 6042
rect 15745 6039 15893 6049
rect 15952 6069 15989 6079
rect 15952 6049 15960 6069
rect 15980 6049 15989 6069
rect 15801 6038 15837 6039
rect 15649 5979 15686 5980
rect 15952 5979 15989 6049
rect 16024 6078 16055 6129
rect 16849 6118 17249 6136
rect 17267 6118 17288 6136
rect 16849 6112 17288 6118
rect 16855 6108 17288 6112
rect 17572 6149 17584 6167
rect 17602 6149 17615 6167
rect 17572 6123 17615 6149
rect 17688 6123 17715 6210
rect 17977 6201 18017 6210
rect 17234 6106 17286 6108
rect 17572 6102 17715 6123
rect 17759 6175 17793 6191
rect 17977 6181 18370 6201
rect 18390 6181 18393 6201
rect 18708 6194 18739 6215
rect 18926 6194 18962 6304
rect 18981 6303 19018 6304
rect 19077 6303 19114 6304
rect 19037 6244 19127 6250
rect 19037 6224 19046 6244
rect 19066 6242 19127 6244
rect 19066 6224 19091 6242
rect 19037 6222 19091 6224
rect 19111 6222 19127 6242
rect 19037 6216 19127 6222
rect 18551 6193 18588 6194
rect 17977 6176 18393 6181
rect 18550 6184 18588 6193
rect 17977 6175 18318 6176
rect 17759 6105 17796 6175
rect 17911 6115 17942 6116
rect 17572 6100 17709 6102
rect 16074 6078 16111 6079
rect 16024 6069 16111 6078
rect 16024 6049 16082 6069
rect 16102 6049 16111 6069
rect 16024 6039 16111 6049
rect 16170 6069 16207 6079
rect 16170 6049 16178 6069
rect 16198 6049 16207 6069
rect 17572 6058 17615 6100
rect 17759 6085 17768 6105
rect 17788 6085 17796 6105
rect 17759 6075 17796 6085
rect 17855 6105 17942 6115
rect 17855 6085 17864 6105
rect 17884 6085 17942 6105
rect 17855 6076 17942 6085
rect 17855 6075 17892 6076
rect 16024 6038 16055 6039
rect 15648 5978 15989 5979
rect 16170 5978 16207 6049
rect 17570 6048 17615 6058
rect 17237 6041 17274 6046
rect 17228 6037 17275 6041
rect 17228 6019 17247 6037
rect 17265 6019 17275 6037
rect 17570 6030 17579 6048
rect 17597 6030 17615 6048
rect 17570 6024 17615 6030
rect 17911 6025 17942 6076
rect 17977 6105 18014 6175
rect 18280 6174 18317 6175
rect 18550 6164 18559 6184
rect 18579 6164 18588 6184
rect 18550 6156 18588 6164
rect 18654 6188 18739 6194
rect 18769 6193 18806 6194
rect 18654 6168 18662 6188
rect 18682 6168 18739 6188
rect 18654 6160 18739 6168
rect 18768 6184 18806 6193
rect 18768 6164 18777 6184
rect 18797 6164 18806 6184
rect 18654 6159 18690 6160
rect 18768 6156 18806 6164
rect 18872 6188 19016 6194
rect 18872 6168 18880 6188
rect 18900 6169 18932 6188
rect 18953 6169 18988 6188
rect 18900 6168 18988 6169
rect 19008 6168 19016 6188
rect 18872 6160 19016 6168
rect 18872 6159 18908 6160
rect 18980 6159 19016 6160
rect 19082 6193 19119 6194
rect 19082 6192 19120 6193
rect 19082 6184 19146 6192
rect 19082 6164 19091 6184
rect 19111 6170 19146 6184
rect 19166 6170 19169 6190
rect 19111 6165 19169 6170
rect 19111 6164 19146 6165
rect 18551 6127 18588 6156
rect 18552 6125 18588 6127
rect 18129 6115 18165 6116
rect 17977 6085 17986 6105
rect 18006 6085 18014 6105
rect 17977 6075 18014 6085
rect 18073 6105 18221 6115
rect 18321 6112 18417 6114
rect 18073 6085 18082 6105
rect 18102 6085 18192 6105
rect 18212 6085 18221 6105
rect 18073 6076 18221 6085
rect 18279 6105 18417 6112
rect 18279 6085 18288 6105
rect 18308 6085 18417 6105
rect 18552 6103 18743 6125
rect 18769 6124 18806 6156
rect 19082 6152 19146 6164
rect 19186 6126 19213 6304
rect 19045 6124 19213 6126
rect 18769 6098 19213 6124
rect 18279 6076 18417 6085
rect 18073 6075 18110 6076
rect 17570 6021 17607 6024
rect 17803 6022 17844 6023
rect 15573 5973 15989 5978
rect 15573 5953 15576 5973
rect 15596 5953 15989 5973
rect 16020 5954 16207 5978
rect 16832 5976 16872 5981
rect 17228 5976 17275 6019
rect 17695 6015 17844 6022
rect 17695 5995 17754 6015
rect 17774 5995 17813 6015
rect 17833 5995 17844 6015
rect 17695 5987 17844 5995
rect 17911 6018 18068 6025
rect 17911 5998 18031 6018
rect 18051 5998 18068 6018
rect 17911 5988 18068 5998
rect 17911 5987 17946 5988
rect 16832 5937 17275 5976
rect 17911 5966 17942 5987
rect 18129 5966 18165 6076
rect 18184 6075 18221 6076
rect 18280 6075 18317 6076
rect 18240 6016 18330 6022
rect 18240 5996 18249 6016
rect 18269 6014 18330 6016
rect 18269 5996 18294 6014
rect 18240 5994 18294 5996
rect 18314 5994 18330 6014
rect 18240 5988 18330 5994
rect 17754 5965 17791 5966
rect 15926 5922 15966 5930
rect 15926 5900 15934 5922
rect 15958 5900 15966 5922
rect 15632 5676 15800 5677
rect 15926 5676 15966 5900
rect 16429 5904 16597 5905
rect 16832 5904 16872 5937
rect 17228 5904 17275 5937
rect 17567 5957 17604 5959
rect 17567 5949 17609 5957
rect 17567 5931 17577 5949
rect 17595 5931 17609 5949
rect 17567 5922 17609 5931
rect 17753 5956 17791 5965
rect 17753 5936 17762 5956
rect 17782 5936 17791 5956
rect 17753 5928 17791 5936
rect 17857 5960 17942 5966
rect 17972 5965 18009 5966
rect 17857 5940 17865 5960
rect 17885 5940 17942 5960
rect 17857 5932 17942 5940
rect 17971 5956 18009 5965
rect 17971 5936 17980 5956
rect 18000 5936 18009 5956
rect 17857 5931 17893 5932
rect 17971 5928 18009 5936
rect 18075 5964 18219 5966
rect 18075 5960 18127 5964
rect 18075 5940 18083 5960
rect 18103 5944 18127 5960
rect 18147 5960 18219 5964
rect 18147 5944 18191 5960
rect 18103 5940 18191 5944
rect 18211 5940 18219 5960
rect 18075 5932 18219 5940
rect 18075 5931 18111 5932
rect 18183 5931 18219 5932
rect 18285 5965 18322 5966
rect 18285 5964 18323 5965
rect 18285 5956 18349 5964
rect 18285 5936 18294 5956
rect 18314 5942 18349 5956
rect 18369 5942 18372 5962
rect 18314 5937 18372 5942
rect 18314 5936 18349 5937
rect 16429 5903 16873 5904
rect 16429 5878 16874 5903
rect 16429 5876 16597 5878
rect 16793 5877 16874 5878
rect 17043 5877 17092 5903
rect 17228 5877 17277 5904
rect 16429 5698 16456 5876
rect 16496 5838 16560 5850
rect 16836 5846 16873 5877
rect 17054 5846 17091 5877
rect 17236 5852 17277 5877
rect 17568 5897 17609 5922
rect 17754 5897 17791 5928
rect 17972 5897 18009 5928
rect 18285 5924 18349 5936
rect 18389 5898 18416 6076
rect 17568 5870 17617 5897
rect 17753 5871 17802 5897
rect 17971 5896 18052 5897
rect 18248 5896 18416 5898
rect 17971 5871 18416 5896
rect 17972 5870 18416 5871
rect 16496 5837 16531 5838
rect 16473 5832 16531 5837
rect 16473 5812 16476 5832
rect 16496 5818 16531 5832
rect 16551 5818 16560 5838
rect 16496 5810 16560 5818
rect 16522 5809 16560 5810
rect 16523 5808 16560 5809
rect 16626 5842 16662 5843
rect 16734 5842 16770 5843
rect 16626 5834 16770 5842
rect 16626 5814 16634 5834
rect 16654 5830 16742 5834
rect 16654 5814 16698 5830
rect 16626 5810 16698 5814
rect 16718 5814 16742 5830
rect 16762 5814 16770 5834
rect 16718 5810 16770 5814
rect 16626 5808 16770 5810
rect 16836 5838 16874 5846
rect 16952 5842 16988 5843
rect 16836 5818 16845 5838
rect 16865 5818 16874 5838
rect 16836 5809 16874 5818
rect 16903 5834 16988 5842
rect 16903 5814 16960 5834
rect 16980 5814 16988 5834
rect 16836 5808 16873 5809
rect 16903 5808 16988 5814
rect 17054 5838 17092 5846
rect 17054 5818 17063 5838
rect 17083 5818 17092 5838
rect 17054 5809 17092 5818
rect 17236 5843 17278 5852
rect 17236 5825 17250 5843
rect 17268 5825 17278 5843
rect 17236 5817 17278 5825
rect 17241 5815 17278 5817
rect 17570 5837 17617 5870
rect 17973 5837 18013 5870
rect 18248 5869 18416 5870
rect 18879 5874 18919 6098
rect 19045 6097 19213 6098
rect 18879 5852 18887 5874
rect 18911 5852 18919 5874
rect 18879 5844 18919 5852
rect 17054 5808 17091 5809
rect 16515 5780 16605 5786
rect 16515 5760 16531 5780
rect 16551 5778 16605 5780
rect 16551 5760 16576 5778
rect 16515 5758 16576 5760
rect 16596 5758 16605 5778
rect 16515 5752 16605 5758
rect 16528 5698 16565 5699
rect 16624 5698 16661 5699
rect 16680 5698 16716 5808
rect 16903 5787 16934 5808
rect 17570 5798 18013 5837
rect 16899 5786 16934 5787
rect 16777 5776 16934 5786
rect 16777 5756 16794 5776
rect 16814 5756 16934 5776
rect 16777 5749 16934 5756
rect 17001 5779 17150 5787
rect 17001 5759 17012 5779
rect 17032 5759 17071 5779
rect 17091 5759 17150 5779
rect 17001 5752 17150 5759
rect 17570 5755 17617 5798
rect 17973 5793 18013 5798
rect 18638 5796 18825 5820
rect 18856 5801 19249 5821
rect 19269 5801 19272 5821
rect 18856 5796 19272 5801
rect 17001 5751 17042 5752
rect 17238 5750 17275 5753
rect 16735 5698 16772 5699
rect 16428 5689 16566 5698
rect 15632 5650 16076 5676
rect 15632 5648 15800 5650
rect 15632 5470 15659 5648
rect 15699 5610 15763 5622
rect 16039 5618 16076 5650
rect 16102 5649 16293 5671
rect 16428 5669 16537 5689
rect 16557 5669 16566 5689
rect 16428 5662 16566 5669
rect 16624 5689 16772 5698
rect 16624 5669 16633 5689
rect 16653 5669 16743 5689
rect 16763 5669 16772 5689
rect 16428 5660 16524 5662
rect 16624 5659 16772 5669
rect 16831 5689 16868 5699
rect 16831 5669 16839 5689
rect 16859 5669 16868 5689
rect 16680 5658 16716 5659
rect 16257 5647 16293 5649
rect 16257 5618 16294 5647
rect 15699 5609 15734 5610
rect 15676 5604 15734 5609
rect 15676 5584 15679 5604
rect 15699 5590 15734 5604
rect 15754 5590 15763 5610
rect 15699 5582 15763 5590
rect 15725 5581 15763 5582
rect 15726 5580 15763 5581
rect 15829 5614 15865 5615
rect 15937 5614 15973 5615
rect 15829 5606 15973 5614
rect 15829 5586 15837 5606
rect 15857 5605 15945 5606
rect 15857 5586 15892 5605
rect 15913 5586 15945 5605
rect 15965 5586 15973 5606
rect 15829 5580 15973 5586
rect 16039 5610 16077 5618
rect 16155 5614 16191 5615
rect 16039 5590 16048 5610
rect 16068 5590 16077 5610
rect 16039 5581 16077 5590
rect 16106 5606 16191 5614
rect 16106 5586 16163 5606
rect 16183 5586 16191 5606
rect 16039 5580 16076 5581
rect 16106 5580 16191 5586
rect 16257 5610 16295 5618
rect 16257 5590 16266 5610
rect 16286 5590 16295 5610
rect 16528 5599 16565 5600
rect 16831 5599 16868 5669
rect 16903 5698 16934 5749
rect 17230 5744 17275 5750
rect 17230 5726 17248 5744
rect 17266 5726 17275 5744
rect 17570 5737 17580 5755
rect 17598 5737 17617 5755
rect 17570 5733 17617 5737
rect 17571 5728 17608 5733
rect 17230 5716 17275 5726
rect 18638 5725 18675 5796
rect 18856 5795 19197 5796
rect 18790 5735 18821 5736
rect 16953 5698 16990 5699
rect 16903 5689 16990 5698
rect 16903 5669 16961 5689
rect 16981 5669 16990 5689
rect 16903 5659 16990 5669
rect 17049 5689 17086 5699
rect 17049 5669 17057 5689
rect 17077 5669 17086 5689
rect 17230 5674 17273 5716
rect 18638 5705 18647 5725
rect 18667 5705 18675 5725
rect 18638 5695 18675 5705
rect 18734 5725 18821 5735
rect 18734 5705 18743 5725
rect 18763 5705 18821 5725
rect 18734 5696 18821 5705
rect 18734 5695 18771 5696
rect 17136 5672 17273 5674
rect 16903 5658 16934 5659
rect 17049 5599 17086 5669
rect 16527 5598 16868 5599
rect 16257 5581 16295 5590
rect 16452 5593 16868 5598
rect 16257 5580 16294 5581
rect 15718 5552 15808 5558
rect 15718 5532 15734 5552
rect 15754 5550 15808 5552
rect 15754 5532 15779 5550
rect 15718 5530 15779 5532
rect 15799 5530 15808 5550
rect 15718 5524 15808 5530
rect 15731 5470 15768 5471
rect 15827 5470 15864 5471
rect 15883 5470 15919 5580
rect 16106 5559 16137 5580
rect 16452 5573 16455 5593
rect 16475 5573 16868 5593
rect 17052 5583 17086 5599
rect 17130 5651 17273 5672
rect 17559 5666 17611 5668
rect 16828 5564 16868 5573
rect 17130 5564 17157 5651
rect 17230 5625 17273 5651
rect 17230 5607 17243 5625
rect 17261 5607 17273 5625
rect 17557 5662 17990 5666
rect 17557 5656 17996 5662
rect 17557 5638 17578 5656
rect 17596 5638 17996 5656
rect 18790 5645 18821 5696
rect 18856 5725 18893 5795
rect 19159 5794 19196 5795
rect 19008 5735 19044 5736
rect 18856 5705 18865 5725
rect 18885 5705 18893 5725
rect 18856 5695 18893 5705
rect 18952 5725 19100 5735
rect 19200 5732 19296 5734
rect 18952 5705 18961 5725
rect 18981 5705 19071 5725
rect 19091 5705 19100 5725
rect 18952 5696 19100 5705
rect 19158 5725 19296 5732
rect 19158 5705 19167 5725
rect 19187 5705 19296 5725
rect 19158 5696 19296 5705
rect 18952 5695 18989 5696
rect 18682 5642 18723 5643
rect 17557 5620 17996 5638
rect 17230 5596 17273 5607
rect 16102 5558 16137 5559
rect 15980 5548 16137 5558
rect 15980 5528 15997 5548
rect 16017 5528 16137 5548
rect 15980 5521 16137 5528
rect 16204 5551 16353 5559
rect 16204 5531 16215 5551
rect 16235 5531 16274 5551
rect 16294 5531 16353 5551
rect 16828 5547 17157 5564
rect 16828 5546 16868 5547
rect 16204 5524 16353 5531
rect 17225 5535 17265 5538
rect 17225 5529 17268 5535
rect 16850 5526 17268 5529
rect 16204 5523 16245 5524
rect 15938 5470 15975 5471
rect 15631 5461 15769 5470
rect 15329 5286 15369 5458
rect 15631 5441 15740 5461
rect 15760 5441 15769 5461
rect 15631 5434 15769 5441
rect 15827 5461 15975 5470
rect 15827 5441 15836 5461
rect 15856 5441 15946 5461
rect 15966 5441 15975 5461
rect 15631 5432 15727 5434
rect 15827 5431 15975 5441
rect 16034 5461 16071 5471
rect 16034 5441 16042 5461
rect 16062 5441 16071 5461
rect 15883 5430 15919 5431
rect 15731 5371 15768 5372
rect 16034 5371 16071 5441
rect 16106 5470 16137 5521
rect 16850 5508 17241 5526
rect 17259 5508 17268 5526
rect 16850 5506 17268 5508
rect 16850 5498 16877 5506
rect 17118 5503 17268 5506
rect 16430 5492 16598 5493
rect 16849 5492 16877 5498
rect 16430 5476 16877 5492
rect 17225 5498 17268 5503
rect 16156 5470 16193 5471
rect 16106 5461 16193 5470
rect 16106 5441 16164 5461
rect 16184 5441 16193 5461
rect 16106 5431 16193 5441
rect 16252 5461 16289 5471
rect 16252 5441 16260 5461
rect 16280 5441 16289 5461
rect 16106 5430 16137 5431
rect 15730 5370 16071 5371
rect 16252 5370 16289 5441
rect 15655 5365 16071 5370
rect 15655 5345 15658 5365
rect 15678 5345 16071 5365
rect 16102 5346 16289 5370
rect 16430 5466 16874 5476
rect 16430 5464 16598 5466
rect 16430 5286 16457 5464
rect 16497 5426 16561 5438
rect 16837 5434 16874 5466
rect 16900 5465 17091 5487
rect 17055 5463 17091 5465
rect 17055 5434 17092 5463
rect 17225 5442 17265 5498
rect 16497 5425 16532 5426
rect 16474 5420 16532 5425
rect 16474 5400 16477 5420
rect 16497 5406 16532 5420
rect 16552 5406 16561 5426
rect 16497 5398 16561 5406
rect 16523 5397 16561 5398
rect 16524 5396 16561 5397
rect 16627 5430 16663 5431
rect 16735 5430 16771 5431
rect 16627 5422 16771 5430
rect 16627 5402 16635 5422
rect 16655 5402 16690 5422
rect 16710 5402 16743 5422
rect 16763 5402 16771 5422
rect 16627 5396 16771 5402
rect 16837 5426 16875 5434
rect 16953 5430 16989 5431
rect 16837 5406 16846 5426
rect 16866 5406 16875 5426
rect 16837 5397 16875 5406
rect 16904 5422 16989 5430
rect 16904 5402 16961 5422
rect 16981 5402 16989 5422
rect 16837 5396 16874 5397
rect 16904 5396 16989 5402
rect 17055 5426 17093 5434
rect 17055 5406 17064 5426
rect 17084 5406 17093 5426
rect 17225 5424 17237 5442
rect 17255 5424 17265 5442
rect 17225 5414 17265 5424
rect 17559 5431 17611 5620
rect 17957 5595 17996 5620
rect 18574 5635 18723 5642
rect 18574 5615 18633 5635
rect 18653 5615 18692 5635
rect 18712 5615 18723 5635
rect 18574 5607 18723 5615
rect 18790 5638 18947 5645
rect 18790 5618 18910 5638
rect 18930 5618 18947 5638
rect 18790 5608 18947 5618
rect 18790 5607 18825 5608
rect 17741 5570 17928 5594
rect 17957 5575 18352 5595
rect 18372 5575 18375 5595
rect 18790 5586 18821 5607
rect 19008 5586 19044 5696
rect 19063 5695 19100 5696
rect 19159 5695 19196 5696
rect 19119 5636 19209 5642
rect 19119 5616 19128 5636
rect 19148 5634 19209 5636
rect 19148 5616 19173 5634
rect 19119 5614 19173 5616
rect 19193 5614 19209 5634
rect 19119 5608 19209 5614
rect 18633 5585 18670 5586
rect 17957 5570 18375 5575
rect 18632 5576 18670 5585
rect 17741 5499 17778 5570
rect 17957 5569 18300 5570
rect 17957 5566 17996 5569
rect 18262 5568 18299 5569
rect 17893 5509 17924 5510
rect 17741 5479 17750 5499
rect 17770 5479 17778 5499
rect 17741 5469 17778 5479
rect 17837 5499 17924 5509
rect 17837 5479 17846 5499
rect 17866 5479 17924 5499
rect 17837 5470 17924 5479
rect 17837 5469 17874 5470
rect 17055 5397 17093 5406
rect 17559 5413 17575 5431
rect 17593 5413 17611 5431
rect 17893 5419 17924 5470
rect 17959 5499 17996 5566
rect 18632 5556 18641 5576
rect 18661 5556 18670 5576
rect 18632 5548 18670 5556
rect 18736 5580 18821 5586
rect 18851 5585 18888 5586
rect 18736 5560 18744 5580
rect 18764 5560 18821 5580
rect 18736 5552 18821 5560
rect 18850 5576 18888 5585
rect 18850 5556 18859 5576
rect 18879 5556 18888 5576
rect 18736 5551 18772 5552
rect 18850 5548 18888 5556
rect 18954 5580 19098 5586
rect 18954 5560 18962 5580
rect 18982 5575 19070 5580
rect 18982 5560 19018 5575
rect 18954 5558 19018 5560
rect 19037 5560 19070 5575
rect 19090 5560 19098 5580
rect 19037 5558 19098 5560
rect 18954 5552 19098 5558
rect 18954 5551 18990 5552
rect 19062 5551 19098 5552
rect 19164 5585 19201 5586
rect 19164 5584 19202 5585
rect 19164 5576 19228 5584
rect 19164 5556 19173 5576
rect 19193 5562 19228 5576
rect 19248 5562 19251 5582
rect 19193 5557 19251 5562
rect 19193 5556 19228 5557
rect 18633 5519 18670 5548
rect 18634 5517 18670 5519
rect 18111 5509 18147 5510
rect 17959 5479 17968 5499
rect 17988 5479 17996 5499
rect 17959 5469 17996 5479
rect 18055 5499 18203 5509
rect 18303 5506 18399 5508
rect 18055 5479 18064 5499
rect 18084 5479 18174 5499
rect 18194 5479 18203 5499
rect 18055 5470 18203 5479
rect 18261 5499 18399 5506
rect 18261 5479 18270 5499
rect 18290 5479 18399 5499
rect 18634 5495 18825 5517
rect 18851 5516 18888 5548
rect 19164 5544 19228 5556
rect 19268 5518 19295 5696
rect 19127 5516 19295 5518
rect 18851 5502 19295 5516
rect 19319 5539 19347 6485
rect 19319 5509 19364 5539
rect 18851 5490 19298 5502
rect 18894 5488 18927 5490
rect 18261 5470 18399 5479
rect 18055 5469 18092 5470
rect 17785 5416 17826 5417
rect 17055 5396 17092 5397
rect 16516 5368 16606 5374
rect 16516 5348 16532 5368
rect 16552 5366 16606 5368
rect 16552 5348 16577 5366
rect 16516 5346 16577 5348
rect 16597 5346 16606 5366
rect 16516 5340 16606 5346
rect 16529 5286 16566 5287
rect 16625 5286 16662 5287
rect 16681 5286 16717 5396
rect 16904 5375 16935 5396
rect 17559 5395 17611 5413
rect 17677 5409 17826 5416
rect 17677 5389 17736 5409
rect 17756 5389 17795 5409
rect 17815 5389 17826 5409
rect 17677 5381 17826 5389
rect 17893 5412 18050 5419
rect 17893 5392 18013 5412
rect 18033 5392 18050 5412
rect 17893 5382 18050 5392
rect 17893 5381 17928 5382
rect 16900 5374 16935 5375
rect 16778 5364 16935 5374
rect 16778 5344 16795 5364
rect 16815 5344 16935 5364
rect 16778 5337 16935 5344
rect 17002 5367 17151 5375
rect 17002 5347 17013 5367
rect 17033 5347 17072 5367
rect 17092 5347 17151 5367
rect 17002 5340 17151 5347
rect 17217 5343 17269 5361
rect 17893 5360 17924 5381
rect 18111 5360 18147 5470
rect 18166 5469 18203 5470
rect 18262 5469 18299 5470
rect 18222 5410 18312 5416
rect 18222 5390 18231 5410
rect 18251 5408 18312 5410
rect 18251 5390 18276 5408
rect 18222 5388 18276 5390
rect 18296 5388 18312 5408
rect 18222 5382 18312 5388
rect 17736 5359 17773 5360
rect 17002 5339 17043 5340
rect 16736 5286 16773 5287
rect 15330 5271 15369 5286
rect 16429 5277 16567 5286
rect 15330 5270 15496 5271
rect 15622 5270 15662 5272
rect 15330 5244 15772 5270
rect 15330 5242 15496 5244
rect 14994 5130 15031 5138
rect 14994 5111 15002 5130
rect 15023 5111 15031 5130
rect 14994 5105 15031 5111
rect 15330 5064 15355 5242
rect 15395 5204 15459 5216
rect 15735 5212 15772 5244
rect 15798 5243 15989 5265
rect 16429 5257 16538 5277
rect 16558 5257 16567 5277
rect 16429 5250 16567 5257
rect 16625 5277 16773 5286
rect 16625 5257 16634 5277
rect 16654 5257 16744 5277
rect 16764 5257 16773 5277
rect 16429 5248 16525 5250
rect 16625 5247 16773 5257
rect 16832 5277 16869 5287
rect 16832 5257 16840 5277
rect 16860 5257 16869 5277
rect 16681 5246 16717 5247
rect 15953 5241 15989 5243
rect 15953 5212 15990 5241
rect 15395 5203 15430 5204
rect 15372 5198 15430 5203
rect 15372 5178 15375 5198
rect 15395 5184 15430 5198
rect 15450 5184 15459 5204
rect 15395 5176 15459 5184
rect 15421 5175 15459 5176
rect 15422 5174 15459 5175
rect 15525 5208 15561 5209
rect 15633 5208 15669 5209
rect 15525 5203 15669 5208
rect 15525 5200 15587 5203
rect 15525 5180 15533 5200
rect 15553 5180 15587 5200
rect 15525 5177 15587 5180
rect 15613 5200 15669 5203
rect 15613 5180 15641 5200
rect 15661 5180 15669 5200
rect 15613 5177 15669 5180
rect 15525 5174 15669 5177
rect 15735 5204 15773 5212
rect 15851 5208 15887 5209
rect 15735 5184 15744 5204
rect 15764 5184 15773 5204
rect 15735 5175 15773 5184
rect 15802 5200 15887 5208
rect 15802 5180 15859 5200
rect 15879 5180 15887 5200
rect 15735 5174 15772 5175
rect 15802 5174 15887 5180
rect 15953 5204 15991 5212
rect 15953 5184 15962 5204
rect 15982 5184 15991 5204
rect 16832 5190 16869 5257
rect 16904 5286 16935 5337
rect 17217 5325 17235 5343
rect 17253 5325 17269 5343
rect 17735 5350 17773 5359
rect 16954 5286 16991 5287
rect 16904 5277 16991 5286
rect 16904 5257 16962 5277
rect 16982 5257 16991 5277
rect 16904 5247 16991 5257
rect 17050 5277 17087 5287
rect 17050 5257 17058 5277
rect 17078 5257 17087 5277
rect 16904 5246 16935 5247
rect 16529 5187 16566 5188
rect 16832 5187 16871 5190
rect 16528 5186 16871 5187
rect 17050 5186 17087 5257
rect 15953 5175 15991 5184
rect 16453 5181 16871 5186
rect 15953 5174 15990 5175
rect 15414 5146 15504 5152
rect 15414 5126 15430 5146
rect 15450 5144 15504 5146
rect 15450 5126 15475 5144
rect 15414 5124 15475 5126
rect 15495 5124 15504 5144
rect 15414 5118 15504 5124
rect 15427 5064 15464 5065
rect 15523 5064 15560 5065
rect 15579 5064 15615 5174
rect 15802 5153 15833 5174
rect 16453 5161 16456 5181
rect 16476 5161 16871 5181
rect 16900 5162 17087 5186
rect 15798 5152 15833 5153
rect 15676 5142 15833 5152
rect 15676 5122 15693 5142
rect 15713 5122 15833 5142
rect 15676 5115 15833 5122
rect 15900 5145 16049 5153
rect 15900 5125 15911 5145
rect 15931 5125 15970 5145
rect 15990 5125 16049 5145
rect 15900 5118 16049 5125
rect 16832 5136 16871 5161
rect 17217 5136 17269 5325
rect 17563 5332 17603 5342
rect 17563 5314 17573 5332
rect 17591 5314 17603 5332
rect 17735 5330 17744 5350
rect 17764 5330 17773 5350
rect 17735 5322 17773 5330
rect 17839 5354 17924 5360
rect 17954 5359 17991 5360
rect 17839 5334 17847 5354
rect 17867 5334 17924 5354
rect 17839 5326 17924 5334
rect 17953 5350 17991 5359
rect 17953 5330 17962 5350
rect 17982 5330 17991 5350
rect 17839 5325 17875 5326
rect 17953 5322 17991 5330
rect 18057 5354 18201 5360
rect 18057 5334 18065 5354
rect 18085 5334 18118 5354
rect 18138 5334 18173 5354
rect 18193 5334 18201 5354
rect 18057 5326 18201 5334
rect 18057 5325 18093 5326
rect 18165 5325 18201 5326
rect 18267 5359 18304 5360
rect 18267 5358 18305 5359
rect 18267 5350 18331 5358
rect 18267 5330 18276 5350
rect 18296 5336 18331 5350
rect 18351 5336 18354 5356
rect 18296 5331 18354 5336
rect 18296 5330 18331 5331
rect 17563 5258 17603 5314
rect 17736 5293 17773 5322
rect 17737 5291 17773 5293
rect 17737 5269 17928 5291
rect 17954 5290 17991 5322
rect 18267 5318 18331 5330
rect 18371 5292 18398 5470
rect 19256 5445 19298 5490
rect 19319 5491 19330 5509
rect 19352 5491 19364 5509
rect 19319 5485 19364 5491
rect 19320 5484 19364 5485
rect 18230 5290 18398 5292
rect 17954 5280 18398 5290
rect 18539 5386 18726 5410
rect 18757 5391 19150 5411
rect 19170 5391 19173 5411
rect 18757 5386 19173 5391
rect 18539 5315 18576 5386
rect 18757 5385 19098 5386
rect 18691 5325 18722 5326
rect 18539 5295 18548 5315
rect 18568 5295 18576 5315
rect 18539 5285 18576 5295
rect 18635 5315 18722 5325
rect 18635 5295 18644 5315
rect 18664 5295 18722 5315
rect 18635 5286 18722 5295
rect 18635 5285 18672 5286
rect 17560 5253 17603 5258
rect 17951 5264 18398 5280
rect 17951 5258 17979 5264
rect 18230 5263 18398 5264
rect 17560 5250 17710 5253
rect 17951 5250 17978 5258
rect 17560 5248 17978 5250
rect 17560 5230 17569 5248
rect 17587 5230 17978 5248
rect 18691 5235 18722 5286
rect 18757 5315 18794 5385
rect 19060 5384 19097 5385
rect 18909 5325 18945 5326
rect 18757 5295 18766 5315
rect 18786 5295 18794 5315
rect 18757 5285 18794 5295
rect 18853 5315 19001 5325
rect 19101 5322 19197 5324
rect 18853 5295 18862 5315
rect 18882 5295 18972 5315
rect 18992 5295 19001 5315
rect 18853 5286 19001 5295
rect 19059 5315 19197 5322
rect 19059 5295 19068 5315
rect 19088 5295 19197 5315
rect 19059 5286 19197 5295
rect 18853 5285 18890 5286
rect 18583 5232 18624 5233
rect 17560 5227 17978 5230
rect 17560 5221 17603 5227
rect 17563 5218 17603 5221
rect 18478 5225 18624 5232
rect 17960 5209 18000 5210
rect 17671 5192 18000 5209
rect 18478 5205 18534 5225
rect 18554 5205 18593 5225
rect 18613 5205 18624 5225
rect 18478 5197 18624 5205
rect 18691 5228 18848 5235
rect 18691 5208 18811 5228
rect 18831 5208 18848 5228
rect 18691 5198 18848 5208
rect 18691 5197 18726 5198
rect 17555 5149 17598 5160
rect 16832 5118 17271 5136
rect 15900 5117 15941 5118
rect 15634 5064 15671 5065
rect 15330 5055 15465 5064
rect 15330 5035 15436 5055
rect 15456 5035 15465 5055
rect 15330 5028 15465 5035
rect 15523 5055 15671 5064
rect 15523 5035 15532 5055
rect 15552 5035 15642 5055
rect 15662 5035 15671 5055
rect 15330 5026 15423 5028
rect 15523 5025 15671 5035
rect 15730 5055 15767 5065
rect 15730 5035 15738 5055
rect 15758 5035 15767 5055
rect 15579 5024 15615 5025
rect 15427 4965 15464 4966
rect 15730 4965 15767 5035
rect 15802 5064 15833 5115
rect 16832 5100 17232 5118
rect 17250 5100 17271 5118
rect 16832 5094 17271 5100
rect 16838 5090 17271 5094
rect 17555 5131 17567 5149
rect 17585 5131 17598 5149
rect 17555 5105 17598 5131
rect 17671 5105 17698 5192
rect 17960 5183 18000 5192
rect 17217 5088 17269 5090
rect 17555 5084 17698 5105
rect 17742 5157 17776 5173
rect 17960 5163 18353 5183
rect 18373 5163 18376 5183
rect 18691 5176 18722 5197
rect 18909 5176 18945 5286
rect 18964 5285 19001 5286
rect 19060 5285 19097 5286
rect 19020 5226 19110 5232
rect 19020 5206 19029 5226
rect 19049 5224 19110 5226
rect 19049 5206 19074 5224
rect 19020 5204 19074 5206
rect 19094 5204 19110 5224
rect 19020 5198 19110 5204
rect 18534 5175 18571 5176
rect 17960 5158 18376 5163
rect 18533 5166 18571 5175
rect 17960 5157 18301 5158
rect 17742 5087 17779 5157
rect 17894 5097 17925 5098
rect 17555 5082 17692 5084
rect 15852 5064 15889 5065
rect 15802 5055 15889 5064
rect 15802 5035 15860 5055
rect 15880 5035 15889 5055
rect 15802 5025 15889 5035
rect 15948 5055 15985 5065
rect 15948 5035 15956 5055
rect 15976 5035 15985 5055
rect 17555 5040 17598 5082
rect 17742 5067 17751 5087
rect 17771 5067 17779 5087
rect 17742 5057 17779 5067
rect 17838 5087 17925 5097
rect 17838 5067 17847 5087
rect 17867 5067 17925 5087
rect 17838 5058 17925 5067
rect 17838 5057 17875 5058
rect 15802 5024 15833 5025
rect 15426 4964 15767 4965
rect 15948 4964 15985 5035
rect 17553 5030 17598 5040
rect 17220 5023 17257 5028
rect 15351 4959 15767 4964
rect 15351 4939 15354 4959
rect 15374 4939 15767 4959
rect 15798 4940 15985 4964
rect 17211 5019 17258 5023
rect 17211 5001 17230 5019
rect 17248 5001 17258 5019
rect 17553 5012 17562 5030
rect 17580 5012 17598 5030
rect 17553 5006 17598 5012
rect 17894 5007 17925 5058
rect 17960 5087 17997 5157
rect 18263 5156 18300 5157
rect 18533 5146 18542 5166
rect 18562 5146 18571 5166
rect 18533 5138 18571 5146
rect 18637 5170 18722 5176
rect 18752 5175 18789 5176
rect 18637 5150 18645 5170
rect 18665 5150 18722 5170
rect 18637 5142 18722 5150
rect 18751 5166 18789 5175
rect 18751 5146 18760 5166
rect 18780 5146 18789 5166
rect 18637 5141 18673 5142
rect 18751 5138 18789 5146
rect 18855 5170 18999 5176
rect 18855 5150 18863 5170
rect 18883 5167 18971 5170
rect 18883 5150 18918 5167
rect 18855 5149 18918 5150
rect 18937 5150 18971 5167
rect 18991 5150 18999 5170
rect 18937 5149 18999 5150
rect 18855 5142 18999 5149
rect 18855 5141 18891 5142
rect 18963 5141 18999 5142
rect 19065 5175 19102 5176
rect 19065 5174 19103 5175
rect 19125 5174 19152 5178
rect 19065 5172 19152 5174
rect 19065 5166 19129 5172
rect 19065 5146 19074 5166
rect 19094 5152 19129 5166
rect 19149 5152 19152 5172
rect 19094 5147 19152 5152
rect 19094 5146 19129 5147
rect 18534 5109 18571 5138
rect 18535 5107 18571 5109
rect 18112 5097 18148 5098
rect 17960 5067 17969 5087
rect 17989 5067 17997 5087
rect 17960 5057 17997 5067
rect 18056 5087 18204 5097
rect 18304 5094 18400 5096
rect 18056 5067 18065 5087
rect 18085 5067 18175 5087
rect 18195 5067 18204 5087
rect 18056 5058 18204 5067
rect 18262 5087 18400 5094
rect 18262 5067 18271 5087
rect 18291 5067 18400 5087
rect 18535 5085 18726 5107
rect 18752 5106 18789 5138
rect 19065 5134 19129 5146
rect 19169 5108 19196 5286
rect 19028 5106 19196 5108
rect 18752 5080 19196 5106
rect 18262 5058 18400 5067
rect 18056 5057 18093 5058
rect 17553 5003 17590 5006
rect 17786 5004 17827 5005
rect 16819 4942 16857 4943
rect 17211 4942 17258 5001
rect 17678 4997 17827 5004
rect 17678 4977 17737 4997
rect 17757 4977 17796 4997
rect 17816 4977 17827 4997
rect 17678 4969 17827 4977
rect 17894 5000 18051 5007
rect 17894 4980 18014 5000
rect 18034 4980 18051 5000
rect 17894 4970 18051 4980
rect 17894 4969 17929 4970
rect 17894 4948 17925 4969
rect 18112 4948 18148 5058
rect 18167 5057 18204 5058
rect 18263 5057 18300 5058
rect 18223 4998 18313 5004
rect 18223 4978 18232 4998
rect 18252 4996 18313 4998
rect 18252 4978 18277 4996
rect 18223 4976 18277 4978
rect 18297 4976 18313 4996
rect 18223 4970 18313 4976
rect 17737 4947 17774 4948
rect 15571 4938 15636 4939
rect 13686 4860 13724 4861
rect 13285 4822 13724 4860
rect 14596 4860 14604 4882
rect 14628 4860 14636 4882
rect 14596 4852 14636 4860
rect 15907 4904 15947 4912
rect 15907 4882 15915 4904
rect 15939 4882 15947 4904
rect 16819 4904 17258 4942
rect 17550 4939 17587 4941
rect 17550 4931 17592 4939
rect 17550 4913 17560 4931
rect 17578 4913 17592 4931
rect 17550 4904 17592 4913
rect 17736 4938 17774 4947
rect 17736 4918 17745 4938
rect 17765 4918 17774 4938
rect 17736 4910 17774 4918
rect 17840 4942 17925 4948
rect 17955 4947 17992 4948
rect 17840 4922 17848 4942
rect 17868 4922 17925 4942
rect 17840 4914 17925 4922
rect 17954 4938 17992 4947
rect 17954 4918 17963 4938
rect 17983 4918 17992 4938
rect 17840 4913 17876 4914
rect 17954 4910 17992 4918
rect 18058 4946 18202 4948
rect 18058 4942 18110 4946
rect 18058 4922 18066 4942
rect 18086 4926 18110 4942
rect 18130 4942 18202 4946
rect 18130 4926 18174 4942
rect 18086 4922 18174 4926
rect 18194 4922 18202 4942
rect 18058 4914 18202 4922
rect 18058 4913 18094 4914
rect 18166 4913 18202 4914
rect 18268 4947 18305 4948
rect 18268 4946 18306 4947
rect 18268 4938 18332 4946
rect 18268 4918 18277 4938
rect 18297 4924 18332 4938
rect 18352 4924 18355 4944
rect 18297 4919 18355 4924
rect 18297 4918 18332 4919
rect 16819 4903 16857 4904
rect 14907 4825 14972 4826
rect 12113 4806 12148 4807
rect 12090 4801 12148 4806
rect 12090 4781 12093 4801
rect 12113 4787 12148 4801
rect 12168 4787 12177 4807
rect 12113 4779 12177 4787
rect 12139 4778 12177 4779
rect 12140 4777 12177 4778
rect 12243 4811 12279 4812
rect 12351 4811 12387 4812
rect 12243 4803 12387 4811
rect 12243 4783 12251 4803
rect 12271 4799 12359 4803
rect 12271 4783 12315 4799
rect 12243 4779 12315 4783
rect 12335 4783 12359 4799
rect 12379 4783 12387 4803
rect 12335 4779 12387 4783
rect 12243 4777 12387 4779
rect 12453 4807 12491 4815
rect 12569 4811 12605 4812
rect 12453 4787 12462 4807
rect 12482 4787 12491 4807
rect 12453 4778 12491 4787
rect 12520 4803 12605 4811
rect 12520 4783 12577 4803
rect 12597 4783 12605 4803
rect 12453 4777 12490 4778
rect 12520 4777 12605 4783
rect 12671 4807 12709 4815
rect 12671 4787 12680 4807
rect 12700 4787 12709 4807
rect 12671 4778 12709 4787
rect 12853 4812 12895 4821
rect 12853 4794 12867 4812
rect 12885 4794 12895 4812
rect 12853 4786 12895 4794
rect 12858 4784 12895 4786
rect 12671 4777 12708 4778
rect 12132 4749 12222 4755
rect 12132 4729 12148 4749
rect 12168 4747 12222 4749
rect 12168 4729 12193 4747
rect 12132 4727 12193 4729
rect 12213 4727 12222 4747
rect 12132 4721 12222 4727
rect 12145 4667 12182 4668
rect 12241 4667 12278 4668
rect 12297 4667 12333 4777
rect 12520 4756 12551 4777
rect 13285 4763 13332 4822
rect 13686 4821 13724 4822
rect 12516 4755 12551 4756
rect 12394 4745 12551 4755
rect 12394 4725 12411 4745
rect 12431 4725 12551 4745
rect 12394 4718 12551 4725
rect 12618 4748 12767 4756
rect 12618 4728 12629 4748
rect 12649 4728 12688 4748
rect 12708 4728 12767 4748
rect 13285 4745 13295 4763
rect 13313 4745 13332 4763
rect 13285 4741 13332 4745
rect 14558 4800 14745 4824
rect 14776 4805 15169 4825
rect 15189 4805 15192 4825
rect 14776 4800 15192 4805
rect 13286 4736 13323 4741
rect 12618 4721 12767 4728
rect 14558 4729 14595 4800
rect 14776 4799 15117 4800
rect 14710 4739 14741 4740
rect 12618 4720 12659 4721
rect 12855 4719 12892 4722
rect 12352 4667 12389 4668
rect 12045 4658 12183 4667
rect 11249 4619 11693 4645
rect 11249 4617 11417 4619
rect 11249 4439 11276 4617
rect 11316 4579 11380 4591
rect 11656 4587 11693 4619
rect 11719 4618 11910 4640
rect 12045 4638 12154 4658
rect 12174 4638 12183 4658
rect 12045 4631 12183 4638
rect 12241 4658 12389 4667
rect 12241 4638 12250 4658
rect 12270 4638 12360 4658
rect 12380 4638 12389 4658
rect 12045 4629 12141 4631
rect 12241 4628 12389 4638
rect 12448 4658 12485 4668
rect 12448 4638 12456 4658
rect 12476 4638 12485 4658
rect 12297 4627 12333 4628
rect 11874 4616 11910 4618
rect 11874 4587 11911 4616
rect 11316 4578 11351 4579
rect 11293 4573 11351 4578
rect 11293 4553 11296 4573
rect 11316 4559 11351 4573
rect 11371 4559 11380 4579
rect 11316 4553 11380 4559
rect 11293 4551 11380 4553
rect 11293 4547 11320 4551
rect 11342 4550 11380 4551
rect 11343 4549 11380 4550
rect 11446 4583 11482 4584
rect 11554 4583 11590 4584
rect 11446 4576 11590 4583
rect 11446 4575 11508 4576
rect 11446 4555 11454 4575
rect 11474 4558 11508 4575
rect 11527 4575 11590 4576
rect 11527 4558 11562 4575
rect 11474 4555 11562 4558
rect 11582 4555 11590 4575
rect 11446 4549 11590 4555
rect 11656 4579 11694 4587
rect 11772 4583 11808 4584
rect 11656 4559 11665 4579
rect 11685 4559 11694 4579
rect 11656 4550 11694 4559
rect 11723 4575 11808 4583
rect 11723 4555 11780 4575
rect 11800 4555 11808 4575
rect 11656 4549 11693 4550
rect 11723 4549 11808 4555
rect 11874 4579 11912 4587
rect 11874 4559 11883 4579
rect 11903 4559 11912 4579
rect 12145 4568 12182 4569
rect 12448 4568 12485 4638
rect 12520 4667 12551 4718
rect 12847 4713 12892 4719
rect 12847 4695 12865 4713
rect 12883 4695 12892 4713
rect 14558 4709 14567 4729
rect 14587 4709 14595 4729
rect 14558 4699 14595 4709
rect 14654 4729 14741 4739
rect 14654 4709 14663 4729
rect 14683 4709 14741 4729
rect 14654 4700 14741 4709
rect 14654 4699 14691 4700
rect 12847 4685 12892 4695
rect 12570 4667 12607 4668
rect 12520 4658 12607 4667
rect 12520 4638 12578 4658
rect 12598 4638 12607 4658
rect 12520 4628 12607 4638
rect 12666 4658 12703 4668
rect 12666 4638 12674 4658
rect 12694 4638 12703 4658
rect 12847 4643 12890 4685
rect 13274 4674 13326 4676
rect 12753 4641 12890 4643
rect 12520 4627 12551 4628
rect 12666 4568 12703 4638
rect 12144 4567 12485 4568
rect 11874 4550 11912 4559
rect 12069 4562 12485 4567
rect 11874 4549 11911 4550
rect 11335 4521 11425 4527
rect 11335 4501 11351 4521
rect 11371 4519 11425 4521
rect 11371 4501 11396 4519
rect 11335 4499 11396 4501
rect 11416 4499 11425 4519
rect 11335 4493 11425 4499
rect 11348 4439 11385 4440
rect 11444 4439 11481 4440
rect 11500 4439 11536 4549
rect 11723 4528 11754 4549
rect 12069 4542 12072 4562
rect 12092 4542 12485 4562
rect 12669 4552 12703 4568
rect 12747 4620 12890 4641
rect 13272 4670 13705 4674
rect 13272 4664 13711 4670
rect 13272 4646 13293 4664
rect 13311 4646 13711 4664
rect 14710 4649 14741 4700
rect 14776 4729 14813 4799
rect 15079 4798 15116 4799
rect 14928 4739 14964 4740
rect 14776 4709 14785 4729
rect 14805 4709 14813 4729
rect 14776 4699 14813 4709
rect 14872 4729 15020 4739
rect 15120 4736 15216 4738
rect 14872 4709 14881 4729
rect 14901 4709 14991 4729
rect 15011 4709 15020 4729
rect 14872 4700 15020 4709
rect 15078 4729 15216 4736
rect 15078 4709 15087 4729
rect 15107 4709 15216 4729
rect 15078 4700 15216 4709
rect 14872 4699 14909 4700
rect 14602 4646 14643 4647
rect 13272 4628 13711 4646
rect 12445 4533 12485 4542
rect 12747 4533 12774 4620
rect 12847 4594 12890 4620
rect 12847 4576 12860 4594
rect 12878 4576 12890 4594
rect 12847 4565 12890 4576
rect 11719 4527 11754 4528
rect 11597 4517 11754 4527
rect 11597 4497 11614 4517
rect 11634 4497 11754 4517
rect 11597 4490 11754 4497
rect 11821 4520 11967 4528
rect 11821 4500 11832 4520
rect 11852 4500 11891 4520
rect 11911 4500 11967 4520
rect 12445 4516 12774 4533
rect 12445 4515 12485 4516
rect 11821 4493 11967 4500
rect 12842 4504 12882 4507
rect 12842 4498 12885 4504
rect 12467 4495 12885 4498
rect 11821 4492 11862 4493
rect 11555 4439 11592 4440
rect 11248 4430 11386 4439
rect 11248 4410 11357 4430
rect 11377 4410 11386 4430
rect 11248 4403 11386 4410
rect 11444 4430 11592 4439
rect 11444 4410 11453 4430
rect 11473 4410 11563 4430
rect 11583 4410 11592 4430
rect 11248 4401 11344 4403
rect 11444 4400 11592 4410
rect 11651 4430 11688 4440
rect 11651 4410 11659 4430
rect 11679 4410 11688 4430
rect 11500 4399 11536 4400
rect 11348 4340 11385 4341
rect 11651 4340 11688 4410
rect 11723 4439 11754 4490
rect 12467 4477 12858 4495
rect 12876 4477 12885 4495
rect 12467 4475 12885 4477
rect 12467 4467 12494 4475
rect 12735 4472 12885 4475
rect 12047 4461 12215 4462
rect 12466 4461 12494 4467
rect 12047 4445 12494 4461
rect 12842 4467 12885 4472
rect 11773 4439 11810 4440
rect 11723 4430 11810 4439
rect 11723 4410 11781 4430
rect 11801 4410 11810 4430
rect 11723 4400 11810 4410
rect 11869 4430 11906 4440
rect 11869 4410 11877 4430
rect 11897 4410 11906 4430
rect 11723 4399 11754 4400
rect 11347 4339 11688 4340
rect 11869 4339 11906 4410
rect 11272 4334 11688 4339
rect 11272 4314 11275 4334
rect 11295 4314 11688 4334
rect 11719 4315 11906 4339
rect 12047 4435 12491 4445
rect 12047 4433 12215 4435
rect 11081 4240 11125 4241
rect 11081 4234 11126 4240
rect 11081 4216 11093 4234
rect 11115 4216 11126 4234
rect 11147 4235 11189 4280
rect 12047 4255 12074 4433
rect 12114 4395 12178 4407
rect 12454 4403 12491 4435
rect 12517 4434 12708 4456
rect 12672 4432 12708 4434
rect 12672 4403 12709 4432
rect 12842 4411 12882 4467
rect 12114 4394 12149 4395
rect 12091 4389 12149 4394
rect 12091 4369 12094 4389
rect 12114 4375 12149 4389
rect 12169 4375 12178 4395
rect 12114 4367 12178 4375
rect 12140 4366 12178 4367
rect 12141 4365 12178 4366
rect 12244 4399 12280 4400
rect 12352 4399 12388 4400
rect 12244 4391 12388 4399
rect 12244 4371 12252 4391
rect 12272 4371 12307 4391
rect 12327 4371 12360 4391
rect 12380 4371 12388 4391
rect 12244 4365 12388 4371
rect 12454 4395 12492 4403
rect 12570 4399 12606 4400
rect 12454 4375 12463 4395
rect 12483 4375 12492 4395
rect 12454 4366 12492 4375
rect 12521 4391 12606 4399
rect 12521 4371 12578 4391
rect 12598 4371 12606 4391
rect 12454 4365 12491 4366
rect 12521 4365 12606 4371
rect 12672 4395 12710 4403
rect 12672 4375 12681 4395
rect 12701 4375 12710 4395
rect 12842 4393 12854 4411
rect 12872 4393 12882 4411
rect 13274 4439 13326 4628
rect 13672 4603 13711 4628
rect 14494 4639 14643 4646
rect 14494 4619 14553 4639
rect 14573 4619 14612 4639
rect 14632 4619 14643 4639
rect 14494 4611 14643 4619
rect 14710 4642 14867 4649
rect 14710 4622 14830 4642
rect 14850 4622 14867 4642
rect 14710 4612 14867 4622
rect 14710 4611 14745 4612
rect 13456 4578 13643 4602
rect 13672 4583 14067 4603
rect 14087 4583 14090 4603
rect 14710 4590 14741 4611
rect 14928 4590 14964 4700
rect 14983 4699 15020 4700
rect 15079 4699 15116 4700
rect 15039 4640 15129 4646
rect 15039 4620 15048 4640
rect 15068 4638 15129 4640
rect 15068 4620 15093 4638
rect 15039 4618 15093 4620
rect 15113 4618 15129 4638
rect 15039 4612 15129 4618
rect 14553 4589 14590 4590
rect 13672 4578 14090 4583
rect 14552 4580 14590 4589
rect 13456 4507 13493 4578
rect 13672 4577 14015 4578
rect 13672 4574 13711 4577
rect 13977 4576 14014 4577
rect 13608 4517 13639 4518
rect 13456 4487 13465 4507
rect 13485 4487 13493 4507
rect 13456 4477 13493 4487
rect 13552 4507 13639 4517
rect 13552 4487 13561 4507
rect 13581 4487 13639 4507
rect 13552 4478 13639 4487
rect 13552 4477 13589 4478
rect 13274 4421 13290 4439
rect 13308 4421 13326 4439
rect 13608 4427 13639 4478
rect 13674 4507 13711 4574
rect 14552 4560 14561 4580
rect 14581 4560 14590 4580
rect 14552 4552 14590 4560
rect 14656 4584 14741 4590
rect 14771 4589 14808 4590
rect 14656 4564 14664 4584
rect 14684 4564 14741 4584
rect 14656 4556 14741 4564
rect 14770 4580 14808 4589
rect 14770 4560 14779 4580
rect 14799 4560 14808 4580
rect 14656 4555 14692 4556
rect 14770 4552 14808 4560
rect 14874 4584 15018 4590
rect 14874 4564 14882 4584
rect 14902 4578 14990 4584
rect 14902 4564 14931 4578
rect 14874 4556 14931 4564
rect 14874 4555 14910 4556
rect 14954 4564 14990 4578
rect 15010 4564 15018 4584
rect 14954 4556 15018 4564
rect 14982 4555 15018 4556
rect 15084 4589 15121 4590
rect 15084 4588 15122 4589
rect 15084 4580 15148 4588
rect 15084 4560 15093 4580
rect 15113 4566 15148 4580
rect 15168 4566 15171 4586
rect 15113 4561 15171 4566
rect 15113 4560 15148 4561
rect 14553 4523 14590 4552
rect 14554 4521 14590 4523
rect 13826 4517 13862 4518
rect 13674 4487 13683 4507
rect 13703 4487 13711 4507
rect 13674 4477 13711 4487
rect 13770 4507 13918 4517
rect 14018 4514 14114 4516
rect 13770 4487 13779 4507
rect 13799 4487 13889 4507
rect 13909 4487 13918 4507
rect 13770 4478 13918 4487
rect 13976 4507 14114 4514
rect 13976 4487 13985 4507
rect 14005 4487 14114 4507
rect 14554 4499 14745 4521
rect 14771 4520 14808 4552
rect 15084 4548 15148 4560
rect 15188 4522 15215 4700
rect 15512 4653 15549 4659
rect 15512 4634 15520 4653
rect 15541 4634 15549 4653
rect 15512 4626 15549 4634
rect 15047 4520 15215 4522
rect 14771 4494 15215 4520
rect 14881 4492 14921 4494
rect 15047 4493 15215 4494
rect 13976 4478 14114 4487
rect 15174 4488 15215 4493
rect 13770 4477 13807 4478
rect 13500 4424 13541 4425
rect 13274 4403 13326 4421
rect 13392 4417 13541 4424
rect 12842 4383 12882 4393
rect 13392 4397 13451 4417
rect 13471 4397 13510 4417
rect 13530 4397 13541 4417
rect 13392 4389 13541 4397
rect 13608 4420 13765 4427
rect 13608 4400 13728 4420
rect 13748 4400 13765 4420
rect 13608 4390 13765 4400
rect 13608 4389 13643 4390
rect 12672 4366 12710 4375
rect 13608 4368 13639 4389
rect 13826 4368 13862 4478
rect 13881 4477 13918 4478
rect 13977 4477 14014 4478
rect 13937 4418 14027 4424
rect 13937 4398 13946 4418
rect 13966 4416 14027 4418
rect 13966 4398 13991 4416
rect 13937 4396 13991 4398
rect 14011 4396 14027 4416
rect 13937 4390 14027 4396
rect 13451 4367 13488 4368
rect 12672 4365 12709 4366
rect 12133 4337 12223 4343
rect 12133 4317 12149 4337
rect 12169 4335 12223 4337
rect 12169 4317 12194 4335
rect 12133 4315 12194 4317
rect 12214 4315 12223 4335
rect 12133 4309 12223 4315
rect 12146 4255 12183 4256
rect 12242 4255 12279 4256
rect 12298 4255 12334 4365
rect 12521 4344 12552 4365
rect 13450 4358 13488 4367
rect 12517 4343 12552 4344
rect 12395 4333 12552 4343
rect 12395 4313 12412 4333
rect 12432 4313 12552 4333
rect 12395 4306 12552 4313
rect 12619 4336 12768 4344
rect 12619 4316 12630 4336
rect 12650 4316 12689 4336
rect 12709 4316 12768 4336
rect 13278 4340 13318 4350
rect 12619 4309 12768 4316
rect 12834 4312 12886 4330
rect 12619 4308 12660 4309
rect 12353 4255 12390 4256
rect 12046 4246 12184 4255
rect 11518 4235 11551 4237
rect 11147 4223 11594 4235
rect 11081 4186 11126 4216
rect 11098 3240 11126 4186
rect 11150 4209 11594 4223
rect 11150 4207 11318 4209
rect 11150 4029 11177 4207
rect 11217 4169 11281 4181
rect 11557 4177 11594 4209
rect 11620 4208 11811 4230
rect 12046 4226 12155 4246
rect 12175 4226 12184 4246
rect 12046 4219 12184 4226
rect 12242 4246 12390 4255
rect 12242 4226 12251 4246
rect 12271 4226 12361 4246
rect 12381 4226 12390 4246
rect 12046 4217 12142 4219
rect 12242 4216 12390 4226
rect 12449 4246 12486 4256
rect 12449 4226 12457 4246
rect 12477 4226 12486 4246
rect 12298 4215 12334 4216
rect 11775 4206 11811 4208
rect 11775 4177 11812 4206
rect 11217 4168 11252 4169
rect 11194 4163 11252 4168
rect 11194 4143 11197 4163
rect 11217 4149 11252 4163
rect 11272 4149 11281 4169
rect 11217 4141 11281 4149
rect 11243 4140 11281 4141
rect 11244 4139 11281 4140
rect 11347 4173 11383 4174
rect 11455 4173 11491 4174
rect 11347 4167 11491 4173
rect 11347 4165 11408 4167
rect 11347 4145 11355 4165
rect 11375 4150 11408 4165
rect 11427 4165 11491 4167
rect 11427 4150 11463 4165
rect 11375 4145 11463 4150
rect 11483 4145 11491 4165
rect 11347 4139 11491 4145
rect 11557 4169 11595 4177
rect 11673 4173 11709 4174
rect 11557 4149 11566 4169
rect 11586 4149 11595 4169
rect 11557 4140 11595 4149
rect 11624 4165 11709 4173
rect 11624 4145 11681 4165
rect 11701 4145 11709 4165
rect 11557 4139 11594 4140
rect 11624 4139 11709 4145
rect 11775 4169 11813 4177
rect 11775 4149 11784 4169
rect 11804 4149 11813 4169
rect 12449 4159 12486 4226
rect 12521 4255 12552 4306
rect 12834 4294 12852 4312
rect 12870 4294 12886 4312
rect 12571 4255 12608 4256
rect 12521 4246 12608 4255
rect 12521 4226 12579 4246
rect 12599 4226 12608 4246
rect 12521 4216 12608 4226
rect 12667 4246 12704 4256
rect 12667 4226 12675 4246
rect 12695 4226 12704 4246
rect 12521 4215 12552 4216
rect 12146 4156 12183 4157
rect 12449 4156 12488 4159
rect 12145 4155 12488 4156
rect 12667 4155 12704 4226
rect 11775 4140 11813 4149
rect 12070 4150 12488 4155
rect 11775 4139 11812 4140
rect 11236 4111 11326 4117
rect 11236 4091 11252 4111
rect 11272 4109 11326 4111
rect 11272 4091 11297 4109
rect 11236 4089 11297 4091
rect 11317 4089 11326 4109
rect 11236 4083 11326 4089
rect 11249 4029 11286 4030
rect 11345 4029 11382 4030
rect 11401 4029 11437 4139
rect 11624 4118 11655 4139
rect 12070 4130 12073 4150
rect 12093 4130 12488 4150
rect 12517 4131 12704 4155
rect 11620 4117 11655 4118
rect 11498 4107 11655 4117
rect 11498 4087 11515 4107
rect 11535 4087 11655 4107
rect 11498 4080 11655 4087
rect 11722 4110 11871 4118
rect 11722 4090 11733 4110
rect 11753 4090 11792 4110
rect 11812 4090 11871 4110
rect 11722 4083 11871 4090
rect 12449 4105 12488 4130
rect 12834 4105 12886 4294
rect 13278 4322 13288 4340
rect 13306 4322 13318 4340
rect 13450 4338 13459 4358
rect 13479 4338 13488 4358
rect 13450 4330 13488 4338
rect 13554 4362 13639 4368
rect 13669 4367 13706 4368
rect 13554 4342 13562 4362
rect 13582 4342 13639 4362
rect 13554 4334 13639 4342
rect 13668 4358 13706 4367
rect 13668 4338 13677 4358
rect 13697 4338 13706 4358
rect 13554 4333 13590 4334
rect 13668 4330 13706 4338
rect 13772 4362 13916 4368
rect 13772 4342 13780 4362
rect 13800 4342 13833 4362
rect 13853 4342 13888 4362
rect 13908 4342 13916 4362
rect 13772 4334 13916 4342
rect 13772 4333 13808 4334
rect 13880 4333 13916 4334
rect 13982 4367 14019 4368
rect 13982 4366 14020 4367
rect 13982 4358 14046 4366
rect 13982 4338 13991 4358
rect 14011 4344 14046 4358
rect 14066 4344 14069 4364
rect 14011 4339 14069 4344
rect 14011 4338 14046 4339
rect 13278 4266 13318 4322
rect 13451 4301 13488 4330
rect 13452 4299 13488 4301
rect 13452 4277 13643 4299
rect 13669 4298 13706 4330
rect 13982 4326 14046 4338
rect 14086 4300 14113 4478
rect 13945 4298 14113 4300
rect 13669 4288 14113 4298
rect 14254 4394 14441 4418
rect 14472 4399 14865 4419
rect 14885 4399 14888 4419
rect 14472 4394 14888 4399
rect 14254 4323 14291 4394
rect 14472 4393 14813 4394
rect 14406 4333 14437 4334
rect 14254 4303 14263 4323
rect 14283 4303 14291 4323
rect 14254 4293 14291 4303
rect 14350 4323 14437 4333
rect 14350 4303 14359 4323
rect 14379 4303 14437 4323
rect 14350 4294 14437 4303
rect 14350 4293 14387 4294
rect 13275 4261 13318 4266
rect 13666 4272 14113 4288
rect 13666 4266 13694 4272
rect 13945 4271 14113 4272
rect 13275 4258 13425 4261
rect 13666 4258 13693 4266
rect 13275 4256 13693 4258
rect 13275 4238 13284 4256
rect 13302 4238 13693 4256
rect 14406 4243 14437 4294
rect 14472 4323 14509 4393
rect 14775 4392 14812 4393
rect 14624 4333 14660 4334
rect 14472 4303 14481 4323
rect 14501 4303 14509 4323
rect 14472 4293 14509 4303
rect 14568 4323 14716 4333
rect 14816 4330 14912 4332
rect 14568 4303 14577 4323
rect 14597 4303 14687 4323
rect 14707 4303 14716 4323
rect 14568 4294 14716 4303
rect 14774 4323 14912 4330
rect 14774 4303 14783 4323
rect 14803 4303 14912 4323
rect 15174 4306 15214 4488
rect 14774 4294 14912 4303
rect 14568 4293 14605 4294
rect 14298 4240 14339 4241
rect 13275 4235 13693 4238
rect 13275 4229 13318 4235
rect 13278 4226 13318 4229
rect 14190 4233 14339 4240
rect 13675 4217 13715 4218
rect 13386 4200 13715 4217
rect 14190 4213 14249 4233
rect 14269 4213 14308 4233
rect 14328 4213 14339 4233
rect 14190 4205 14339 4213
rect 14406 4236 14563 4243
rect 14406 4216 14526 4236
rect 14546 4216 14563 4236
rect 14406 4206 14563 4216
rect 14406 4205 14441 4206
rect 13270 4157 13313 4168
rect 13270 4139 13282 4157
rect 13300 4139 13313 4157
rect 13270 4113 13313 4139
rect 13386 4113 13413 4200
rect 13675 4191 13715 4200
rect 12449 4087 12888 4105
rect 11722 4082 11763 4083
rect 11456 4029 11493 4030
rect 11149 4020 11287 4029
rect 11149 4000 11258 4020
rect 11278 4000 11287 4020
rect 11149 3993 11287 4000
rect 11345 4020 11493 4029
rect 11345 4000 11354 4020
rect 11374 4000 11464 4020
rect 11484 4000 11493 4020
rect 11149 3991 11245 3993
rect 11345 3990 11493 4000
rect 11552 4020 11589 4030
rect 11552 4000 11560 4020
rect 11580 4000 11589 4020
rect 11401 3989 11437 3990
rect 11249 3930 11286 3931
rect 11552 3930 11589 4000
rect 11624 4029 11655 4080
rect 12449 4069 12849 4087
rect 12867 4069 12888 4087
rect 12449 4063 12888 4069
rect 12455 4059 12888 4063
rect 13270 4092 13413 4113
rect 13457 4165 13491 4181
rect 13675 4171 14068 4191
rect 14088 4171 14091 4191
rect 14406 4184 14437 4205
rect 14624 4184 14660 4294
rect 14679 4293 14716 4294
rect 14775 4293 14812 4294
rect 14735 4234 14825 4240
rect 14735 4214 14744 4234
rect 14764 4232 14825 4234
rect 14764 4214 14789 4232
rect 14735 4212 14789 4214
rect 14809 4212 14825 4232
rect 14735 4206 14825 4212
rect 14249 4183 14286 4184
rect 13675 4166 14091 4171
rect 14248 4174 14286 4183
rect 13675 4165 14016 4166
rect 13457 4095 13494 4165
rect 13609 4105 13640 4106
rect 13270 4090 13407 4092
rect 12834 4057 12886 4059
rect 13270 4048 13313 4090
rect 13457 4075 13466 4095
rect 13486 4075 13494 4095
rect 13457 4065 13494 4075
rect 13553 4095 13640 4105
rect 13553 4075 13562 4095
rect 13582 4075 13640 4095
rect 13553 4066 13640 4075
rect 13553 4065 13590 4066
rect 13268 4038 13313 4048
rect 11674 4029 11711 4030
rect 11624 4020 11711 4029
rect 11624 4000 11682 4020
rect 11702 4000 11711 4020
rect 11624 3990 11711 4000
rect 11770 4020 11807 4030
rect 11770 4000 11778 4020
rect 11798 4000 11807 4020
rect 13268 4020 13277 4038
rect 13295 4020 13313 4038
rect 13268 4014 13313 4020
rect 13609 4015 13640 4066
rect 13675 4095 13712 4165
rect 13978 4164 14015 4165
rect 14248 4154 14257 4174
rect 14277 4154 14286 4174
rect 14248 4146 14286 4154
rect 14352 4178 14437 4184
rect 14467 4183 14504 4184
rect 14352 4158 14360 4178
rect 14380 4158 14437 4178
rect 14352 4150 14437 4158
rect 14466 4174 14504 4183
rect 14466 4154 14475 4174
rect 14495 4154 14504 4174
rect 14352 4149 14388 4150
rect 14466 4146 14504 4154
rect 14570 4178 14714 4184
rect 14570 4158 14578 4178
rect 14598 4159 14630 4178
rect 14651 4159 14686 4178
rect 14598 4158 14686 4159
rect 14706 4158 14714 4178
rect 14570 4150 14714 4158
rect 14570 4149 14606 4150
rect 14678 4149 14714 4150
rect 14780 4183 14817 4184
rect 14780 4182 14818 4183
rect 14780 4174 14844 4182
rect 14780 4154 14789 4174
rect 14809 4160 14844 4174
rect 14864 4160 14867 4180
rect 14809 4155 14867 4160
rect 14809 4154 14844 4155
rect 14249 4117 14286 4146
rect 14250 4115 14286 4117
rect 13827 4105 13863 4106
rect 13675 4075 13684 4095
rect 13704 4075 13712 4095
rect 13675 4065 13712 4075
rect 13771 4095 13919 4105
rect 14019 4102 14115 4104
rect 13771 4075 13780 4095
rect 13800 4075 13890 4095
rect 13910 4075 13919 4095
rect 13771 4066 13919 4075
rect 13977 4095 14115 4102
rect 13977 4075 13986 4095
rect 14006 4075 14115 4095
rect 14250 4093 14441 4115
rect 14467 4114 14504 4146
rect 14780 4142 14844 4154
rect 14884 4116 14911 4294
rect 14743 4114 14911 4116
rect 14467 4088 14911 4114
rect 13977 4066 14115 4075
rect 13771 4065 13808 4066
rect 13268 4011 13305 4014
rect 13501 4012 13542 4013
rect 11624 3989 11655 3990
rect 11248 3929 11589 3930
rect 11770 3929 11807 4000
rect 13393 4005 13542 4012
rect 12837 3992 12874 3997
rect 12828 3988 12875 3992
rect 12828 3970 12847 3988
rect 12865 3970 12875 3988
rect 13393 3985 13452 4005
rect 13472 3985 13511 4005
rect 13531 3985 13542 4005
rect 13393 3977 13542 3985
rect 13609 4008 13766 4015
rect 13609 3988 13729 4008
rect 13749 3988 13766 4008
rect 13609 3978 13766 3988
rect 13609 3977 13644 3978
rect 11173 3924 11589 3929
rect 11173 3904 11176 3924
rect 11196 3904 11589 3924
rect 11620 3905 11807 3929
rect 12432 3927 12472 3932
rect 12828 3927 12875 3970
rect 13609 3956 13640 3977
rect 13827 3956 13863 4066
rect 13882 4065 13919 4066
rect 13978 4065 14015 4066
rect 13938 4006 14028 4012
rect 13938 3986 13947 4006
rect 13967 4004 14028 4006
rect 13967 3986 13992 4004
rect 13938 3984 13992 3986
rect 14012 3984 14028 4004
rect 13938 3978 14028 3984
rect 13452 3955 13489 3956
rect 12432 3888 12875 3927
rect 13265 3947 13302 3949
rect 13265 3939 13307 3947
rect 13265 3921 13275 3939
rect 13293 3921 13307 3939
rect 13265 3912 13307 3921
rect 13451 3946 13489 3955
rect 13451 3926 13460 3946
rect 13480 3926 13489 3946
rect 13451 3918 13489 3926
rect 13555 3950 13640 3956
rect 13670 3955 13707 3956
rect 13555 3930 13563 3950
rect 13583 3930 13640 3950
rect 13555 3922 13640 3930
rect 13669 3946 13707 3955
rect 13669 3926 13678 3946
rect 13698 3926 13707 3946
rect 13555 3921 13591 3922
rect 13669 3918 13707 3926
rect 13773 3954 13917 3956
rect 13773 3950 13825 3954
rect 13773 3930 13781 3950
rect 13801 3934 13825 3950
rect 13845 3950 13917 3954
rect 13845 3934 13889 3950
rect 13801 3930 13889 3934
rect 13909 3930 13917 3950
rect 13773 3922 13917 3930
rect 13773 3921 13809 3922
rect 13881 3921 13917 3922
rect 13983 3955 14020 3956
rect 13983 3954 14021 3955
rect 13983 3946 14047 3954
rect 13983 3926 13992 3946
rect 14012 3932 14047 3946
rect 14067 3932 14070 3952
rect 14012 3927 14070 3932
rect 14012 3926 14047 3927
rect 11526 3873 11566 3881
rect 11526 3851 11534 3873
rect 11558 3851 11566 3873
rect 11232 3627 11400 3628
rect 11526 3627 11566 3851
rect 12029 3855 12197 3856
rect 12432 3855 12472 3888
rect 12828 3855 12875 3888
rect 13266 3887 13307 3912
rect 13452 3887 13489 3918
rect 13670 3887 13707 3918
rect 13983 3914 14047 3926
rect 14087 3888 14114 4066
rect 13266 3860 13315 3887
rect 13451 3861 13500 3887
rect 13669 3886 13750 3887
rect 13946 3886 14114 3888
rect 13669 3861 14114 3886
rect 13670 3860 14114 3861
rect 12029 3854 12473 3855
rect 12029 3829 12474 3854
rect 12029 3827 12197 3829
rect 12393 3828 12474 3829
rect 12643 3828 12692 3854
rect 12828 3828 12877 3855
rect 12029 3649 12056 3827
rect 12096 3789 12160 3801
rect 12436 3797 12473 3828
rect 12654 3797 12691 3828
rect 12836 3803 12877 3828
rect 13268 3827 13315 3860
rect 13671 3827 13711 3860
rect 13946 3859 14114 3860
rect 14577 3864 14617 4088
rect 14743 4087 14911 4088
rect 14577 3842 14585 3864
rect 14609 3842 14617 3864
rect 14577 3834 14617 3842
rect 12096 3788 12131 3789
rect 12073 3783 12131 3788
rect 12073 3763 12076 3783
rect 12096 3769 12131 3783
rect 12151 3769 12160 3789
rect 12096 3761 12160 3769
rect 12122 3760 12160 3761
rect 12123 3759 12160 3760
rect 12226 3793 12262 3794
rect 12334 3793 12370 3794
rect 12226 3785 12370 3793
rect 12226 3765 12234 3785
rect 12254 3781 12342 3785
rect 12254 3765 12298 3781
rect 12226 3761 12298 3765
rect 12318 3765 12342 3781
rect 12362 3765 12370 3785
rect 12318 3761 12370 3765
rect 12226 3759 12370 3761
rect 12436 3789 12474 3797
rect 12552 3793 12588 3794
rect 12436 3769 12445 3789
rect 12465 3769 12474 3789
rect 12436 3760 12474 3769
rect 12503 3785 12588 3793
rect 12503 3765 12560 3785
rect 12580 3765 12588 3785
rect 12436 3759 12473 3760
rect 12503 3759 12588 3765
rect 12654 3789 12692 3797
rect 12654 3769 12663 3789
rect 12683 3769 12692 3789
rect 12654 3760 12692 3769
rect 12836 3794 12878 3803
rect 12836 3776 12850 3794
rect 12868 3776 12878 3794
rect 12836 3768 12878 3776
rect 12841 3766 12878 3768
rect 13268 3788 13711 3827
rect 12654 3759 12691 3760
rect 12115 3731 12205 3737
rect 12115 3711 12131 3731
rect 12151 3729 12205 3731
rect 12151 3711 12176 3729
rect 12115 3709 12176 3711
rect 12196 3709 12205 3729
rect 12115 3703 12205 3709
rect 12128 3649 12165 3650
rect 12224 3649 12261 3650
rect 12280 3649 12316 3759
rect 12503 3738 12534 3759
rect 13268 3745 13315 3788
rect 13671 3783 13711 3788
rect 14336 3786 14523 3810
rect 14554 3791 14947 3811
rect 14967 3791 14970 3811
rect 14554 3786 14970 3791
rect 12499 3737 12534 3738
rect 12377 3727 12534 3737
rect 12377 3707 12394 3727
rect 12414 3707 12534 3727
rect 12377 3700 12534 3707
rect 12601 3730 12750 3738
rect 12601 3710 12612 3730
rect 12632 3710 12671 3730
rect 12691 3710 12750 3730
rect 13268 3727 13278 3745
rect 13296 3727 13315 3745
rect 13268 3723 13315 3727
rect 13269 3718 13306 3723
rect 12601 3703 12750 3710
rect 14336 3715 14373 3786
rect 14554 3785 14895 3786
rect 14488 3725 14519 3726
rect 12601 3702 12642 3703
rect 12838 3701 12875 3704
rect 12335 3649 12372 3650
rect 12028 3640 12166 3649
rect 11232 3601 11676 3627
rect 11232 3599 11400 3601
rect 11232 3421 11259 3599
rect 11299 3561 11363 3573
rect 11639 3569 11676 3601
rect 11702 3600 11893 3622
rect 12028 3620 12137 3640
rect 12157 3620 12166 3640
rect 12028 3613 12166 3620
rect 12224 3640 12372 3649
rect 12224 3620 12233 3640
rect 12253 3620 12343 3640
rect 12363 3620 12372 3640
rect 12028 3611 12124 3613
rect 12224 3610 12372 3620
rect 12431 3640 12468 3650
rect 12431 3620 12439 3640
rect 12459 3620 12468 3640
rect 12280 3609 12316 3610
rect 11857 3598 11893 3600
rect 11857 3569 11894 3598
rect 11299 3560 11334 3561
rect 11276 3555 11334 3560
rect 11276 3535 11279 3555
rect 11299 3541 11334 3555
rect 11354 3541 11363 3561
rect 11299 3533 11363 3541
rect 11325 3532 11363 3533
rect 11326 3531 11363 3532
rect 11429 3565 11465 3566
rect 11537 3565 11573 3566
rect 11429 3557 11573 3565
rect 11429 3537 11437 3557
rect 11457 3556 11545 3557
rect 11457 3537 11492 3556
rect 11513 3537 11545 3556
rect 11565 3537 11573 3557
rect 11429 3531 11573 3537
rect 11639 3561 11677 3569
rect 11755 3565 11791 3566
rect 11639 3541 11648 3561
rect 11668 3541 11677 3561
rect 11639 3532 11677 3541
rect 11706 3557 11791 3565
rect 11706 3537 11763 3557
rect 11783 3537 11791 3557
rect 11639 3531 11676 3532
rect 11706 3531 11791 3537
rect 11857 3561 11895 3569
rect 11857 3541 11866 3561
rect 11886 3541 11895 3561
rect 12128 3550 12165 3551
rect 12431 3550 12468 3620
rect 12503 3649 12534 3700
rect 12830 3695 12875 3701
rect 12830 3677 12848 3695
rect 12866 3677 12875 3695
rect 14336 3695 14345 3715
rect 14365 3695 14373 3715
rect 14336 3685 14373 3695
rect 14432 3715 14519 3725
rect 14432 3695 14441 3715
rect 14461 3695 14519 3715
rect 14432 3686 14519 3695
rect 14432 3685 14469 3686
rect 12830 3667 12875 3677
rect 12553 3649 12590 3650
rect 12503 3640 12590 3649
rect 12503 3620 12561 3640
rect 12581 3620 12590 3640
rect 12503 3610 12590 3620
rect 12649 3640 12686 3650
rect 12649 3620 12657 3640
rect 12677 3620 12686 3640
rect 12830 3625 12873 3667
rect 13257 3656 13309 3658
rect 12736 3623 12873 3625
rect 12503 3609 12534 3610
rect 12649 3550 12686 3620
rect 12127 3549 12468 3550
rect 11857 3532 11895 3541
rect 12052 3544 12468 3549
rect 11857 3531 11894 3532
rect 11318 3503 11408 3509
rect 11318 3483 11334 3503
rect 11354 3501 11408 3503
rect 11354 3483 11379 3501
rect 11318 3481 11379 3483
rect 11399 3481 11408 3501
rect 11318 3475 11408 3481
rect 11331 3421 11368 3422
rect 11427 3421 11464 3422
rect 11483 3421 11519 3531
rect 11706 3510 11737 3531
rect 12052 3524 12055 3544
rect 12075 3524 12468 3544
rect 12652 3534 12686 3550
rect 12730 3602 12873 3623
rect 13255 3652 13688 3656
rect 13255 3646 13694 3652
rect 13255 3628 13276 3646
rect 13294 3628 13694 3646
rect 14488 3635 14519 3686
rect 14554 3715 14591 3785
rect 14857 3784 14894 3785
rect 14706 3725 14742 3726
rect 14554 3695 14563 3715
rect 14583 3695 14591 3715
rect 14554 3685 14591 3695
rect 14650 3715 14798 3725
rect 14898 3722 14994 3724
rect 14650 3695 14659 3715
rect 14679 3695 14769 3715
rect 14789 3695 14798 3715
rect 14650 3686 14798 3695
rect 14856 3715 14994 3722
rect 14856 3695 14865 3715
rect 14885 3695 14994 3715
rect 14856 3686 14994 3695
rect 14650 3685 14687 3686
rect 14380 3632 14421 3633
rect 13255 3610 13694 3628
rect 12428 3515 12468 3524
rect 12730 3515 12757 3602
rect 12830 3576 12873 3602
rect 12830 3558 12843 3576
rect 12861 3558 12873 3576
rect 12830 3547 12873 3558
rect 11702 3509 11737 3510
rect 11580 3499 11737 3509
rect 11580 3479 11597 3499
rect 11617 3479 11737 3499
rect 11580 3472 11737 3479
rect 11804 3502 11953 3510
rect 11804 3482 11815 3502
rect 11835 3482 11874 3502
rect 11894 3482 11953 3502
rect 12428 3498 12757 3515
rect 12428 3497 12468 3498
rect 11804 3475 11953 3482
rect 12825 3486 12865 3489
rect 12825 3480 12868 3486
rect 12450 3477 12868 3480
rect 11804 3474 11845 3475
rect 11538 3421 11575 3422
rect 11231 3412 11369 3421
rect 11231 3392 11340 3412
rect 11360 3392 11369 3412
rect 11231 3385 11369 3392
rect 11427 3412 11575 3421
rect 11427 3392 11436 3412
rect 11456 3392 11546 3412
rect 11566 3392 11575 3412
rect 11231 3383 11327 3385
rect 11427 3382 11575 3392
rect 11634 3412 11671 3422
rect 11634 3392 11642 3412
rect 11662 3392 11671 3412
rect 11483 3381 11519 3382
rect 11331 3322 11368 3323
rect 11634 3322 11671 3392
rect 11706 3421 11737 3472
rect 12450 3459 12841 3477
rect 12859 3459 12868 3477
rect 12450 3457 12868 3459
rect 12450 3449 12477 3457
rect 12718 3454 12868 3457
rect 12030 3443 12198 3444
rect 12449 3443 12477 3449
rect 12030 3427 12477 3443
rect 12825 3449 12868 3454
rect 11756 3421 11793 3422
rect 11706 3412 11793 3421
rect 11706 3392 11764 3412
rect 11784 3392 11793 3412
rect 11706 3382 11793 3392
rect 11852 3412 11889 3422
rect 11852 3392 11860 3412
rect 11880 3392 11889 3412
rect 11706 3381 11737 3382
rect 11330 3321 11671 3322
rect 11852 3321 11889 3392
rect 11255 3316 11671 3321
rect 11255 3296 11258 3316
rect 11278 3296 11671 3316
rect 11702 3297 11889 3321
rect 12030 3417 12474 3427
rect 12030 3415 12198 3417
rect 11097 3222 11126 3240
rect 12030 3237 12057 3415
rect 12097 3377 12161 3389
rect 12437 3385 12474 3417
rect 12500 3416 12691 3438
rect 12655 3414 12691 3416
rect 12655 3385 12692 3414
rect 12825 3393 12865 3449
rect 12097 3376 12132 3377
rect 12074 3371 12132 3376
rect 12074 3351 12077 3371
rect 12097 3357 12132 3371
rect 12152 3357 12161 3377
rect 12097 3349 12161 3357
rect 12123 3348 12161 3349
rect 12124 3347 12161 3348
rect 12227 3381 12263 3382
rect 12335 3381 12371 3382
rect 12227 3373 12371 3381
rect 12227 3353 12235 3373
rect 12255 3353 12290 3373
rect 12310 3353 12343 3373
rect 12363 3353 12371 3373
rect 12227 3347 12371 3353
rect 12437 3377 12475 3385
rect 12553 3381 12589 3382
rect 12437 3357 12446 3377
rect 12466 3357 12475 3377
rect 12437 3348 12475 3357
rect 12504 3373 12589 3381
rect 12504 3353 12561 3373
rect 12581 3353 12589 3373
rect 12437 3347 12474 3348
rect 12504 3347 12589 3353
rect 12655 3377 12693 3385
rect 12655 3357 12664 3377
rect 12684 3357 12693 3377
rect 12825 3375 12837 3393
rect 12855 3375 12865 3393
rect 13257 3421 13309 3610
rect 13655 3585 13694 3610
rect 14272 3625 14421 3632
rect 14272 3605 14331 3625
rect 14351 3605 14390 3625
rect 14410 3605 14421 3625
rect 14272 3597 14421 3605
rect 14488 3628 14645 3635
rect 14488 3608 14608 3628
rect 14628 3608 14645 3628
rect 14488 3598 14645 3608
rect 14488 3597 14523 3598
rect 13439 3560 13626 3584
rect 13655 3565 14050 3585
rect 14070 3565 14073 3585
rect 14488 3576 14519 3597
rect 14706 3576 14742 3686
rect 14761 3685 14798 3686
rect 14857 3685 14894 3686
rect 14817 3626 14907 3632
rect 14817 3606 14826 3626
rect 14846 3624 14907 3626
rect 14846 3606 14871 3624
rect 14817 3604 14871 3606
rect 14891 3604 14907 3624
rect 14817 3598 14907 3604
rect 14331 3575 14368 3576
rect 13655 3560 14073 3565
rect 14330 3566 14368 3575
rect 13439 3489 13476 3560
rect 13655 3559 13998 3560
rect 13655 3556 13694 3559
rect 13960 3558 13997 3559
rect 13591 3499 13622 3500
rect 13439 3469 13448 3489
rect 13468 3469 13476 3489
rect 13439 3459 13476 3469
rect 13535 3489 13622 3499
rect 13535 3469 13544 3489
rect 13564 3469 13622 3489
rect 13535 3460 13622 3469
rect 13535 3459 13572 3460
rect 13257 3403 13273 3421
rect 13291 3403 13309 3421
rect 13591 3409 13622 3460
rect 13657 3489 13694 3556
rect 14330 3546 14339 3566
rect 14359 3546 14368 3566
rect 14330 3538 14368 3546
rect 14434 3570 14519 3576
rect 14549 3575 14586 3576
rect 14434 3550 14442 3570
rect 14462 3550 14519 3570
rect 14434 3542 14519 3550
rect 14548 3566 14586 3575
rect 14548 3546 14557 3566
rect 14577 3546 14586 3566
rect 14434 3541 14470 3542
rect 14548 3538 14586 3546
rect 14652 3571 14796 3576
rect 14652 3570 14714 3571
rect 14652 3550 14660 3570
rect 14680 3552 14714 3570
rect 14735 3570 14796 3571
rect 14735 3552 14768 3570
rect 14680 3550 14768 3552
rect 14788 3550 14796 3570
rect 14652 3542 14796 3550
rect 14652 3541 14688 3542
rect 14760 3541 14796 3542
rect 14862 3575 14899 3576
rect 14862 3574 14900 3575
rect 14862 3566 14926 3574
rect 14862 3546 14871 3566
rect 14891 3552 14926 3566
rect 14946 3552 14949 3572
rect 14891 3547 14949 3552
rect 14891 3546 14926 3547
rect 14331 3509 14368 3538
rect 14332 3507 14368 3509
rect 13809 3499 13845 3500
rect 13657 3469 13666 3489
rect 13686 3469 13694 3489
rect 13657 3459 13694 3469
rect 13753 3489 13901 3499
rect 14001 3496 14097 3498
rect 13753 3469 13762 3489
rect 13782 3469 13872 3489
rect 13892 3469 13901 3489
rect 13753 3460 13901 3469
rect 13959 3489 14097 3496
rect 13959 3469 13968 3489
rect 13988 3469 14097 3489
rect 14332 3485 14523 3507
rect 14549 3506 14586 3538
rect 14862 3534 14926 3546
rect 14966 3508 14993 3686
rect 14825 3506 14993 3508
rect 14549 3492 14993 3506
rect 14549 3480 14996 3492
rect 14592 3478 14625 3480
rect 13959 3460 14097 3469
rect 13753 3459 13790 3460
rect 13483 3406 13524 3407
rect 13257 3385 13309 3403
rect 13375 3399 13524 3406
rect 12825 3365 12865 3375
rect 13375 3379 13434 3399
rect 13454 3379 13493 3399
rect 13513 3379 13524 3399
rect 13375 3371 13524 3379
rect 13591 3402 13748 3409
rect 13591 3382 13711 3402
rect 13731 3382 13748 3402
rect 13591 3372 13748 3382
rect 13591 3371 13626 3372
rect 12655 3348 12693 3357
rect 13591 3350 13622 3371
rect 13809 3350 13845 3460
rect 13864 3459 13901 3460
rect 13960 3459 13997 3460
rect 13920 3400 14010 3406
rect 13920 3380 13929 3400
rect 13949 3398 14010 3400
rect 13949 3380 13974 3398
rect 13920 3378 13974 3380
rect 13994 3378 14010 3398
rect 13920 3372 14010 3378
rect 13434 3349 13471 3350
rect 12655 3347 12692 3348
rect 12116 3319 12206 3325
rect 12116 3299 12132 3319
rect 12152 3317 12206 3319
rect 12152 3299 12177 3317
rect 12116 3297 12177 3299
rect 12197 3297 12206 3317
rect 12116 3291 12206 3297
rect 12129 3237 12166 3238
rect 12225 3237 12262 3238
rect 12281 3237 12317 3347
rect 12504 3326 12535 3347
rect 13433 3340 13471 3349
rect 12500 3325 12535 3326
rect 12378 3315 12535 3325
rect 12378 3295 12395 3315
rect 12415 3295 12535 3315
rect 12378 3288 12535 3295
rect 12602 3318 12751 3326
rect 12602 3298 12613 3318
rect 12633 3298 12672 3318
rect 12692 3298 12751 3318
rect 13261 3322 13301 3332
rect 12602 3291 12751 3298
rect 12817 3294 12869 3312
rect 12602 3290 12643 3291
rect 12336 3237 12373 3238
rect 11067 3220 11126 3222
rect 12029 3228 12167 3237
rect 11067 3219 11235 3220
rect 11361 3219 11401 3221
rect 11067 3193 11511 3219
rect 11067 3191 11235 3193
rect 11067 3189 11148 3191
rect 11067 3013 11094 3189
rect 11134 3153 11198 3165
rect 11474 3161 11511 3193
rect 11537 3192 11728 3214
rect 12029 3208 12138 3228
rect 12158 3208 12167 3228
rect 12029 3201 12167 3208
rect 12225 3228 12373 3237
rect 12225 3208 12234 3228
rect 12254 3208 12344 3228
rect 12364 3208 12373 3228
rect 12029 3199 12125 3201
rect 12225 3198 12373 3208
rect 12432 3228 12469 3238
rect 12432 3208 12440 3228
rect 12460 3208 12469 3228
rect 12281 3197 12317 3198
rect 11692 3190 11728 3192
rect 11692 3161 11729 3190
rect 11134 3152 11169 3153
rect 11111 3147 11169 3152
rect 11111 3127 11114 3147
rect 11134 3133 11169 3147
rect 11189 3133 11198 3153
rect 11134 3125 11198 3133
rect 11160 3124 11198 3125
rect 11161 3123 11198 3124
rect 11264 3157 11300 3158
rect 11372 3157 11408 3158
rect 11264 3149 11408 3157
rect 11264 3129 11272 3149
rect 11292 3148 11380 3149
rect 11292 3130 11327 3148
rect 11345 3130 11380 3148
rect 11292 3129 11380 3130
rect 11400 3129 11408 3149
rect 11264 3123 11408 3129
rect 11474 3153 11512 3161
rect 11590 3157 11626 3158
rect 11474 3133 11483 3153
rect 11503 3133 11512 3153
rect 11474 3124 11512 3133
rect 11541 3149 11626 3157
rect 11541 3129 11598 3149
rect 11618 3129 11626 3149
rect 11474 3123 11511 3124
rect 11541 3123 11626 3129
rect 11692 3153 11730 3161
rect 11692 3133 11701 3153
rect 11721 3133 11730 3153
rect 12432 3141 12469 3208
rect 12504 3237 12535 3288
rect 12817 3276 12835 3294
rect 12853 3276 12869 3294
rect 12554 3237 12591 3238
rect 12504 3228 12591 3237
rect 12504 3208 12562 3228
rect 12582 3208 12591 3228
rect 12504 3198 12591 3208
rect 12650 3228 12687 3238
rect 12650 3208 12658 3228
rect 12678 3208 12687 3228
rect 12504 3197 12535 3198
rect 12129 3138 12166 3139
rect 12432 3138 12471 3141
rect 12128 3137 12471 3138
rect 12650 3137 12687 3208
rect 11692 3124 11730 3133
rect 12053 3132 12471 3137
rect 11692 3123 11729 3124
rect 11153 3095 11243 3101
rect 11153 3075 11169 3095
rect 11189 3093 11243 3095
rect 11189 3075 11214 3093
rect 11153 3073 11214 3075
rect 11234 3073 11243 3093
rect 11153 3067 11243 3073
rect 11166 3013 11203 3014
rect 11262 3013 11299 3014
rect 11318 3013 11354 3123
rect 11541 3102 11572 3123
rect 12053 3112 12056 3132
rect 12076 3112 12471 3132
rect 12500 3113 12687 3137
rect 11537 3101 11572 3102
rect 11415 3091 11572 3101
rect 11415 3071 11432 3091
rect 11452 3071 11572 3091
rect 11415 3064 11572 3071
rect 11639 3094 11788 3102
rect 11639 3074 11650 3094
rect 11670 3074 11709 3094
rect 11729 3074 11788 3094
rect 11639 3067 11788 3074
rect 12432 3087 12471 3112
rect 12817 3087 12869 3276
rect 13261 3304 13271 3322
rect 13289 3304 13301 3322
rect 13433 3320 13442 3340
rect 13462 3320 13471 3340
rect 13433 3312 13471 3320
rect 13537 3344 13622 3350
rect 13652 3349 13689 3350
rect 13537 3324 13545 3344
rect 13565 3324 13622 3344
rect 13537 3316 13622 3324
rect 13651 3340 13689 3349
rect 13651 3320 13660 3340
rect 13680 3320 13689 3340
rect 13537 3315 13573 3316
rect 13651 3312 13689 3320
rect 13755 3344 13899 3350
rect 13755 3324 13763 3344
rect 13783 3324 13816 3344
rect 13836 3324 13871 3344
rect 13891 3324 13899 3344
rect 13755 3316 13899 3324
rect 13755 3315 13791 3316
rect 13863 3315 13899 3316
rect 13965 3349 14002 3350
rect 13965 3348 14003 3349
rect 13965 3340 14029 3348
rect 13965 3320 13974 3340
rect 13994 3326 14029 3340
rect 14049 3326 14052 3346
rect 13994 3321 14052 3326
rect 13994 3320 14029 3321
rect 13261 3248 13301 3304
rect 13434 3283 13471 3312
rect 13435 3281 13471 3283
rect 13435 3259 13626 3281
rect 13652 3280 13689 3312
rect 13965 3308 14029 3320
rect 14069 3282 14096 3460
rect 14954 3435 14996 3480
rect 13928 3280 14096 3282
rect 13652 3270 14096 3280
rect 14237 3376 14424 3400
rect 14455 3381 14848 3401
rect 14868 3381 14871 3401
rect 14455 3376 14871 3381
rect 14237 3305 14274 3376
rect 14455 3375 14796 3376
rect 14389 3315 14420 3316
rect 14237 3285 14246 3305
rect 14266 3285 14274 3305
rect 14237 3275 14274 3285
rect 14333 3305 14420 3315
rect 14333 3285 14342 3305
rect 14362 3285 14420 3305
rect 14333 3276 14420 3285
rect 14333 3275 14370 3276
rect 13258 3243 13301 3248
rect 13649 3254 14096 3270
rect 13649 3248 13677 3254
rect 13928 3253 14096 3254
rect 13258 3240 13408 3243
rect 13649 3240 13676 3248
rect 13258 3238 13676 3240
rect 13258 3220 13267 3238
rect 13285 3220 13676 3238
rect 14389 3225 14420 3276
rect 14455 3305 14492 3375
rect 14758 3374 14795 3375
rect 14607 3315 14643 3316
rect 14455 3285 14464 3305
rect 14484 3285 14492 3305
rect 14455 3275 14492 3285
rect 14551 3305 14699 3315
rect 14799 3312 14895 3314
rect 14551 3285 14560 3305
rect 14580 3285 14670 3305
rect 14690 3285 14699 3305
rect 14551 3276 14699 3285
rect 14757 3305 14895 3312
rect 14757 3285 14766 3305
rect 14786 3285 14895 3305
rect 14757 3276 14895 3285
rect 14551 3275 14588 3276
rect 14281 3222 14322 3223
rect 13258 3217 13676 3220
rect 13258 3211 13301 3217
rect 13261 3208 13301 3211
rect 14176 3215 14322 3222
rect 13658 3199 13698 3200
rect 13369 3182 13698 3199
rect 14176 3195 14232 3215
rect 14252 3195 14291 3215
rect 14311 3195 14322 3215
rect 14176 3187 14322 3195
rect 14389 3218 14546 3225
rect 14389 3198 14509 3218
rect 14529 3198 14546 3218
rect 14389 3188 14546 3198
rect 14389 3187 14424 3188
rect 13253 3139 13296 3150
rect 13253 3121 13265 3139
rect 13283 3121 13296 3139
rect 13253 3095 13296 3121
rect 13369 3095 13396 3182
rect 13658 3173 13698 3182
rect 12432 3069 12871 3087
rect 11639 3066 11680 3067
rect 11373 3013 11410 3014
rect 11066 3004 11204 3013
rect 11066 2984 11175 3004
rect 11195 2984 11204 3004
rect 11066 2977 11204 2984
rect 11262 3004 11410 3013
rect 11262 2984 11271 3004
rect 11291 2984 11381 3004
rect 11401 2984 11410 3004
rect 11066 2975 11162 2977
rect 11262 2974 11410 2984
rect 11469 3004 11506 3014
rect 11469 2984 11477 3004
rect 11497 2984 11506 3004
rect 11318 2973 11354 2974
rect 11166 2914 11203 2915
rect 11469 2914 11506 2984
rect 11541 3013 11572 3064
rect 12432 3051 12832 3069
rect 12850 3051 12871 3069
rect 12432 3045 12871 3051
rect 12438 3041 12871 3045
rect 13253 3074 13396 3095
rect 13440 3147 13474 3163
rect 13658 3153 14051 3173
rect 14071 3153 14074 3173
rect 14389 3166 14420 3187
rect 14607 3166 14643 3276
rect 14662 3275 14699 3276
rect 14758 3275 14795 3276
rect 14718 3216 14808 3222
rect 14718 3196 14727 3216
rect 14747 3214 14808 3216
rect 14747 3196 14772 3214
rect 14718 3194 14772 3196
rect 14792 3194 14808 3214
rect 14718 3188 14808 3194
rect 14232 3165 14269 3166
rect 13658 3148 14074 3153
rect 14231 3156 14269 3165
rect 13658 3147 13999 3148
rect 13440 3077 13477 3147
rect 13592 3087 13623 3088
rect 13253 3072 13390 3074
rect 12817 3039 12869 3041
rect 13253 3030 13296 3072
rect 13440 3057 13449 3077
rect 13469 3057 13477 3077
rect 13440 3047 13477 3057
rect 13536 3077 13623 3087
rect 13536 3057 13545 3077
rect 13565 3057 13623 3077
rect 13536 3048 13623 3057
rect 13536 3047 13573 3048
rect 13251 3020 13296 3030
rect 11591 3013 11628 3014
rect 11541 3004 11628 3013
rect 11541 2984 11599 3004
rect 11619 2984 11628 3004
rect 11541 2974 11628 2984
rect 11687 3004 11724 3014
rect 11687 2984 11695 3004
rect 11715 2984 11724 3004
rect 13251 3002 13260 3020
rect 13278 3002 13296 3020
rect 13251 2996 13296 3002
rect 13592 2997 13623 3048
rect 13658 3077 13695 3147
rect 13961 3146 13998 3147
rect 14231 3136 14240 3156
rect 14260 3136 14269 3156
rect 14231 3128 14269 3136
rect 14335 3160 14420 3166
rect 14450 3165 14487 3166
rect 14335 3140 14343 3160
rect 14363 3140 14420 3160
rect 14335 3132 14420 3140
rect 14449 3156 14487 3165
rect 14449 3136 14458 3156
rect 14478 3136 14487 3156
rect 14335 3131 14371 3132
rect 14449 3128 14487 3136
rect 14553 3160 14697 3166
rect 14553 3140 14561 3160
rect 14581 3157 14669 3160
rect 14581 3140 14616 3157
rect 14553 3139 14616 3140
rect 14635 3140 14669 3157
rect 14689 3140 14697 3160
rect 14635 3139 14697 3140
rect 14553 3132 14697 3139
rect 14553 3131 14589 3132
rect 14661 3131 14697 3132
rect 14763 3165 14800 3166
rect 14763 3164 14801 3165
rect 14823 3164 14850 3168
rect 14763 3162 14850 3164
rect 14763 3156 14827 3162
rect 14763 3136 14772 3156
rect 14792 3142 14827 3156
rect 14847 3142 14850 3162
rect 14792 3137 14850 3142
rect 14792 3136 14827 3137
rect 14232 3099 14269 3128
rect 14233 3097 14269 3099
rect 13810 3087 13846 3088
rect 13658 3057 13667 3077
rect 13687 3057 13695 3077
rect 13658 3047 13695 3057
rect 13754 3077 13902 3087
rect 14002 3084 14098 3086
rect 13754 3057 13763 3077
rect 13783 3057 13873 3077
rect 13893 3057 13902 3077
rect 13754 3048 13902 3057
rect 13960 3077 14098 3084
rect 13960 3057 13969 3077
rect 13989 3057 14098 3077
rect 14233 3075 14424 3097
rect 14450 3096 14487 3128
rect 14763 3124 14827 3136
rect 14867 3098 14894 3276
rect 14726 3096 14894 3098
rect 14450 3070 14894 3096
rect 13960 3048 14098 3057
rect 13754 3047 13791 3048
rect 13251 2993 13288 2996
rect 13484 2994 13525 2995
rect 11541 2973 11572 2974
rect 11165 2913 11506 2914
rect 11687 2913 11724 2984
rect 13376 2987 13525 2994
rect 12820 2974 12857 2979
rect 11090 2908 11506 2913
rect 11090 2888 11093 2908
rect 11113 2888 11506 2908
rect 11537 2889 11724 2913
rect 12811 2970 12858 2974
rect 12811 2952 12830 2970
rect 12848 2952 12858 2970
rect 13376 2967 13435 2987
rect 13455 2967 13494 2987
rect 13514 2967 13525 2987
rect 13376 2959 13525 2967
rect 13592 2990 13749 2997
rect 13592 2970 13712 2990
rect 13732 2970 13749 2990
rect 13592 2960 13749 2970
rect 13592 2959 13627 2960
rect 12811 2904 12858 2952
rect 13592 2938 13623 2959
rect 13810 2938 13846 3048
rect 13865 3047 13902 3048
rect 13961 3047 13998 3048
rect 13921 2988 14011 2994
rect 13921 2968 13930 2988
rect 13950 2986 14011 2988
rect 13950 2968 13975 2986
rect 13921 2966 13975 2968
rect 13995 2966 14011 2986
rect 13921 2960 14011 2966
rect 13435 2937 13472 2938
rect 12435 2901 12858 2904
rect 11310 2887 11375 2888
rect 12413 2871 12858 2901
rect 13247 2929 13285 2931
rect 13247 2921 13290 2929
rect 13247 2903 13258 2921
rect 13276 2903 13290 2921
rect 13247 2876 13290 2903
rect 13434 2928 13472 2937
rect 13434 2908 13443 2928
rect 13463 2908 13472 2928
rect 13434 2900 13472 2908
rect 13538 2932 13623 2938
rect 13653 2937 13690 2938
rect 13538 2912 13546 2932
rect 13566 2912 13623 2932
rect 13538 2904 13623 2912
rect 13652 2928 13690 2937
rect 13652 2908 13661 2928
rect 13681 2908 13690 2928
rect 13538 2903 13574 2904
rect 13652 2900 13690 2908
rect 13756 2936 13900 2938
rect 13756 2932 13808 2936
rect 13756 2912 13764 2932
rect 13784 2916 13808 2932
rect 13828 2932 13900 2936
rect 13828 2916 13872 2932
rect 13784 2912 13872 2916
rect 13892 2912 13900 2932
rect 13756 2904 13900 2912
rect 13756 2903 13792 2904
rect 13864 2903 13900 2904
rect 13966 2937 14003 2938
rect 13966 2936 14004 2937
rect 13966 2928 14030 2936
rect 13966 2908 13975 2928
rect 13995 2914 14030 2928
rect 14050 2914 14053 2934
rect 13995 2909 14053 2914
rect 13995 2908 14030 2909
rect 11506 2855 11546 2863
rect 11506 2833 11514 2855
rect 11538 2833 11546 2855
rect 11111 2604 11148 2610
rect 11111 2585 11119 2604
rect 11140 2585 11148 2604
rect 11111 2577 11148 2585
rect 10811 2456 10818 2478
rect 10842 2456 10850 2478
rect 10811 2450 10850 2456
rect 10341 2445 10381 2447
rect 10507 2446 10675 2447
rect 10609 2445 10646 2446
rect 9575 2429 9713 2438
rect 9369 2428 9406 2429
rect 9099 2375 9140 2376
rect 8873 2354 8925 2372
rect 8991 2368 9140 2375
rect 8428 2335 8468 2345
rect 8991 2348 9050 2368
rect 9070 2348 9109 2368
rect 9129 2348 9140 2368
rect 8991 2340 9140 2348
rect 9207 2371 9364 2378
rect 9207 2351 9327 2371
rect 9347 2351 9364 2371
rect 9207 2341 9364 2351
rect 9207 2340 9242 2341
rect 8258 2318 8296 2327
rect 9207 2319 9238 2340
rect 9425 2319 9461 2429
rect 9480 2428 9517 2429
rect 9576 2428 9613 2429
rect 9536 2369 9626 2375
rect 9536 2349 9545 2369
rect 9565 2367 9626 2369
rect 9565 2349 9590 2367
rect 9536 2347 9590 2349
rect 9610 2347 9626 2367
rect 9536 2341 9626 2347
rect 9050 2318 9087 2319
rect 8258 2317 8295 2318
rect 7719 2289 7809 2295
rect 7719 2269 7735 2289
rect 7755 2287 7809 2289
rect 7755 2269 7780 2287
rect 7719 2267 7780 2269
rect 7800 2267 7809 2287
rect 7719 2261 7809 2267
rect 7732 2207 7769 2208
rect 7828 2207 7865 2208
rect 7884 2207 7920 2317
rect 8107 2296 8138 2317
rect 9049 2309 9087 2318
rect 8103 2295 8138 2296
rect 7981 2285 8138 2295
rect 7981 2265 7998 2285
rect 8018 2265 8138 2285
rect 7981 2258 8138 2265
rect 8205 2288 8354 2296
rect 8205 2268 8216 2288
rect 8236 2268 8275 2288
rect 8295 2268 8354 2288
rect 8877 2291 8917 2301
rect 8205 2261 8354 2268
rect 8420 2264 8472 2282
rect 8205 2260 8246 2261
rect 7939 2207 7976 2208
rect 7632 2198 7770 2207
rect 7104 2187 7137 2189
rect 6733 2175 7180 2187
rect 5965 2053 6133 2055
rect 5689 2027 6133 2053
rect 5199 2005 5337 2014
rect 4993 2004 5030 2005
rect 4490 1950 4527 1953
rect 4723 1951 4764 1952
rect 2846 1928 2877 1929
rect 2470 1868 2811 1869
rect 2992 1868 3029 1939
rect 4615 1944 4764 1951
rect 4059 1931 4096 1936
rect 4050 1927 4097 1931
rect 4050 1909 4069 1927
rect 4087 1909 4097 1927
rect 4615 1924 4674 1944
rect 4694 1924 4733 1944
rect 4753 1924 4764 1944
rect 4615 1916 4764 1924
rect 4831 1947 4988 1954
rect 4831 1927 4951 1947
rect 4971 1927 4988 1947
rect 4831 1917 4988 1927
rect 4831 1916 4866 1917
rect 2395 1863 2811 1868
rect 2395 1843 2398 1863
rect 2418 1843 2811 1863
rect 2842 1844 3029 1868
rect 3654 1866 3694 1871
rect 4050 1866 4097 1909
rect 4831 1895 4862 1916
rect 5049 1895 5085 2005
rect 5104 2004 5141 2005
rect 5200 2004 5237 2005
rect 5160 1945 5250 1951
rect 5160 1925 5169 1945
rect 5189 1943 5250 1945
rect 5189 1925 5214 1943
rect 5160 1923 5214 1925
rect 5234 1923 5250 1943
rect 5160 1917 5250 1923
rect 4674 1894 4711 1895
rect 3654 1827 4097 1866
rect 4487 1886 4524 1888
rect 4487 1878 4529 1886
rect 4487 1860 4497 1878
rect 4515 1860 4529 1878
rect 4487 1851 4529 1860
rect 4673 1885 4711 1894
rect 4673 1865 4682 1885
rect 4702 1865 4711 1885
rect 4673 1857 4711 1865
rect 4777 1889 4862 1895
rect 4892 1894 4929 1895
rect 4777 1869 4785 1889
rect 4805 1869 4862 1889
rect 4777 1861 4862 1869
rect 4891 1885 4929 1894
rect 4891 1865 4900 1885
rect 4920 1865 4929 1885
rect 4777 1860 4813 1861
rect 4891 1857 4929 1865
rect 4995 1893 5139 1895
rect 4995 1889 5047 1893
rect 4995 1869 5003 1889
rect 5023 1873 5047 1889
rect 5067 1889 5139 1893
rect 5067 1873 5111 1889
rect 5023 1869 5111 1873
rect 5131 1869 5139 1889
rect 4995 1861 5139 1869
rect 4995 1860 5031 1861
rect 5103 1860 5139 1861
rect 5205 1894 5242 1895
rect 5205 1893 5243 1894
rect 5205 1885 5269 1893
rect 5205 1865 5214 1885
rect 5234 1871 5269 1885
rect 5289 1871 5292 1891
rect 5234 1866 5292 1871
rect 5234 1865 5269 1866
rect 1435 1768 1443 1790
rect 1467 1768 1475 1790
rect 1435 1760 1475 1768
rect 2748 1812 2788 1820
rect 2748 1790 2756 1812
rect 2780 1790 2788 1812
rect 126 1714 569 1753
rect 126 1671 173 1714
rect 529 1709 569 1714
rect 1194 1712 1381 1736
rect 1412 1717 1805 1737
rect 1825 1717 1828 1737
rect 1412 1712 1828 1717
rect 126 1653 136 1671
rect 154 1653 173 1671
rect 126 1649 173 1653
rect 127 1644 164 1649
rect 1194 1641 1231 1712
rect 1412 1711 1753 1712
rect 1346 1651 1377 1652
rect 1194 1621 1203 1641
rect 1223 1621 1231 1641
rect 1194 1611 1231 1621
rect 1290 1641 1377 1651
rect 1290 1621 1299 1641
rect 1319 1621 1377 1641
rect 1290 1612 1377 1621
rect 1290 1611 1327 1612
rect 115 1582 167 1584
rect 113 1578 546 1582
rect 113 1572 552 1578
rect 113 1554 134 1572
rect 152 1554 552 1572
rect 1346 1561 1377 1612
rect 1412 1641 1449 1711
rect 1715 1710 1752 1711
rect 1564 1651 1600 1652
rect 1412 1621 1421 1641
rect 1441 1621 1449 1641
rect 1412 1611 1449 1621
rect 1508 1641 1656 1651
rect 1756 1648 1852 1650
rect 1508 1621 1517 1641
rect 1537 1621 1627 1641
rect 1647 1621 1656 1641
rect 1508 1612 1656 1621
rect 1714 1641 1852 1648
rect 1714 1621 1723 1641
rect 1743 1621 1852 1641
rect 1714 1612 1852 1621
rect 1508 1611 1545 1612
rect 1238 1558 1279 1559
rect 113 1536 552 1554
rect 115 1347 167 1536
rect 513 1511 552 1536
rect 1130 1551 1279 1558
rect 1130 1531 1189 1551
rect 1209 1531 1248 1551
rect 1268 1531 1279 1551
rect 1130 1523 1279 1531
rect 1346 1554 1503 1561
rect 1346 1534 1466 1554
rect 1486 1534 1503 1554
rect 1346 1524 1503 1534
rect 1346 1523 1381 1524
rect 297 1486 484 1510
rect 513 1491 908 1511
rect 928 1491 931 1511
rect 1346 1502 1377 1523
rect 1564 1502 1600 1612
rect 1619 1611 1656 1612
rect 1715 1611 1752 1612
rect 1675 1552 1765 1558
rect 1675 1532 1684 1552
rect 1704 1550 1765 1552
rect 1704 1532 1729 1550
rect 1675 1530 1729 1532
rect 1749 1530 1765 1550
rect 1675 1524 1765 1530
rect 1189 1501 1226 1502
rect 513 1486 931 1491
rect 1188 1492 1226 1501
rect 297 1415 334 1486
rect 513 1485 856 1486
rect 513 1482 552 1485
rect 818 1484 855 1485
rect 449 1425 480 1426
rect 297 1395 306 1415
rect 326 1395 334 1415
rect 297 1385 334 1395
rect 393 1415 480 1425
rect 393 1395 402 1415
rect 422 1395 480 1415
rect 393 1386 480 1395
rect 393 1385 430 1386
rect 115 1329 131 1347
rect 149 1329 167 1347
rect 449 1335 480 1386
rect 515 1415 552 1482
rect 1188 1472 1197 1492
rect 1217 1472 1226 1492
rect 1188 1464 1226 1472
rect 1292 1496 1377 1502
rect 1407 1501 1444 1502
rect 1292 1476 1300 1496
rect 1320 1476 1377 1496
rect 1292 1468 1377 1476
rect 1406 1492 1444 1501
rect 1406 1472 1415 1492
rect 1435 1472 1444 1492
rect 1292 1467 1328 1468
rect 1406 1464 1444 1472
rect 1510 1496 1654 1502
rect 1510 1476 1518 1496
rect 1538 1491 1626 1496
rect 1538 1476 1574 1491
rect 1510 1474 1574 1476
rect 1593 1476 1626 1491
rect 1646 1476 1654 1496
rect 1593 1474 1654 1476
rect 1510 1468 1654 1474
rect 1510 1467 1546 1468
rect 1618 1467 1654 1468
rect 1720 1501 1757 1502
rect 1720 1500 1758 1501
rect 1720 1492 1784 1500
rect 1720 1472 1729 1492
rect 1749 1478 1784 1492
rect 1804 1478 1807 1498
rect 1749 1473 1807 1478
rect 1749 1472 1784 1473
rect 1189 1435 1226 1464
rect 1190 1433 1226 1435
rect 667 1425 703 1426
rect 515 1395 524 1415
rect 544 1395 552 1415
rect 515 1385 552 1395
rect 611 1415 759 1425
rect 859 1422 955 1424
rect 611 1395 620 1415
rect 640 1395 730 1415
rect 750 1395 759 1415
rect 611 1386 759 1395
rect 817 1415 955 1422
rect 817 1395 826 1415
rect 846 1395 955 1415
rect 1190 1411 1381 1433
rect 1407 1432 1444 1464
rect 1720 1460 1784 1472
rect 1824 1434 1851 1612
rect 1683 1432 1851 1434
rect 1407 1418 1851 1432
rect 2454 1566 2622 1567
rect 2748 1566 2788 1790
rect 3251 1794 3419 1795
rect 3654 1794 3694 1827
rect 4050 1794 4097 1827
rect 4488 1826 4529 1851
rect 4674 1826 4711 1857
rect 4892 1826 4929 1857
rect 5205 1853 5269 1865
rect 5309 1827 5336 2005
rect 4488 1799 4537 1826
rect 4673 1800 4722 1826
rect 4891 1825 4972 1826
rect 5168 1825 5336 1827
rect 4891 1800 5336 1825
rect 4892 1799 5336 1800
rect 3251 1793 3695 1794
rect 3251 1768 3696 1793
rect 3251 1766 3419 1768
rect 3615 1767 3696 1768
rect 3865 1767 3914 1793
rect 4050 1767 4099 1794
rect 3251 1588 3278 1766
rect 3318 1728 3382 1740
rect 3658 1736 3695 1767
rect 3876 1736 3913 1767
rect 4058 1742 4099 1767
rect 4490 1766 4537 1799
rect 4893 1766 4933 1799
rect 5168 1798 5336 1799
rect 5799 1803 5839 2027
rect 5965 2026 6133 2027
rect 6736 2161 7180 2175
rect 6736 2159 6904 2161
rect 6736 1981 6763 2159
rect 6803 2121 6867 2133
rect 7143 2129 7180 2161
rect 7206 2160 7397 2182
rect 7632 2178 7741 2198
rect 7761 2178 7770 2198
rect 7632 2171 7770 2178
rect 7828 2198 7976 2207
rect 7828 2178 7837 2198
rect 7857 2178 7947 2198
rect 7967 2178 7976 2198
rect 7632 2169 7728 2171
rect 7828 2168 7976 2178
rect 8035 2198 8072 2208
rect 8035 2178 8043 2198
rect 8063 2178 8072 2198
rect 7884 2167 7920 2168
rect 7361 2158 7397 2160
rect 7361 2129 7398 2158
rect 6803 2120 6838 2121
rect 6780 2115 6838 2120
rect 6780 2095 6783 2115
rect 6803 2101 6838 2115
rect 6858 2101 6867 2121
rect 6803 2093 6867 2101
rect 6829 2092 6867 2093
rect 6830 2091 6867 2092
rect 6933 2125 6969 2126
rect 7041 2125 7077 2126
rect 6933 2117 7077 2125
rect 6933 2097 6941 2117
rect 6961 2115 7049 2117
rect 6961 2097 6994 2115
rect 6933 2096 6994 2097
rect 7015 2097 7049 2115
rect 7069 2097 7077 2117
rect 7015 2096 7077 2097
rect 6933 2091 7077 2096
rect 7143 2121 7181 2129
rect 7259 2125 7295 2126
rect 7143 2101 7152 2121
rect 7172 2101 7181 2121
rect 7143 2092 7181 2101
rect 7210 2117 7295 2125
rect 7210 2097 7267 2117
rect 7287 2097 7295 2117
rect 7143 2091 7180 2092
rect 7210 2091 7295 2097
rect 7361 2121 7399 2129
rect 7361 2101 7370 2121
rect 7390 2101 7399 2121
rect 8035 2111 8072 2178
rect 8107 2207 8138 2258
rect 8420 2246 8438 2264
rect 8456 2246 8472 2264
rect 8157 2207 8194 2208
rect 8107 2198 8194 2207
rect 8107 2178 8165 2198
rect 8185 2178 8194 2198
rect 8107 2168 8194 2178
rect 8253 2198 8290 2208
rect 8253 2178 8261 2198
rect 8281 2178 8290 2198
rect 8107 2167 8138 2168
rect 7732 2108 7769 2109
rect 8035 2108 8074 2111
rect 7731 2107 8074 2108
rect 8253 2107 8290 2178
rect 7361 2092 7399 2101
rect 7656 2102 8074 2107
rect 7361 2091 7398 2092
rect 6822 2063 6912 2069
rect 6822 2043 6838 2063
rect 6858 2061 6912 2063
rect 6858 2043 6883 2061
rect 6822 2041 6883 2043
rect 6903 2041 6912 2061
rect 6822 2035 6912 2041
rect 6835 1981 6872 1982
rect 6931 1981 6968 1982
rect 6987 1981 7023 2091
rect 7210 2070 7241 2091
rect 7656 2082 7659 2102
rect 7679 2082 8074 2102
rect 8103 2083 8290 2107
rect 7206 2069 7241 2070
rect 7084 2059 7241 2069
rect 7084 2039 7101 2059
rect 7121 2039 7241 2059
rect 7084 2032 7241 2039
rect 7308 2062 7457 2070
rect 7308 2042 7319 2062
rect 7339 2042 7378 2062
rect 7398 2042 7457 2062
rect 7308 2035 7457 2042
rect 8035 2057 8074 2082
rect 8420 2057 8472 2246
rect 8877 2273 8887 2291
rect 8905 2273 8917 2291
rect 9049 2289 9058 2309
rect 9078 2289 9087 2309
rect 9049 2281 9087 2289
rect 9153 2313 9238 2319
rect 9268 2318 9305 2319
rect 9153 2293 9161 2313
rect 9181 2293 9238 2313
rect 9153 2285 9238 2293
rect 9267 2309 9305 2318
rect 9267 2289 9276 2309
rect 9296 2289 9305 2309
rect 9153 2284 9189 2285
rect 9267 2281 9305 2289
rect 9371 2313 9515 2319
rect 9371 2293 9379 2313
rect 9399 2293 9432 2313
rect 9452 2293 9487 2313
rect 9507 2293 9515 2313
rect 9371 2285 9515 2293
rect 9371 2284 9407 2285
rect 9479 2284 9515 2285
rect 9581 2318 9618 2319
rect 9581 2317 9619 2318
rect 9581 2309 9645 2317
rect 9581 2289 9590 2309
rect 9610 2295 9645 2309
rect 9665 2295 9668 2315
rect 9610 2290 9668 2295
rect 9610 2289 9645 2290
rect 8877 2217 8917 2273
rect 9050 2252 9087 2281
rect 9051 2250 9087 2252
rect 9051 2228 9242 2250
rect 9268 2249 9305 2281
rect 9581 2277 9645 2289
rect 9685 2251 9712 2429
rect 9544 2249 9712 2251
rect 9268 2239 9712 2249
rect 9853 2345 10040 2369
rect 10071 2350 10464 2370
rect 10484 2350 10487 2370
rect 10071 2345 10487 2350
rect 9853 2274 9890 2345
rect 10071 2344 10412 2345
rect 10005 2284 10036 2285
rect 9853 2254 9862 2274
rect 9882 2254 9890 2274
rect 9853 2244 9890 2254
rect 9949 2274 10036 2284
rect 9949 2254 9958 2274
rect 9978 2254 10036 2274
rect 9949 2245 10036 2254
rect 9949 2244 9986 2245
rect 8874 2212 8917 2217
rect 9265 2223 9712 2239
rect 9265 2217 9293 2223
rect 9544 2222 9712 2223
rect 8874 2209 9024 2212
rect 9265 2209 9292 2217
rect 8874 2207 9292 2209
rect 8874 2189 8883 2207
rect 8901 2189 9292 2207
rect 10005 2194 10036 2245
rect 10071 2274 10108 2344
rect 10374 2343 10411 2344
rect 10612 2286 10645 2445
rect 10223 2284 10259 2285
rect 10071 2254 10080 2274
rect 10100 2254 10108 2274
rect 10071 2244 10108 2254
rect 10167 2274 10315 2284
rect 10415 2281 10511 2283
rect 10167 2254 10176 2274
rect 10196 2254 10286 2274
rect 10306 2254 10315 2274
rect 10167 2245 10315 2254
rect 10373 2274 10511 2281
rect 10373 2254 10382 2274
rect 10402 2254 10511 2274
rect 10612 2282 10648 2286
rect 10612 2264 10621 2282
rect 10643 2264 10648 2282
rect 10612 2258 10648 2264
rect 10373 2245 10511 2254
rect 10167 2244 10204 2245
rect 9897 2191 9938 2192
rect 8874 2186 9292 2189
rect 8874 2180 8917 2186
rect 8877 2177 8917 2180
rect 9789 2184 9938 2191
rect 9274 2168 9314 2169
rect 8985 2151 9314 2168
rect 9789 2164 9848 2184
rect 9868 2164 9907 2184
rect 9927 2164 9938 2184
rect 9789 2156 9938 2164
rect 10005 2187 10162 2194
rect 10005 2167 10125 2187
rect 10145 2167 10162 2187
rect 10005 2157 10162 2167
rect 10005 2156 10040 2157
rect 8869 2108 8912 2119
rect 8869 2090 8881 2108
rect 8899 2090 8912 2108
rect 8869 2064 8912 2090
rect 8985 2064 9012 2151
rect 9274 2142 9314 2151
rect 8035 2039 8474 2057
rect 7308 2034 7349 2035
rect 7042 1981 7079 1982
rect 6735 1972 6873 1981
rect 6735 1952 6844 1972
rect 6864 1952 6873 1972
rect 6735 1945 6873 1952
rect 6931 1972 7079 1981
rect 6931 1952 6940 1972
rect 6960 1952 7050 1972
rect 7070 1952 7079 1972
rect 6735 1943 6831 1945
rect 6931 1942 7079 1952
rect 7138 1972 7175 1982
rect 7138 1952 7146 1972
rect 7166 1952 7175 1972
rect 6987 1941 7023 1942
rect 6835 1882 6872 1883
rect 7138 1882 7175 1952
rect 7210 1981 7241 2032
rect 8035 2021 8435 2039
rect 8453 2021 8474 2039
rect 8035 2015 8474 2021
rect 8041 2011 8474 2015
rect 8869 2043 9012 2064
rect 9056 2116 9090 2132
rect 9274 2122 9667 2142
rect 9687 2122 9690 2142
rect 10005 2135 10036 2156
rect 10223 2135 10259 2245
rect 10278 2244 10315 2245
rect 10374 2244 10411 2245
rect 10334 2185 10424 2191
rect 10334 2165 10343 2185
rect 10363 2183 10424 2185
rect 10363 2165 10388 2183
rect 10334 2163 10388 2165
rect 10408 2163 10424 2183
rect 10334 2157 10424 2163
rect 9848 2134 9885 2135
rect 9274 2117 9690 2122
rect 9847 2125 9885 2134
rect 9274 2116 9615 2117
rect 9056 2046 9093 2116
rect 9208 2056 9239 2057
rect 8869 2041 9006 2043
rect 8420 2009 8472 2011
rect 8869 1999 8912 2041
rect 9056 2026 9065 2046
rect 9085 2026 9093 2046
rect 9056 2016 9093 2026
rect 9152 2046 9239 2056
rect 9152 2026 9161 2046
rect 9181 2026 9239 2046
rect 9152 2017 9239 2026
rect 9152 2016 9189 2017
rect 8867 1989 8912 1999
rect 7260 1981 7297 1982
rect 7210 1972 7297 1981
rect 7210 1952 7268 1972
rect 7288 1952 7297 1972
rect 7210 1942 7297 1952
rect 7356 1972 7393 1982
rect 7356 1952 7364 1972
rect 7384 1952 7393 1972
rect 8867 1971 8876 1989
rect 8894 1971 8912 1989
rect 8867 1965 8912 1971
rect 9208 1966 9239 2017
rect 9274 2046 9311 2116
rect 9577 2115 9614 2116
rect 9847 2105 9856 2125
rect 9876 2105 9885 2125
rect 9847 2097 9885 2105
rect 9951 2129 10036 2135
rect 10066 2134 10103 2135
rect 9951 2109 9959 2129
rect 9979 2109 10036 2129
rect 9951 2101 10036 2109
rect 10065 2125 10103 2134
rect 10065 2105 10074 2125
rect 10094 2105 10103 2125
rect 9951 2100 9987 2101
rect 10065 2097 10103 2105
rect 10169 2129 10313 2135
rect 10169 2109 10177 2129
rect 10197 2110 10229 2129
rect 10250 2110 10285 2129
rect 10197 2109 10285 2110
rect 10305 2109 10313 2129
rect 10169 2101 10313 2109
rect 10169 2100 10205 2101
rect 10277 2100 10313 2101
rect 10379 2134 10416 2135
rect 10379 2133 10417 2134
rect 10379 2125 10443 2133
rect 10379 2105 10388 2125
rect 10408 2111 10443 2125
rect 10463 2111 10466 2131
rect 10408 2106 10466 2111
rect 10408 2105 10443 2106
rect 9848 2068 9885 2097
rect 9849 2066 9885 2068
rect 9426 2056 9462 2057
rect 9274 2026 9283 2046
rect 9303 2026 9311 2046
rect 9274 2016 9311 2026
rect 9370 2046 9518 2056
rect 9618 2053 9714 2055
rect 9370 2026 9379 2046
rect 9399 2026 9489 2046
rect 9509 2026 9518 2046
rect 9370 2017 9518 2026
rect 9576 2046 9714 2053
rect 9576 2026 9585 2046
rect 9605 2026 9714 2046
rect 9849 2044 10040 2066
rect 10066 2065 10103 2097
rect 10379 2093 10443 2105
rect 10483 2067 10510 2245
rect 11115 2244 11148 2577
rect 11212 2609 11380 2610
rect 11506 2609 11546 2833
rect 12009 2837 12177 2838
rect 12413 2837 12454 2871
rect 12811 2850 12858 2871
rect 12009 2827 12454 2837
rect 12526 2835 12669 2836
rect 12009 2811 12453 2827
rect 12009 2809 12177 2811
rect 12373 2810 12453 2811
rect 12526 2810 12671 2835
rect 12813 2810 12858 2850
rect 12009 2631 12036 2809
rect 12076 2771 12140 2783
rect 12416 2779 12453 2810
rect 12634 2779 12671 2810
rect 12816 2803 12858 2810
rect 13248 2869 13290 2876
rect 13435 2869 13472 2900
rect 13653 2869 13690 2900
rect 13966 2896 14030 2908
rect 14070 2870 14097 3048
rect 13248 2829 13293 2869
rect 13435 2844 13580 2869
rect 13653 2868 13733 2869
rect 13929 2868 14097 2870
rect 13653 2852 14097 2868
rect 13437 2843 13580 2844
rect 13652 2842 14097 2852
rect 13248 2808 13295 2829
rect 13652 2808 13693 2842
rect 13929 2841 14097 2842
rect 14560 2846 14600 3070
rect 14726 3069 14894 3070
rect 14958 3102 14991 3435
rect 14958 3094 14995 3102
rect 14958 3075 14966 3094
rect 14987 3075 14995 3094
rect 14958 3069 14995 3075
rect 14560 2824 14568 2846
rect 14592 2824 14600 2846
rect 14560 2816 14600 2824
rect 12076 2770 12111 2771
rect 12053 2765 12111 2770
rect 12053 2745 12056 2765
rect 12076 2751 12111 2765
rect 12131 2751 12140 2771
rect 12076 2743 12140 2751
rect 12102 2742 12140 2743
rect 12103 2741 12140 2742
rect 12206 2775 12242 2776
rect 12314 2775 12350 2776
rect 12206 2767 12350 2775
rect 12206 2747 12214 2767
rect 12234 2763 12322 2767
rect 12234 2747 12278 2763
rect 12206 2743 12278 2747
rect 12298 2747 12322 2763
rect 12342 2747 12350 2767
rect 12298 2743 12350 2747
rect 12206 2741 12350 2743
rect 12416 2771 12454 2779
rect 12532 2775 12568 2776
rect 12416 2751 12425 2771
rect 12445 2751 12454 2771
rect 12416 2742 12454 2751
rect 12483 2767 12568 2775
rect 12483 2747 12540 2767
rect 12560 2747 12568 2767
rect 12416 2741 12453 2742
rect 12483 2741 12568 2747
rect 12634 2771 12672 2779
rect 12634 2751 12643 2771
rect 12663 2751 12672 2771
rect 12634 2742 12672 2751
rect 12816 2776 12859 2803
rect 12816 2758 12830 2776
rect 12848 2758 12859 2776
rect 12816 2750 12859 2758
rect 12821 2748 12859 2750
rect 13248 2778 13693 2808
rect 14731 2791 14796 2792
rect 13248 2775 13671 2778
rect 12634 2741 12671 2742
rect 12095 2713 12185 2719
rect 12095 2693 12111 2713
rect 12131 2711 12185 2713
rect 12131 2693 12156 2711
rect 12095 2691 12156 2693
rect 12176 2691 12185 2711
rect 12095 2685 12185 2691
rect 12108 2631 12145 2632
rect 12204 2631 12241 2632
rect 12260 2631 12296 2741
rect 12483 2720 12514 2741
rect 13248 2727 13295 2775
rect 12479 2719 12514 2720
rect 12357 2709 12514 2719
rect 12357 2689 12374 2709
rect 12394 2689 12514 2709
rect 12357 2682 12514 2689
rect 12581 2712 12730 2720
rect 12581 2692 12592 2712
rect 12612 2692 12651 2712
rect 12671 2692 12730 2712
rect 13248 2709 13258 2727
rect 13276 2709 13295 2727
rect 13248 2705 13295 2709
rect 14382 2766 14569 2790
rect 14600 2771 14993 2791
rect 15013 2771 15016 2791
rect 14600 2766 15016 2771
rect 13249 2700 13286 2705
rect 12581 2685 12730 2692
rect 14382 2695 14419 2766
rect 14600 2765 14941 2766
rect 14534 2705 14565 2706
rect 12581 2684 12622 2685
rect 12818 2683 12855 2686
rect 12315 2631 12352 2632
rect 12008 2622 12146 2631
rect 11212 2583 11656 2609
rect 11212 2581 11380 2583
rect 11212 2403 11239 2581
rect 11279 2543 11343 2555
rect 11619 2551 11656 2583
rect 11682 2582 11873 2604
rect 12008 2602 12117 2622
rect 12137 2602 12146 2622
rect 12008 2595 12146 2602
rect 12204 2622 12352 2631
rect 12204 2602 12213 2622
rect 12233 2602 12323 2622
rect 12343 2602 12352 2622
rect 12008 2593 12104 2595
rect 12204 2592 12352 2602
rect 12411 2622 12448 2632
rect 12411 2602 12419 2622
rect 12439 2602 12448 2622
rect 12260 2591 12296 2592
rect 11837 2580 11873 2582
rect 11837 2551 11874 2580
rect 11279 2542 11314 2543
rect 11256 2537 11314 2542
rect 11256 2517 11259 2537
rect 11279 2523 11314 2537
rect 11334 2523 11343 2543
rect 11279 2517 11343 2523
rect 11256 2515 11343 2517
rect 11256 2511 11283 2515
rect 11305 2514 11343 2515
rect 11306 2513 11343 2514
rect 11409 2547 11445 2548
rect 11517 2547 11553 2548
rect 11409 2540 11553 2547
rect 11409 2539 11471 2540
rect 11409 2519 11417 2539
rect 11437 2522 11471 2539
rect 11490 2539 11553 2540
rect 11490 2522 11525 2539
rect 11437 2519 11525 2522
rect 11545 2519 11553 2539
rect 11409 2513 11553 2519
rect 11619 2543 11657 2551
rect 11735 2547 11771 2548
rect 11619 2523 11628 2543
rect 11648 2523 11657 2543
rect 11619 2514 11657 2523
rect 11686 2539 11771 2547
rect 11686 2519 11743 2539
rect 11763 2519 11771 2539
rect 11619 2513 11656 2514
rect 11686 2513 11771 2519
rect 11837 2543 11875 2551
rect 11837 2523 11846 2543
rect 11866 2523 11875 2543
rect 12108 2532 12145 2533
rect 12411 2532 12448 2602
rect 12483 2631 12514 2682
rect 12810 2677 12855 2683
rect 12810 2659 12828 2677
rect 12846 2659 12855 2677
rect 14382 2675 14391 2695
rect 14411 2675 14419 2695
rect 14382 2665 14419 2675
rect 14478 2695 14565 2705
rect 14478 2675 14487 2695
rect 14507 2675 14565 2695
rect 14478 2666 14565 2675
rect 14478 2665 14515 2666
rect 12810 2649 12855 2659
rect 12533 2631 12570 2632
rect 12483 2622 12570 2631
rect 12483 2602 12541 2622
rect 12561 2602 12570 2622
rect 12483 2592 12570 2602
rect 12629 2622 12666 2632
rect 12629 2602 12637 2622
rect 12657 2602 12666 2622
rect 12810 2607 12853 2649
rect 13237 2638 13289 2640
rect 12716 2605 12853 2607
rect 12483 2591 12514 2592
rect 12629 2532 12666 2602
rect 12107 2531 12448 2532
rect 11837 2514 11875 2523
rect 12032 2526 12448 2531
rect 11837 2513 11874 2514
rect 11298 2485 11388 2491
rect 11298 2465 11314 2485
rect 11334 2483 11388 2485
rect 11334 2465 11359 2483
rect 11298 2463 11359 2465
rect 11379 2463 11388 2483
rect 11298 2457 11388 2463
rect 11311 2403 11348 2404
rect 11407 2403 11444 2404
rect 11463 2403 11499 2513
rect 11686 2492 11717 2513
rect 12032 2506 12035 2526
rect 12055 2506 12448 2526
rect 12632 2516 12666 2532
rect 12710 2584 12853 2605
rect 13235 2634 13668 2638
rect 13235 2628 13674 2634
rect 13235 2610 13256 2628
rect 13274 2610 13674 2628
rect 14534 2615 14565 2666
rect 14600 2695 14637 2765
rect 14903 2764 14940 2765
rect 14752 2705 14788 2706
rect 14600 2675 14609 2695
rect 14629 2675 14637 2695
rect 14600 2665 14637 2675
rect 14696 2695 14844 2705
rect 14944 2702 15040 2704
rect 14696 2675 14705 2695
rect 14725 2675 14815 2695
rect 14835 2675 14844 2695
rect 14696 2666 14844 2675
rect 14902 2695 15040 2702
rect 14902 2675 14911 2695
rect 14931 2675 15040 2695
rect 14902 2666 15040 2675
rect 14696 2665 14733 2666
rect 14426 2612 14467 2613
rect 13235 2592 13674 2610
rect 12408 2497 12448 2506
rect 12710 2497 12737 2584
rect 12810 2558 12853 2584
rect 12810 2540 12823 2558
rect 12841 2540 12853 2558
rect 12810 2529 12853 2540
rect 11682 2491 11717 2492
rect 11560 2481 11717 2491
rect 11560 2461 11577 2481
rect 11597 2461 11717 2481
rect 11560 2454 11717 2461
rect 11784 2484 11930 2492
rect 11784 2464 11795 2484
rect 11815 2464 11854 2484
rect 11874 2464 11930 2484
rect 12408 2480 12737 2497
rect 12408 2479 12448 2480
rect 11784 2457 11930 2464
rect 12805 2468 12845 2471
rect 12805 2462 12848 2468
rect 12430 2459 12848 2462
rect 11784 2456 11825 2457
rect 11518 2403 11555 2404
rect 11211 2394 11349 2403
rect 11211 2374 11320 2394
rect 11340 2374 11349 2394
rect 11211 2367 11349 2374
rect 11407 2394 11555 2403
rect 11407 2374 11416 2394
rect 11436 2374 11526 2394
rect 11546 2374 11555 2394
rect 11211 2365 11307 2367
rect 11407 2364 11555 2374
rect 11614 2394 11651 2404
rect 11614 2374 11622 2394
rect 11642 2374 11651 2394
rect 11463 2363 11499 2364
rect 11311 2304 11348 2305
rect 11614 2304 11651 2374
rect 11686 2403 11717 2454
rect 12430 2441 12821 2459
rect 12839 2441 12848 2459
rect 12430 2439 12848 2441
rect 12430 2431 12457 2439
rect 12698 2436 12848 2439
rect 12010 2425 12178 2426
rect 12429 2425 12457 2431
rect 12010 2409 12457 2425
rect 12805 2431 12848 2436
rect 11736 2403 11773 2404
rect 11686 2394 11773 2403
rect 11686 2374 11744 2394
rect 11764 2374 11773 2394
rect 11686 2364 11773 2374
rect 11832 2394 11869 2404
rect 11832 2374 11840 2394
rect 11860 2374 11869 2394
rect 11686 2363 11717 2364
rect 11310 2303 11651 2304
rect 11832 2303 11869 2374
rect 11235 2298 11651 2303
rect 11235 2278 11238 2298
rect 11258 2278 11651 2298
rect 11682 2279 11869 2303
rect 12010 2399 12454 2409
rect 12010 2397 12178 2399
rect 11110 2199 11152 2244
rect 12010 2219 12037 2397
rect 12077 2359 12141 2371
rect 12417 2367 12454 2399
rect 12480 2398 12671 2420
rect 12635 2396 12671 2398
rect 12635 2367 12672 2396
rect 12805 2375 12845 2431
rect 12077 2358 12112 2359
rect 12054 2353 12112 2358
rect 12054 2333 12057 2353
rect 12077 2339 12112 2353
rect 12132 2339 12141 2359
rect 12077 2331 12141 2339
rect 12103 2330 12141 2331
rect 12104 2329 12141 2330
rect 12207 2363 12243 2364
rect 12315 2363 12351 2364
rect 12207 2355 12351 2363
rect 12207 2335 12215 2355
rect 12235 2335 12270 2355
rect 12290 2335 12323 2355
rect 12343 2335 12351 2355
rect 12207 2329 12351 2335
rect 12417 2359 12455 2367
rect 12533 2363 12569 2364
rect 12417 2339 12426 2359
rect 12446 2339 12455 2359
rect 12417 2330 12455 2339
rect 12484 2355 12569 2363
rect 12484 2335 12541 2355
rect 12561 2335 12569 2355
rect 12417 2329 12454 2330
rect 12484 2329 12569 2335
rect 12635 2359 12673 2367
rect 12635 2339 12644 2359
rect 12664 2339 12673 2359
rect 12805 2357 12817 2375
rect 12835 2357 12845 2375
rect 13237 2403 13289 2592
rect 13635 2567 13674 2592
rect 14318 2605 14467 2612
rect 14318 2585 14377 2605
rect 14397 2585 14436 2605
rect 14456 2585 14467 2605
rect 14318 2577 14467 2585
rect 14534 2608 14691 2615
rect 14534 2588 14654 2608
rect 14674 2588 14691 2608
rect 14534 2578 14691 2588
rect 14534 2577 14569 2578
rect 13419 2542 13606 2566
rect 13635 2547 14030 2567
rect 14050 2547 14053 2567
rect 14534 2556 14565 2577
rect 14752 2556 14788 2666
rect 14807 2665 14844 2666
rect 14903 2665 14940 2666
rect 14863 2606 14953 2612
rect 14863 2586 14872 2606
rect 14892 2604 14953 2606
rect 14892 2586 14917 2604
rect 14863 2584 14917 2586
rect 14937 2584 14953 2604
rect 14863 2578 14953 2584
rect 14377 2555 14414 2556
rect 13635 2542 14053 2547
rect 14376 2546 14414 2555
rect 13419 2471 13456 2542
rect 13635 2541 13978 2542
rect 13635 2538 13674 2541
rect 13940 2540 13977 2541
rect 13571 2481 13602 2482
rect 13419 2451 13428 2471
rect 13448 2451 13456 2471
rect 13419 2441 13456 2451
rect 13515 2471 13602 2481
rect 13515 2451 13524 2471
rect 13544 2451 13602 2471
rect 13515 2442 13602 2451
rect 13515 2441 13552 2442
rect 13237 2385 13253 2403
rect 13271 2385 13289 2403
rect 13571 2391 13602 2442
rect 13637 2471 13674 2538
rect 14376 2526 14385 2546
rect 14405 2526 14414 2546
rect 14376 2518 14414 2526
rect 14480 2550 14565 2556
rect 14595 2555 14632 2556
rect 14480 2530 14488 2550
rect 14508 2530 14565 2550
rect 14480 2522 14565 2530
rect 14594 2546 14632 2555
rect 14594 2526 14603 2546
rect 14623 2526 14632 2546
rect 14480 2521 14516 2522
rect 14594 2518 14632 2526
rect 14698 2554 14842 2556
rect 14698 2550 14758 2554
rect 14698 2530 14706 2550
rect 14726 2532 14758 2550
rect 14781 2550 14842 2554
rect 14781 2532 14814 2550
rect 14726 2530 14814 2532
rect 14834 2530 14842 2550
rect 14698 2522 14842 2530
rect 14698 2521 14734 2522
rect 14806 2521 14842 2522
rect 14908 2555 14945 2556
rect 14908 2554 14946 2555
rect 14908 2546 14972 2554
rect 14908 2526 14917 2546
rect 14937 2532 14972 2546
rect 14992 2532 14995 2552
rect 14937 2527 14995 2532
rect 14937 2526 14972 2527
rect 14377 2489 14414 2518
rect 14378 2487 14414 2489
rect 13789 2481 13825 2482
rect 13637 2451 13646 2471
rect 13666 2451 13674 2471
rect 13637 2441 13674 2451
rect 13733 2471 13881 2481
rect 13981 2478 14077 2480
rect 13733 2451 13742 2471
rect 13762 2451 13852 2471
rect 13872 2451 13881 2471
rect 13733 2442 13881 2451
rect 13939 2471 14077 2478
rect 13939 2451 13948 2471
rect 13968 2451 14077 2471
rect 14378 2465 14569 2487
rect 14595 2486 14632 2518
rect 14908 2514 14972 2526
rect 14595 2485 14870 2486
rect 15012 2485 15039 2666
rect 14595 2460 15039 2485
rect 15175 2491 15214 4306
rect 15516 4293 15549 4626
rect 15613 4658 15781 4659
rect 15907 4658 15947 4882
rect 16410 4886 16578 4887
rect 16819 4886 16854 4903
rect 17211 4893 17258 4904
rect 16410 4860 16854 4886
rect 16410 4858 16578 4860
rect 16774 4859 16854 4860
rect 17009 4859 17076 4885
rect 17215 4859 17258 4893
rect 16410 4680 16437 4858
rect 16477 4820 16541 4832
rect 16817 4828 16854 4859
rect 17035 4828 17072 4859
rect 17217 4834 17258 4859
rect 17551 4879 17592 4904
rect 17737 4879 17774 4910
rect 17955 4879 17992 4910
rect 18268 4906 18332 4918
rect 18372 4880 18399 5058
rect 17551 4845 17594 4879
rect 17733 4853 17800 4879
rect 17955 4878 18035 4879
rect 18231 4878 18399 4880
rect 17955 4852 18399 4878
rect 17551 4834 17598 4845
rect 17955 4835 17990 4852
rect 18231 4851 18399 4852
rect 18862 4856 18902 5080
rect 19028 5079 19196 5080
rect 19260 5112 19293 5445
rect 19595 5432 19634 7247
rect 19770 7253 20214 7278
rect 19770 7072 19797 7253
rect 19939 7252 20214 7253
rect 19837 7212 19901 7224
rect 20177 7220 20214 7252
rect 20240 7251 20431 7273
rect 20732 7267 20841 7287
rect 20861 7267 20870 7287
rect 20732 7260 20870 7267
rect 20928 7287 21076 7296
rect 20928 7267 20937 7287
rect 20957 7267 21047 7287
rect 21067 7267 21076 7287
rect 20732 7258 20828 7260
rect 20928 7257 21076 7267
rect 21135 7287 21172 7297
rect 21135 7267 21143 7287
rect 21163 7267 21172 7287
rect 20984 7256 21020 7257
rect 20395 7249 20431 7251
rect 20395 7220 20432 7249
rect 19837 7211 19872 7212
rect 19814 7206 19872 7211
rect 19814 7186 19817 7206
rect 19837 7192 19872 7206
rect 19892 7192 19901 7212
rect 19837 7184 19901 7192
rect 19863 7183 19901 7184
rect 19864 7182 19901 7183
rect 19967 7216 20003 7217
rect 20075 7216 20111 7217
rect 19967 7208 20111 7216
rect 19967 7188 19975 7208
rect 19995 7206 20083 7208
rect 19995 7188 20028 7206
rect 19967 7184 20028 7188
rect 20051 7188 20083 7206
rect 20103 7188 20111 7208
rect 20051 7184 20111 7188
rect 19967 7182 20111 7184
rect 20177 7212 20215 7220
rect 20293 7216 20329 7217
rect 20177 7192 20186 7212
rect 20206 7192 20215 7212
rect 20177 7183 20215 7192
rect 20244 7208 20329 7216
rect 20244 7188 20301 7208
rect 20321 7188 20329 7208
rect 20177 7182 20214 7183
rect 20244 7182 20329 7188
rect 20395 7212 20433 7220
rect 20395 7192 20404 7212
rect 20424 7192 20433 7212
rect 21135 7200 21172 7267
rect 21207 7296 21238 7347
rect 21520 7335 21538 7353
rect 21556 7335 21572 7353
rect 21257 7296 21294 7297
rect 21207 7287 21294 7296
rect 21207 7267 21265 7287
rect 21285 7267 21294 7287
rect 21207 7257 21294 7267
rect 21353 7287 21390 7297
rect 21353 7267 21361 7287
rect 21381 7267 21390 7287
rect 21207 7256 21238 7257
rect 20832 7197 20869 7198
rect 21135 7197 21174 7200
rect 20831 7196 21174 7197
rect 21353 7196 21390 7267
rect 20395 7183 20433 7192
rect 20756 7191 21174 7196
rect 20395 7182 20432 7183
rect 19856 7154 19946 7160
rect 19856 7134 19872 7154
rect 19892 7152 19946 7154
rect 19892 7134 19917 7152
rect 19856 7132 19917 7134
rect 19937 7132 19946 7152
rect 19856 7126 19946 7132
rect 19869 7072 19906 7073
rect 19965 7072 20002 7073
rect 20021 7072 20057 7182
rect 20244 7161 20275 7182
rect 20756 7171 20759 7191
rect 20779 7171 21174 7191
rect 21203 7172 21390 7196
rect 20240 7160 20275 7161
rect 20118 7150 20275 7160
rect 20118 7130 20135 7150
rect 20155 7130 20275 7150
rect 20118 7123 20275 7130
rect 20342 7153 20491 7161
rect 20342 7133 20353 7153
rect 20373 7133 20412 7153
rect 20432 7133 20491 7153
rect 20342 7126 20491 7133
rect 21135 7146 21174 7171
rect 21520 7146 21572 7335
rect 21964 7363 21974 7381
rect 21992 7363 22004 7381
rect 22136 7379 22145 7399
rect 22165 7379 22174 7399
rect 22136 7371 22174 7379
rect 22240 7403 22325 7409
rect 22355 7408 22392 7409
rect 22240 7383 22248 7403
rect 22268 7383 22325 7403
rect 22240 7375 22325 7383
rect 22354 7399 22392 7408
rect 22354 7379 22363 7399
rect 22383 7379 22392 7399
rect 22240 7374 22276 7375
rect 22354 7371 22392 7379
rect 22458 7403 22602 7409
rect 22458 7383 22466 7403
rect 22486 7383 22519 7403
rect 22539 7383 22574 7403
rect 22594 7383 22602 7403
rect 22458 7375 22602 7383
rect 22458 7374 22494 7375
rect 22566 7374 22602 7375
rect 22668 7408 22705 7409
rect 22668 7407 22706 7408
rect 22668 7399 22732 7407
rect 22668 7379 22677 7399
rect 22697 7385 22732 7399
rect 22752 7385 22755 7405
rect 22697 7380 22755 7385
rect 22697 7379 22732 7380
rect 21964 7307 22004 7363
rect 22137 7342 22174 7371
rect 22138 7340 22174 7342
rect 22138 7318 22329 7340
rect 22355 7339 22392 7371
rect 22668 7367 22732 7379
rect 22772 7341 22799 7519
rect 23657 7494 23699 7539
rect 22631 7339 22799 7341
rect 22355 7329 22799 7339
rect 22940 7435 23127 7459
rect 23158 7440 23551 7460
rect 23571 7440 23574 7460
rect 23158 7435 23574 7440
rect 22940 7364 22977 7435
rect 23158 7434 23499 7435
rect 23092 7374 23123 7375
rect 22940 7344 22949 7364
rect 22969 7344 22977 7364
rect 22940 7334 22977 7344
rect 23036 7364 23123 7374
rect 23036 7344 23045 7364
rect 23065 7344 23123 7364
rect 23036 7335 23123 7344
rect 23036 7334 23073 7335
rect 21961 7302 22004 7307
rect 22352 7313 22799 7329
rect 22352 7307 22380 7313
rect 22631 7312 22799 7313
rect 21961 7299 22111 7302
rect 22352 7299 22379 7307
rect 21961 7297 22379 7299
rect 21961 7279 21970 7297
rect 21988 7279 22379 7297
rect 23092 7284 23123 7335
rect 23158 7364 23195 7434
rect 23461 7433 23498 7434
rect 23310 7374 23346 7375
rect 23158 7344 23167 7364
rect 23187 7344 23195 7364
rect 23158 7334 23195 7344
rect 23254 7364 23402 7374
rect 23502 7371 23598 7373
rect 23254 7344 23263 7364
rect 23283 7344 23373 7364
rect 23393 7344 23402 7364
rect 23254 7335 23402 7344
rect 23460 7364 23598 7371
rect 23460 7344 23469 7364
rect 23489 7344 23598 7364
rect 23460 7335 23598 7344
rect 23254 7334 23291 7335
rect 22984 7281 23025 7282
rect 21961 7276 22379 7279
rect 21961 7270 22004 7276
rect 21964 7267 22004 7270
rect 22879 7274 23025 7281
rect 22361 7258 22401 7259
rect 22072 7241 22401 7258
rect 22879 7254 22935 7274
rect 22955 7254 22994 7274
rect 23014 7254 23025 7274
rect 22879 7246 23025 7254
rect 23092 7277 23249 7284
rect 23092 7257 23212 7277
rect 23232 7257 23249 7277
rect 23092 7247 23249 7257
rect 23092 7246 23127 7247
rect 21956 7198 21999 7209
rect 21956 7180 21968 7198
rect 21986 7180 21999 7198
rect 21956 7154 21999 7180
rect 22072 7154 22099 7241
rect 22361 7232 22401 7241
rect 21135 7128 21574 7146
rect 20342 7125 20383 7126
rect 20076 7072 20113 7073
rect 19769 7063 19907 7072
rect 19769 7043 19878 7063
rect 19898 7043 19907 7063
rect 19769 7036 19907 7043
rect 19965 7063 20113 7072
rect 19965 7043 19974 7063
rect 19994 7043 20084 7063
rect 20104 7043 20113 7063
rect 19769 7034 19865 7036
rect 19965 7033 20113 7043
rect 20172 7063 20209 7073
rect 20172 7043 20180 7063
rect 20200 7043 20209 7063
rect 20021 7032 20057 7033
rect 19869 6973 19906 6974
rect 20172 6973 20209 7043
rect 20244 7072 20275 7123
rect 21135 7110 21535 7128
rect 21553 7110 21574 7128
rect 21135 7104 21574 7110
rect 21141 7100 21574 7104
rect 21956 7133 22099 7154
rect 22143 7206 22177 7222
rect 22361 7212 22754 7232
rect 22774 7212 22777 7232
rect 23092 7225 23123 7246
rect 23310 7225 23346 7335
rect 23365 7334 23402 7335
rect 23461 7334 23498 7335
rect 23421 7275 23511 7281
rect 23421 7255 23430 7275
rect 23450 7273 23511 7275
rect 23450 7255 23475 7273
rect 23421 7253 23475 7255
rect 23495 7253 23511 7273
rect 23421 7247 23511 7253
rect 22935 7224 22972 7225
rect 22361 7207 22777 7212
rect 22934 7215 22972 7224
rect 22361 7206 22702 7207
rect 22143 7136 22180 7206
rect 22295 7146 22326 7147
rect 21956 7131 22093 7133
rect 21520 7098 21572 7100
rect 21956 7089 21999 7131
rect 22143 7116 22152 7136
rect 22172 7116 22180 7136
rect 22143 7106 22180 7116
rect 22239 7136 22326 7146
rect 22239 7116 22248 7136
rect 22268 7116 22326 7136
rect 22239 7107 22326 7116
rect 22239 7106 22276 7107
rect 21954 7079 21999 7089
rect 20294 7072 20331 7073
rect 20244 7063 20331 7072
rect 20244 7043 20302 7063
rect 20322 7043 20331 7063
rect 20244 7033 20331 7043
rect 20390 7063 20427 7073
rect 20390 7043 20398 7063
rect 20418 7043 20427 7063
rect 21954 7061 21963 7079
rect 21981 7061 21999 7079
rect 21954 7055 21999 7061
rect 22295 7056 22326 7107
rect 22361 7136 22398 7206
rect 22664 7205 22701 7206
rect 22934 7195 22943 7215
rect 22963 7195 22972 7215
rect 22934 7187 22972 7195
rect 23038 7219 23123 7225
rect 23153 7224 23190 7225
rect 23038 7199 23046 7219
rect 23066 7199 23123 7219
rect 23038 7191 23123 7199
rect 23152 7215 23190 7224
rect 23152 7195 23161 7215
rect 23181 7195 23190 7215
rect 23038 7190 23074 7191
rect 23152 7187 23190 7195
rect 23256 7219 23400 7225
rect 23256 7199 23264 7219
rect 23284 7216 23372 7219
rect 23284 7199 23319 7216
rect 23256 7198 23319 7199
rect 23338 7199 23372 7216
rect 23392 7199 23400 7219
rect 23338 7198 23400 7199
rect 23256 7191 23400 7198
rect 23256 7190 23292 7191
rect 23364 7190 23400 7191
rect 23466 7224 23503 7225
rect 23466 7223 23504 7224
rect 23526 7223 23553 7227
rect 23466 7221 23553 7223
rect 23466 7215 23530 7221
rect 23466 7195 23475 7215
rect 23495 7201 23530 7215
rect 23550 7201 23553 7221
rect 23495 7196 23553 7201
rect 23495 7195 23530 7196
rect 22935 7158 22972 7187
rect 22936 7156 22972 7158
rect 22513 7146 22549 7147
rect 22361 7116 22370 7136
rect 22390 7116 22398 7136
rect 22361 7106 22398 7116
rect 22457 7136 22605 7146
rect 22705 7143 22801 7145
rect 22457 7116 22466 7136
rect 22486 7116 22576 7136
rect 22596 7116 22605 7136
rect 22457 7107 22605 7116
rect 22663 7136 22801 7143
rect 22663 7116 22672 7136
rect 22692 7116 22801 7136
rect 22936 7134 23127 7156
rect 23153 7155 23190 7187
rect 23466 7183 23530 7195
rect 23570 7157 23597 7335
rect 23429 7155 23597 7157
rect 23153 7129 23597 7155
rect 22663 7107 22801 7116
rect 22457 7106 22494 7107
rect 21954 7052 21991 7055
rect 22187 7053 22228 7054
rect 20244 7032 20275 7033
rect 19868 6972 20209 6973
rect 20390 6972 20427 7043
rect 22079 7046 22228 7053
rect 21523 7033 21560 7038
rect 19793 6967 20209 6972
rect 19793 6947 19796 6967
rect 19816 6947 20209 6967
rect 20240 6948 20427 6972
rect 21514 7029 21561 7033
rect 21514 7011 21533 7029
rect 21551 7011 21561 7029
rect 22079 7026 22138 7046
rect 22158 7026 22197 7046
rect 22217 7026 22228 7046
rect 22079 7018 22228 7026
rect 22295 7049 22452 7056
rect 22295 7029 22415 7049
rect 22435 7029 22452 7049
rect 22295 7019 22452 7029
rect 22295 7018 22330 7019
rect 21514 6963 21561 7011
rect 22295 6997 22326 7018
rect 22513 6997 22549 7107
rect 22568 7106 22605 7107
rect 22664 7106 22701 7107
rect 22624 7047 22714 7053
rect 22624 7027 22633 7047
rect 22653 7045 22714 7047
rect 22653 7027 22678 7045
rect 22624 7025 22678 7027
rect 22698 7025 22714 7045
rect 22624 7019 22714 7025
rect 22138 6996 22175 6997
rect 21138 6960 21561 6963
rect 20013 6946 20078 6947
rect 21116 6930 21561 6960
rect 21950 6988 21988 6990
rect 21950 6980 21993 6988
rect 21950 6962 21961 6980
rect 21979 6962 21993 6980
rect 21950 6935 21993 6962
rect 22137 6987 22175 6996
rect 22137 6967 22146 6987
rect 22166 6967 22175 6987
rect 22137 6959 22175 6967
rect 22241 6991 22326 6997
rect 22356 6996 22393 6997
rect 22241 6971 22249 6991
rect 22269 6971 22326 6991
rect 22241 6963 22326 6971
rect 22355 6987 22393 6996
rect 22355 6967 22364 6987
rect 22384 6967 22393 6987
rect 22241 6962 22277 6963
rect 22355 6959 22393 6967
rect 22459 6995 22603 6997
rect 22459 6991 22511 6995
rect 22459 6971 22467 6991
rect 22487 6975 22511 6991
rect 22531 6991 22603 6995
rect 22531 6975 22575 6991
rect 22487 6971 22575 6975
rect 22595 6971 22603 6991
rect 22459 6963 22603 6971
rect 22459 6962 22495 6963
rect 22567 6962 22603 6963
rect 22669 6996 22706 6997
rect 22669 6995 22707 6996
rect 22669 6987 22733 6995
rect 22669 6967 22678 6987
rect 22698 6973 22733 6987
rect 22753 6973 22756 6993
rect 22698 6968 22756 6973
rect 22698 6967 22733 6968
rect 20209 6914 20249 6922
rect 20209 6892 20217 6914
rect 20241 6892 20249 6914
rect 19814 6663 19851 6669
rect 19814 6644 19822 6663
rect 19843 6644 19851 6663
rect 19814 6636 19851 6644
rect 19818 6303 19851 6636
rect 19915 6668 20083 6669
rect 20209 6668 20249 6892
rect 20712 6896 20880 6897
rect 21116 6896 21157 6930
rect 21514 6909 21561 6930
rect 20712 6886 21157 6896
rect 21229 6894 21372 6895
rect 20712 6870 21156 6886
rect 20712 6868 20880 6870
rect 21076 6869 21156 6870
rect 21229 6869 21374 6894
rect 21516 6869 21561 6909
rect 20712 6690 20739 6868
rect 20779 6830 20843 6842
rect 21119 6838 21156 6869
rect 21337 6838 21374 6869
rect 21519 6862 21561 6869
rect 21951 6928 21993 6935
rect 22138 6928 22175 6959
rect 22356 6928 22393 6959
rect 22669 6955 22733 6967
rect 22773 6929 22800 7107
rect 21951 6888 21996 6928
rect 22138 6903 22283 6928
rect 22356 6927 22436 6928
rect 22632 6927 22800 6929
rect 22356 6911 22800 6927
rect 22140 6902 22283 6903
rect 22355 6901 22800 6911
rect 21951 6867 21998 6888
rect 22355 6867 22396 6901
rect 22632 6900 22800 6901
rect 23263 6905 23303 7129
rect 23429 7128 23597 7129
rect 23661 7161 23694 7494
rect 24299 7493 24326 7671
rect 24366 7633 24430 7645
rect 24706 7641 24743 7673
rect 24769 7672 24960 7694
rect 25095 7692 25204 7712
rect 25224 7692 25233 7712
rect 25095 7685 25233 7692
rect 25291 7712 25439 7721
rect 25291 7692 25300 7712
rect 25320 7692 25410 7712
rect 25430 7692 25439 7712
rect 25095 7683 25191 7685
rect 25291 7682 25439 7692
rect 25498 7712 25535 7722
rect 25498 7692 25506 7712
rect 25526 7692 25535 7712
rect 25347 7681 25383 7682
rect 24924 7670 24960 7672
rect 24924 7641 24961 7670
rect 24366 7632 24401 7633
rect 24343 7627 24401 7632
rect 24343 7607 24346 7627
rect 24366 7613 24401 7627
rect 24421 7613 24430 7633
rect 24366 7605 24430 7613
rect 24392 7604 24430 7605
rect 24393 7603 24430 7604
rect 24496 7637 24532 7638
rect 24604 7637 24640 7638
rect 24496 7629 24640 7637
rect 24496 7609 24504 7629
rect 24524 7628 24612 7629
rect 24524 7609 24559 7628
rect 24580 7609 24612 7628
rect 24632 7609 24640 7629
rect 24496 7603 24640 7609
rect 24706 7633 24744 7641
rect 24822 7637 24858 7638
rect 24706 7613 24715 7633
rect 24735 7613 24744 7633
rect 24706 7604 24744 7613
rect 24773 7629 24858 7637
rect 24773 7609 24830 7629
rect 24850 7609 24858 7629
rect 24706 7603 24743 7604
rect 24773 7603 24858 7609
rect 24924 7633 24962 7641
rect 24924 7613 24933 7633
rect 24953 7613 24962 7633
rect 25195 7622 25232 7623
rect 25498 7622 25535 7692
rect 25570 7721 25601 7772
rect 25897 7767 25942 7773
rect 25897 7749 25915 7767
rect 25933 7749 25942 7767
rect 27416 7766 27425 7786
rect 27445 7766 27453 7786
rect 27416 7756 27453 7766
rect 27512 7786 27599 7796
rect 27512 7766 27521 7786
rect 27541 7766 27599 7786
rect 27512 7757 27599 7766
rect 27512 7756 27549 7757
rect 25897 7739 25942 7749
rect 25620 7721 25657 7722
rect 25570 7712 25657 7721
rect 25570 7692 25628 7712
rect 25648 7692 25657 7712
rect 25570 7682 25657 7692
rect 25716 7712 25753 7722
rect 25716 7692 25724 7712
rect 25744 7692 25753 7712
rect 25897 7697 25940 7739
rect 26337 7727 26389 7729
rect 25803 7695 25940 7697
rect 25570 7681 25601 7682
rect 25716 7622 25753 7692
rect 25194 7621 25535 7622
rect 24924 7604 24962 7613
rect 25119 7616 25535 7621
rect 24924 7603 24961 7604
rect 24385 7575 24475 7581
rect 24385 7555 24401 7575
rect 24421 7573 24475 7575
rect 24421 7555 24446 7573
rect 24385 7553 24446 7555
rect 24466 7553 24475 7573
rect 24385 7547 24475 7553
rect 24398 7493 24435 7494
rect 24494 7493 24531 7494
rect 24550 7493 24586 7603
rect 24773 7582 24804 7603
rect 25119 7596 25122 7616
rect 25142 7596 25535 7616
rect 25719 7606 25753 7622
rect 25797 7674 25940 7695
rect 26335 7723 26768 7727
rect 26335 7717 26774 7723
rect 26335 7699 26356 7717
rect 26374 7699 26774 7717
rect 27568 7706 27599 7757
rect 27634 7786 27671 7856
rect 27937 7855 27974 7856
rect 27786 7796 27822 7797
rect 27634 7766 27643 7786
rect 27663 7766 27671 7786
rect 27634 7756 27671 7766
rect 27730 7786 27878 7796
rect 27978 7793 28074 7795
rect 27730 7766 27739 7786
rect 27759 7766 27849 7786
rect 27869 7766 27878 7786
rect 27730 7757 27878 7766
rect 27936 7786 28074 7793
rect 27936 7766 27945 7786
rect 27965 7766 28074 7786
rect 27936 7757 28074 7766
rect 27730 7756 27767 7757
rect 27460 7703 27501 7704
rect 26335 7681 26774 7699
rect 25495 7587 25535 7596
rect 25797 7587 25824 7674
rect 25897 7648 25940 7674
rect 25897 7630 25910 7648
rect 25928 7630 25940 7648
rect 25897 7619 25940 7630
rect 24769 7581 24804 7582
rect 24647 7571 24804 7581
rect 24647 7551 24664 7571
rect 24684 7551 24804 7571
rect 24647 7544 24804 7551
rect 24871 7574 25020 7582
rect 24871 7554 24882 7574
rect 24902 7554 24941 7574
rect 24961 7554 25020 7574
rect 25495 7570 25824 7587
rect 25495 7569 25535 7570
rect 24871 7547 25020 7554
rect 25892 7558 25932 7561
rect 25892 7552 25935 7558
rect 25517 7549 25935 7552
rect 24871 7546 24912 7547
rect 24605 7493 24642 7494
rect 24298 7484 24436 7493
rect 24161 7474 24197 7480
rect 24161 7456 24166 7474
rect 24188 7456 24197 7474
rect 24161 7452 24197 7456
rect 24298 7464 24407 7484
rect 24427 7464 24436 7484
rect 24298 7457 24436 7464
rect 24494 7484 24642 7493
rect 24494 7464 24503 7484
rect 24523 7464 24613 7484
rect 24633 7464 24642 7484
rect 24298 7455 24394 7457
rect 24494 7454 24642 7464
rect 24701 7484 24738 7494
rect 24701 7464 24709 7484
rect 24729 7464 24738 7484
rect 24550 7453 24586 7454
rect 24164 7293 24197 7452
rect 24398 7394 24435 7395
rect 24701 7394 24738 7464
rect 24773 7493 24804 7544
rect 25517 7531 25908 7549
rect 25926 7531 25935 7549
rect 25517 7529 25935 7531
rect 25517 7521 25544 7529
rect 25785 7526 25935 7529
rect 25097 7515 25265 7516
rect 25516 7515 25544 7521
rect 25097 7499 25544 7515
rect 25892 7521 25935 7526
rect 24823 7493 24860 7494
rect 24773 7484 24860 7493
rect 24773 7464 24831 7484
rect 24851 7464 24860 7484
rect 24773 7454 24860 7464
rect 24919 7484 24956 7494
rect 24919 7464 24927 7484
rect 24947 7464 24956 7484
rect 24773 7453 24804 7454
rect 24397 7393 24738 7394
rect 24919 7393 24956 7464
rect 24322 7388 24738 7393
rect 24322 7368 24325 7388
rect 24345 7368 24738 7388
rect 24769 7369 24956 7393
rect 25097 7489 25541 7499
rect 25097 7487 25265 7489
rect 25097 7309 25124 7487
rect 25164 7449 25228 7461
rect 25504 7457 25541 7489
rect 25567 7488 25758 7510
rect 25722 7486 25758 7488
rect 25722 7457 25759 7486
rect 25892 7465 25932 7521
rect 25164 7448 25199 7449
rect 25141 7443 25199 7448
rect 25141 7423 25144 7443
rect 25164 7429 25199 7443
rect 25219 7429 25228 7449
rect 25164 7421 25228 7429
rect 25190 7420 25228 7421
rect 25191 7419 25228 7420
rect 25294 7453 25330 7454
rect 25402 7453 25438 7454
rect 25294 7445 25438 7453
rect 25294 7425 25302 7445
rect 25322 7425 25357 7445
rect 25377 7425 25410 7445
rect 25430 7425 25438 7445
rect 25294 7419 25438 7425
rect 25504 7449 25542 7457
rect 25620 7453 25656 7454
rect 25504 7429 25513 7449
rect 25533 7429 25542 7449
rect 25504 7420 25542 7429
rect 25571 7445 25656 7453
rect 25571 7425 25628 7445
rect 25648 7425 25656 7445
rect 25504 7419 25541 7420
rect 25571 7419 25656 7425
rect 25722 7449 25760 7457
rect 25722 7429 25731 7449
rect 25751 7429 25760 7449
rect 25892 7447 25904 7465
rect 25922 7447 25932 7465
rect 26337 7492 26389 7681
rect 26735 7656 26774 7681
rect 27352 7696 27501 7703
rect 27352 7676 27411 7696
rect 27431 7676 27470 7696
rect 27490 7676 27501 7696
rect 27352 7668 27501 7676
rect 27568 7699 27725 7706
rect 27568 7679 27688 7699
rect 27708 7679 27725 7699
rect 27568 7669 27725 7679
rect 27568 7668 27603 7669
rect 26519 7631 26706 7655
rect 26735 7636 27130 7656
rect 27150 7636 27153 7656
rect 27568 7647 27599 7668
rect 27786 7647 27822 7757
rect 27841 7756 27878 7757
rect 27937 7756 27974 7757
rect 27897 7697 27987 7703
rect 27897 7677 27906 7697
rect 27926 7695 27987 7697
rect 27926 7677 27951 7695
rect 27897 7675 27951 7677
rect 27971 7675 27987 7695
rect 27897 7669 27987 7675
rect 27411 7646 27448 7647
rect 26735 7631 27153 7636
rect 27410 7637 27448 7646
rect 26519 7560 26556 7631
rect 26735 7630 27078 7631
rect 26735 7627 26774 7630
rect 27040 7629 27077 7630
rect 26671 7570 26702 7571
rect 26519 7540 26528 7560
rect 26548 7540 26556 7560
rect 26519 7530 26556 7540
rect 26615 7560 26702 7570
rect 26615 7540 26624 7560
rect 26644 7540 26702 7560
rect 26615 7531 26702 7540
rect 26615 7530 26652 7531
rect 26337 7474 26353 7492
rect 26371 7474 26389 7492
rect 26671 7480 26702 7531
rect 26737 7560 26774 7627
rect 27410 7617 27419 7637
rect 27439 7617 27448 7637
rect 27410 7609 27448 7617
rect 27514 7641 27599 7647
rect 27629 7646 27666 7647
rect 27514 7621 27522 7641
rect 27542 7621 27599 7641
rect 27514 7613 27599 7621
rect 27628 7637 27666 7646
rect 27628 7617 27637 7637
rect 27657 7617 27666 7637
rect 27514 7612 27550 7613
rect 27628 7609 27666 7617
rect 27732 7642 27876 7647
rect 27732 7641 27794 7642
rect 27732 7621 27740 7641
rect 27760 7623 27794 7641
rect 27815 7641 27876 7642
rect 27815 7623 27848 7641
rect 27760 7621 27848 7623
rect 27868 7621 27876 7641
rect 27732 7613 27876 7621
rect 27732 7612 27768 7613
rect 27840 7612 27876 7613
rect 27942 7646 27979 7647
rect 27942 7645 27980 7646
rect 27942 7637 28006 7645
rect 27942 7617 27951 7637
rect 27971 7623 28006 7637
rect 28026 7623 28029 7643
rect 27971 7618 28029 7623
rect 27971 7617 28006 7618
rect 27411 7580 27448 7609
rect 27412 7578 27448 7580
rect 26889 7570 26925 7571
rect 26737 7540 26746 7560
rect 26766 7540 26774 7560
rect 26737 7530 26774 7540
rect 26833 7560 26981 7570
rect 27081 7567 27177 7569
rect 26833 7540 26842 7560
rect 26862 7540 26952 7560
rect 26972 7540 26981 7560
rect 26833 7531 26981 7540
rect 27039 7560 27177 7567
rect 27039 7540 27048 7560
rect 27068 7540 27177 7560
rect 27412 7556 27603 7578
rect 27629 7577 27666 7609
rect 27942 7605 28006 7617
rect 28046 7579 28073 7757
rect 27905 7577 28073 7579
rect 27629 7563 28073 7577
rect 28676 7711 28844 7712
rect 28970 7711 29010 7935
rect 29473 7939 29641 7940
rect 29876 7939 29916 7972
rect 30272 7939 30319 7972
rect 30710 7971 30751 7996
rect 30896 7971 30933 8002
rect 31114 7971 31151 8002
rect 31427 7998 31491 8010
rect 31531 7972 31558 8150
rect 30710 7944 30759 7971
rect 30895 7945 30944 7971
rect 31113 7970 31194 7971
rect 31390 7970 31558 7972
rect 31113 7945 31558 7970
rect 31114 7944 31558 7945
rect 29473 7938 29917 7939
rect 29473 7913 29918 7938
rect 29473 7911 29641 7913
rect 29837 7912 29918 7913
rect 30087 7912 30136 7938
rect 30272 7912 30321 7939
rect 29473 7733 29500 7911
rect 29540 7873 29604 7885
rect 29880 7881 29917 7912
rect 30098 7881 30135 7912
rect 30280 7887 30321 7912
rect 30712 7911 30759 7944
rect 31115 7911 31155 7944
rect 31390 7943 31558 7944
rect 32021 7948 32061 8172
rect 32187 8171 32355 8172
rect 32958 8306 33402 8320
rect 32958 8304 33126 8306
rect 32958 8126 32985 8304
rect 33025 8266 33089 8278
rect 33365 8274 33402 8306
rect 33428 8305 33619 8327
rect 33854 8323 33963 8343
rect 33983 8323 33992 8343
rect 33854 8316 33992 8323
rect 34050 8343 34198 8352
rect 34050 8323 34059 8343
rect 34079 8323 34169 8343
rect 34189 8323 34198 8343
rect 33854 8314 33950 8316
rect 34050 8313 34198 8323
rect 34257 8343 34294 8353
rect 34257 8323 34265 8343
rect 34285 8323 34294 8343
rect 34106 8312 34142 8313
rect 33583 8303 33619 8305
rect 33583 8274 33620 8303
rect 33025 8265 33060 8266
rect 33002 8260 33060 8265
rect 33002 8240 33005 8260
rect 33025 8246 33060 8260
rect 33080 8246 33089 8266
rect 33025 8238 33089 8246
rect 33051 8237 33089 8238
rect 33052 8236 33089 8237
rect 33155 8270 33191 8271
rect 33263 8270 33299 8271
rect 33155 8264 33299 8270
rect 33155 8262 33216 8264
rect 33155 8242 33163 8262
rect 33183 8247 33216 8262
rect 33235 8262 33299 8264
rect 33235 8247 33271 8262
rect 33183 8242 33271 8247
rect 33291 8242 33299 8262
rect 33155 8236 33299 8242
rect 33365 8266 33403 8274
rect 33481 8270 33517 8271
rect 33365 8246 33374 8266
rect 33394 8246 33403 8266
rect 33365 8237 33403 8246
rect 33432 8262 33517 8270
rect 33432 8242 33489 8262
rect 33509 8242 33517 8262
rect 33365 8236 33402 8237
rect 33432 8236 33517 8242
rect 33583 8266 33621 8274
rect 33583 8246 33592 8266
rect 33612 8246 33621 8266
rect 34257 8256 34294 8323
rect 34329 8352 34360 8403
rect 34642 8391 34660 8409
rect 34678 8391 34694 8409
rect 34379 8352 34416 8353
rect 34329 8343 34416 8352
rect 34329 8323 34387 8343
rect 34407 8323 34416 8343
rect 34329 8313 34416 8323
rect 34475 8343 34512 8353
rect 34475 8323 34483 8343
rect 34503 8323 34512 8343
rect 34329 8312 34360 8313
rect 33954 8253 33991 8254
rect 34257 8253 34296 8256
rect 33953 8252 34296 8253
rect 34475 8252 34512 8323
rect 33583 8237 33621 8246
rect 33878 8247 34296 8252
rect 33583 8236 33620 8237
rect 33044 8208 33134 8214
rect 33044 8188 33060 8208
rect 33080 8206 33134 8208
rect 33080 8188 33105 8206
rect 33044 8186 33105 8188
rect 33125 8186 33134 8206
rect 33044 8180 33134 8186
rect 33057 8126 33094 8127
rect 33153 8126 33190 8127
rect 33209 8126 33245 8236
rect 33432 8215 33463 8236
rect 33878 8227 33881 8247
rect 33901 8227 34296 8247
rect 34325 8228 34512 8252
rect 33428 8214 33463 8215
rect 33306 8204 33463 8214
rect 33306 8184 33323 8204
rect 33343 8184 33463 8204
rect 33306 8177 33463 8184
rect 33530 8207 33679 8215
rect 33530 8187 33541 8207
rect 33561 8187 33600 8207
rect 33620 8187 33679 8207
rect 33530 8180 33679 8187
rect 34257 8202 34296 8227
rect 34642 8202 34694 8391
rect 34257 8184 34696 8202
rect 33530 8179 33571 8180
rect 33264 8126 33301 8127
rect 32957 8117 33095 8126
rect 32957 8097 33066 8117
rect 33086 8097 33095 8117
rect 32957 8090 33095 8097
rect 33153 8117 33301 8126
rect 33153 8097 33162 8117
rect 33182 8097 33272 8117
rect 33292 8097 33301 8117
rect 32957 8088 33053 8090
rect 33153 8087 33301 8097
rect 33360 8117 33397 8127
rect 33360 8097 33368 8117
rect 33388 8097 33397 8117
rect 33209 8086 33245 8087
rect 33057 8027 33094 8028
rect 33360 8027 33397 8097
rect 33432 8126 33463 8177
rect 34257 8166 34657 8184
rect 34675 8166 34696 8184
rect 34257 8160 34696 8166
rect 34263 8156 34696 8160
rect 34642 8154 34694 8156
rect 33482 8126 33519 8127
rect 33432 8117 33519 8126
rect 33432 8097 33490 8117
rect 33510 8097 33519 8117
rect 33432 8087 33519 8097
rect 33578 8117 33615 8127
rect 33578 8097 33586 8117
rect 33606 8097 33615 8117
rect 33432 8086 33463 8087
rect 33056 8026 33397 8027
rect 33578 8026 33615 8097
rect 34645 8089 34682 8094
rect 34636 8085 34683 8089
rect 34636 8067 34655 8085
rect 34673 8067 34683 8085
rect 32981 8021 33397 8026
rect 32981 8001 32984 8021
rect 33004 8001 33397 8021
rect 33428 8002 33615 8026
rect 34240 8024 34280 8029
rect 34636 8024 34683 8067
rect 34240 7985 34683 8024
rect 32021 7926 32029 7948
rect 32053 7926 32061 7948
rect 32021 7918 32061 7926
rect 33334 7970 33374 7978
rect 33334 7948 33342 7970
rect 33366 7948 33374 7970
rect 29540 7872 29575 7873
rect 29517 7867 29575 7872
rect 29517 7847 29520 7867
rect 29540 7853 29575 7867
rect 29595 7853 29604 7873
rect 29540 7845 29604 7853
rect 29566 7844 29604 7845
rect 29567 7843 29604 7844
rect 29670 7877 29706 7878
rect 29778 7877 29814 7878
rect 29670 7869 29814 7877
rect 29670 7849 29678 7869
rect 29698 7865 29786 7869
rect 29698 7849 29742 7865
rect 29670 7845 29742 7849
rect 29762 7849 29786 7865
rect 29806 7849 29814 7869
rect 29762 7845 29814 7849
rect 29670 7843 29814 7845
rect 29880 7873 29918 7881
rect 29996 7877 30032 7878
rect 29880 7853 29889 7873
rect 29909 7853 29918 7873
rect 29880 7844 29918 7853
rect 29947 7869 30032 7877
rect 29947 7849 30004 7869
rect 30024 7849 30032 7869
rect 29880 7843 29917 7844
rect 29947 7843 30032 7849
rect 30098 7873 30136 7881
rect 30098 7853 30107 7873
rect 30127 7853 30136 7873
rect 30098 7844 30136 7853
rect 30280 7878 30322 7887
rect 30280 7860 30294 7878
rect 30312 7860 30322 7878
rect 30280 7852 30322 7860
rect 30285 7850 30322 7852
rect 30712 7872 31155 7911
rect 30098 7843 30135 7844
rect 29559 7815 29649 7821
rect 29559 7795 29575 7815
rect 29595 7813 29649 7815
rect 29595 7795 29620 7813
rect 29559 7793 29620 7795
rect 29640 7793 29649 7813
rect 29559 7787 29649 7793
rect 29572 7733 29609 7734
rect 29668 7733 29705 7734
rect 29724 7733 29760 7843
rect 29947 7822 29978 7843
rect 30712 7829 30759 7872
rect 31115 7867 31155 7872
rect 31780 7870 31967 7894
rect 31998 7875 32391 7895
rect 32411 7875 32414 7895
rect 31998 7870 32414 7875
rect 29943 7821 29978 7822
rect 29821 7811 29978 7821
rect 29821 7791 29838 7811
rect 29858 7791 29978 7811
rect 29821 7784 29978 7791
rect 30045 7814 30194 7822
rect 30045 7794 30056 7814
rect 30076 7794 30115 7814
rect 30135 7794 30194 7814
rect 30712 7811 30722 7829
rect 30740 7811 30759 7829
rect 30712 7807 30759 7811
rect 30713 7802 30750 7807
rect 30045 7787 30194 7794
rect 31780 7799 31817 7870
rect 31998 7869 32339 7870
rect 31932 7809 31963 7810
rect 30045 7786 30086 7787
rect 30282 7785 30319 7788
rect 29779 7733 29816 7734
rect 29472 7724 29610 7733
rect 28676 7685 29120 7711
rect 28676 7683 28844 7685
rect 27629 7551 28076 7563
rect 27672 7549 27705 7551
rect 27039 7531 27177 7540
rect 26833 7530 26870 7531
rect 26563 7477 26604 7478
rect 26337 7456 26389 7474
rect 26455 7470 26604 7477
rect 25892 7437 25932 7447
rect 26455 7450 26514 7470
rect 26534 7450 26573 7470
rect 26593 7450 26604 7470
rect 26455 7442 26604 7450
rect 26671 7473 26828 7480
rect 26671 7453 26791 7473
rect 26811 7453 26828 7473
rect 26671 7443 26828 7453
rect 26671 7442 26706 7443
rect 25722 7420 25760 7429
rect 26671 7421 26702 7442
rect 26889 7421 26925 7531
rect 26944 7530 26981 7531
rect 27040 7530 27077 7531
rect 27000 7471 27090 7477
rect 27000 7451 27009 7471
rect 27029 7469 27090 7471
rect 27029 7451 27054 7469
rect 27000 7449 27054 7451
rect 27074 7449 27090 7469
rect 27000 7443 27090 7449
rect 26514 7420 26551 7421
rect 25722 7419 25759 7420
rect 25183 7391 25273 7397
rect 25183 7371 25199 7391
rect 25219 7389 25273 7391
rect 25219 7371 25244 7389
rect 25183 7369 25244 7371
rect 25264 7369 25273 7389
rect 25183 7363 25273 7369
rect 25196 7309 25233 7310
rect 25292 7309 25329 7310
rect 25348 7309 25384 7419
rect 25571 7398 25602 7419
rect 26513 7411 26551 7420
rect 25567 7397 25602 7398
rect 25445 7387 25602 7397
rect 25445 7367 25462 7387
rect 25482 7367 25602 7387
rect 25445 7360 25602 7367
rect 25669 7390 25818 7398
rect 25669 7370 25680 7390
rect 25700 7370 25739 7390
rect 25759 7370 25818 7390
rect 26341 7393 26381 7403
rect 25669 7363 25818 7370
rect 25884 7366 25936 7384
rect 25669 7362 25710 7363
rect 25403 7309 25440 7310
rect 25096 7300 25234 7309
rect 24163 7292 24200 7293
rect 24134 7291 24302 7292
rect 24428 7291 24468 7293
rect 23959 7282 23998 7288
rect 23959 7260 23967 7282
rect 23991 7260 23998 7282
rect 23661 7153 23698 7161
rect 23661 7134 23669 7153
rect 23690 7134 23698 7153
rect 23661 7128 23698 7134
rect 23263 6883 23271 6905
rect 23295 6883 23303 6905
rect 23263 6875 23303 6883
rect 20779 6829 20814 6830
rect 20756 6824 20814 6829
rect 20756 6804 20759 6824
rect 20779 6810 20814 6824
rect 20834 6810 20843 6830
rect 20779 6802 20843 6810
rect 20805 6801 20843 6802
rect 20806 6800 20843 6801
rect 20909 6834 20945 6835
rect 21017 6834 21053 6835
rect 20909 6826 21053 6834
rect 20909 6806 20917 6826
rect 20937 6822 21025 6826
rect 20937 6806 20981 6822
rect 20909 6802 20981 6806
rect 21001 6806 21025 6822
rect 21045 6806 21053 6826
rect 21001 6802 21053 6806
rect 20909 6800 21053 6802
rect 21119 6830 21157 6838
rect 21235 6834 21271 6835
rect 21119 6810 21128 6830
rect 21148 6810 21157 6830
rect 21119 6801 21157 6810
rect 21186 6826 21271 6834
rect 21186 6806 21243 6826
rect 21263 6806 21271 6826
rect 21119 6800 21156 6801
rect 21186 6800 21271 6806
rect 21337 6830 21375 6838
rect 21337 6810 21346 6830
rect 21366 6810 21375 6830
rect 21337 6801 21375 6810
rect 21519 6835 21562 6862
rect 21519 6817 21533 6835
rect 21551 6817 21562 6835
rect 21519 6809 21562 6817
rect 21524 6807 21562 6809
rect 21951 6837 22396 6867
rect 23434 6850 23499 6851
rect 21951 6834 22374 6837
rect 21337 6800 21374 6801
rect 20798 6772 20888 6778
rect 20798 6752 20814 6772
rect 20834 6770 20888 6772
rect 20834 6752 20859 6770
rect 20798 6750 20859 6752
rect 20879 6750 20888 6770
rect 20798 6744 20888 6750
rect 20811 6690 20848 6691
rect 20907 6690 20944 6691
rect 20963 6690 20999 6800
rect 21186 6779 21217 6800
rect 21951 6786 21998 6834
rect 21182 6778 21217 6779
rect 21060 6768 21217 6778
rect 21060 6748 21077 6768
rect 21097 6748 21217 6768
rect 21060 6741 21217 6748
rect 21284 6771 21433 6779
rect 21284 6751 21295 6771
rect 21315 6751 21354 6771
rect 21374 6751 21433 6771
rect 21951 6768 21961 6786
rect 21979 6768 21998 6786
rect 21951 6764 21998 6768
rect 23085 6825 23272 6849
rect 23303 6830 23696 6850
rect 23716 6830 23719 6850
rect 23303 6825 23719 6830
rect 21952 6759 21989 6764
rect 21284 6744 21433 6751
rect 23085 6754 23122 6825
rect 23303 6824 23644 6825
rect 23237 6764 23268 6765
rect 21284 6743 21325 6744
rect 21521 6742 21558 6745
rect 21018 6690 21055 6691
rect 20711 6681 20849 6690
rect 19915 6642 20359 6668
rect 19915 6640 20083 6642
rect 19915 6462 19942 6640
rect 19982 6602 20046 6614
rect 20322 6610 20359 6642
rect 20385 6641 20576 6663
rect 20711 6661 20820 6681
rect 20840 6661 20849 6681
rect 20711 6654 20849 6661
rect 20907 6681 21055 6690
rect 20907 6661 20916 6681
rect 20936 6661 21026 6681
rect 21046 6661 21055 6681
rect 20711 6652 20807 6654
rect 20907 6651 21055 6661
rect 21114 6681 21151 6691
rect 21114 6661 21122 6681
rect 21142 6661 21151 6681
rect 20963 6650 20999 6651
rect 20540 6639 20576 6641
rect 20540 6610 20577 6639
rect 19982 6601 20017 6602
rect 19959 6596 20017 6601
rect 19959 6576 19962 6596
rect 19982 6582 20017 6596
rect 20037 6582 20046 6602
rect 19982 6576 20046 6582
rect 19959 6574 20046 6576
rect 19959 6570 19986 6574
rect 20008 6573 20046 6574
rect 20009 6572 20046 6573
rect 20112 6606 20148 6607
rect 20220 6606 20256 6607
rect 20112 6599 20256 6606
rect 20112 6598 20174 6599
rect 20112 6578 20120 6598
rect 20140 6581 20174 6598
rect 20193 6598 20256 6599
rect 20193 6581 20228 6598
rect 20140 6578 20228 6581
rect 20248 6578 20256 6598
rect 20112 6572 20256 6578
rect 20322 6602 20360 6610
rect 20438 6606 20474 6607
rect 20322 6582 20331 6602
rect 20351 6582 20360 6602
rect 20322 6573 20360 6582
rect 20389 6598 20474 6606
rect 20389 6578 20446 6598
rect 20466 6578 20474 6598
rect 20322 6572 20359 6573
rect 20389 6572 20474 6578
rect 20540 6602 20578 6610
rect 20540 6582 20549 6602
rect 20569 6582 20578 6602
rect 20811 6591 20848 6592
rect 21114 6591 21151 6661
rect 21186 6690 21217 6741
rect 21513 6736 21558 6742
rect 21513 6718 21531 6736
rect 21549 6718 21558 6736
rect 23085 6734 23094 6754
rect 23114 6734 23122 6754
rect 23085 6724 23122 6734
rect 23181 6754 23268 6764
rect 23181 6734 23190 6754
rect 23210 6734 23268 6754
rect 23181 6725 23268 6734
rect 23181 6724 23218 6725
rect 21513 6708 21558 6718
rect 21236 6690 21273 6691
rect 21186 6681 21273 6690
rect 21186 6661 21244 6681
rect 21264 6661 21273 6681
rect 21186 6651 21273 6661
rect 21332 6681 21369 6691
rect 21332 6661 21340 6681
rect 21360 6661 21369 6681
rect 21513 6666 21556 6708
rect 21940 6697 21992 6699
rect 21419 6664 21556 6666
rect 21186 6650 21217 6651
rect 21332 6591 21369 6661
rect 20810 6590 21151 6591
rect 20540 6573 20578 6582
rect 20735 6585 21151 6590
rect 20540 6572 20577 6573
rect 20001 6544 20091 6550
rect 20001 6524 20017 6544
rect 20037 6542 20091 6544
rect 20037 6524 20062 6542
rect 20001 6522 20062 6524
rect 20082 6522 20091 6542
rect 20001 6516 20091 6522
rect 20014 6462 20051 6463
rect 20110 6462 20147 6463
rect 20166 6462 20202 6572
rect 20389 6551 20420 6572
rect 20735 6565 20738 6585
rect 20758 6565 21151 6585
rect 21335 6575 21369 6591
rect 21413 6643 21556 6664
rect 21938 6693 22371 6697
rect 21938 6687 22377 6693
rect 21938 6669 21959 6687
rect 21977 6669 22377 6687
rect 23237 6674 23268 6725
rect 23303 6754 23340 6824
rect 23606 6823 23643 6824
rect 23455 6764 23491 6765
rect 23303 6734 23312 6754
rect 23332 6734 23340 6754
rect 23303 6724 23340 6734
rect 23399 6754 23547 6764
rect 23647 6761 23743 6763
rect 23399 6734 23408 6754
rect 23428 6734 23518 6754
rect 23538 6734 23547 6754
rect 23399 6725 23547 6734
rect 23605 6754 23743 6761
rect 23605 6734 23614 6754
rect 23634 6734 23743 6754
rect 23605 6725 23743 6734
rect 23399 6724 23436 6725
rect 23129 6671 23170 6672
rect 21938 6651 22377 6669
rect 21111 6556 21151 6565
rect 21413 6556 21440 6643
rect 21513 6617 21556 6643
rect 21513 6599 21526 6617
rect 21544 6599 21556 6617
rect 21513 6588 21556 6599
rect 20385 6550 20420 6551
rect 20263 6540 20420 6550
rect 20263 6520 20280 6540
rect 20300 6520 20420 6540
rect 20263 6513 20420 6520
rect 20487 6543 20633 6551
rect 20487 6523 20498 6543
rect 20518 6523 20557 6543
rect 20577 6523 20633 6543
rect 21111 6539 21440 6556
rect 21111 6538 21151 6539
rect 20487 6516 20633 6523
rect 21508 6527 21548 6530
rect 21508 6521 21551 6527
rect 21133 6518 21551 6521
rect 20487 6515 20528 6516
rect 20221 6462 20258 6463
rect 19914 6453 20052 6462
rect 19914 6433 20023 6453
rect 20043 6433 20052 6453
rect 19914 6426 20052 6433
rect 20110 6453 20258 6462
rect 20110 6433 20119 6453
rect 20139 6433 20229 6453
rect 20249 6433 20258 6453
rect 19914 6424 20010 6426
rect 20110 6423 20258 6433
rect 20317 6453 20354 6463
rect 20317 6433 20325 6453
rect 20345 6433 20354 6453
rect 20166 6422 20202 6423
rect 20014 6363 20051 6364
rect 20317 6363 20354 6433
rect 20389 6462 20420 6513
rect 21133 6500 21524 6518
rect 21542 6500 21551 6518
rect 21133 6498 21551 6500
rect 21133 6490 21160 6498
rect 21401 6495 21551 6498
rect 20713 6484 20881 6485
rect 21132 6484 21160 6490
rect 20713 6468 21160 6484
rect 21508 6490 21551 6495
rect 20439 6462 20476 6463
rect 20389 6453 20476 6462
rect 20389 6433 20447 6453
rect 20467 6433 20476 6453
rect 20389 6423 20476 6433
rect 20535 6453 20572 6463
rect 20535 6433 20543 6453
rect 20563 6433 20572 6453
rect 20389 6422 20420 6423
rect 20013 6362 20354 6363
rect 20535 6362 20572 6433
rect 19938 6357 20354 6362
rect 19938 6337 19941 6357
rect 19961 6337 20354 6357
rect 20385 6338 20572 6362
rect 20713 6458 21157 6468
rect 20713 6456 20881 6458
rect 19813 6258 19855 6303
rect 20713 6278 20740 6456
rect 20780 6418 20844 6430
rect 21120 6426 21157 6458
rect 21183 6457 21374 6479
rect 21338 6455 21374 6457
rect 21338 6426 21375 6455
rect 21508 6434 21548 6490
rect 20780 6417 20815 6418
rect 20757 6412 20815 6417
rect 20757 6392 20760 6412
rect 20780 6398 20815 6412
rect 20835 6398 20844 6418
rect 20780 6390 20844 6398
rect 20806 6389 20844 6390
rect 20807 6388 20844 6389
rect 20910 6422 20946 6423
rect 21018 6422 21054 6423
rect 20910 6414 21054 6422
rect 20910 6394 20918 6414
rect 20938 6394 20973 6414
rect 20993 6394 21026 6414
rect 21046 6394 21054 6414
rect 20910 6388 21054 6394
rect 21120 6418 21158 6426
rect 21236 6422 21272 6423
rect 21120 6398 21129 6418
rect 21149 6398 21158 6418
rect 21120 6389 21158 6398
rect 21187 6414 21272 6422
rect 21187 6394 21244 6414
rect 21264 6394 21272 6414
rect 21120 6388 21157 6389
rect 21187 6388 21272 6394
rect 21338 6418 21376 6426
rect 21338 6398 21347 6418
rect 21367 6398 21376 6418
rect 21508 6416 21520 6434
rect 21538 6416 21548 6434
rect 21940 6462 21992 6651
rect 22338 6626 22377 6651
rect 23021 6664 23170 6671
rect 23021 6644 23080 6664
rect 23100 6644 23139 6664
rect 23159 6644 23170 6664
rect 23021 6636 23170 6644
rect 23237 6667 23394 6674
rect 23237 6647 23357 6667
rect 23377 6647 23394 6667
rect 23237 6637 23394 6647
rect 23237 6636 23272 6637
rect 22122 6601 22309 6625
rect 22338 6606 22733 6626
rect 22753 6606 22756 6626
rect 23237 6615 23268 6636
rect 23455 6615 23491 6725
rect 23510 6724 23547 6725
rect 23606 6724 23643 6725
rect 23566 6665 23656 6671
rect 23566 6645 23575 6665
rect 23595 6663 23656 6665
rect 23595 6645 23620 6663
rect 23566 6643 23620 6645
rect 23640 6643 23656 6663
rect 23566 6637 23656 6643
rect 23080 6614 23117 6615
rect 22338 6601 22756 6606
rect 23079 6605 23117 6614
rect 22122 6530 22159 6601
rect 22338 6600 22681 6601
rect 22338 6597 22377 6600
rect 22643 6599 22680 6600
rect 22274 6540 22305 6541
rect 22122 6510 22131 6530
rect 22151 6510 22159 6530
rect 22122 6500 22159 6510
rect 22218 6530 22305 6540
rect 22218 6510 22227 6530
rect 22247 6510 22305 6530
rect 22218 6501 22305 6510
rect 22218 6500 22255 6501
rect 21940 6444 21956 6462
rect 21974 6444 21992 6462
rect 22274 6450 22305 6501
rect 22340 6530 22377 6597
rect 23079 6585 23088 6605
rect 23108 6585 23117 6605
rect 23079 6577 23117 6585
rect 23183 6609 23268 6615
rect 23298 6614 23335 6615
rect 23183 6589 23191 6609
rect 23211 6589 23268 6609
rect 23183 6581 23268 6589
rect 23297 6605 23335 6614
rect 23297 6585 23306 6605
rect 23326 6585 23335 6605
rect 23183 6580 23219 6581
rect 23297 6577 23335 6585
rect 23401 6609 23545 6615
rect 23401 6589 23409 6609
rect 23429 6608 23517 6609
rect 23429 6590 23464 6608
rect 23482 6590 23517 6608
rect 23429 6589 23517 6590
rect 23537 6589 23545 6609
rect 23401 6581 23545 6589
rect 23401 6580 23437 6581
rect 23509 6580 23545 6581
rect 23611 6614 23648 6615
rect 23611 6613 23649 6614
rect 23611 6605 23675 6613
rect 23611 6585 23620 6605
rect 23640 6591 23675 6605
rect 23695 6591 23698 6611
rect 23640 6586 23698 6591
rect 23640 6585 23675 6586
rect 23080 6548 23117 6577
rect 23081 6546 23117 6548
rect 22492 6540 22528 6541
rect 22340 6510 22349 6530
rect 22369 6510 22377 6530
rect 22340 6500 22377 6510
rect 22436 6530 22584 6540
rect 22684 6537 22780 6539
rect 22436 6510 22445 6530
rect 22465 6510 22555 6530
rect 22575 6510 22584 6530
rect 22436 6501 22584 6510
rect 22642 6530 22780 6537
rect 22642 6510 22651 6530
rect 22671 6510 22780 6530
rect 23081 6524 23272 6546
rect 23298 6545 23335 6577
rect 23611 6573 23675 6585
rect 23715 6549 23742 6725
rect 23661 6547 23742 6549
rect 23574 6545 23742 6547
rect 23298 6519 23742 6545
rect 23408 6517 23448 6519
rect 23574 6518 23742 6519
rect 22642 6501 22780 6510
rect 23683 6516 23742 6518
rect 22436 6500 22473 6501
rect 22166 6447 22207 6448
rect 21940 6426 21992 6444
rect 22058 6440 22207 6447
rect 21508 6406 21548 6416
rect 22058 6420 22117 6440
rect 22137 6420 22176 6440
rect 22196 6420 22207 6440
rect 22058 6412 22207 6420
rect 22274 6443 22431 6450
rect 22274 6423 22394 6443
rect 22414 6423 22431 6443
rect 22274 6413 22431 6423
rect 22274 6412 22309 6413
rect 21338 6389 21376 6398
rect 22274 6391 22305 6412
rect 22492 6391 22528 6501
rect 22547 6500 22584 6501
rect 22643 6500 22680 6501
rect 22603 6441 22693 6447
rect 22603 6421 22612 6441
rect 22632 6439 22693 6441
rect 22632 6421 22657 6439
rect 22603 6419 22657 6421
rect 22677 6419 22693 6439
rect 22603 6413 22693 6419
rect 22117 6390 22154 6391
rect 21338 6388 21375 6389
rect 20799 6360 20889 6366
rect 20799 6340 20815 6360
rect 20835 6358 20889 6360
rect 20835 6340 20860 6358
rect 20799 6338 20860 6340
rect 20880 6338 20889 6358
rect 20799 6332 20889 6338
rect 20812 6278 20849 6279
rect 20908 6278 20945 6279
rect 20964 6278 21000 6388
rect 21187 6367 21218 6388
rect 22116 6381 22154 6390
rect 21183 6366 21218 6367
rect 21061 6356 21218 6366
rect 21061 6336 21078 6356
rect 21098 6336 21218 6356
rect 21061 6329 21218 6336
rect 21285 6359 21434 6367
rect 21285 6339 21296 6359
rect 21316 6339 21355 6359
rect 21375 6339 21434 6359
rect 21944 6363 21984 6373
rect 21285 6332 21434 6339
rect 21500 6335 21552 6353
rect 21285 6331 21326 6332
rect 21019 6278 21056 6279
rect 20712 6269 20850 6278
rect 20184 6258 20217 6260
rect 19813 6246 20260 6258
rect 19816 6232 20260 6246
rect 19816 6230 19984 6232
rect 19816 6052 19843 6230
rect 19883 6192 19947 6204
rect 20223 6200 20260 6232
rect 20286 6231 20477 6253
rect 20712 6249 20821 6269
rect 20841 6249 20850 6269
rect 20712 6242 20850 6249
rect 20908 6269 21056 6278
rect 20908 6249 20917 6269
rect 20937 6249 21027 6269
rect 21047 6249 21056 6269
rect 20712 6240 20808 6242
rect 20908 6239 21056 6249
rect 21115 6269 21152 6279
rect 21115 6249 21123 6269
rect 21143 6249 21152 6269
rect 20964 6238 21000 6239
rect 20441 6229 20477 6231
rect 20441 6200 20478 6229
rect 19883 6191 19918 6192
rect 19860 6186 19918 6191
rect 19860 6166 19863 6186
rect 19883 6172 19918 6186
rect 19938 6172 19947 6192
rect 19883 6164 19947 6172
rect 19909 6163 19947 6164
rect 19910 6162 19947 6163
rect 20013 6196 20049 6197
rect 20121 6196 20157 6197
rect 20013 6188 20157 6196
rect 20013 6168 20021 6188
rect 20041 6186 20129 6188
rect 20041 6168 20074 6186
rect 20013 6167 20074 6168
rect 20095 6168 20129 6186
rect 20149 6168 20157 6188
rect 20095 6167 20157 6168
rect 20013 6162 20157 6167
rect 20223 6192 20261 6200
rect 20339 6196 20375 6197
rect 20223 6172 20232 6192
rect 20252 6172 20261 6192
rect 20223 6163 20261 6172
rect 20290 6188 20375 6196
rect 20290 6168 20347 6188
rect 20367 6168 20375 6188
rect 20223 6162 20260 6163
rect 20290 6162 20375 6168
rect 20441 6192 20479 6200
rect 20441 6172 20450 6192
rect 20470 6172 20479 6192
rect 21115 6182 21152 6249
rect 21187 6278 21218 6329
rect 21500 6317 21518 6335
rect 21536 6317 21552 6335
rect 21237 6278 21274 6279
rect 21187 6269 21274 6278
rect 21187 6249 21245 6269
rect 21265 6249 21274 6269
rect 21187 6239 21274 6249
rect 21333 6269 21370 6279
rect 21333 6249 21341 6269
rect 21361 6249 21370 6269
rect 21187 6238 21218 6239
rect 20812 6179 20849 6180
rect 21115 6179 21154 6182
rect 20811 6178 21154 6179
rect 21333 6178 21370 6249
rect 20441 6163 20479 6172
rect 20736 6173 21154 6178
rect 20441 6162 20478 6163
rect 19902 6134 19992 6140
rect 19902 6114 19918 6134
rect 19938 6132 19992 6134
rect 19938 6114 19963 6132
rect 19902 6112 19963 6114
rect 19983 6112 19992 6132
rect 19902 6106 19992 6112
rect 19915 6052 19952 6053
rect 20011 6052 20048 6053
rect 20067 6052 20103 6162
rect 20290 6141 20321 6162
rect 20736 6153 20739 6173
rect 20759 6153 21154 6173
rect 21183 6154 21370 6178
rect 20286 6140 20321 6141
rect 20164 6130 20321 6140
rect 20164 6110 20181 6130
rect 20201 6110 20321 6130
rect 20164 6103 20321 6110
rect 20388 6133 20537 6141
rect 20388 6113 20399 6133
rect 20419 6113 20458 6133
rect 20478 6113 20537 6133
rect 20388 6106 20537 6113
rect 21115 6128 21154 6153
rect 21500 6128 21552 6317
rect 21944 6345 21954 6363
rect 21972 6345 21984 6363
rect 22116 6361 22125 6381
rect 22145 6361 22154 6381
rect 22116 6353 22154 6361
rect 22220 6385 22305 6391
rect 22335 6390 22372 6391
rect 22220 6365 22228 6385
rect 22248 6365 22305 6385
rect 22220 6357 22305 6365
rect 22334 6381 22372 6390
rect 22334 6361 22343 6381
rect 22363 6361 22372 6381
rect 22220 6356 22256 6357
rect 22334 6353 22372 6361
rect 22438 6385 22582 6391
rect 22438 6365 22446 6385
rect 22466 6365 22499 6385
rect 22519 6365 22554 6385
rect 22574 6365 22582 6385
rect 22438 6357 22582 6365
rect 22438 6356 22474 6357
rect 22546 6356 22582 6357
rect 22648 6390 22685 6391
rect 22648 6389 22686 6390
rect 22648 6381 22712 6389
rect 22648 6361 22657 6381
rect 22677 6367 22712 6381
rect 22732 6367 22735 6387
rect 22677 6362 22735 6367
rect 22677 6361 22712 6362
rect 21944 6289 21984 6345
rect 22117 6324 22154 6353
rect 22118 6322 22154 6324
rect 22118 6300 22309 6322
rect 22335 6321 22372 6353
rect 22648 6349 22712 6361
rect 22752 6323 22779 6501
rect 23683 6498 23712 6516
rect 22611 6321 22779 6323
rect 22335 6311 22779 6321
rect 22920 6417 23107 6441
rect 23138 6422 23531 6442
rect 23551 6422 23554 6442
rect 23138 6417 23554 6422
rect 22920 6346 22957 6417
rect 23138 6416 23479 6417
rect 23072 6356 23103 6357
rect 22920 6326 22929 6346
rect 22949 6326 22957 6346
rect 22920 6316 22957 6326
rect 23016 6346 23103 6356
rect 23016 6326 23025 6346
rect 23045 6326 23103 6346
rect 23016 6317 23103 6326
rect 23016 6316 23053 6317
rect 21941 6284 21984 6289
rect 22332 6295 22779 6311
rect 22332 6289 22360 6295
rect 22611 6294 22779 6295
rect 21941 6281 22091 6284
rect 22332 6281 22359 6289
rect 21941 6279 22359 6281
rect 21941 6261 21950 6279
rect 21968 6261 22359 6279
rect 23072 6266 23103 6317
rect 23138 6346 23175 6416
rect 23441 6415 23478 6416
rect 23290 6356 23326 6357
rect 23138 6326 23147 6346
rect 23167 6326 23175 6346
rect 23138 6316 23175 6326
rect 23234 6346 23382 6356
rect 23482 6353 23578 6355
rect 23234 6326 23243 6346
rect 23263 6326 23353 6346
rect 23373 6326 23382 6346
rect 23234 6317 23382 6326
rect 23440 6346 23578 6353
rect 23440 6326 23449 6346
rect 23469 6326 23578 6346
rect 23440 6317 23578 6326
rect 23234 6316 23271 6317
rect 22964 6263 23005 6264
rect 21941 6258 22359 6261
rect 21941 6252 21984 6258
rect 21944 6249 21984 6252
rect 22856 6256 23005 6263
rect 22341 6240 22381 6241
rect 22052 6223 22381 6240
rect 22856 6236 22915 6256
rect 22935 6236 22974 6256
rect 22994 6236 23005 6256
rect 22856 6228 23005 6236
rect 23072 6259 23229 6266
rect 23072 6239 23192 6259
rect 23212 6239 23229 6259
rect 23072 6229 23229 6239
rect 23072 6228 23107 6229
rect 21936 6180 21979 6191
rect 21936 6162 21948 6180
rect 21966 6162 21979 6180
rect 21936 6136 21979 6162
rect 22052 6136 22079 6223
rect 22341 6214 22381 6223
rect 21115 6110 21554 6128
rect 20388 6105 20429 6106
rect 20122 6052 20159 6053
rect 19815 6043 19953 6052
rect 19815 6023 19924 6043
rect 19944 6023 19953 6043
rect 19815 6016 19953 6023
rect 20011 6043 20159 6052
rect 20011 6023 20020 6043
rect 20040 6023 20130 6043
rect 20150 6023 20159 6043
rect 19815 6014 19911 6016
rect 20011 6013 20159 6023
rect 20218 6043 20255 6053
rect 20218 6023 20226 6043
rect 20246 6023 20255 6043
rect 20067 6012 20103 6013
rect 19915 5953 19952 5954
rect 20218 5953 20255 6023
rect 20290 6052 20321 6103
rect 21115 6092 21515 6110
rect 21533 6092 21554 6110
rect 21115 6086 21554 6092
rect 21121 6082 21554 6086
rect 21936 6115 22079 6136
rect 22123 6188 22157 6204
rect 22341 6194 22734 6214
rect 22754 6194 22757 6214
rect 23072 6207 23103 6228
rect 23290 6207 23326 6317
rect 23345 6316 23382 6317
rect 23441 6316 23478 6317
rect 23401 6257 23491 6263
rect 23401 6237 23410 6257
rect 23430 6255 23491 6257
rect 23430 6237 23455 6255
rect 23401 6235 23455 6237
rect 23475 6235 23491 6255
rect 23401 6229 23491 6235
rect 22915 6206 22952 6207
rect 22341 6189 22757 6194
rect 22914 6197 22952 6206
rect 22341 6188 22682 6189
rect 22123 6118 22160 6188
rect 22275 6128 22306 6129
rect 21936 6113 22073 6115
rect 21500 6080 21552 6082
rect 21936 6071 21979 6113
rect 22123 6098 22132 6118
rect 22152 6098 22160 6118
rect 22123 6088 22160 6098
rect 22219 6118 22306 6128
rect 22219 6098 22228 6118
rect 22248 6098 22306 6118
rect 22219 6089 22306 6098
rect 22219 6088 22256 6089
rect 21934 6061 21979 6071
rect 20340 6052 20377 6053
rect 20290 6043 20377 6052
rect 20290 6023 20348 6043
rect 20368 6023 20377 6043
rect 20290 6013 20377 6023
rect 20436 6043 20473 6053
rect 20436 6023 20444 6043
rect 20464 6023 20473 6043
rect 21934 6043 21943 6061
rect 21961 6043 21979 6061
rect 21934 6037 21979 6043
rect 22275 6038 22306 6089
rect 22341 6118 22378 6188
rect 22644 6187 22681 6188
rect 22914 6177 22923 6197
rect 22943 6177 22952 6197
rect 22914 6169 22952 6177
rect 23018 6201 23103 6207
rect 23133 6206 23170 6207
rect 23018 6181 23026 6201
rect 23046 6181 23103 6201
rect 23018 6173 23103 6181
rect 23132 6197 23170 6206
rect 23132 6177 23141 6197
rect 23161 6177 23170 6197
rect 23018 6172 23054 6173
rect 23132 6169 23170 6177
rect 23236 6201 23380 6207
rect 23236 6181 23244 6201
rect 23264 6182 23296 6201
rect 23317 6182 23352 6201
rect 23264 6181 23352 6182
rect 23372 6181 23380 6201
rect 23236 6173 23380 6181
rect 23236 6172 23272 6173
rect 23344 6172 23380 6173
rect 23446 6206 23483 6207
rect 23446 6205 23484 6206
rect 23446 6197 23510 6205
rect 23446 6177 23455 6197
rect 23475 6183 23510 6197
rect 23530 6183 23533 6203
rect 23475 6178 23533 6183
rect 23475 6177 23510 6178
rect 22915 6140 22952 6169
rect 22916 6138 22952 6140
rect 22493 6128 22529 6129
rect 22341 6098 22350 6118
rect 22370 6098 22378 6118
rect 22341 6088 22378 6098
rect 22437 6118 22585 6128
rect 22685 6125 22781 6127
rect 22437 6098 22446 6118
rect 22466 6098 22556 6118
rect 22576 6098 22585 6118
rect 22437 6089 22585 6098
rect 22643 6118 22781 6125
rect 22643 6098 22652 6118
rect 22672 6098 22781 6118
rect 22916 6116 23107 6138
rect 23133 6137 23170 6169
rect 23446 6165 23510 6177
rect 23550 6139 23577 6317
rect 23409 6137 23577 6139
rect 23133 6111 23577 6137
rect 22643 6089 22781 6098
rect 22437 6088 22474 6089
rect 21934 6034 21971 6037
rect 22167 6035 22208 6036
rect 20290 6012 20321 6013
rect 19914 5952 20255 5953
rect 20436 5952 20473 6023
rect 22059 6028 22208 6035
rect 21503 6015 21540 6020
rect 21494 6011 21541 6015
rect 21494 5993 21513 6011
rect 21531 5993 21541 6011
rect 22059 6008 22118 6028
rect 22138 6008 22177 6028
rect 22197 6008 22208 6028
rect 22059 6000 22208 6008
rect 22275 6031 22432 6038
rect 22275 6011 22395 6031
rect 22415 6011 22432 6031
rect 22275 6001 22432 6011
rect 22275 6000 22310 6001
rect 19839 5947 20255 5952
rect 19839 5927 19842 5947
rect 19862 5927 20255 5947
rect 20286 5928 20473 5952
rect 21098 5950 21138 5955
rect 21494 5950 21541 5993
rect 22275 5979 22306 6000
rect 22493 5979 22529 6089
rect 22548 6088 22585 6089
rect 22644 6088 22681 6089
rect 22604 6029 22694 6035
rect 22604 6009 22613 6029
rect 22633 6027 22694 6029
rect 22633 6009 22658 6027
rect 22604 6007 22658 6009
rect 22678 6007 22694 6027
rect 22604 6001 22694 6007
rect 22118 5978 22155 5979
rect 21098 5911 21541 5950
rect 21931 5970 21968 5972
rect 21931 5962 21973 5970
rect 21931 5944 21941 5962
rect 21959 5944 21973 5962
rect 21931 5935 21973 5944
rect 22117 5969 22155 5978
rect 22117 5949 22126 5969
rect 22146 5949 22155 5969
rect 22117 5941 22155 5949
rect 22221 5973 22306 5979
rect 22336 5978 22373 5979
rect 22221 5953 22229 5973
rect 22249 5953 22306 5973
rect 22221 5945 22306 5953
rect 22335 5969 22373 5978
rect 22335 5949 22344 5969
rect 22364 5949 22373 5969
rect 22221 5944 22257 5945
rect 22335 5941 22373 5949
rect 22439 5977 22583 5979
rect 22439 5973 22491 5977
rect 22439 5953 22447 5973
rect 22467 5957 22491 5973
rect 22511 5973 22583 5977
rect 22511 5957 22555 5973
rect 22467 5953 22555 5957
rect 22575 5953 22583 5973
rect 22439 5945 22583 5953
rect 22439 5944 22475 5945
rect 22547 5944 22583 5945
rect 22649 5978 22686 5979
rect 22649 5977 22687 5978
rect 22649 5969 22713 5977
rect 22649 5949 22658 5969
rect 22678 5955 22713 5969
rect 22733 5955 22736 5975
rect 22678 5950 22736 5955
rect 22678 5949 22713 5950
rect 20192 5896 20232 5904
rect 20192 5874 20200 5896
rect 20224 5874 20232 5896
rect 19898 5650 20066 5651
rect 20192 5650 20232 5874
rect 20695 5878 20863 5879
rect 21098 5878 21138 5911
rect 21494 5878 21541 5911
rect 21932 5910 21973 5935
rect 22118 5910 22155 5941
rect 22336 5910 22373 5941
rect 22649 5937 22713 5949
rect 22753 5911 22780 6089
rect 21932 5883 21981 5910
rect 22117 5884 22166 5910
rect 22335 5909 22416 5910
rect 22612 5909 22780 5911
rect 22335 5884 22780 5909
rect 22336 5883 22780 5884
rect 20695 5877 21139 5878
rect 20695 5852 21140 5877
rect 20695 5850 20863 5852
rect 21059 5851 21140 5852
rect 21309 5851 21358 5877
rect 21494 5851 21543 5878
rect 20695 5672 20722 5850
rect 20762 5812 20826 5824
rect 21102 5820 21139 5851
rect 21320 5820 21357 5851
rect 21502 5826 21543 5851
rect 21934 5850 21981 5883
rect 22337 5850 22377 5883
rect 22612 5882 22780 5883
rect 23243 5887 23283 6111
rect 23409 6110 23577 6111
rect 23243 5865 23251 5887
rect 23275 5865 23283 5887
rect 23243 5857 23283 5865
rect 20762 5811 20797 5812
rect 20739 5806 20797 5811
rect 20739 5786 20742 5806
rect 20762 5792 20797 5806
rect 20817 5792 20826 5812
rect 20762 5784 20826 5792
rect 20788 5783 20826 5784
rect 20789 5782 20826 5783
rect 20892 5816 20928 5817
rect 21000 5816 21036 5817
rect 20892 5808 21036 5816
rect 20892 5788 20900 5808
rect 20920 5804 21008 5808
rect 20920 5788 20964 5804
rect 20892 5784 20964 5788
rect 20984 5788 21008 5804
rect 21028 5788 21036 5808
rect 20984 5784 21036 5788
rect 20892 5782 21036 5784
rect 21102 5812 21140 5820
rect 21218 5816 21254 5817
rect 21102 5792 21111 5812
rect 21131 5792 21140 5812
rect 21102 5783 21140 5792
rect 21169 5808 21254 5816
rect 21169 5788 21226 5808
rect 21246 5788 21254 5808
rect 21102 5782 21139 5783
rect 21169 5782 21254 5788
rect 21320 5812 21358 5820
rect 21320 5792 21329 5812
rect 21349 5792 21358 5812
rect 21320 5783 21358 5792
rect 21502 5817 21544 5826
rect 21502 5799 21516 5817
rect 21534 5799 21544 5817
rect 21502 5791 21544 5799
rect 21507 5789 21544 5791
rect 21934 5811 22377 5850
rect 21320 5782 21357 5783
rect 20781 5754 20871 5760
rect 20781 5734 20797 5754
rect 20817 5752 20871 5754
rect 20817 5734 20842 5752
rect 20781 5732 20842 5734
rect 20862 5732 20871 5752
rect 20781 5726 20871 5732
rect 20794 5672 20831 5673
rect 20890 5672 20927 5673
rect 20946 5672 20982 5782
rect 21169 5761 21200 5782
rect 21934 5768 21981 5811
rect 22337 5806 22377 5811
rect 23002 5809 23189 5833
rect 23220 5814 23613 5834
rect 23633 5814 23636 5834
rect 23220 5809 23636 5814
rect 21165 5760 21200 5761
rect 21043 5750 21200 5760
rect 21043 5730 21060 5750
rect 21080 5730 21200 5750
rect 21043 5723 21200 5730
rect 21267 5753 21416 5761
rect 21267 5733 21278 5753
rect 21298 5733 21337 5753
rect 21357 5733 21416 5753
rect 21934 5750 21944 5768
rect 21962 5750 21981 5768
rect 21934 5746 21981 5750
rect 21935 5741 21972 5746
rect 21267 5726 21416 5733
rect 23002 5738 23039 5809
rect 23220 5808 23561 5809
rect 23154 5748 23185 5749
rect 21267 5725 21308 5726
rect 21504 5724 21541 5727
rect 21001 5672 21038 5673
rect 20694 5663 20832 5672
rect 19898 5624 20342 5650
rect 19898 5622 20066 5624
rect 19898 5444 19925 5622
rect 19965 5584 20029 5596
rect 20305 5592 20342 5624
rect 20368 5623 20559 5645
rect 20694 5643 20803 5663
rect 20823 5643 20832 5663
rect 20694 5636 20832 5643
rect 20890 5663 21038 5672
rect 20890 5643 20899 5663
rect 20919 5643 21009 5663
rect 21029 5643 21038 5663
rect 20694 5634 20790 5636
rect 20890 5633 21038 5643
rect 21097 5663 21134 5673
rect 21097 5643 21105 5663
rect 21125 5643 21134 5663
rect 20946 5632 20982 5633
rect 20523 5621 20559 5623
rect 20523 5592 20560 5621
rect 19965 5583 20000 5584
rect 19942 5578 20000 5583
rect 19942 5558 19945 5578
rect 19965 5564 20000 5578
rect 20020 5564 20029 5584
rect 19965 5556 20029 5564
rect 19991 5555 20029 5556
rect 19992 5554 20029 5555
rect 20095 5588 20131 5589
rect 20203 5588 20239 5589
rect 20095 5580 20239 5588
rect 20095 5560 20103 5580
rect 20123 5579 20211 5580
rect 20123 5560 20158 5579
rect 20179 5560 20211 5579
rect 20231 5560 20239 5580
rect 20095 5554 20239 5560
rect 20305 5584 20343 5592
rect 20421 5588 20457 5589
rect 20305 5564 20314 5584
rect 20334 5564 20343 5584
rect 20305 5555 20343 5564
rect 20372 5580 20457 5588
rect 20372 5560 20429 5580
rect 20449 5560 20457 5580
rect 20305 5554 20342 5555
rect 20372 5554 20457 5560
rect 20523 5584 20561 5592
rect 20523 5564 20532 5584
rect 20552 5564 20561 5584
rect 20794 5573 20831 5574
rect 21097 5573 21134 5643
rect 21169 5672 21200 5723
rect 21496 5718 21541 5724
rect 21496 5700 21514 5718
rect 21532 5700 21541 5718
rect 23002 5718 23011 5738
rect 23031 5718 23039 5738
rect 23002 5708 23039 5718
rect 23098 5738 23185 5748
rect 23098 5718 23107 5738
rect 23127 5718 23185 5738
rect 23098 5709 23185 5718
rect 23098 5708 23135 5709
rect 21496 5690 21541 5700
rect 21219 5672 21256 5673
rect 21169 5663 21256 5672
rect 21169 5643 21227 5663
rect 21247 5643 21256 5663
rect 21169 5633 21256 5643
rect 21315 5663 21352 5673
rect 21315 5643 21323 5663
rect 21343 5643 21352 5663
rect 21496 5648 21539 5690
rect 21923 5679 21975 5681
rect 21402 5646 21539 5648
rect 21169 5632 21200 5633
rect 21315 5573 21352 5643
rect 20793 5572 21134 5573
rect 20523 5555 20561 5564
rect 20718 5567 21134 5572
rect 20523 5554 20560 5555
rect 19984 5526 20074 5532
rect 19984 5506 20000 5526
rect 20020 5524 20074 5526
rect 20020 5506 20045 5524
rect 19984 5504 20045 5506
rect 20065 5504 20074 5524
rect 19984 5498 20074 5504
rect 19997 5444 20034 5445
rect 20093 5444 20130 5445
rect 20149 5444 20185 5554
rect 20372 5533 20403 5554
rect 20718 5547 20721 5567
rect 20741 5547 21134 5567
rect 21318 5557 21352 5573
rect 21396 5625 21539 5646
rect 21921 5675 22354 5679
rect 21921 5669 22360 5675
rect 21921 5651 21942 5669
rect 21960 5651 22360 5669
rect 23154 5658 23185 5709
rect 23220 5738 23257 5808
rect 23523 5807 23560 5808
rect 23372 5748 23408 5749
rect 23220 5718 23229 5738
rect 23249 5718 23257 5738
rect 23220 5708 23257 5718
rect 23316 5738 23464 5748
rect 23564 5745 23660 5747
rect 23316 5718 23325 5738
rect 23345 5718 23435 5738
rect 23455 5718 23464 5738
rect 23316 5709 23464 5718
rect 23522 5738 23660 5745
rect 23522 5718 23531 5738
rect 23551 5718 23660 5738
rect 23522 5709 23660 5718
rect 23316 5708 23353 5709
rect 23046 5655 23087 5656
rect 21921 5633 22360 5651
rect 21094 5538 21134 5547
rect 21396 5538 21423 5625
rect 21496 5599 21539 5625
rect 21496 5581 21509 5599
rect 21527 5581 21539 5599
rect 21496 5570 21539 5581
rect 20368 5532 20403 5533
rect 20246 5522 20403 5532
rect 20246 5502 20263 5522
rect 20283 5502 20403 5522
rect 20246 5495 20403 5502
rect 20470 5525 20619 5533
rect 20470 5505 20481 5525
rect 20501 5505 20540 5525
rect 20560 5505 20619 5525
rect 21094 5521 21423 5538
rect 21094 5520 21134 5521
rect 20470 5498 20619 5505
rect 21491 5509 21531 5512
rect 21491 5503 21534 5509
rect 21116 5500 21534 5503
rect 20470 5497 20511 5498
rect 20204 5444 20241 5445
rect 19897 5435 20035 5444
rect 19595 5260 19635 5432
rect 19897 5415 20006 5435
rect 20026 5415 20035 5435
rect 19897 5408 20035 5415
rect 20093 5435 20241 5444
rect 20093 5415 20102 5435
rect 20122 5415 20212 5435
rect 20232 5415 20241 5435
rect 19897 5406 19993 5408
rect 20093 5405 20241 5415
rect 20300 5435 20337 5445
rect 20300 5415 20308 5435
rect 20328 5415 20337 5435
rect 20149 5404 20185 5405
rect 19997 5345 20034 5346
rect 20300 5345 20337 5415
rect 20372 5444 20403 5495
rect 21116 5482 21507 5500
rect 21525 5482 21534 5500
rect 21116 5480 21534 5482
rect 21116 5472 21143 5480
rect 21384 5477 21534 5480
rect 20696 5466 20864 5467
rect 21115 5466 21143 5472
rect 20696 5450 21143 5466
rect 21491 5472 21534 5477
rect 20422 5444 20459 5445
rect 20372 5435 20459 5444
rect 20372 5415 20430 5435
rect 20450 5415 20459 5435
rect 20372 5405 20459 5415
rect 20518 5435 20555 5445
rect 20518 5415 20526 5435
rect 20546 5415 20555 5435
rect 20372 5404 20403 5405
rect 19996 5344 20337 5345
rect 20518 5344 20555 5415
rect 19921 5339 20337 5344
rect 19921 5319 19924 5339
rect 19944 5319 20337 5339
rect 20368 5320 20555 5344
rect 20696 5440 21140 5450
rect 20696 5438 20864 5440
rect 20696 5260 20723 5438
rect 20763 5400 20827 5412
rect 21103 5408 21140 5440
rect 21166 5439 21357 5461
rect 21321 5437 21357 5439
rect 21321 5408 21358 5437
rect 21491 5416 21531 5472
rect 20763 5399 20798 5400
rect 20740 5394 20798 5399
rect 20740 5374 20743 5394
rect 20763 5380 20798 5394
rect 20818 5380 20827 5400
rect 20763 5372 20827 5380
rect 20789 5371 20827 5372
rect 20790 5370 20827 5371
rect 20893 5404 20929 5405
rect 21001 5404 21037 5405
rect 20893 5396 21037 5404
rect 20893 5376 20901 5396
rect 20921 5376 20956 5396
rect 20976 5376 21009 5396
rect 21029 5376 21037 5396
rect 20893 5370 21037 5376
rect 21103 5400 21141 5408
rect 21219 5404 21255 5405
rect 21103 5380 21112 5400
rect 21132 5380 21141 5400
rect 21103 5371 21141 5380
rect 21170 5396 21255 5404
rect 21170 5376 21227 5396
rect 21247 5376 21255 5396
rect 21103 5370 21140 5371
rect 21170 5370 21255 5376
rect 21321 5400 21359 5408
rect 21321 5380 21330 5400
rect 21350 5380 21359 5400
rect 21491 5398 21503 5416
rect 21521 5398 21531 5416
rect 21923 5444 21975 5633
rect 22321 5608 22360 5633
rect 22938 5648 23087 5655
rect 22938 5628 22997 5648
rect 23017 5628 23056 5648
rect 23076 5628 23087 5648
rect 22938 5620 23087 5628
rect 23154 5651 23311 5658
rect 23154 5631 23274 5651
rect 23294 5631 23311 5651
rect 23154 5621 23311 5631
rect 23154 5620 23189 5621
rect 22105 5583 22292 5607
rect 22321 5588 22716 5608
rect 22736 5588 22739 5608
rect 23154 5599 23185 5620
rect 23372 5599 23408 5709
rect 23427 5708 23464 5709
rect 23523 5708 23560 5709
rect 23483 5649 23573 5655
rect 23483 5629 23492 5649
rect 23512 5647 23573 5649
rect 23512 5629 23537 5647
rect 23483 5627 23537 5629
rect 23557 5627 23573 5647
rect 23483 5621 23573 5627
rect 22997 5598 23034 5599
rect 22321 5583 22739 5588
rect 22996 5589 23034 5598
rect 22105 5512 22142 5583
rect 22321 5582 22664 5583
rect 22321 5579 22360 5582
rect 22626 5581 22663 5582
rect 22257 5522 22288 5523
rect 22105 5492 22114 5512
rect 22134 5492 22142 5512
rect 22105 5482 22142 5492
rect 22201 5512 22288 5522
rect 22201 5492 22210 5512
rect 22230 5492 22288 5512
rect 22201 5483 22288 5492
rect 22201 5482 22238 5483
rect 21923 5426 21939 5444
rect 21957 5426 21975 5444
rect 22257 5432 22288 5483
rect 22323 5512 22360 5579
rect 22996 5569 23005 5589
rect 23025 5569 23034 5589
rect 22996 5561 23034 5569
rect 23100 5593 23185 5599
rect 23215 5598 23252 5599
rect 23100 5573 23108 5593
rect 23128 5573 23185 5593
rect 23100 5565 23185 5573
rect 23214 5589 23252 5598
rect 23214 5569 23223 5589
rect 23243 5569 23252 5589
rect 23100 5564 23136 5565
rect 23214 5561 23252 5569
rect 23318 5593 23462 5599
rect 23318 5573 23326 5593
rect 23346 5588 23434 5593
rect 23346 5573 23382 5588
rect 23318 5571 23382 5573
rect 23401 5573 23434 5588
rect 23454 5573 23462 5593
rect 23401 5571 23462 5573
rect 23318 5565 23462 5571
rect 23318 5564 23354 5565
rect 23426 5564 23462 5565
rect 23528 5598 23565 5599
rect 23528 5597 23566 5598
rect 23528 5589 23592 5597
rect 23528 5569 23537 5589
rect 23557 5575 23592 5589
rect 23612 5575 23615 5595
rect 23557 5570 23615 5575
rect 23557 5569 23592 5570
rect 22997 5532 23034 5561
rect 22998 5530 23034 5532
rect 22475 5522 22511 5523
rect 22323 5492 22332 5512
rect 22352 5492 22360 5512
rect 22323 5482 22360 5492
rect 22419 5512 22567 5522
rect 22667 5519 22763 5521
rect 22419 5492 22428 5512
rect 22448 5492 22538 5512
rect 22558 5492 22567 5512
rect 22419 5483 22567 5492
rect 22625 5512 22763 5519
rect 22625 5492 22634 5512
rect 22654 5492 22763 5512
rect 22998 5508 23189 5530
rect 23215 5529 23252 5561
rect 23528 5557 23592 5569
rect 23632 5531 23659 5709
rect 23491 5529 23659 5531
rect 23215 5515 23659 5529
rect 23683 5552 23711 6498
rect 23683 5522 23728 5552
rect 23215 5503 23662 5515
rect 23258 5501 23291 5503
rect 22625 5483 22763 5492
rect 22419 5482 22456 5483
rect 22149 5429 22190 5430
rect 21923 5408 21975 5426
rect 22041 5422 22190 5429
rect 21491 5388 21531 5398
rect 22041 5402 22100 5422
rect 22120 5402 22159 5422
rect 22179 5402 22190 5422
rect 22041 5394 22190 5402
rect 22257 5425 22414 5432
rect 22257 5405 22377 5425
rect 22397 5405 22414 5425
rect 22257 5395 22414 5405
rect 22257 5394 22292 5395
rect 21321 5371 21359 5380
rect 22257 5373 22288 5394
rect 22475 5373 22511 5483
rect 22530 5482 22567 5483
rect 22626 5482 22663 5483
rect 22586 5423 22676 5429
rect 22586 5403 22595 5423
rect 22615 5421 22676 5423
rect 22615 5403 22640 5421
rect 22586 5401 22640 5403
rect 22660 5401 22676 5421
rect 22586 5395 22676 5401
rect 22100 5372 22137 5373
rect 21321 5370 21358 5371
rect 20782 5342 20872 5348
rect 20782 5322 20798 5342
rect 20818 5340 20872 5342
rect 20818 5322 20843 5340
rect 20782 5320 20843 5322
rect 20863 5320 20872 5340
rect 20782 5314 20872 5320
rect 20795 5260 20832 5261
rect 20891 5260 20928 5261
rect 20947 5260 20983 5370
rect 21170 5349 21201 5370
rect 22099 5363 22137 5372
rect 21166 5348 21201 5349
rect 21044 5338 21201 5348
rect 21044 5318 21061 5338
rect 21081 5318 21201 5338
rect 21044 5311 21201 5318
rect 21268 5341 21417 5349
rect 21268 5321 21279 5341
rect 21299 5321 21338 5341
rect 21358 5321 21417 5341
rect 21927 5345 21967 5355
rect 21268 5314 21417 5321
rect 21483 5317 21535 5335
rect 21268 5313 21309 5314
rect 21002 5260 21039 5261
rect 19596 5245 19635 5260
rect 20695 5251 20833 5260
rect 19596 5244 19762 5245
rect 19888 5244 19928 5246
rect 19596 5218 20038 5244
rect 19596 5216 19762 5218
rect 19260 5104 19297 5112
rect 19260 5085 19268 5104
rect 19289 5085 19297 5104
rect 19260 5079 19297 5085
rect 19596 5038 19621 5216
rect 19661 5178 19725 5190
rect 20001 5186 20038 5218
rect 20064 5217 20255 5239
rect 20695 5231 20804 5251
rect 20824 5231 20833 5251
rect 20695 5224 20833 5231
rect 20891 5251 21039 5260
rect 20891 5231 20900 5251
rect 20920 5231 21010 5251
rect 21030 5231 21039 5251
rect 20695 5222 20791 5224
rect 20891 5221 21039 5231
rect 21098 5251 21135 5261
rect 21098 5231 21106 5251
rect 21126 5231 21135 5251
rect 20947 5220 20983 5221
rect 20219 5215 20255 5217
rect 20219 5186 20256 5215
rect 19661 5177 19696 5178
rect 19638 5172 19696 5177
rect 19638 5152 19641 5172
rect 19661 5158 19696 5172
rect 19716 5158 19725 5178
rect 19661 5150 19725 5158
rect 19687 5149 19725 5150
rect 19688 5148 19725 5149
rect 19791 5182 19827 5183
rect 19899 5182 19935 5183
rect 19791 5177 19935 5182
rect 19791 5174 19853 5177
rect 19791 5154 19799 5174
rect 19819 5154 19853 5174
rect 19791 5151 19853 5154
rect 19879 5174 19935 5177
rect 19879 5154 19907 5174
rect 19927 5154 19935 5174
rect 19879 5151 19935 5154
rect 19791 5148 19935 5151
rect 20001 5178 20039 5186
rect 20117 5182 20153 5183
rect 20001 5158 20010 5178
rect 20030 5158 20039 5178
rect 20001 5149 20039 5158
rect 20068 5174 20153 5182
rect 20068 5154 20125 5174
rect 20145 5154 20153 5174
rect 20001 5148 20038 5149
rect 20068 5148 20153 5154
rect 20219 5178 20257 5186
rect 20219 5158 20228 5178
rect 20248 5158 20257 5178
rect 21098 5164 21135 5231
rect 21170 5260 21201 5311
rect 21483 5299 21501 5317
rect 21519 5299 21535 5317
rect 21220 5260 21257 5261
rect 21170 5251 21257 5260
rect 21170 5231 21228 5251
rect 21248 5231 21257 5251
rect 21170 5221 21257 5231
rect 21316 5251 21353 5261
rect 21316 5231 21324 5251
rect 21344 5231 21353 5251
rect 21170 5220 21201 5221
rect 20795 5161 20832 5162
rect 21098 5161 21137 5164
rect 20794 5160 21137 5161
rect 21316 5160 21353 5231
rect 20219 5149 20257 5158
rect 20719 5155 21137 5160
rect 20219 5148 20256 5149
rect 19680 5120 19770 5126
rect 19680 5100 19696 5120
rect 19716 5118 19770 5120
rect 19716 5100 19741 5118
rect 19680 5098 19741 5100
rect 19761 5098 19770 5118
rect 19680 5092 19770 5098
rect 19693 5038 19730 5039
rect 19789 5038 19826 5039
rect 19845 5038 19881 5148
rect 20068 5127 20099 5148
rect 20719 5135 20722 5155
rect 20742 5135 21137 5155
rect 21166 5136 21353 5160
rect 20064 5126 20099 5127
rect 19942 5116 20099 5126
rect 19942 5096 19959 5116
rect 19979 5096 20099 5116
rect 19942 5089 20099 5096
rect 20166 5119 20315 5127
rect 20166 5099 20177 5119
rect 20197 5099 20236 5119
rect 20256 5099 20315 5119
rect 20166 5092 20315 5099
rect 21098 5110 21137 5135
rect 21483 5110 21535 5299
rect 21927 5327 21937 5345
rect 21955 5327 21967 5345
rect 22099 5343 22108 5363
rect 22128 5343 22137 5363
rect 22099 5335 22137 5343
rect 22203 5367 22288 5373
rect 22318 5372 22355 5373
rect 22203 5347 22211 5367
rect 22231 5347 22288 5367
rect 22203 5339 22288 5347
rect 22317 5363 22355 5372
rect 22317 5343 22326 5363
rect 22346 5343 22355 5363
rect 22203 5338 22239 5339
rect 22317 5335 22355 5343
rect 22421 5367 22565 5373
rect 22421 5347 22429 5367
rect 22449 5347 22482 5367
rect 22502 5347 22537 5367
rect 22557 5347 22565 5367
rect 22421 5339 22565 5347
rect 22421 5338 22457 5339
rect 22529 5338 22565 5339
rect 22631 5372 22668 5373
rect 22631 5371 22669 5372
rect 22631 5363 22695 5371
rect 22631 5343 22640 5363
rect 22660 5349 22695 5363
rect 22715 5349 22718 5369
rect 22660 5344 22718 5349
rect 22660 5343 22695 5344
rect 21927 5271 21967 5327
rect 22100 5306 22137 5335
rect 22101 5304 22137 5306
rect 22101 5282 22292 5304
rect 22318 5303 22355 5335
rect 22631 5331 22695 5343
rect 22735 5305 22762 5483
rect 23620 5458 23662 5503
rect 23683 5504 23694 5522
rect 23716 5504 23728 5522
rect 23683 5498 23728 5504
rect 23684 5497 23728 5498
rect 22594 5303 22762 5305
rect 22318 5293 22762 5303
rect 22903 5399 23090 5423
rect 23121 5404 23514 5424
rect 23534 5404 23537 5424
rect 23121 5399 23537 5404
rect 22903 5328 22940 5399
rect 23121 5398 23462 5399
rect 23055 5338 23086 5339
rect 22903 5308 22912 5328
rect 22932 5308 22940 5328
rect 22903 5298 22940 5308
rect 22999 5328 23086 5338
rect 22999 5308 23008 5328
rect 23028 5308 23086 5328
rect 22999 5299 23086 5308
rect 22999 5298 23036 5299
rect 21924 5266 21967 5271
rect 22315 5277 22762 5293
rect 22315 5271 22343 5277
rect 22594 5276 22762 5277
rect 21924 5263 22074 5266
rect 22315 5263 22342 5271
rect 21924 5261 22342 5263
rect 21924 5243 21933 5261
rect 21951 5243 22342 5261
rect 23055 5248 23086 5299
rect 23121 5328 23158 5398
rect 23424 5397 23461 5398
rect 23273 5338 23309 5339
rect 23121 5308 23130 5328
rect 23150 5308 23158 5328
rect 23121 5298 23158 5308
rect 23217 5328 23365 5338
rect 23465 5335 23561 5337
rect 23217 5308 23226 5328
rect 23246 5308 23336 5328
rect 23356 5308 23365 5328
rect 23217 5299 23365 5308
rect 23423 5328 23561 5335
rect 23423 5308 23432 5328
rect 23452 5308 23561 5328
rect 23423 5299 23561 5308
rect 23217 5298 23254 5299
rect 22947 5245 22988 5246
rect 21924 5240 22342 5243
rect 21924 5234 21967 5240
rect 21927 5231 21967 5234
rect 22842 5238 22988 5245
rect 22324 5222 22364 5223
rect 22035 5205 22364 5222
rect 22842 5218 22898 5238
rect 22918 5218 22957 5238
rect 22977 5218 22988 5238
rect 22842 5210 22988 5218
rect 23055 5241 23212 5248
rect 23055 5221 23175 5241
rect 23195 5221 23212 5241
rect 23055 5211 23212 5221
rect 23055 5210 23090 5211
rect 21919 5162 21962 5173
rect 21919 5144 21931 5162
rect 21949 5144 21962 5162
rect 21919 5118 21962 5144
rect 22035 5118 22062 5205
rect 22324 5196 22364 5205
rect 21098 5092 21537 5110
rect 20166 5091 20207 5092
rect 19900 5038 19937 5039
rect 19596 5029 19731 5038
rect 19596 5009 19702 5029
rect 19722 5009 19731 5029
rect 19596 5002 19731 5009
rect 19789 5029 19937 5038
rect 19789 5009 19798 5029
rect 19818 5009 19908 5029
rect 19928 5009 19937 5029
rect 19596 5000 19689 5002
rect 19789 4999 19937 5009
rect 19996 5029 20033 5039
rect 19996 5009 20004 5029
rect 20024 5009 20033 5029
rect 19845 4998 19881 4999
rect 19693 4939 19730 4940
rect 19996 4939 20033 5009
rect 20068 5038 20099 5089
rect 21098 5074 21498 5092
rect 21516 5074 21537 5092
rect 21098 5068 21537 5074
rect 21104 5064 21537 5068
rect 21919 5097 22062 5118
rect 22106 5170 22140 5186
rect 22324 5176 22717 5196
rect 22737 5176 22740 5196
rect 23055 5189 23086 5210
rect 23273 5189 23309 5299
rect 23328 5298 23365 5299
rect 23424 5298 23461 5299
rect 23384 5239 23474 5245
rect 23384 5219 23393 5239
rect 23413 5237 23474 5239
rect 23413 5219 23438 5237
rect 23384 5217 23438 5219
rect 23458 5217 23474 5237
rect 23384 5211 23474 5217
rect 22898 5188 22935 5189
rect 22324 5171 22740 5176
rect 22897 5179 22935 5188
rect 22324 5170 22665 5171
rect 22106 5100 22143 5170
rect 22258 5110 22289 5111
rect 21919 5095 22056 5097
rect 21483 5062 21535 5064
rect 21919 5053 21962 5095
rect 22106 5080 22115 5100
rect 22135 5080 22143 5100
rect 22106 5070 22143 5080
rect 22202 5100 22289 5110
rect 22202 5080 22211 5100
rect 22231 5080 22289 5100
rect 22202 5071 22289 5080
rect 22202 5070 22239 5071
rect 21917 5043 21962 5053
rect 20118 5038 20155 5039
rect 20068 5029 20155 5038
rect 20068 5009 20126 5029
rect 20146 5009 20155 5029
rect 20068 4999 20155 5009
rect 20214 5029 20251 5039
rect 20214 5009 20222 5029
rect 20242 5009 20251 5029
rect 21917 5025 21926 5043
rect 21944 5025 21962 5043
rect 21917 5019 21962 5025
rect 22258 5020 22289 5071
rect 22324 5100 22361 5170
rect 22627 5169 22664 5170
rect 22897 5159 22906 5179
rect 22926 5159 22935 5179
rect 22897 5151 22935 5159
rect 23001 5183 23086 5189
rect 23116 5188 23153 5189
rect 23001 5163 23009 5183
rect 23029 5163 23086 5183
rect 23001 5155 23086 5163
rect 23115 5179 23153 5188
rect 23115 5159 23124 5179
rect 23144 5159 23153 5179
rect 23001 5154 23037 5155
rect 23115 5151 23153 5159
rect 23219 5183 23363 5189
rect 23219 5163 23227 5183
rect 23247 5180 23335 5183
rect 23247 5163 23282 5180
rect 23219 5162 23282 5163
rect 23301 5163 23335 5180
rect 23355 5163 23363 5183
rect 23301 5162 23363 5163
rect 23219 5155 23363 5162
rect 23219 5154 23255 5155
rect 23327 5154 23363 5155
rect 23429 5188 23466 5189
rect 23429 5187 23467 5188
rect 23489 5187 23516 5191
rect 23429 5185 23516 5187
rect 23429 5179 23493 5185
rect 23429 5159 23438 5179
rect 23458 5165 23493 5179
rect 23513 5165 23516 5185
rect 23458 5160 23516 5165
rect 23458 5159 23493 5160
rect 22898 5122 22935 5151
rect 22899 5120 22935 5122
rect 22476 5110 22512 5111
rect 22324 5080 22333 5100
rect 22353 5080 22361 5100
rect 22324 5070 22361 5080
rect 22420 5100 22568 5110
rect 22668 5107 22764 5109
rect 22420 5080 22429 5100
rect 22449 5080 22539 5100
rect 22559 5080 22568 5100
rect 22420 5071 22568 5080
rect 22626 5100 22764 5107
rect 22626 5080 22635 5100
rect 22655 5080 22764 5100
rect 22899 5098 23090 5120
rect 23116 5119 23153 5151
rect 23429 5147 23493 5159
rect 23533 5121 23560 5299
rect 23392 5119 23560 5121
rect 23116 5093 23560 5119
rect 22626 5071 22764 5080
rect 22420 5070 22457 5071
rect 21917 5016 21954 5019
rect 22150 5017 22191 5018
rect 20068 4998 20099 4999
rect 19692 4938 20033 4939
rect 20214 4938 20251 5009
rect 22042 5010 22191 5017
rect 21486 4997 21523 5002
rect 19617 4933 20033 4938
rect 19617 4913 19620 4933
rect 19640 4913 20033 4933
rect 20064 4914 20251 4938
rect 21477 4993 21524 4997
rect 21477 4975 21496 4993
rect 21514 4975 21524 4993
rect 22042 4990 22101 5010
rect 22121 4990 22160 5010
rect 22180 4990 22191 5010
rect 22042 4982 22191 4990
rect 22258 5013 22415 5020
rect 22258 4993 22378 5013
rect 22398 4993 22415 5013
rect 22258 4983 22415 4993
rect 22258 4982 22293 4983
rect 21085 4916 21123 4917
rect 21477 4916 21524 4975
rect 22258 4961 22289 4982
rect 22476 4961 22512 5071
rect 22531 5070 22568 5071
rect 22627 5070 22664 5071
rect 22587 5011 22677 5017
rect 22587 4991 22596 5011
rect 22616 5009 22677 5011
rect 22616 4991 22641 5009
rect 22587 4989 22641 4991
rect 22661 4989 22677 5009
rect 22587 4983 22677 4989
rect 22101 4960 22138 4961
rect 21914 4952 21951 4954
rect 21914 4944 21956 4952
rect 21914 4926 21924 4944
rect 21942 4926 21956 4944
rect 21914 4917 21956 4926
rect 22100 4951 22138 4960
rect 22100 4931 22109 4951
rect 22129 4931 22138 4951
rect 22100 4923 22138 4931
rect 22204 4955 22289 4961
rect 22319 4960 22356 4961
rect 22204 4935 22212 4955
rect 22232 4935 22289 4955
rect 22204 4927 22289 4935
rect 22318 4951 22356 4960
rect 22318 4931 22327 4951
rect 22347 4931 22356 4951
rect 22204 4926 22240 4927
rect 22318 4923 22356 4931
rect 22422 4959 22566 4961
rect 22422 4955 22474 4959
rect 22422 4935 22430 4955
rect 22450 4939 22474 4955
rect 22494 4955 22566 4959
rect 22494 4939 22538 4955
rect 22450 4935 22538 4939
rect 22558 4935 22566 4955
rect 22422 4927 22566 4935
rect 22422 4926 22458 4927
rect 22530 4926 22566 4927
rect 22632 4960 22669 4961
rect 22632 4959 22670 4960
rect 22632 4951 22696 4959
rect 22632 4931 22641 4951
rect 22661 4937 22696 4951
rect 22716 4937 22719 4957
rect 22661 4932 22719 4937
rect 22661 4931 22696 4932
rect 19837 4912 19902 4913
rect 17952 4834 17990 4835
rect 16477 4819 16512 4820
rect 16454 4814 16512 4819
rect 16454 4794 16457 4814
rect 16477 4800 16512 4814
rect 16532 4800 16541 4820
rect 16477 4792 16541 4800
rect 16503 4791 16541 4792
rect 16504 4790 16541 4791
rect 16607 4824 16643 4825
rect 16715 4824 16751 4825
rect 16607 4816 16751 4824
rect 16607 4796 16615 4816
rect 16635 4812 16723 4816
rect 16635 4796 16679 4812
rect 16607 4792 16679 4796
rect 16699 4796 16723 4812
rect 16743 4796 16751 4816
rect 16699 4792 16751 4796
rect 16607 4790 16751 4792
rect 16817 4820 16855 4828
rect 16933 4824 16969 4825
rect 16817 4800 16826 4820
rect 16846 4800 16855 4820
rect 16817 4791 16855 4800
rect 16884 4816 16969 4824
rect 16884 4796 16941 4816
rect 16961 4796 16969 4816
rect 16817 4790 16854 4791
rect 16884 4790 16969 4796
rect 17035 4820 17073 4828
rect 17035 4800 17044 4820
rect 17064 4800 17073 4820
rect 17035 4791 17073 4800
rect 17217 4825 17259 4834
rect 17217 4807 17231 4825
rect 17249 4807 17259 4825
rect 17217 4799 17259 4807
rect 17222 4797 17259 4799
rect 17551 4796 17990 4834
rect 18862 4834 18870 4856
rect 18894 4834 18902 4856
rect 18862 4826 18902 4834
rect 20173 4878 20213 4886
rect 20173 4856 20181 4878
rect 20205 4856 20213 4878
rect 21085 4878 21524 4916
rect 21085 4877 21123 4878
rect 19173 4799 19238 4800
rect 17035 4790 17072 4791
rect 16496 4762 16586 4768
rect 16496 4742 16512 4762
rect 16532 4760 16586 4762
rect 16532 4742 16557 4760
rect 16496 4740 16557 4742
rect 16577 4740 16586 4760
rect 16496 4734 16586 4740
rect 16509 4680 16546 4681
rect 16605 4680 16642 4681
rect 16661 4680 16697 4790
rect 16884 4769 16915 4790
rect 16880 4768 16915 4769
rect 16758 4758 16915 4768
rect 16758 4738 16775 4758
rect 16795 4738 16915 4758
rect 16758 4731 16915 4738
rect 16982 4761 17131 4769
rect 16982 4741 16993 4761
rect 17013 4741 17052 4761
rect 17072 4741 17131 4761
rect 16982 4734 17131 4741
rect 17551 4737 17598 4796
rect 17952 4795 17990 4796
rect 16982 4733 17023 4734
rect 17219 4732 17256 4735
rect 16716 4680 16753 4681
rect 16409 4671 16547 4680
rect 15613 4632 16057 4658
rect 15613 4630 15781 4632
rect 15613 4452 15640 4630
rect 15680 4592 15744 4604
rect 16020 4600 16057 4632
rect 16083 4631 16274 4653
rect 16409 4651 16518 4671
rect 16538 4651 16547 4671
rect 16409 4644 16547 4651
rect 16605 4671 16753 4680
rect 16605 4651 16614 4671
rect 16634 4651 16724 4671
rect 16744 4651 16753 4671
rect 16409 4642 16505 4644
rect 16605 4641 16753 4651
rect 16812 4671 16849 4681
rect 16812 4651 16820 4671
rect 16840 4651 16849 4671
rect 16661 4640 16697 4641
rect 16238 4629 16274 4631
rect 16238 4600 16275 4629
rect 15680 4591 15715 4592
rect 15657 4586 15715 4591
rect 15657 4566 15660 4586
rect 15680 4572 15715 4586
rect 15735 4572 15744 4592
rect 15680 4566 15744 4572
rect 15657 4564 15744 4566
rect 15657 4560 15684 4564
rect 15706 4563 15744 4564
rect 15707 4562 15744 4563
rect 15810 4596 15846 4597
rect 15918 4596 15954 4597
rect 15810 4589 15954 4596
rect 15810 4588 15872 4589
rect 15810 4568 15818 4588
rect 15838 4571 15872 4588
rect 15891 4588 15954 4589
rect 15891 4571 15926 4588
rect 15838 4568 15926 4571
rect 15946 4568 15954 4588
rect 15810 4562 15954 4568
rect 16020 4592 16058 4600
rect 16136 4596 16172 4597
rect 16020 4572 16029 4592
rect 16049 4572 16058 4592
rect 16020 4563 16058 4572
rect 16087 4588 16172 4596
rect 16087 4568 16144 4588
rect 16164 4568 16172 4588
rect 16020 4562 16057 4563
rect 16087 4562 16172 4568
rect 16238 4592 16276 4600
rect 16238 4572 16247 4592
rect 16267 4572 16276 4592
rect 16509 4581 16546 4582
rect 16812 4581 16849 4651
rect 16884 4680 16915 4731
rect 17211 4726 17256 4732
rect 17211 4708 17229 4726
rect 17247 4708 17256 4726
rect 17551 4719 17561 4737
rect 17579 4719 17598 4737
rect 17551 4715 17598 4719
rect 18824 4774 19011 4798
rect 19042 4779 19435 4799
rect 19455 4779 19458 4799
rect 19042 4774 19458 4779
rect 17552 4710 17589 4715
rect 17211 4698 17256 4708
rect 18824 4703 18861 4774
rect 19042 4773 19383 4774
rect 18976 4713 19007 4714
rect 16934 4680 16971 4681
rect 16884 4671 16971 4680
rect 16884 4651 16942 4671
rect 16962 4651 16971 4671
rect 16884 4641 16971 4651
rect 17030 4671 17067 4681
rect 17030 4651 17038 4671
rect 17058 4651 17067 4671
rect 17211 4656 17254 4698
rect 18824 4683 18833 4703
rect 18853 4683 18861 4703
rect 18824 4673 18861 4683
rect 18920 4703 19007 4713
rect 18920 4683 18929 4703
rect 18949 4683 19007 4703
rect 18920 4674 19007 4683
rect 18920 4673 18957 4674
rect 17117 4654 17254 4656
rect 16884 4640 16915 4641
rect 17030 4581 17067 4651
rect 16508 4580 16849 4581
rect 16238 4563 16276 4572
rect 16433 4575 16849 4580
rect 16238 4562 16275 4563
rect 15699 4534 15789 4540
rect 15699 4514 15715 4534
rect 15735 4532 15789 4534
rect 15735 4514 15760 4532
rect 15699 4512 15760 4514
rect 15780 4512 15789 4532
rect 15699 4506 15789 4512
rect 15712 4452 15749 4453
rect 15808 4452 15845 4453
rect 15864 4452 15900 4562
rect 16087 4541 16118 4562
rect 16433 4555 16436 4575
rect 16456 4555 16849 4575
rect 17033 4565 17067 4581
rect 17111 4633 17254 4654
rect 17540 4648 17592 4650
rect 16809 4546 16849 4555
rect 17111 4546 17138 4633
rect 17211 4607 17254 4633
rect 17211 4589 17224 4607
rect 17242 4589 17254 4607
rect 17538 4644 17971 4648
rect 17538 4638 17977 4644
rect 17538 4620 17559 4638
rect 17577 4620 17977 4638
rect 18976 4623 19007 4674
rect 19042 4703 19079 4773
rect 19345 4772 19382 4773
rect 19194 4713 19230 4714
rect 19042 4683 19051 4703
rect 19071 4683 19079 4703
rect 19042 4673 19079 4683
rect 19138 4703 19286 4713
rect 19386 4710 19482 4712
rect 19138 4683 19147 4703
rect 19167 4683 19257 4703
rect 19277 4683 19286 4703
rect 19138 4674 19286 4683
rect 19344 4703 19482 4710
rect 19344 4683 19353 4703
rect 19373 4683 19482 4703
rect 19344 4674 19482 4683
rect 19138 4673 19175 4674
rect 18868 4620 18909 4621
rect 17538 4602 17977 4620
rect 17211 4578 17254 4589
rect 16083 4540 16118 4541
rect 15961 4530 16118 4540
rect 15961 4510 15978 4530
rect 15998 4510 16118 4530
rect 15961 4503 16118 4510
rect 16185 4533 16331 4541
rect 16185 4513 16196 4533
rect 16216 4513 16255 4533
rect 16275 4513 16331 4533
rect 16809 4529 17138 4546
rect 16809 4528 16849 4529
rect 16185 4506 16331 4513
rect 17206 4517 17246 4520
rect 17206 4511 17249 4517
rect 16831 4508 17249 4511
rect 16185 4505 16226 4506
rect 15919 4452 15956 4453
rect 15612 4443 15750 4452
rect 15612 4423 15721 4443
rect 15741 4423 15750 4443
rect 15612 4416 15750 4423
rect 15808 4443 15956 4452
rect 15808 4423 15817 4443
rect 15837 4423 15927 4443
rect 15947 4423 15956 4443
rect 15612 4414 15708 4416
rect 15808 4413 15956 4423
rect 16015 4443 16052 4453
rect 16015 4423 16023 4443
rect 16043 4423 16052 4443
rect 15864 4412 15900 4413
rect 15712 4353 15749 4354
rect 16015 4353 16052 4423
rect 16087 4452 16118 4503
rect 16831 4490 17222 4508
rect 17240 4490 17249 4508
rect 16831 4488 17249 4490
rect 16831 4480 16858 4488
rect 17099 4485 17249 4488
rect 16411 4474 16579 4475
rect 16830 4474 16858 4480
rect 16411 4458 16858 4474
rect 17206 4480 17249 4485
rect 16137 4452 16174 4453
rect 16087 4443 16174 4452
rect 16087 4423 16145 4443
rect 16165 4423 16174 4443
rect 16087 4413 16174 4423
rect 16233 4443 16270 4453
rect 16233 4423 16241 4443
rect 16261 4423 16270 4443
rect 16087 4412 16118 4413
rect 15711 4352 16052 4353
rect 16233 4352 16270 4423
rect 15636 4347 16052 4352
rect 15636 4327 15639 4347
rect 15659 4327 16052 4347
rect 16083 4328 16270 4352
rect 16411 4448 16855 4458
rect 16411 4446 16579 4448
rect 15445 4253 15489 4254
rect 15445 4247 15490 4253
rect 15445 4229 15457 4247
rect 15479 4229 15490 4247
rect 15511 4248 15553 4293
rect 16411 4268 16438 4446
rect 16478 4408 16542 4420
rect 16818 4416 16855 4448
rect 16881 4447 17072 4469
rect 17036 4445 17072 4447
rect 17036 4416 17073 4445
rect 17206 4424 17246 4480
rect 16478 4407 16513 4408
rect 16455 4402 16513 4407
rect 16455 4382 16458 4402
rect 16478 4388 16513 4402
rect 16533 4388 16542 4408
rect 16478 4380 16542 4388
rect 16504 4379 16542 4380
rect 16505 4378 16542 4379
rect 16608 4412 16644 4413
rect 16716 4412 16752 4413
rect 16608 4404 16752 4412
rect 16608 4384 16616 4404
rect 16636 4384 16671 4404
rect 16691 4384 16724 4404
rect 16744 4384 16752 4404
rect 16608 4378 16752 4384
rect 16818 4408 16856 4416
rect 16934 4412 16970 4413
rect 16818 4388 16827 4408
rect 16847 4388 16856 4408
rect 16818 4379 16856 4388
rect 16885 4404 16970 4412
rect 16885 4384 16942 4404
rect 16962 4384 16970 4404
rect 16818 4378 16855 4379
rect 16885 4378 16970 4384
rect 17036 4408 17074 4416
rect 17036 4388 17045 4408
rect 17065 4388 17074 4408
rect 17206 4406 17218 4424
rect 17236 4406 17246 4424
rect 17206 4396 17246 4406
rect 17540 4413 17592 4602
rect 17938 4577 17977 4602
rect 18760 4613 18909 4620
rect 18760 4593 18819 4613
rect 18839 4593 18878 4613
rect 18898 4593 18909 4613
rect 18760 4585 18909 4593
rect 18976 4616 19133 4623
rect 18976 4596 19096 4616
rect 19116 4596 19133 4616
rect 18976 4586 19133 4596
rect 18976 4585 19011 4586
rect 17722 4552 17909 4576
rect 17938 4557 18333 4577
rect 18353 4557 18356 4577
rect 18976 4564 19007 4585
rect 19194 4564 19230 4674
rect 19249 4673 19286 4674
rect 19345 4673 19382 4674
rect 19305 4614 19395 4620
rect 19305 4594 19314 4614
rect 19334 4612 19395 4614
rect 19334 4594 19359 4612
rect 19305 4592 19359 4594
rect 19379 4592 19395 4612
rect 19305 4586 19395 4592
rect 18819 4563 18856 4564
rect 17938 4552 18356 4557
rect 18818 4554 18856 4563
rect 17722 4481 17759 4552
rect 17938 4551 18281 4552
rect 17938 4548 17977 4551
rect 18243 4550 18280 4551
rect 17874 4491 17905 4492
rect 17722 4461 17731 4481
rect 17751 4461 17759 4481
rect 17722 4451 17759 4461
rect 17818 4481 17905 4491
rect 17818 4461 17827 4481
rect 17847 4461 17905 4481
rect 17818 4452 17905 4461
rect 17818 4451 17855 4452
rect 17036 4379 17074 4388
rect 17540 4395 17556 4413
rect 17574 4395 17592 4413
rect 17874 4401 17905 4452
rect 17940 4481 17977 4548
rect 18818 4534 18827 4554
rect 18847 4534 18856 4554
rect 18818 4526 18856 4534
rect 18922 4558 19007 4564
rect 19037 4563 19074 4564
rect 18922 4538 18930 4558
rect 18950 4538 19007 4558
rect 18922 4530 19007 4538
rect 19036 4554 19074 4563
rect 19036 4534 19045 4554
rect 19065 4534 19074 4554
rect 18922 4529 18958 4530
rect 19036 4526 19074 4534
rect 19140 4558 19284 4564
rect 19140 4538 19148 4558
rect 19168 4552 19256 4558
rect 19168 4538 19197 4552
rect 19140 4530 19197 4538
rect 19140 4529 19176 4530
rect 19220 4538 19256 4552
rect 19276 4538 19284 4558
rect 19220 4530 19284 4538
rect 19248 4529 19284 4530
rect 19350 4563 19387 4564
rect 19350 4562 19388 4563
rect 19350 4554 19414 4562
rect 19350 4534 19359 4554
rect 19379 4540 19414 4554
rect 19434 4540 19437 4560
rect 19379 4535 19437 4540
rect 19379 4534 19414 4535
rect 18819 4497 18856 4526
rect 18820 4495 18856 4497
rect 18092 4491 18128 4492
rect 17940 4461 17949 4481
rect 17969 4461 17977 4481
rect 17940 4451 17977 4461
rect 18036 4481 18184 4491
rect 18284 4488 18380 4490
rect 18036 4461 18045 4481
rect 18065 4461 18155 4481
rect 18175 4461 18184 4481
rect 18036 4452 18184 4461
rect 18242 4481 18380 4488
rect 18242 4461 18251 4481
rect 18271 4461 18380 4481
rect 18820 4473 19011 4495
rect 19037 4494 19074 4526
rect 19350 4522 19414 4534
rect 19454 4496 19481 4674
rect 19778 4627 19815 4633
rect 19778 4608 19786 4627
rect 19807 4608 19815 4627
rect 19778 4600 19815 4608
rect 19313 4494 19481 4496
rect 19037 4468 19481 4494
rect 19147 4466 19187 4468
rect 19313 4467 19481 4468
rect 18242 4452 18380 4461
rect 19440 4462 19481 4467
rect 18036 4451 18073 4452
rect 17766 4398 17807 4399
rect 17036 4378 17073 4379
rect 16497 4350 16587 4356
rect 16497 4330 16513 4350
rect 16533 4348 16587 4350
rect 16533 4330 16558 4348
rect 16497 4328 16558 4330
rect 16578 4328 16587 4348
rect 16497 4322 16587 4328
rect 16510 4268 16547 4269
rect 16606 4268 16643 4269
rect 16662 4268 16698 4378
rect 16885 4357 16916 4378
rect 17540 4377 17592 4395
rect 17658 4391 17807 4398
rect 17658 4371 17717 4391
rect 17737 4371 17776 4391
rect 17796 4371 17807 4391
rect 17658 4363 17807 4371
rect 17874 4394 18031 4401
rect 17874 4374 17994 4394
rect 18014 4374 18031 4394
rect 17874 4364 18031 4374
rect 17874 4363 17909 4364
rect 16881 4356 16916 4357
rect 16759 4346 16916 4356
rect 16759 4326 16776 4346
rect 16796 4326 16916 4346
rect 16759 4319 16916 4326
rect 16983 4349 17132 4357
rect 16983 4329 16994 4349
rect 17014 4329 17053 4349
rect 17073 4329 17132 4349
rect 16983 4322 17132 4329
rect 17198 4325 17250 4343
rect 17874 4342 17905 4363
rect 18092 4342 18128 4452
rect 18147 4451 18184 4452
rect 18243 4451 18280 4452
rect 18203 4392 18293 4398
rect 18203 4372 18212 4392
rect 18232 4390 18293 4392
rect 18232 4372 18257 4390
rect 18203 4370 18257 4372
rect 18277 4370 18293 4390
rect 18203 4364 18293 4370
rect 17717 4341 17754 4342
rect 16983 4321 17024 4322
rect 16717 4268 16754 4269
rect 16410 4259 16548 4268
rect 15882 4248 15915 4250
rect 15511 4236 15958 4248
rect 15445 4199 15490 4229
rect 15462 3253 15490 4199
rect 15514 4222 15958 4236
rect 15514 4220 15682 4222
rect 15514 4042 15541 4220
rect 15581 4182 15645 4194
rect 15921 4190 15958 4222
rect 15984 4221 16175 4243
rect 16410 4239 16519 4259
rect 16539 4239 16548 4259
rect 16410 4232 16548 4239
rect 16606 4259 16754 4268
rect 16606 4239 16615 4259
rect 16635 4239 16725 4259
rect 16745 4239 16754 4259
rect 16410 4230 16506 4232
rect 16606 4229 16754 4239
rect 16813 4259 16850 4269
rect 16813 4239 16821 4259
rect 16841 4239 16850 4259
rect 16662 4228 16698 4229
rect 16139 4219 16175 4221
rect 16139 4190 16176 4219
rect 15581 4181 15616 4182
rect 15558 4176 15616 4181
rect 15558 4156 15561 4176
rect 15581 4162 15616 4176
rect 15636 4162 15645 4182
rect 15581 4154 15645 4162
rect 15607 4153 15645 4154
rect 15608 4152 15645 4153
rect 15711 4186 15747 4187
rect 15819 4186 15855 4187
rect 15711 4180 15855 4186
rect 15711 4178 15772 4180
rect 15711 4158 15719 4178
rect 15739 4163 15772 4178
rect 15791 4178 15855 4180
rect 15791 4163 15827 4178
rect 15739 4158 15827 4163
rect 15847 4158 15855 4178
rect 15711 4152 15855 4158
rect 15921 4182 15959 4190
rect 16037 4186 16073 4187
rect 15921 4162 15930 4182
rect 15950 4162 15959 4182
rect 15921 4153 15959 4162
rect 15988 4178 16073 4186
rect 15988 4158 16045 4178
rect 16065 4158 16073 4178
rect 15921 4152 15958 4153
rect 15988 4152 16073 4158
rect 16139 4182 16177 4190
rect 16139 4162 16148 4182
rect 16168 4162 16177 4182
rect 16813 4172 16850 4239
rect 16885 4268 16916 4319
rect 17198 4307 17216 4325
rect 17234 4307 17250 4325
rect 17716 4332 17754 4341
rect 16935 4268 16972 4269
rect 16885 4259 16972 4268
rect 16885 4239 16943 4259
rect 16963 4239 16972 4259
rect 16885 4229 16972 4239
rect 17031 4259 17068 4269
rect 17031 4239 17039 4259
rect 17059 4239 17068 4259
rect 16885 4228 16916 4229
rect 16510 4169 16547 4170
rect 16813 4169 16852 4172
rect 16509 4168 16852 4169
rect 17031 4168 17068 4239
rect 16139 4153 16177 4162
rect 16434 4163 16852 4168
rect 16139 4152 16176 4153
rect 15600 4124 15690 4130
rect 15600 4104 15616 4124
rect 15636 4122 15690 4124
rect 15636 4104 15661 4122
rect 15600 4102 15661 4104
rect 15681 4102 15690 4122
rect 15600 4096 15690 4102
rect 15613 4042 15650 4043
rect 15709 4042 15746 4043
rect 15765 4042 15801 4152
rect 15988 4131 16019 4152
rect 16434 4143 16437 4163
rect 16457 4143 16852 4163
rect 16881 4144 17068 4168
rect 15984 4130 16019 4131
rect 15862 4120 16019 4130
rect 15862 4100 15879 4120
rect 15899 4100 16019 4120
rect 15862 4093 16019 4100
rect 16086 4123 16235 4131
rect 16086 4103 16097 4123
rect 16117 4103 16156 4123
rect 16176 4103 16235 4123
rect 16086 4096 16235 4103
rect 16813 4118 16852 4143
rect 17198 4118 17250 4307
rect 17544 4314 17584 4324
rect 17544 4296 17554 4314
rect 17572 4296 17584 4314
rect 17716 4312 17725 4332
rect 17745 4312 17754 4332
rect 17716 4304 17754 4312
rect 17820 4336 17905 4342
rect 17935 4341 17972 4342
rect 17820 4316 17828 4336
rect 17848 4316 17905 4336
rect 17820 4308 17905 4316
rect 17934 4332 17972 4341
rect 17934 4312 17943 4332
rect 17963 4312 17972 4332
rect 17820 4307 17856 4308
rect 17934 4304 17972 4312
rect 18038 4336 18182 4342
rect 18038 4316 18046 4336
rect 18066 4316 18099 4336
rect 18119 4316 18154 4336
rect 18174 4316 18182 4336
rect 18038 4308 18182 4316
rect 18038 4307 18074 4308
rect 18146 4307 18182 4308
rect 18248 4341 18285 4342
rect 18248 4340 18286 4341
rect 18248 4332 18312 4340
rect 18248 4312 18257 4332
rect 18277 4318 18312 4332
rect 18332 4318 18335 4338
rect 18277 4313 18335 4318
rect 18277 4312 18312 4313
rect 17544 4240 17584 4296
rect 17717 4275 17754 4304
rect 17718 4273 17754 4275
rect 17718 4251 17909 4273
rect 17935 4272 17972 4304
rect 18248 4300 18312 4312
rect 18352 4274 18379 4452
rect 18211 4272 18379 4274
rect 17935 4262 18379 4272
rect 18520 4368 18707 4392
rect 18738 4373 19131 4393
rect 19151 4373 19154 4393
rect 18738 4368 19154 4373
rect 18520 4297 18557 4368
rect 18738 4367 19079 4368
rect 18672 4307 18703 4308
rect 18520 4277 18529 4297
rect 18549 4277 18557 4297
rect 18520 4267 18557 4277
rect 18616 4297 18703 4307
rect 18616 4277 18625 4297
rect 18645 4277 18703 4297
rect 18616 4268 18703 4277
rect 18616 4267 18653 4268
rect 17541 4235 17584 4240
rect 17932 4246 18379 4262
rect 17932 4240 17960 4246
rect 18211 4245 18379 4246
rect 17541 4232 17691 4235
rect 17932 4232 17959 4240
rect 17541 4230 17959 4232
rect 17541 4212 17550 4230
rect 17568 4212 17959 4230
rect 18672 4217 18703 4268
rect 18738 4297 18775 4367
rect 19041 4366 19078 4367
rect 18890 4307 18926 4308
rect 18738 4277 18747 4297
rect 18767 4277 18775 4297
rect 18738 4267 18775 4277
rect 18834 4297 18982 4307
rect 19082 4304 19178 4306
rect 18834 4277 18843 4297
rect 18863 4277 18953 4297
rect 18973 4277 18982 4297
rect 18834 4268 18982 4277
rect 19040 4297 19178 4304
rect 19040 4277 19049 4297
rect 19069 4277 19178 4297
rect 19440 4280 19480 4462
rect 19040 4268 19178 4277
rect 18834 4267 18871 4268
rect 18564 4214 18605 4215
rect 17541 4209 17959 4212
rect 17541 4203 17584 4209
rect 17544 4200 17584 4203
rect 18456 4207 18605 4214
rect 17941 4191 17981 4192
rect 17652 4174 17981 4191
rect 18456 4187 18515 4207
rect 18535 4187 18574 4207
rect 18594 4187 18605 4207
rect 18456 4179 18605 4187
rect 18672 4210 18829 4217
rect 18672 4190 18792 4210
rect 18812 4190 18829 4210
rect 18672 4180 18829 4190
rect 18672 4179 18707 4180
rect 17536 4131 17579 4142
rect 16813 4100 17252 4118
rect 16086 4095 16127 4096
rect 15820 4042 15857 4043
rect 15513 4033 15651 4042
rect 15513 4013 15622 4033
rect 15642 4013 15651 4033
rect 15513 4006 15651 4013
rect 15709 4033 15857 4042
rect 15709 4013 15718 4033
rect 15738 4013 15828 4033
rect 15848 4013 15857 4033
rect 15513 4004 15609 4006
rect 15709 4003 15857 4013
rect 15916 4033 15953 4043
rect 15916 4013 15924 4033
rect 15944 4013 15953 4033
rect 15765 4002 15801 4003
rect 15613 3943 15650 3944
rect 15916 3943 15953 4013
rect 15988 4042 16019 4093
rect 16813 4082 17213 4100
rect 17231 4082 17252 4100
rect 16813 4076 17252 4082
rect 16819 4072 17252 4076
rect 17536 4113 17548 4131
rect 17566 4113 17579 4131
rect 17536 4087 17579 4113
rect 17652 4087 17679 4174
rect 17941 4165 17981 4174
rect 17198 4070 17250 4072
rect 17536 4066 17679 4087
rect 17723 4139 17757 4155
rect 17941 4145 18334 4165
rect 18354 4145 18357 4165
rect 18672 4158 18703 4179
rect 18890 4158 18926 4268
rect 18945 4267 18982 4268
rect 19041 4267 19078 4268
rect 19001 4208 19091 4214
rect 19001 4188 19010 4208
rect 19030 4206 19091 4208
rect 19030 4188 19055 4206
rect 19001 4186 19055 4188
rect 19075 4186 19091 4206
rect 19001 4180 19091 4186
rect 18515 4157 18552 4158
rect 17941 4140 18357 4145
rect 18514 4148 18552 4157
rect 17941 4139 18282 4140
rect 17723 4069 17760 4139
rect 17875 4079 17906 4080
rect 17536 4064 17673 4066
rect 16038 4042 16075 4043
rect 15988 4033 16075 4042
rect 15988 4013 16046 4033
rect 16066 4013 16075 4033
rect 15988 4003 16075 4013
rect 16134 4033 16171 4043
rect 16134 4013 16142 4033
rect 16162 4013 16171 4033
rect 17536 4022 17579 4064
rect 17723 4049 17732 4069
rect 17752 4049 17760 4069
rect 17723 4039 17760 4049
rect 17819 4069 17906 4079
rect 17819 4049 17828 4069
rect 17848 4049 17906 4069
rect 17819 4040 17906 4049
rect 17819 4039 17856 4040
rect 15988 4002 16019 4003
rect 15612 3942 15953 3943
rect 16134 3942 16171 4013
rect 17534 4012 17579 4022
rect 17201 4005 17238 4010
rect 17192 4001 17239 4005
rect 17192 3983 17211 4001
rect 17229 3983 17239 4001
rect 17534 3994 17543 4012
rect 17561 3994 17579 4012
rect 17534 3988 17579 3994
rect 17875 3989 17906 4040
rect 17941 4069 17978 4139
rect 18244 4138 18281 4139
rect 18514 4128 18523 4148
rect 18543 4128 18552 4148
rect 18514 4120 18552 4128
rect 18618 4152 18703 4158
rect 18733 4157 18770 4158
rect 18618 4132 18626 4152
rect 18646 4132 18703 4152
rect 18618 4124 18703 4132
rect 18732 4148 18770 4157
rect 18732 4128 18741 4148
rect 18761 4128 18770 4148
rect 18618 4123 18654 4124
rect 18732 4120 18770 4128
rect 18836 4152 18980 4158
rect 18836 4132 18844 4152
rect 18864 4133 18896 4152
rect 18917 4133 18952 4152
rect 18864 4132 18952 4133
rect 18972 4132 18980 4152
rect 18836 4124 18980 4132
rect 18836 4123 18872 4124
rect 18944 4123 18980 4124
rect 19046 4157 19083 4158
rect 19046 4156 19084 4157
rect 19046 4148 19110 4156
rect 19046 4128 19055 4148
rect 19075 4134 19110 4148
rect 19130 4134 19133 4154
rect 19075 4129 19133 4134
rect 19075 4128 19110 4129
rect 18515 4091 18552 4120
rect 18516 4089 18552 4091
rect 18093 4079 18129 4080
rect 17941 4049 17950 4069
rect 17970 4049 17978 4069
rect 17941 4039 17978 4049
rect 18037 4069 18185 4079
rect 18285 4076 18381 4078
rect 18037 4049 18046 4069
rect 18066 4049 18156 4069
rect 18176 4049 18185 4069
rect 18037 4040 18185 4049
rect 18243 4069 18381 4076
rect 18243 4049 18252 4069
rect 18272 4049 18381 4069
rect 18516 4067 18707 4089
rect 18733 4088 18770 4120
rect 19046 4116 19110 4128
rect 19150 4090 19177 4268
rect 19009 4088 19177 4090
rect 18733 4062 19177 4088
rect 18243 4040 18381 4049
rect 18037 4039 18074 4040
rect 17534 3985 17571 3988
rect 17767 3986 17808 3987
rect 15537 3937 15953 3942
rect 15537 3917 15540 3937
rect 15560 3917 15953 3937
rect 15984 3918 16171 3942
rect 16796 3940 16836 3945
rect 17192 3940 17239 3983
rect 17659 3979 17808 3986
rect 17659 3959 17718 3979
rect 17738 3959 17777 3979
rect 17797 3959 17808 3979
rect 17659 3951 17808 3959
rect 17875 3982 18032 3989
rect 17875 3962 17995 3982
rect 18015 3962 18032 3982
rect 17875 3952 18032 3962
rect 17875 3951 17910 3952
rect 16796 3901 17239 3940
rect 17875 3930 17906 3951
rect 18093 3930 18129 4040
rect 18148 4039 18185 4040
rect 18244 4039 18281 4040
rect 18204 3980 18294 3986
rect 18204 3960 18213 3980
rect 18233 3978 18294 3980
rect 18233 3960 18258 3978
rect 18204 3958 18258 3960
rect 18278 3958 18294 3978
rect 18204 3952 18294 3958
rect 17718 3929 17755 3930
rect 15890 3886 15930 3894
rect 15890 3864 15898 3886
rect 15922 3864 15930 3886
rect 15596 3640 15764 3641
rect 15890 3640 15930 3864
rect 16393 3868 16561 3869
rect 16796 3868 16836 3901
rect 17192 3868 17239 3901
rect 17531 3921 17568 3923
rect 17531 3913 17573 3921
rect 17531 3895 17541 3913
rect 17559 3895 17573 3913
rect 17531 3886 17573 3895
rect 17717 3920 17755 3929
rect 17717 3900 17726 3920
rect 17746 3900 17755 3920
rect 17717 3892 17755 3900
rect 17821 3924 17906 3930
rect 17936 3929 17973 3930
rect 17821 3904 17829 3924
rect 17849 3904 17906 3924
rect 17821 3896 17906 3904
rect 17935 3920 17973 3929
rect 17935 3900 17944 3920
rect 17964 3900 17973 3920
rect 17821 3895 17857 3896
rect 17935 3892 17973 3900
rect 18039 3928 18183 3930
rect 18039 3924 18091 3928
rect 18039 3904 18047 3924
rect 18067 3908 18091 3924
rect 18111 3924 18183 3928
rect 18111 3908 18155 3924
rect 18067 3904 18155 3908
rect 18175 3904 18183 3924
rect 18039 3896 18183 3904
rect 18039 3895 18075 3896
rect 18147 3895 18183 3896
rect 18249 3929 18286 3930
rect 18249 3928 18287 3929
rect 18249 3920 18313 3928
rect 18249 3900 18258 3920
rect 18278 3906 18313 3920
rect 18333 3906 18336 3926
rect 18278 3901 18336 3906
rect 18278 3900 18313 3901
rect 16393 3867 16837 3868
rect 16393 3842 16838 3867
rect 16393 3840 16561 3842
rect 16757 3841 16838 3842
rect 17007 3841 17056 3867
rect 17192 3841 17241 3868
rect 16393 3662 16420 3840
rect 16460 3802 16524 3814
rect 16800 3810 16837 3841
rect 17018 3810 17055 3841
rect 17200 3816 17241 3841
rect 17532 3861 17573 3886
rect 17718 3861 17755 3892
rect 17936 3861 17973 3892
rect 18249 3888 18313 3900
rect 18353 3862 18380 4040
rect 17532 3834 17581 3861
rect 17717 3835 17766 3861
rect 17935 3860 18016 3861
rect 18212 3860 18380 3862
rect 17935 3835 18380 3860
rect 17936 3834 18380 3835
rect 16460 3801 16495 3802
rect 16437 3796 16495 3801
rect 16437 3776 16440 3796
rect 16460 3782 16495 3796
rect 16515 3782 16524 3802
rect 16460 3774 16524 3782
rect 16486 3773 16524 3774
rect 16487 3772 16524 3773
rect 16590 3806 16626 3807
rect 16698 3806 16734 3807
rect 16590 3798 16734 3806
rect 16590 3778 16598 3798
rect 16618 3794 16706 3798
rect 16618 3778 16662 3794
rect 16590 3774 16662 3778
rect 16682 3778 16706 3794
rect 16726 3778 16734 3798
rect 16682 3774 16734 3778
rect 16590 3772 16734 3774
rect 16800 3802 16838 3810
rect 16916 3806 16952 3807
rect 16800 3782 16809 3802
rect 16829 3782 16838 3802
rect 16800 3773 16838 3782
rect 16867 3798 16952 3806
rect 16867 3778 16924 3798
rect 16944 3778 16952 3798
rect 16800 3772 16837 3773
rect 16867 3772 16952 3778
rect 17018 3802 17056 3810
rect 17018 3782 17027 3802
rect 17047 3782 17056 3802
rect 17018 3773 17056 3782
rect 17200 3807 17242 3816
rect 17200 3789 17214 3807
rect 17232 3789 17242 3807
rect 17200 3781 17242 3789
rect 17205 3779 17242 3781
rect 17534 3801 17581 3834
rect 17937 3801 17977 3834
rect 18212 3833 18380 3834
rect 18843 3838 18883 4062
rect 19009 4061 19177 4062
rect 18843 3816 18851 3838
rect 18875 3816 18883 3838
rect 18843 3808 18883 3816
rect 17018 3772 17055 3773
rect 16479 3744 16569 3750
rect 16479 3724 16495 3744
rect 16515 3742 16569 3744
rect 16515 3724 16540 3742
rect 16479 3722 16540 3724
rect 16560 3722 16569 3742
rect 16479 3716 16569 3722
rect 16492 3662 16529 3663
rect 16588 3662 16625 3663
rect 16644 3662 16680 3772
rect 16867 3751 16898 3772
rect 17534 3762 17977 3801
rect 16863 3750 16898 3751
rect 16741 3740 16898 3750
rect 16741 3720 16758 3740
rect 16778 3720 16898 3740
rect 16741 3713 16898 3720
rect 16965 3743 17114 3751
rect 16965 3723 16976 3743
rect 16996 3723 17035 3743
rect 17055 3723 17114 3743
rect 16965 3716 17114 3723
rect 17534 3719 17581 3762
rect 17937 3757 17977 3762
rect 18602 3760 18789 3784
rect 18820 3765 19213 3785
rect 19233 3765 19236 3785
rect 18820 3760 19236 3765
rect 16965 3715 17006 3716
rect 17202 3714 17239 3717
rect 16699 3662 16736 3663
rect 16392 3653 16530 3662
rect 15596 3614 16040 3640
rect 15596 3612 15764 3614
rect 15596 3434 15623 3612
rect 15663 3574 15727 3586
rect 16003 3582 16040 3614
rect 16066 3613 16257 3635
rect 16392 3633 16501 3653
rect 16521 3633 16530 3653
rect 16392 3626 16530 3633
rect 16588 3653 16736 3662
rect 16588 3633 16597 3653
rect 16617 3633 16707 3653
rect 16727 3633 16736 3653
rect 16392 3624 16488 3626
rect 16588 3623 16736 3633
rect 16795 3653 16832 3663
rect 16795 3633 16803 3653
rect 16823 3633 16832 3653
rect 16644 3622 16680 3623
rect 16221 3611 16257 3613
rect 16221 3582 16258 3611
rect 15663 3573 15698 3574
rect 15640 3568 15698 3573
rect 15640 3548 15643 3568
rect 15663 3554 15698 3568
rect 15718 3554 15727 3574
rect 15663 3546 15727 3554
rect 15689 3545 15727 3546
rect 15690 3544 15727 3545
rect 15793 3578 15829 3579
rect 15901 3578 15937 3579
rect 15793 3570 15937 3578
rect 15793 3550 15801 3570
rect 15821 3569 15909 3570
rect 15821 3550 15856 3569
rect 15877 3550 15909 3569
rect 15929 3550 15937 3570
rect 15793 3544 15937 3550
rect 16003 3574 16041 3582
rect 16119 3578 16155 3579
rect 16003 3554 16012 3574
rect 16032 3554 16041 3574
rect 16003 3545 16041 3554
rect 16070 3570 16155 3578
rect 16070 3550 16127 3570
rect 16147 3550 16155 3570
rect 16003 3544 16040 3545
rect 16070 3544 16155 3550
rect 16221 3574 16259 3582
rect 16221 3554 16230 3574
rect 16250 3554 16259 3574
rect 16492 3563 16529 3564
rect 16795 3563 16832 3633
rect 16867 3662 16898 3713
rect 17194 3708 17239 3714
rect 17194 3690 17212 3708
rect 17230 3690 17239 3708
rect 17534 3701 17544 3719
rect 17562 3701 17581 3719
rect 17534 3697 17581 3701
rect 17535 3692 17572 3697
rect 17194 3680 17239 3690
rect 18602 3689 18639 3760
rect 18820 3759 19161 3760
rect 18754 3699 18785 3700
rect 16917 3662 16954 3663
rect 16867 3653 16954 3662
rect 16867 3633 16925 3653
rect 16945 3633 16954 3653
rect 16867 3623 16954 3633
rect 17013 3653 17050 3663
rect 17013 3633 17021 3653
rect 17041 3633 17050 3653
rect 17194 3638 17237 3680
rect 18602 3669 18611 3689
rect 18631 3669 18639 3689
rect 18602 3659 18639 3669
rect 18698 3689 18785 3699
rect 18698 3669 18707 3689
rect 18727 3669 18785 3689
rect 18698 3660 18785 3669
rect 18698 3659 18735 3660
rect 17100 3636 17237 3638
rect 16867 3622 16898 3623
rect 17013 3563 17050 3633
rect 16491 3562 16832 3563
rect 16221 3545 16259 3554
rect 16416 3557 16832 3562
rect 16221 3544 16258 3545
rect 15682 3516 15772 3522
rect 15682 3496 15698 3516
rect 15718 3514 15772 3516
rect 15718 3496 15743 3514
rect 15682 3494 15743 3496
rect 15763 3494 15772 3514
rect 15682 3488 15772 3494
rect 15695 3434 15732 3435
rect 15791 3434 15828 3435
rect 15847 3434 15883 3544
rect 16070 3523 16101 3544
rect 16416 3537 16419 3557
rect 16439 3537 16832 3557
rect 17016 3547 17050 3563
rect 17094 3615 17237 3636
rect 17523 3630 17575 3632
rect 16792 3528 16832 3537
rect 17094 3528 17121 3615
rect 17194 3589 17237 3615
rect 17194 3571 17207 3589
rect 17225 3571 17237 3589
rect 17521 3626 17954 3630
rect 17521 3620 17960 3626
rect 17521 3602 17542 3620
rect 17560 3602 17960 3620
rect 18754 3609 18785 3660
rect 18820 3689 18857 3759
rect 19123 3758 19160 3759
rect 18972 3699 19008 3700
rect 18820 3669 18829 3689
rect 18849 3669 18857 3689
rect 18820 3659 18857 3669
rect 18916 3689 19064 3699
rect 19164 3696 19260 3698
rect 18916 3669 18925 3689
rect 18945 3669 19035 3689
rect 19055 3669 19064 3689
rect 18916 3660 19064 3669
rect 19122 3689 19260 3696
rect 19122 3669 19131 3689
rect 19151 3669 19260 3689
rect 19122 3660 19260 3669
rect 18916 3659 18953 3660
rect 18646 3606 18687 3607
rect 17521 3584 17960 3602
rect 17194 3560 17237 3571
rect 16066 3522 16101 3523
rect 15944 3512 16101 3522
rect 15944 3492 15961 3512
rect 15981 3492 16101 3512
rect 15944 3485 16101 3492
rect 16168 3515 16317 3523
rect 16168 3495 16179 3515
rect 16199 3495 16238 3515
rect 16258 3495 16317 3515
rect 16792 3511 17121 3528
rect 16792 3510 16832 3511
rect 16168 3488 16317 3495
rect 17189 3499 17229 3502
rect 17189 3493 17232 3499
rect 16814 3490 17232 3493
rect 16168 3487 16209 3488
rect 15902 3434 15939 3435
rect 15595 3425 15733 3434
rect 15595 3405 15704 3425
rect 15724 3405 15733 3425
rect 15595 3398 15733 3405
rect 15791 3425 15939 3434
rect 15791 3405 15800 3425
rect 15820 3405 15910 3425
rect 15930 3405 15939 3425
rect 15595 3396 15691 3398
rect 15791 3395 15939 3405
rect 15998 3425 16035 3435
rect 15998 3405 16006 3425
rect 16026 3405 16035 3425
rect 15847 3394 15883 3395
rect 15695 3335 15732 3336
rect 15998 3335 16035 3405
rect 16070 3434 16101 3485
rect 16814 3472 17205 3490
rect 17223 3472 17232 3490
rect 16814 3470 17232 3472
rect 16814 3462 16841 3470
rect 17082 3467 17232 3470
rect 16394 3456 16562 3457
rect 16813 3456 16841 3462
rect 16394 3440 16841 3456
rect 17189 3462 17232 3467
rect 16120 3434 16157 3435
rect 16070 3425 16157 3434
rect 16070 3405 16128 3425
rect 16148 3405 16157 3425
rect 16070 3395 16157 3405
rect 16216 3425 16253 3435
rect 16216 3405 16224 3425
rect 16244 3405 16253 3425
rect 16070 3394 16101 3395
rect 15694 3334 16035 3335
rect 16216 3334 16253 3405
rect 15619 3329 16035 3334
rect 15619 3309 15622 3329
rect 15642 3309 16035 3329
rect 16066 3310 16253 3334
rect 16394 3430 16838 3440
rect 16394 3428 16562 3430
rect 15461 3235 15490 3253
rect 16394 3250 16421 3428
rect 16461 3390 16525 3402
rect 16801 3398 16838 3430
rect 16864 3429 17055 3451
rect 17019 3427 17055 3429
rect 17019 3398 17056 3427
rect 17189 3406 17229 3462
rect 16461 3389 16496 3390
rect 16438 3384 16496 3389
rect 16438 3364 16441 3384
rect 16461 3370 16496 3384
rect 16516 3370 16525 3390
rect 16461 3362 16525 3370
rect 16487 3361 16525 3362
rect 16488 3360 16525 3361
rect 16591 3394 16627 3395
rect 16699 3394 16735 3395
rect 16591 3386 16735 3394
rect 16591 3366 16599 3386
rect 16619 3366 16654 3386
rect 16674 3366 16707 3386
rect 16727 3366 16735 3386
rect 16591 3360 16735 3366
rect 16801 3390 16839 3398
rect 16917 3394 16953 3395
rect 16801 3370 16810 3390
rect 16830 3370 16839 3390
rect 16801 3361 16839 3370
rect 16868 3386 16953 3394
rect 16868 3366 16925 3386
rect 16945 3366 16953 3386
rect 16801 3360 16838 3361
rect 16868 3360 16953 3366
rect 17019 3390 17057 3398
rect 17019 3370 17028 3390
rect 17048 3370 17057 3390
rect 17189 3388 17201 3406
rect 17219 3388 17229 3406
rect 17189 3378 17229 3388
rect 17523 3395 17575 3584
rect 17921 3559 17960 3584
rect 18538 3599 18687 3606
rect 18538 3579 18597 3599
rect 18617 3579 18656 3599
rect 18676 3579 18687 3599
rect 18538 3571 18687 3579
rect 18754 3602 18911 3609
rect 18754 3582 18874 3602
rect 18894 3582 18911 3602
rect 18754 3572 18911 3582
rect 18754 3571 18789 3572
rect 17705 3534 17892 3558
rect 17921 3539 18316 3559
rect 18336 3539 18339 3559
rect 18754 3550 18785 3571
rect 18972 3550 19008 3660
rect 19027 3659 19064 3660
rect 19123 3659 19160 3660
rect 19083 3600 19173 3606
rect 19083 3580 19092 3600
rect 19112 3598 19173 3600
rect 19112 3580 19137 3598
rect 19083 3578 19137 3580
rect 19157 3578 19173 3598
rect 19083 3572 19173 3578
rect 18597 3549 18634 3550
rect 17921 3534 18339 3539
rect 18596 3540 18634 3549
rect 17705 3463 17742 3534
rect 17921 3533 18264 3534
rect 17921 3530 17960 3533
rect 18226 3532 18263 3533
rect 17857 3473 17888 3474
rect 17705 3443 17714 3463
rect 17734 3443 17742 3463
rect 17705 3433 17742 3443
rect 17801 3463 17888 3473
rect 17801 3443 17810 3463
rect 17830 3443 17888 3463
rect 17801 3434 17888 3443
rect 17801 3433 17838 3434
rect 17019 3361 17057 3370
rect 17523 3377 17539 3395
rect 17557 3377 17575 3395
rect 17857 3383 17888 3434
rect 17923 3463 17960 3530
rect 18596 3520 18605 3540
rect 18625 3520 18634 3540
rect 18596 3512 18634 3520
rect 18700 3544 18785 3550
rect 18815 3549 18852 3550
rect 18700 3524 18708 3544
rect 18728 3524 18785 3544
rect 18700 3516 18785 3524
rect 18814 3540 18852 3549
rect 18814 3520 18823 3540
rect 18843 3520 18852 3540
rect 18700 3515 18736 3516
rect 18814 3512 18852 3520
rect 18918 3545 19062 3550
rect 18918 3544 18980 3545
rect 18918 3524 18926 3544
rect 18946 3526 18980 3544
rect 19001 3544 19062 3545
rect 19001 3526 19034 3544
rect 18946 3524 19034 3526
rect 19054 3524 19062 3544
rect 18918 3516 19062 3524
rect 18918 3515 18954 3516
rect 19026 3515 19062 3516
rect 19128 3549 19165 3550
rect 19128 3548 19166 3549
rect 19128 3540 19192 3548
rect 19128 3520 19137 3540
rect 19157 3526 19192 3540
rect 19212 3526 19215 3546
rect 19157 3521 19215 3526
rect 19157 3520 19192 3521
rect 18597 3483 18634 3512
rect 18598 3481 18634 3483
rect 18075 3473 18111 3474
rect 17923 3443 17932 3463
rect 17952 3443 17960 3463
rect 17923 3433 17960 3443
rect 18019 3463 18167 3473
rect 18267 3470 18363 3472
rect 18019 3443 18028 3463
rect 18048 3443 18138 3463
rect 18158 3443 18167 3463
rect 18019 3434 18167 3443
rect 18225 3463 18363 3470
rect 18225 3443 18234 3463
rect 18254 3443 18363 3463
rect 18598 3459 18789 3481
rect 18815 3480 18852 3512
rect 19128 3508 19192 3520
rect 19232 3482 19259 3660
rect 19091 3480 19259 3482
rect 18815 3466 19259 3480
rect 18815 3454 19262 3466
rect 18858 3452 18891 3454
rect 18225 3434 18363 3443
rect 18019 3433 18056 3434
rect 17749 3380 17790 3381
rect 17019 3360 17056 3361
rect 16480 3332 16570 3338
rect 16480 3312 16496 3332
rect 16516 3330 16570 3332
rect 16516 3312 16541 3330
rect 16480 3310 16541 3312
rect 16561 3310 16570 3330
rect 16480 3304 16570 3310
rect 16493 3250 16530 3251
rect 16589 3250 16626 3251
rect 16645 3250 16681 3360
rect 16868 3339 16899 3360
rect 17523 3359 17575 3377
rect 17641 3373 17790 3380
rect 17641 3353 17700 3373
rect 17720 3353 17759 3373
rect 17779 3353 17790 3373
rect 17641 3345 17790 3353
rect 17857 3376 18014 3383
rect 17857 3356 17977 3376
rect 17997 3356 18014 3376
rect 17857 3346 18014 3356
rect 17857 3345 17892 3346
rect 16864 3338 16899 3339
rect 16742 3328 16899 3338
rect 16742 3308 16759 3328
rect 16779 3308 16899 3328
rect 16742 3301 16899 3308
rect 16966 3331 17115 3339
rect 16966 3311 16977 3331
rect 16997 3311 17036 3331
rect 17056 3311 17115 3331
rect 16966 3304 17115 3311
rect 17181 3307 17233 3325
rect 17857 3324 17888 3345
rect 18075 3324 18111 3434
rect 18130 3433 18167 3434
rect 18226 3433 18263 3434
rect 18186 3374 18276 3380
rect 18186 3354 18195 3374
rect 18215 3372 18276 3374
rect 18215 3354 18240 3372
rect 18186 3352 18240 3354
rect 18260 3352 18276 3372
rect 18186 3346 18276 3352
rect 17700 3323 17737 3324
rect 16966 3303 17007 3304
rect 16700 3250 16737 3251
rect 15431 3233 15490 3235
rect 16393 3241 16531 3250
rect 15431 3232 15599 3233
rect 15725 3232 15765 3234
rect 15431 3206 15875 3232
rect 15431 3204 15599 3206
rect 15431 3202 15512 3204
rect 15431 3026 15458 3202
rect 15498 3166 15562 3178
rect 15838 3174 15875 3206
rect 15901 3205 16092 3227
rect 16393 3221 16502 3241
rect 16522 3221 16531 3241
rect 16393 3214 16531 3221
rect 16589 3241 16737 3250
rect 16589 3221 16598 3241
rect 16618 3221 16708 3241
rect 16728 3221 16737 3241
rect 16393 3212 16489 3214
rect 16589 3211 16737 3221
rect 16796 3241 16833 3251
rect 16796 3221 16804 3241
rect 16824 3221 16833 3241
rect 16645 3210 16681 3211
rect 16056 3203 16092 3205
rect 16056 3174 16093 3203
rect 15498 3165 15533 3166
rect 15475 3160 15533 3165
rect 15475 3140 15478 3160
rect 15498 3146 15533 3160
rect 15553 3146 15562 3166
rect 15498 3138 15562 3146
rect 15524 3137 15562 3138
rect 15525 3136 15562 3137
rect 15628 3170 15664 3171
rect 15736 3170 15772 3171
rect 15628 3162 15772 3170
rect 15628 3142 15636 3162
rect 15656 3161 15744 3162
rect 15656 3143 15691 3161
rect 15709 3143 15744 3161
rect 15656 3142 15744 3143
rect 15764 3142 15772 3162
rect 15628 3136 15772 3142
rect 15838 3166 15876 3174
rect 15954 3170 15990 3171
rect 15838 3146 15847 3166
rect 15867 3146 15876 3166
rect 15838 3137 15876 3146
rect 15905 3162 15990 3170
rect 15905 3142 15962 3162
rect 15982 3142 15990 3162
rect 15838 3136 15875 3137
rect 15905 3136 15990 3142
rect 16056 3166 16094 3174
rect 16056 3146 16065 3166
rect 16085 3146 16094 3166
rect 16796 3154 16833 3221
rect 16868 3250 16899 3301
rect 17181 3289 17199 3307
rect 17217 3289 17233 3307
rect 17699 3314 17737 3323
rect 16918 3250 16955 3251
rect 16868 3241 16955 3250
rect 16868 3221 16926 3241
rect 16946 3221 16955 3241
rect 16868 3211 16955 3221
rect 17014 3241 17051 3251
rect 17014 3221 17022 3241
rect 17042 3221 17051 3241
rect 16868 3210 16899 3211
rect 16493 3151 16530 3152
rect 16796 3151 16835 3154
rect 16492 3150 16835 3151
rect 17014 3150 17051 3221
rect 16056 3137 16094 3146
rect 16417 3145 16835 3150
rect 16056 3136 16093 3137
rect 15517 3108 15607 3114
rect 15517 3088 15533 3108
rect 15553 3106 15607 3108
rect 15553 3088 15578 3106
rect 15517 3086 15578 3088
rect 15598 3086 15607 3106
rect 15517 3080 15607 3086
rect 15530 3026 15567 3027
rect 15626 3026 15663 3027
rect 15682 3026 15718 3136
rect 15905 3115 15936 3136
rect 16417 3125 16420 3145
rect 16440 3125 16835 3145
rect 16864 3126 17051 3150
rect 15901 3114 15936 3115
rect 15779 3104 15936 3114
rect 15779 3084 15796 3104
rect 15816 3084 15936 3104
rect 15779 3077 15936 3084
rect 16003 3107 16152 3115
rect 16003 3087 16014 3107
rect 16034 3087 16073 3107
rect 16093 3087 16152 3107
rect 16003 3080 16152 3087
rect 16796 3100 16835 3125
rect 17181 3100 17233 3289
rect 17527 3296 17567 3306
rect 17527 3278 17537 3296
rect 17555 3278 17567 3296
rect 17699 3294 17708 3314
rect 17728 3294 17737 3314
rect 17699 3286 17737 3294
rect 17803 3318 17888 3324
rect 17918 3323 17955 3324
rect 17803 3298 17811 3318
rect 17831 3298 17888 3318
rect 17803 3290 17888 3298
rect 17917 3314 17955 3323
rect 17917 3294 17926 3314
rect 17946 3294 17955 3314
rect 17803 3289 17839 3290
rect 17917 3286 17955 3294
rect 18021 3318 18165 3324
rect 18021 3298 18029 3318
rect 18049 3298 18082 3318
rect 18102 3298 18137 3318
rect 18157 3298 18165 3318
rect 18021 3290 18165 3298
rect 18021 3289 18057 3290
rect 18129 3289 18165 3290
rect 18231 3323 18268 3324
rect 18231 3322 18269 3323
rect 18231 3314 18295 3322
rect 18231 3294 18240 3314
rect 18260 3300 18295 3314
rect 18315 3300 18318 3320
rect 18260 3295 18318 3300
rect 18260 3294 18295 3295
rect 17527 3222 17567 3278
rect 17700 3257 17737 3286
rect 17701 3255 17737 3257
rect 17701 3233 17892 3255
rect 17918 3254 17955 3286
rect 18231 3282 18295 3294
rect 18335 3256 18362 3434
rect 19220 3409 19262 3454
rect 18194 3254 18362 3256
rect 17918 3244 18362 3254
rect 18503 3350 18690 3374
rect 18721 3355 19114 3375
rect 19134 3355 19137 3375
rect 18721 3350 19137 3355
rect 18503 3279 18540 3350
rect 18721 3349 19062 3350
rect 18655 3289 18686 3290
rect 18503 3259 18512 3279
rect 18532 3259 18540 3279
rect 18503 3249 18540 3259
rect 18599 3279 18686 3289
rect 18599 3259 18608 3279
rect 18628 3259 18686 3279
rect 18599 3250 18686 3259
rect 18599 3249 18636 3250
rect 17524 3217 17567 3222
rect 17915 3228 18362 3244
rect 17915 3222 17943 3228
rect 18194 3227 18362 3228
rect 17524 3214 17674 3217
rect 17915 3214 17942 3222
rect 17524 3212 17942 3214
rect 17524 3194 17533 3212
rect 17551 3194 17942 3212
rect 18655 3199 18686 3250
rect 18721 3279 18758 3349
rect 19024 3348 19061 3349
rect 18873 3289 18909 3290
rect 18721 3259 18730 3279
rect 18750 3259 18758 3279
rect 18721 3249 18758 3259
rect 18817 3279 18965 3289
rect 19065 3286 19161 3288
rect 18817 3259 18826 3279
rect 18846 3259 18936 3279
rect 18956 3259 18965 3279
rect 18817 3250 18965 3259
rect 19023 3279 19161 3286
rect 19023 3259 19032 3279
rect 19052 3259 19161 3279
rect 19023 3250 19161 3259
rect 18817 3249 18854 3250
rect 18547 3196 18588 3197
rect 17524 3191 17942 3194
rect 17524 3185 17567 3191
rect 17527 3182 17567 3185
rect 18442 3189 18588 3196
rect 17924 3173 17964 3174
rect 17635 3156 17964 3173
rect 18442 3169 18498 3189
rect 18518 3169 18557 3189
rect 18577 3169 18588 3189
rect 18442 3161 18588 3169
rect 18655 3192 18812 3199
rect 18655 3172 18775 3192
rect 18795 3172 18812 3192
rect 18655 3162 18812 3172
rect 18655 3161 18690 3162
rect 17519 3113 17562 3124
rect 16796 3082 17235 3100
rect 16003 3079 16044 3080
rect 15737 3026 15774 3027
rect 15430 3017 15568 3026
rect 15430 2997 15539 3017
rect 15559 2997 15568 3017
rect 15430 2990 15568 2997
rect 15626 3017 15774 3026
rect 15626 2997 15635 3017
rect 15655 2997 15745 3017
rect 15765 2997 15774 3017
rect 15430 2988 15526 2990
rect 15626 2987 15774 2997
rect 15833 3017 15870 3027
rect 15833 2997 15841 3017
rect 15861 2997 15870 3017
rect 15682 2986 15718 2987
rect 15530 2927 15567 2928
rect 15833 2927 15870 2997
rect 15905 3026 15936 3077
rect 16796 3064 17196 3082
rect 17214 3064 17235 3082
rect 16796 3058 17235 3064
rect 16802 3054 17235 3058
rect 17519 3095 17531 3113
rect 17549 3095 17562 3113
rect 17519 3069 17562 3095
rect 17635 3069 17662 3156
rect 17924 3147 17964 3156
rect 17181 3052 17233 3054
rect 17519 3048 17662 3069
rect 17706 3121 17740 3137
rect 17924 3127 18317 3147
rect 18337 3127 18340 3147
rect 18655 3140 18686 3161
rect 18873 3140 18909 3250
rect 18928 3249 18965 3250
rect 19024 3249 19061 3250
rect 18984 3190 19074 3196
rect 18984 3170 18993 3190
rect 19013 3188 19074 3190
rect 19013 3170 19038 3188
rect 18984 3168 19038 3170
rect 19058 3168 19074 3188
rect 18984 3162 19074 3168
rect 18498 3139 18535 3140
rect 17924 3122 18340 3127
rect 18497 3130 18535 3139
rect 17924 3121 18265 3122
rect 17706 3051 17743 3121
rect 17858 3061 17889 3062
rect 17519 3046 17656 3048
rect 15955 3026 15992 3027
rect 15905 3017 15992 3026
rect 15905 2997 15963 3017
rect 15983 2997 15992 3017
rect 15905 2987 15992 2997
rect 16051 3017 16088 3027
rect 16051 2997 16059 3017
rect 16079 2997 16088 3017
rect 17519 3004 17562 3046
rect 17706 3031 17715 3051
rect 17735 3031 17743 3051
rect 17706 3021 17743 3031
rect 17802 3051 17889 3061
rect 17802 3031 17811 3051
rect 17831 3031 17889 3051
rect 17802 3022 17889 3031
rect 17802 3021 17839 3022
rect 15905 2986 15936 2987
rect 15529 2926 15870 2927
rect 16051 2926 16088 2997
rect 17517 2994 17562 3004
rect 17184 2987 17221 2992
rect 15454 2921 15870 2926
rect 15454 2901 15457 2921
rect 15477 2901 15870 2921
rect 15901 2902 16088 2926
rect 17175 2983 17222 2987
rect 17175 2965 17194 2983
rect 17212 2965 17222 2983
rect 17517 2976 17526 2994
rect 17544 2976 17562 2994
rect 17517 2970 17562 2976
rect 17858 2971 17889 3022
rect 17924 3051 17961 3121
rect 18227 3120 18264 3121
rect 18497 3110 18506 3130
rect 18526 3110 18535 3130
rect 18497 3102 18535 3110
rect 18601 3134 18686 3140
rect 18716 3139 18753 3140
rect 18601 3114 18609 3134
rect 18629 3114 18686 3134
rect 18601 3106 18686 3114
rect 18715 3130 18753 3139
rect 18715 3110 18724 3130
rect 18744 3110 18753 3130
rect 18601 3105 18637 3106
rect 18715 3102 18753 3110
rect 18819 3134 18963 3140
rect 18819 3114 18827 3134
rect 18847 3131 18935 3134
rect 18847 3114 18882 3131
rect 18819 3113 18882 3114
rect 18901 3114 18935 3131
rect 18955 3114 18963 3134
rect 18901 3113 18963 3114
rect 18819 3106 18963 3113
rect 18819 3105 18855 3106
rect 18927 3105 18963 3106
rect 19029 3139 19066 3140
rect 19029 3138 19067 3139
rect 19089 3138 19116 3142
rect 19029 3136 19116 3138
rect 19029 3130 19093 3136
rect 19029 3110 19038 3130
rect 19058 3116 19093 3130
rect 19113 3116 19116 3136
rect 19058 3111 19116 3116
rect 19058 3110 19093 3111
rect 18498 3073 18535 3102
rect 18499 3071 18535 3073
rect 18076 3061 18112 3062
rect 17924 3031 17933 3051
rect 17953 3031 17961 3051
rect 17924 3021 17961 3031
rect 18020 3051 18168 3061
rect 18268 3058 18364 3060
rect 18020 3031 18029 3051
rect 18049 3031 18139 3051
rect 18159 3031 18168 3051
rect 18020 3022 18168 3031
rect 18226 3051 18364 3058
rect 18226 3031 18235 3051
rect 18255 3031 18364 3051
rect 18499 3049 18690 3071
rect 18716 3070 18753 3102
rect 19029 3098 19093 3110
rect 19133 3072 19160 3250
rect 18992 3070 19160 3072
rect 18716 3044 19160 3070
rect 18226 3022 18364 3031
rect 18020 3021 18057 3022
rect 17517 2967 17554 2970
rect 17750 2968 17791 2969
rect 17175 2917 17222 2965
rect 17642 2961 17791 2968
rect 17642 2941 17701 2961
rect 17721 2941 17760 2961
rect 17780 2941 17791 2961
rect 17642 2933 17791 2941
rect 17858 2964 18015 2971
rect 17858 2944 17978 2964
rect 17998 2944 18015 2964
rect 17858 2934 18015 2944
rect 17858 2933 17893 2934
rect 16799 2914 17222 2917
rect 15674 2900 15739 2901
rect 16777 2884 17222 2914
rect 17858 2912 17889 2933
rect 18076 2912 18112 3022
rect 18131 3021 18168 3022
rect 18227 3021 18264 3022
rect 18187 2962 18277 2968
rect 18187 2942 18196 2962
rect 18216 2960 18277 2962
rect 18216 2942 18241 2960
rect 18187 2940 18241 2942
rect 18261 2940 18277 2960
rect 18187 2934 18277 2940
rect 17701 2911 17738 2912
rect 15870 2868 15910 2876
rect 15870 2846 15878 2868
rect 15902 2846 15910 2868
rect 15475 2617 15512 2623
rect 15475 2598 15483 2617
rect 15504 2598 15512 2617
rect 15475 2590 15512 2598
rect 15175 2469 15182 2491
rect 15206 2469 15214 2491
rect 15175 2463 15214 2469
rect 14705 2458 14745 2460
rect 14871 2459 15039 2460
rect 14973 2458 15010 2459
rect 13939 2442 14077 2451
rect 13733 2441 13770 2442
rect 13463 2388 13504 2389
rect 13237 2367 13289 2385
rect 13355 2381 13504 2388
rect 12805 2347 12845 2357
rect 13355 2361 13414 2381
rect 13434 2361 13473 2381
rect 13493 2361 13504 2381
rect 13355 2353 13504 2361
rect 13571 2384 13728 2391
rect 13571 2364 13691 2384
rect 13711 2364 13728 2384
rect 13571 2354 13728 2364
rect 13571 2353 13606 2354
rect 12635 2330 12673 2339
rect 13571 2332 13602 2353
rect 13789 2332 13825 2442
rect 13844 2441 13881 2442
rect 13940 2441 13977 2442
rect 13900 2382 13990 2388
rect 13900 2362 13909 2382
rect 13929 2380 13990 2382
rect 13929 2362 13954 2380
rect 13900 2360 13954 2362
rect 13974 2360 13990 2380
rect 13900 2354 13990 2360
rect 13414 2331 13451 2332
rect 12635 2329 12672 2330
rect 12096 2301 12186 2307
rect 12096 2281 12112 2301
rect 12132 2299 12186 2301
rect 12132 2281 12157 2299
rect 12096 2279 12157 2281
rect 12177 2279 12186 2299
rect 12096 2273 12186 2279
rect 12109 2219 12146 2220
rect 12205 2219 12242 2220
rect 12261 2219 12297 2329
rect 12484 2308 12515 2329
rect 13413 2322 13451 2331
rect 12480 2307 12515 2308
rect 12358 2297 12515 2307
rect 12358 2277 12375 2297
rect 12395 2277 12515 2297
rect 12358 2270 12515 2277
rect 12582 2300 12731 2308
rect 12582 2280 12593 2300
rect 12613 2280 12652 2300
rect 12672 2280 12731 2300
rect 13241 2304 13281 2314
rect 12582 2273 12731 2280
rect 12797 2276 12849 2294
rect 12582 2272 12623 2273
rect 12316 2219 12353 2220
rect 12009 2210 12147 2219
rect 11481 2199 11514 2201
rect 11110 2187 11557 2199
rect 10342 2065 10510 2067
rect 10066 2039 10510 2065
rect 9576 2017 9714 2026
rect 9370 2016 9407 2017
rect 8867 1962 8904 1965
rect 9100 1963 9141 1964
rect 7210 1941 7241 1942
rect 6834 1881 7175 1882
rect 7356 1881 7393 1952
rect 8992 1956 9141 1963
rect 8423 1944 8460 1949
rect 8414 1940 8461 1944
rect 8414 1922 8433 1940
rect 8451 1922 8461 1940
rect 8992 1936 9051 1956
rect 9071 1936 9110 1956
rect 9130 1936 9141 1956
rect 8992 1928 9141 1936
rect 9208 1959 9365 1966
rect 9208 1939 9328 1959
rect 9348 1939 9365 1959
rect 9208 1929 9365 1939
rect 9208 1928 9243 1929
rect 6759 1876 7175 1881
rect 6759 1856 6762 1876
rect 6782 1856 7175 1876
rect 7206 1857 7393 1881
rect 8018 1879 8058 1884
rect 8414 1879 8461 1922
rect 9208 1907 9239 1928
rect 9426 1907 9462 2017
rect 9481 2016 9518 2017
rect 9577 2016 9614 2017
rect 9537 1957 9627 1963
rect 9537 1937 9546 1957
rect 9566 1955 9627 1957
rect 9566 1937 9591 1955
rect 9537 1935 9591 1937
rect 9611 1935 9627 1955
rect 9537 1929 9627 1935
rect 9051 1906 9088 1907
rect 8018 1840 8461 1879
rect 8864 1898 8901 1900
rect 8864 1890 8906 1898
rect 8864 1872 8874 1890
rect 8892 1872 8906 1890
rect 8864 1863 8906 1872
rect 9050 1897 9088 1906
rect 9050 1877 9059 1897
rect 9079 1877 9088 1897
rect 9050 1869 9088 1877
rect 9154 1901 9239 1907
rect 9269 1906 9306 1907
rect 9154 1881 9162 1901
rect 9182 1881 9239 1901
rect 9154 1873 9239 1881
rect 9268 1897 9306 1906
rect 9268 1877 9277 1897
rect 9297 1877 9306 1897
rect 9154 1872 9190 1873
rect 9268 1869 9306 1877
rect 9372 1905 9516 1907
rect 9372 1901 9424 1905
rect 9372 1881 9380 1901
rect 9400 1885 9424 1901
rect 9444 1901 9516 1905
rect 9444 1885 9488 1901
rect 9400 1881 9488 1885
rect 9508 1881 9516 1901
rect 9372 1873 9516 1881
rect 9372 1872 9408 1873
rect 9480 1872 9516 1873
rect 9582 1906 9619 1907
rect 9582 1905 9620 1906
rect 9582 1897 9646 1905
rect 9582 1877 9591 1897
rect 9611 1883 9646 1897
rect 9666 1883 9669 1903
rect 9611 1878 9669 1883
rect 9611 1877 9646 1878
rect 5799 1781 5807 1803
rect 5831 1781 5839 1803
rect 5799 1773 5839 1781
rect 7112 1825 7152 1833
rect 7112 1803 7120 1825
rect 7144 1803 7152 1825
rect 3318 1727 3353 1728
rect 3295 1722 3353 1727
rect 3295 1702 3298 1722
rect 3318 1708 3353 1722
rect 3373 1708 3382 1728
rect 3318 1700 3382 1708
rect 3344 1699 3382 1700
rect 3345 1698 3382 1699
rect 3448 1732 3484 1733
rect 3556 1732 3592 1733
rect 3448 1724 3592 1732
rect 3448 1704 3456 1724
rect 3476 1720 3564 1724
rect 3476 1704 3520 1720
rect 3448 1700 3520 1704
rect 3540 1704 3564 1720
rect 3584 1704 3592 1724
rect 3540 1700 3592 1704
rect 3448 1698 3592 1700
rect 3658 1728 3696 1736
rect 3774 1732 3810 1733
rect 3658 1708 3667 1728
rect 3687 1708 3696 1728
rect 3658 1699 3696 1708
rect 3725 1724 3810 1732
rect 3725 1704 3782 1724
rect 3802 1704 3810 1724
rect 3658 1698 3695 1699
rect 3725 1698 3810 1704
rect 3876 1728 3914 1736
rect 3876 1708 3885 1728
rect 3905 1708 3914 1728
rect 3876 1699 3914 1708
rect 4058 1733 4100 1742
rect 4058 1715 4072 1733
rect 4090 1715 4100 1733
rect 4058 1707 4100 1715
rect 4063 1705 4100 1707
rect 4490 1727 4933 1766
rect 3876 1698 3913 1699
rect 3337 1670 3427 1676
rect 3337 1650 3353 1670
rect 3373 1668 3427 1670
rect 3373 1650 3398 1668
rect 3337 1648 3398 1650
rect 3418 1648 3427 1668
rect 3337 1642 3427 1648
rect 3350 1588 3387 1589
rect 3446 1588 3483 1589
rect 3502 1588 3538 1698
rect 3725 1677 3756 1698
rect 4490 1684 4537 1727
rect 4893 1722 4933 1727
rect 5558 1725 5745 1749
rect 5776 1730 6169 1750
rect 6189 1730 6192 1750
rect 5776 1725 6192 1730
rect 3721 1676 3756 1677
rect 3599 1666 3756 1676
rect 3599 1646 3616 1666
rect 3636 1646 3756 1666
rect 3599 1639 3756 1646
rect 3823 1669 3972 1677
rect 3823 1649 3834 1669
rect 3854 1649 3893 1669
rect 3913 1649 3972 1669
rect 4490 1666 4500 1684
rect 4518 1666 4537 1684
rect 4490 1662 4537 1666
rect 4491 1657 4528 1662
rect 3823 1642 3972 1649
rect 5558 1654 5595 1725
rect 5776 1724 6117 1725
rect 5710 1664 5741 1665
rect 3823 1641 3864 1642
rect 4060 1640 4097 1643
rect 3557 1588 3594 1589
rect 3250 1579 3388 1588
rect 2454 1540 2898 1566
rect 2454 1538 2622 1540
rect 1407 1406 1854 1418
rect 1450 1404 1483 1406
rect 817 1386 955 1395
rect 611 1385 648 1386
rect 341 1332 382 1333
rect 115 1311 167 1329
rect 233 1325 382 1332
rect 233 1305 292 1325
rect 312 1305 351 1325
rect 371 1305 382 1325
rect 233 1297 382 1305
rect 449 1328 606 1335
rect 449 1308 569 1328
rect 589 1308 606 1328
rect 449 1298 606 1308
rect 449 1297 484 1298
rect 449 1276 480 1297
rect 667 1276 703 1386
rect 722 1385 759 1386
rect 818 1385 855 1386
rect 778 1326 868 1332
rect 778 1306 787 1326
rect 807 1324 868 1326
rect 807 1306 832 1324
rect 778 1304 832 1306
rect 852 1304 868 1324
rect 778 1298 868 1304
rect 292 1275 329 1276
rect 291 1266 329 1275
rect 119 1248 159 1258
rect 119 1230 129 1248
rect 147 1230 159 1248
rect 291 1246 300 1266
rect 320 1246 329 1266
rect 291 1238 329 1246
rect 395 1270 480 1276
rect 510 1275 547 1276
rect 395 1250 403 1270
rect 423 1250 480 1270
rect 395 1242 480 1250
rect 509 1266 547 1275
rect 509 1246 518 1266
rect 538 1246 547 1266
rect 395 1241 431 1242
rect 509 1238 547 1246
rect 613 1270 757 1276
rect 613 1250 621 1270
rect 641 1250 674 1270
rect 694 1250 729 1270
rect 749 1250 757 1270
rect 613 1242 757 1250
rect 613 1241 649 1242
rect 721 1241 757 1242
rect 823 1275 860 1276
rect 823 1274 861 1275
rect 823 1266 887 1274
rect 823 1246 832 1266
rect 852 1252 887 1266
rect 907 1252 910 1272
rect 852 1247 910 1252
rect 852 1246 887 1247
rect 119 1174 159 1230
rect 292 1209 329 1238
rect 293 1207 329 1209
rect 293 1185 484 1207
rect 510 1206 547 1238
rect 823 1234 887 1246
rect 927 1208 954 1386
rect 1812 1361 1854 1406
rect 786 1206 954 1208
rect 510 1196 954 1206
rect 1095 1302 1282 1326
rect 1313 1307 1706 1327
rect 1726 1307 1729 1327
rect 1313 1302 1729 1307
rect 1095 1231 1132 1302
rect 1313 1301 1654 1302
rect 1247 1241 1278 1242
rect 1095 1211 1104 1231
rect 1124 1211 1132 1231
rect 1095 1201 1132 1211
rect 1191 1231 1278 1241
rect 1191 1211 1200 1231
rect 1220 1211 1278 1231
rect 1191 1202 1278 1211
rect 1191 1201 1228 1202
rect 116 1169 159 1174
rect 507 1180 954 1196
rect 507 1174 535 1180
rect 786 1179 954 1180
rect 116 1166 266 1169
rect 507 1166 534 1174
rect 116 1164 534 1166
rect 116 1146 125 1164
rect 143 1146 534 1164
rect 1247 1151 1278 1202
rect 1313 1231 1350 1301
rect 1616 1300 1653 1301
rect 1465 1241 1501 1242
rect 1313 1211 1322 1231
rect 1342 1211 1350 1231
rect 1313 1201 1350 1211
rect 1409 1231 1557 1241
rect 1657 1238 1753 1240
rect 1409 1211 1418 1231
rect 1438 1211 1528 1231
rect 1548 1211 1557 1231
rect 1409 1202 1557 1211
rect 1615 1231 1753 1238
rect 1615 1211 1624 1231
rect 1644 1211 1753 1231
rect 1615 1202 1753 1211
rect 1409 1201 1446 1202
rect 1139 1148 1180 1149
rect 116 1143 534 1146
rect 116 1137 159 1143
rect 119 1134 159 1137
rect 1034 1141 1180 1148
rect 516 1125 556 1126
rect 227 1108 556 1125
rect 1034 1121 1090 1141
rect 1110 1121 1149 1141
rect 1169 1121 1180 1141
rect 1034 1113 1180 1121
rect 1247 1144 1404 1151
rect 1247 1124 1367 1144
rect 1387 1124 1404 1144
rect 1247 1114 1404 1124
rect 1247 1113 1282 1114
rect 111 1065 154 1076
rect 111 1047 123 1065
rect 141 1047 154 1065
rect 111 1021 154 1047
rect 227 1021 254 1108
rect 516 1099 556 1108
rect 111 1000 254 1021
rect 298 1073 332 1089
rect 516 1079 909 1099
rect 929 1079 932 1099
rect 1247 1092 1278 1113
rect 1465 1092 1501 1202
rect 1520 1201 1557 1202
rect 1616 1201 1653 1202
rect 1576 1142 1666 1148
rect 1576 1122 1585 1142
rect 1605 1140 1666 1142
rect 1605 1122 1630 1140
rect 1576 1120 1630 1122
rect 1650 1120 1666 1140
rect 1576 1114 1666 1120
rect 1090 1091 1127 1092
rect 516 1074 932 1079
rect 1089 1082 1127 1091
rect 516 1073 857 1074
rect 298 1003 335 1073
rect 450 1013 481 1014
rect 111 998 248 1000
rect 111 956 154 998
rect 298 983 307 1003
rect 327 983 335 1003
rect 298 973 335 983
rect 394 1003 481 1013
rect 394 983 403 1003
rect 423 983 481 1003
rect 394 974 481 983
rect 394 973 431 974
rect 109 946 154 956
rect 109 928 118 946
rect 136 928 154 946
rect 109 922 154 928
rect 450 923 481 974
rect 516 1003 553 1073
rect 819 1072 856 1073
rect 1089 1062 1098 1082
rect 1118 1062 1127 1082
rect 1089 1054 1127 1062
rect 1193 1086 1278 1092
rect 1308 1091 1345 1092
rect 1193 1066 1201 1086
rect 1221 1066 1278 1086
rect 1193 1058 1278 1066
rect 1307 1082 1345 1091
rect 1307 1062 1316 1082
rect 1336 1062 1345 1082
rect 1193 1057 1229 1058
rect 1307 1054 1345 1062
rect 1411 1086 1555 1092
rect 1411 1066 1419 1086
rect 1439 1083 1527 1086
rect 1439 1066 1474 1083
rect 1411 1065 1474 1066
rect 1493 1066 1527 1083
rect 1547 1066 1555 1086
rect 1493 1065 1555 1066
rect 1411 1058 1555 1065
rect 1411 1057 1447 1058
rect 1519 1057 1555 1058
rect 1621 1091 1658 1092
rect 1621 1090 1659 1091
rect 1681 1090 1708 1094
rect 1621 1088 1708 1090
rect 1621 1082 1685 1088
rect 1621 1062 1630 1082
rect 1650 1068 1685 1082
rect 1705 1068 1708 1088
rect 1650 1063 1708 1068
rect 1650 1062 1685 1063
rect 1090 1025 1127 1054
rect 1091 1023 1127 1025
rect 668 1013 704 1014
rect 516 983 525 1003
rect 545 983 553 1003
rect 516 973 553 983
rect 612 1003 760 1013
rect 860 1010 956 1012
rect 612 983 621 1003
rect 641 983 731 1003
rect 751 983 760 1003
rect 612 974 760 983
rect 818 1003 956 1010
rect 818 983 827 1003
rect 847 983 956 1003
rect 1091 1001 1282 1023
rect 1308 1022 1345 1054
rect 1621 1050 1685 1062
rect 1725 1024 1752 1202
rect 1584 1022 1752 1024
rect 1308 996 1752 1022
rect 818 974 956 983
rect 612 973 649 974
rect 109 919 146 922
rect 342 920 383 921
rect 234 913 383 920
rect 234 893 293 913
rect 313 893 352 913
rect 372 893 383 913
rect 234 885 383 893
rect 450 916 607 923
rect 450 896 570 916
rect 590 896 607 916
rect 450 886 607 896
rect 450 885 485 886
rect 450 864 481 885
rect 668 864 704 974
rect 723 973 760 974
rect 819 973 856 974
rect 779 914 869 920
rect 779 894 788 914
rect 808 912 869 914
rect 808 894 833 912
rect 779 892 833 894
rect 853 892 869 912
rect 779 886 869 892
rect 293 863 330 864
rect 106 855 143 857
rect 106 847 148 855
rect 106 829 116 847
rect 134 829 148 847
rect 106 820 148 829
rect 292 854 330 863
rect 292 834 301 854
rect 321 834 330 854
rect 292 826 330 834
rect 396 858 481 864
rect 511 863 548 864
rect 396 838 404 858
rect 424 838 481 858
rect 396 830 481 838
rect 510 854 548 863
rect 510 834 519 854
rect 539 834 548 854
rect 396 829 432 830
rect 510 826 548 834
rect 614 862 758 864
rect 614 858 666 862
rect 614 838 622 858
rect 642 842 666 858
rect 686 858 758 862
rect 686 842 730 858
rect 642 838 730 842
rect 750 838 758 858
rect 614 830 758 838
rect 614 829 650 830
rect 722 829 758 830
rect 824 863 861 864
rect 824 862 862 863
rect 824 854 888 862
rect 824 834 833 854
rect 853 840 888 854
rect 908 840 911 860
rect 853 835 911 840
rect 853 834 888 835
rect 107 795 148 820
rect 293 795 330 826
rect 511 804 548 826
rect 824 822 888 834
rect 506 795 548 804
rect 928 796 955 974
rect 107 783 152 795
rect 103 725 152 783
rect 293 769 355 795
rect 506 794 591 795
rect 787 794 955 796
rect 506 768 955 794
rect 506 725 545 768
rect 787 767 955 768
rect 1418 772 1458 996
rect 1584 995 1752 996
rect 1816 1028 1849 1361
rect 2454 1360 2481 1538
rect 2521 1500 2585 1512
rect 2861 1508 2898 1540
rect 2924 1539 3115 1561
rect 3250 1559 3359 1579
rect 3379 1559 3388 1579
rect 3250 1552 3388 1559
rect 3446 1579 3594 1588
rect 3446 1559 3455 1579
rect 3475 1559 3565 1579
rect 3585 1559 3594 1579
rect 3250 1550 3346 1552
rect 3446 1549 3594 1559
rect 3653 1579 3690 1589
rect 3653 1559 3661 1579
rect 3681 1559 3690 1579
rect 3502 1548 3538 1549
rect 3079 1537 3115 1539
rect 3079 1508 3116 1537
rect 2521 1499 2556 1500
rect 2498 1494 2556 1499
rect 2498 1474 2501 1494
rect 2521 1480 2556 1494
rect 2576 1480 2585 1500
rect 2521 1472 2585 1480
rect 2547 1471 2585 1472
rect 2548 1470 2585 1471
rect 2651 1504 2687 1505
rect 2759 1504 2795 1505
rect 2651 1496 2795 1504
rect 2651 1476 2659 1496
rect 2679 1495 2767 1496
rect 2679 1476 2714 1495
rect 2735 1476 2767 1495
rect 2787 1476 2795 1496
rect 2651 1470 2795 1476
rect 2861 1500 2899 1508
rect 2977 1504 3013 1505
rect 2861 1480 2870 1500
rect 2890 1480 2899 1500
rect 2861 1471 2899 1480
rect 2928 1496 3013 1504
rect 2928 1476 2985 1496
rect 3005 1476 3013 1496
rect 2861 1470 2898 1471
rect 2928 1470 3013 1476
rect 3079 1500 3117 1508
rect 3079 1480 3088 1500
rect 3108 1480 3117 1500
rect 3350 1489 3387 1490
rect 3653 1489 3690 1559
rect 3725 1588 3756 1639
rect 4052 1634 4097 1640
rect 4052 1616 4070 1634
rect 4088 1616 4097 1634
rect 5558 1634 5567 1654
rect 5587 1634 5595 1654
rect 5558 1624 5595 1634
rect 5654 1654 5741 1664
rect 5654 1634 5663 1654
rect 5683 1634 5741 1654
rect 5654 1625 5741 1634
rect 5654 1624 5691 1625
rect 4052 1606 4097 1616
rect 3775 1588 3812 1589
rect 3725 1579 3812 1588
rect 3725 1559 3783 1579
rect 3803 1559 3812 1579
rect 3725 1549 3812 1559
rect 3871 1579 3908 1589
rect 3871 1559 3879 1579
rect 3899 1559 3908 1579
rect 4052 1564 4095 1606
rect 4479 1595 4531 1597
rect 3958 1562 4095 1564
rect 3725 1548 3756 1549
rect 3871 1489 3908 1559
rect 3349 1488 3690 1489
rect 3079 1471 3117 1480
rect 3274 1483 3690 1488
rect 3079 1470 3116 1471
rect 2540 1442 2630 1448
rect 2540 1422 2556 1442
rect 2576 1440 2630 1442
rect 2576 1422 2601 1440
rect 2540 1420 2601 1422
rect 2621 1420 2630 1440
rect 2540 1414 2630 1420
rect 2553 1360 2590 1361
rect 2649 1360 2686 1361
rect 2705 1360 2741 1470
rect 2928 1449 2959 1470
rect 3274 1463 3277 1483
rect 3297 1463 3690 1483
rect 3874 1473 3908 1489
rect 3952 1541 4095 1562
rect 4477 1591 4910 1595
rect 4477 1585 4916 1591
rect 4477 1567 4498 1585
rect 4516 1567 4916 1585
rect 5710 1574 5741 1625
rect 5776 1654 5813 1724
rect 6079 1723 6116 1724
rect 5928 1664 5964 1665
rect 5776 1634 5785 1654
rect 5805 1634 5813 1654
rect 5776 1624 5813 1634
rect 5872 1654 6020 1664
rect 6120 1661 6216 1663
rect 5872 1634 5881 1654
rect 5901 1634 5991 1654
rect 6011 1634 6020 1654
rect 5872 1625 6020 1634
rect 6078 1654 6216 1661
rect 6078 1634 6087 1654
rect 6107 1634 6216 1654
rect 6078 1625 6216 1634
rect 5872 1624 5909 1625
rect 5602 1571 5643 1572
rect 4477 1549 4916 1567
rect 3650 1454 3690 1463
rect 3952 1454 3979 1541
rect 4052 1515 4095 1541
rect 4052 1497 4065 1515
rect 4083 1497 4095 1515
rect 4052 1486 4095 1497
rect 2924 1448 2959 1449
rect 2802 1438 2959 1448
rect 2802 1418 2819 1438
rect 2839 1418 2959 1438
rect 2802 1411 2959 1418
rect 3026 1441 3175 1449
rect 3026 1421 3037 1441
rect 3057 1421 3096 1441
rect 3116 1421 3175 1441
rect 3650 1437 3979 1454
rect 3650 1436 3690 1437
rect 3026 1414 3175 1421
rect 4047 1425 4087 1428
rect 4047 1419 4090 1425
rect 3672 1416 4090 1419
rect 3026 1413 3067 1414
rect 2760 1360 2797 1361
rect 2453 1351 2591 1360
rect 2453 1331 2562 1351
rect 2582 1331 2591 1351
rect 2453 1324 2591 1331
rect 2649 1351 2797 1360
rect 2649 1331 2658 1351
rect 2678 1331 2768 1351
rect 2788 1331 2797 1351
rect 2453 1322 2549 1324
rect 2649 1321 2797 1331
rect 2856 1351 2893 1361
rect 2856 1331 2864 1351
rect 2884 1331 2893 1351
rect 2705 1320 2741 1321
rect 2553 1261 2590 1262
rect 2856 1261 2893 1331
rect 2928 1360 2959 1411
rect 3672 1398 4063 1416
rect 4081 1398 4090 1416
rect 3672 1396 4090 1398
rect 3672 1388 3699 1396
rect 3940 1393 4090 1396
rect 3252 1382 3420 1383
rect 3671 1382 3699 1388
rect 3252 1366 3699 1382
rect 4047 1388 4090 1393
rect 2978 1360 3015 1361
rect 2928 1351 3015 1360
rect 2928 1331 2986 1351
rect 3006 1331 3015 1351
rect 2928 1321 3015 1331
rect 3074 1351 3111 1361
rect 3074 1331 3082 1351
rect 3102 1331 3111 1351
rect 2928 1320 2959 1321
rect 2552 1260 2893 1261
rect 3074 1260 3111 1331
rect 2477 1255 2893 1260
rect 2477 1235 2480 1255
rect 2500 1235 2893 1255
rect 2924 1236 3111 1260
rect 3252 1356 3696 1366
rect 3252 1354 3420 1356
rect 3252 1176 3279 1354
rect 3319 1316 3383 1328
rect 3659 1324 3696 1356
rect 3722 1355 3913 1377
rect 3877 1353 3913 1355
rect 3877 1324 3914 1353
rect 4047 1332 4087 1388
rect 3319 1315 3354 1316
rect 3296 1310 3354 1315
rect 3296 1290 3299 1310
rect 3319 1296 3354 1310
rect 3374 1296 3383 1316
rect 3319 1288 3383 1296
rect 3345 1287 3383 1288
rect 3346 1286 3383 1287
rect 3449 1320 3485 1321
rect 3557 1320 3593 1321
rect 3449 1312 3593 1320
rect 3449 1292 3457 1312
rect 3477 1292 3512 1312
rect 3532 1292 3565 1312
rect 3585 1292 3593 1312
rect 3449 1286 3593 1292
rect 3659 1316 3697 1324
rect 3775 1320 3811 1321
rect 3659 1296 3668 1316
rect 3688 1296 3697 1316
rect 3659 1287 3697 1296
rect 3726 1312 3811 1320
rect 3726 1292 3783 1312
rect 3803 1292 3811 1312
rect 3659 1286 3696 1287
rect 3726 1286 3811 1292
rect 3877 1316 3915 1324
rect 3877 1296 3886 1316
rect 3906 1296 3915 1316
rect 4047 1314 4059 1332
rect 4077 1314 4087 1332
rect 4479 1360 4531 1549
rect 4877 1524 4916 1549
rect 5494 1564 5643 1571
rect 5494 1544 5553 1564
rect 5573 1544 5612 1564
rect 5632 1544 5643 1564
rect 5494 1536 5643 1544
rect 5710 1567 5867 1574
rect 5710 1547 5830 1567
rect 5850 1547 5867 1567
rect 5710 1537 5867 1547
rect 5710 1536 5745 1537
rect 4661 1499 4848 1523
rect 4877 1504 5272 1524
rect 5292 1504 5295 1524
rect 5710 1515 5741 1536
rect 5928 1515 5964 1625
rect 5983 1624 6020 1625
rect 6079 1624 6116 1625
rect 6039 1565 6129 1571
rect 6039 1545 6048 1565
rect 6068 1563 6129 1565
rect 6068 1545 6093 1563
rect 6039 1543 6093 1545
rect 6113 1543 6129 1563
rect 6039 1537 6129 1543
rect 5553 1514 5590 1515
rect 4877 1499 5295 1504
rect 5552 1505 5590 1514
rect 4661 1428 4698 1499
rect 4877 1498 5220 1499
rect 4877 1495 4916 1498
rect 5182 1497 5219 1498
rect 4813 1438 4844 1439
rect 4661 1408 4670 1428
rect 4690 1408 4698 1428
rect 4661 1398 4698 1408
rect 4757 1428 4844 1438
rect 4757 1408 4766 1428
rect 4786 1408 4844 1428
rect 4757 1399 4844 1408
rect 4757 1398 4794 1399
rect 4479 1342 4495 1360
rect 4513 1342 4531 1360
rect 4813 1348 4844 1399
rect 4879 1428 4916 1495
rect 5552 1485 5561 1505
rect 5581 1485 5590 1505
rect 5552 1477 5590 1485
rect 5656 1509 5741 1515
rect 5771 1514 5808 1515
rect 5656 1489 5664 1509
rect 5684 1489 5741 1509
rect 5656 1481 5741 1489
rect 5770 1505 5808 1514
rect 5770 1485 5779 1505
rect 5799 1485 5808 1505
rect 5656 1480 5692 1481
rect 5770 1477 5808 1485
rect 5874 1509 6018 1515
rect 5874 1489 5882 1509
rect 5902 1504 5990 1509
rect 5902 1489 5938 1504
rect 5874 1487 5938 1489
rect 5957 1489 5990 1504
rect 6010 1489 6018 1509
rect 5957 1487 6018 1489
rect 5874 1481 6018 1487
rect 5874 1480 5910 1481
rect 5982 1480 6018 1481
rect 6084 1514 6121 1515
rect 6084 1513 6122 1514
rect 6084 1505 6148 1513
rect 6084 1485 6093 1505
rect 6113 1491 6148 1505
rect 6168 1491 6171 1511
rect 6113 1486 6171 1491
rect 6113 1485 6148 1486
rect 5553 1448 5590 1477
rect 5554 1446 5590 1448
rect 5031 1438 5067 1439
rect 4879 1408 4888 1428
rect 4908 1408 4916 1428
rect 4879 1398 4916 1408
rect 4975 1428 5123 1438
rect 5223 1435 5319 1437
rect 4975 1408 4984 1428
rect 5004 1408 5094 1428
rect 5114 1408 5123 1428
rect 4975 1399 5123 1408
rect 5181 1428 5319 1435
rect 5181 1408 5190 1428
rect 5210 1408 5319 1428
rect 5554 1424 5745 1446
rect 5771 1445 5808 1477
rect 6084 1473 6148 1485
rect 6188 1447 6215 1625
rect 6047 1445 6215 1447
rect 5771 1431 6215 1445
rect 6818 1579 6986 1580
rect 7112 1579 7152 1803
rect 7615 1807 7783 1808
rect 8018 1807 8058 1840
rect 8414 1807 8461 1840
rect 8865 1838 8906 1863
rect 9051 1838 9088 1869
rect 9269 1838 9306 1869
rect 9582 1865 9646 1877
rect 9686 1839 9713 2017
rect 8865 1811 8914 1838
rect 9050 1812 9099 1838
rect 9268 1837 9349 1838
rect 9545 1837 9713 1839
rect 9268 1812 9713 1837
rect 9269 1811 9713 1812
rect 7615 1806 8059 1807
rect 7615 1781 8060 1806
rect 7615 1779 7783 1781
rect 7979 1780 8060 1781
rect 8229 1780 8278 1806
rect 8414 1780 8463 1807
rect 7615 1601 7642 1779
rect 7682 1741 7746 1753
rect 8022 1749 8059 1780
rect 8240 1749 8277 1780
rect 8422 1755 8463 1780
rect 8867 1778 8914 1811
rect 9270 1778 9310 1811
rect 9545 1810 9713 1811
rect 10176 1815 10216 2039
rect 10342 2038 10510 2039
rect 11113 2173 11557 2187
rect 11113 2171 11281 2173
rect 11113 1993 11140 2171
rect 11180 2133 11244 2145
rect 11520 2141 11557 2173
rect 11583 2172 11774 2194
rect 12009 2190 12118 2210
rect 12138 2190 12147 2210
rect 12009 2183 12147 2190
rect 12205 2210 12353 2219
rect 12205 2190 12214 2210
rect 12234 2190 12324 2210
rect 12344 2190 12353 2210
rect 12009 2181 12105 2183
rect 12205 2180 12353 2190
rect 12412 2210 12449 2220
rect 12412 2190 12420 2210
rect 12440 2190 12449 2210
rect 12261 2179 12297 2180
rect 11738 2170 11774 2172
rect 11738 2141 11775 2170
rect 11180 2132 11215 2133
rect 11157 2127 11215 2132
rect 11157 2107 11160 2127
rect 11180 2113 11215 2127
rect 11235 2113 11244 2133
rect 11180 2105 11244 2113
rect 11206 2104 11244 2105
rect 11207 2103 11244 2104
rect 11310 2137 11346 2138
rect 11418 2137 11454 2138
rect 11310 2129 11454 2137
rect 11310 2109 11318 2129
rect 11338 2127 11426 2129
rect 11338 2109 11371 2127
rect 11310 2108 11371 2109
rect 11392 2109 11426 2127
rect 11446 2109 11454 2129
rect 11392 2108 11454 2109
rect 11310 2103 11454 2108
rect 11520 2133 11558 2141
rect 11636 2137 11672 2138
rect 11520 2113 11529 2133
rect 11549 2113 11558 2133
rect 11520 2104 11558 2113
rect 11587 2129 11672 2137
rect 11587 2109 11644 2129
rect 11664 2109 11672 2129
rect 11520 2103 11557 2104
rect 11587 2103 11672 2109
rect 11738 2133 11776 2141
rect 11738 2113 11747 2133
rect 11767 2113 11776 2133
rect 12412 2123 12449 2190
rect 12484 2219 12515 2270
rect 12797 2258 12815 2276
rect 12833 2258 12849 2276
rect 12534 2219 12571 2220
rect 12484 2210 12571 2219
rect 12484 2190 12542 2210
rect 12562 2190 12571 2210
rect 12484 2180 12571 2190
rect 12630 2210 12667 2220
rect 12630 2190 12638 2210
rect 12658 2190 12667 2210
rect 12484 2179 12515 2180
rect 12109 2120 12146 2121
rect 12412 2120 12451 2123
rect 12108 2119 12451 2120
rect 12630 2119 12667 2190
rect 11738 2104 11776 2113
rect 12033 2114 12451 2119
rect 11738 2103 11775 2104
rect 11199 2075 11289 2081
rect 11199 2055 11215 2075
rect 11235 2073 11289 2075
rect 11235 2055 11260 2073
rect 11199 2053 11260 2055
rect 11280 2053 11289 2073
rect 11199 2047 11289 2053
rect 11212 1993 11249 1994
rect 11308 1993 11345 1994
rect 11364 1993 11400 2103
rect 11587 2082 11618 2103
rect 12033 2094 12036 2114
rect 12056 2094 12451 2114
rect 12480 2095 12667 2119
rect 11583 2081 11618 2082
rect 11461 2071 11618 2081
rect 11461 2051 11478 2071
rect 11498 2051 11618 2071
rect 11461 2044 11618 2051
rect 11685 2074 11834 2082
rect 11685 2054 11696 2074
rect 11716 2054 11755 2074
rect 11775 2054 11834 2074
rect 11685 2047 11834 2054
rect 12412 2069 12451 2094
rect 12797 2069 12849 2258
rect 13241 2286 13251 2304
rect 13269 2286 13281 2304
rect 13413 2302 13422 2322
rect 13442 2302 13451 2322
rect 13413 2294 13451 2302
rect 13517 2326 13602 2332
rect 13632 2331 13669 2332
rect 13517 2306 13525 2326
rect 13545 2306 13602 2326
rect 13517 2298 13602 2306
rect 13631 2322 13669 2331
rect 13631 2302 13640 2322
rect 13660 2302 13669 2322
rect 13517 2297 13553 2298
rect 13631 2294 13669 2302
rect 13735 2326 13879 2332
rect 13735 2306 13743 2326
rect 13763 2306 13796 2326
rect 13816 2306 13851 2326
rect 13871 2306 13879 2326
rect 13735 2298 13879 2306
rect 13735 2297 13771 2298
rect 13843 2297 13879 2298
rect 13945 2331 13982 2332
rect 13945 2330 13983 2331
rect 13945 2322 14009 2330
rect 13945 2302 13954 2322
rect 13974 2308 14009 2322
rect 14029 2308 14032 2328
rect 13974 2303 14032 2308
rect 13974 2302 14009 2303
rect 13241 2230 13281 2286
rect 13414 2265 13451 2294
rect 13415 2263 13451 2265
rect 13415 2241 13606 2263
rect 13632 2262 13669 2294
rect 13945 2290 14009 2302
rect 14049 2264 14076 2442
rect 13908 2262 14076 2264
rect 13632 2252 14076 2262
rect 14217 2358 14404 2382
rect 14435 2363 14828 2383
rect 14848 2363 14851 2383
rect 14435 2358 14851 2363
rect 14217 2287 14254 2358
rect 14435 2357 14776 2358
rect 14369 2297 14400 2298
rect 14217 2267 14226 2287
rect 14246 2267 14254 2287
rect 14217 2257 14254 2267
rect 14313 2287 14400 2297
rect 14313 2267 14322 2287
rect 14342 2267 14400 2287
rect 14313 2258 14400 2267
rect 14313 2257 14350 2258
rect 13238 2225 13281 2230
rect 13629 2236 14076 2252
rect 13629 2230 13657 2236
rect 13908 2235 14076 2236
rect 13238 2222 13388 2225
rect 13629 2222 13656 2230
rect 13238 2220 13656 2222
rect 13238 2202 13247 2220
rect 13265 2202 13656 2220
rect 14369 2207 14400 2258
rect 14435 2287 14472 2357
rect 14738 2356 14775 2357
rect 14976 2299 15009 2458
rect 14587 2297 14623 2298
rect 14435 2267 14444 2287
rect 14464 2267 14472 2287
rect 14435 2257 14472 2267
rect 14531 2287 14679 2297
rect 14779 2294 14875 2296
rect 14531 2267 14540 2287
rect 14560 2267 14650 2287
rect 14670 2267 14679 2287
rect 14531 2258 14679 2267
rect 14737 2287 14875 2294
rect 14737 2267 14746 2287
rect 14766 2267 14875 2287
rect 14976 2295 15012 2299
rect 14976 2277 14985 2295
rect 15007 2277 15012 2295
rect 14976 2271 15012 2277
rect 14737 2258 14875 2267
rect 14531 2257 14568 2258
rect 14261 2204 14302 2205
rect 13238 2199 13656 2202
rect 13238 2193 13281 2199
rect 13241 2190 13281 2193
rect 14153 2197 14302 2204
rect 13638 2181 13678 2182
rect 13349 2164 13678 2181
rect 14153 2177 14212 2197
rect 14232 2177 14271 2197
rect 14291 2177 14302 2197
rect 14153 2169 14302 2177
rect 14369 2200 14526 2207
rect 14369 2180 14489 2200
rect 14509 2180 14526 2200
rect 14369 2170 14526 2180
rect 14369 2169 14404 2170
rect 13233 2121 13276 2132
rect 13233 2103 13245 2121
rect 13263 2103 13276 2121
rect 13233 2077 13276 2103
rect 13349 2077 13376 2164
rect 13638 2155 13678 2164
rect 12412 2051 12851 2069
rect 11685 2046 11726 2047
rect 11419 1993 11456 1994
rect 11112 1984 11250 1993
rect 11112 1964 11221 1984
rect 11241 1964 11250 1984
rect 11112 1957 11250 1964
rect 11308 1984 11456 1993
rect 11308 1964 11317 1984
rect 11337 1964 11427 1984
rect 11447 1964 11456 1984
rect 11112 1955 11208 1957
rect 11308 1954 11456 1964
rect 11515 1984 11552 1994
rect 11515 1964 11523 1984
rect 11543 1964 11552 1984
rect 11364 1953 11400 1954
rect 11212 1894 11249 1895
rect 11515 1894 11552 1964
rect 11587 1993 11618 2044
rect 12412 2033 12812 2051
rect 12830 2033 12851 2051
rect 12412 2027 12851 2033
rect 12418 2023 12851 2027
rect 13233 2056 13376 2077
rect 13420 2129 13454 2145
rect 13638 2135 14031 2155
rect 14051 2135 14054 2155
rect 14369 2148 14400 2169
rect 14587 2148 14623 2258
rect 14642 2257 14679 2258
rect 14738 2257 14775 2258
rect 14698 2198 14788 2204
rect 14698 2178 14707 2198
rect 14727 2196 14788 2198
rect 14727 2178 14752 2196
rect 14698 2176 14752 2178
rect 14772 2176 14788 2196
rect 14698 2170 14788 2176
rect 14212 2147 14249 2148
rect 13638 2130 14054 2135
rect 14211 2138 14249 2147
rect 13638 2129 13979 2130
rect 13420 2059 13457 2129
rect 13572 2069 13603 2070
rect 13233 2054 13370 2056
rect 12797 2021 12849 2023
rect 13233 2012 13276 2054
rect 13420 2039 13429 2059
rect 13449 2039 13457 2059
rect 13420 2029 13457 2039
rect 13516 2059 13603 2069
rect 13516 2039 13525 2059
rect 13545 2039 13603 2059
rect 13516 2030 13603 2039
rect 13516 2029 13553 2030
rect 13231 2002 13276 2012
rect 11637 1993 11674 1994
rect 11587 1984 11674 1993
rect 11587 1964 11645 1984
rect 11665 1964 11674 1984
rect 11587 1954 11674 1964
rect 11733 1984 11770 1994
rect 11733 1964 11741 1984
rect 11761 1964 11770 1984
rect 13231 1984 13240 2002
rect 13258 1984 13276 2002
rect 13231 1978 13276 1984
rect 13572 1979 13603 2030
rect 13638 2059 13675 2129
rect 13941 2128 13978 2129
rect 14211 2118 14220 2138
rect 14240 2118 14249 2138
rect 14211 2110 14249 2118
rect 14315 2142 14400 2148
rect 14430 2147 14467 2148
rect 14315 2122 14323 2142
rect 14343 2122 14400 2142
rect 14315 2114 14400 2122
rect 14429 2138 14467 2147
rect 14429 2118 14438 2138
rect 14458 2118 14467 2138
rect 14315 2113 14351 2114
rect 14429 2110 14467 2118
rect 14533 2142 14677 2148
rect 14533 2122 14541 2142
rect 14561 2123 14593 2142
rect 14614 2123 14649 2142
rect 14561 2122 14649 2123
rect 14669 2122 14677 2142
rect 14533 2114 14677 2122
rect 14533 2113 14569 2114
rect 14641 2113 14677 2114
rect 14743 2147 14780 2148
rect 14743 2146 14781 2147
rect 14743 2138 14807 2146
rect 14743 2118 14752 2138
rect 14772 2124 14807 2138
rect 14827 2124 14830 2144
rect 14772 2119 14830 2124
rect 14772 2118 14807 2119
rect 14212 2081 14249 2110
rect 14213 2079 14249 2081
rect 13790 2069 13826 2070
rect 13638 2039 13647 2059
rect 13667 2039 13675 2059
rect 13638 2029 13675 2039
rect 13734 2059 13882 2069
rect 13982 2066 14078 2068
rect 13734 2039 13743 2059
rect 13763 2039 13853 2059
rect 13873 2039 13882 2059
rect 13734 2030 13882 2039
rect 13940 2059 14078 2066
rect 13940 2039 13949 2059
rect 13969 2039 14078 2059
rect 14213 2057 14404 2079
rect 14430 2078 14467 2110
rect 14743 2106 14807 2118
rect 14847 2080 14874 2258
rect 15479 2257 15512 2590
rect 15576 2622 15744 2623
rect 15870 2622 15910 2846
rect 16373 2850 16541 2851
rect 16777 2850 16818 2884
rect 17175 2863 17222 2884
rect 16373 2840 16818 2850
rect 16890 2848 17033 2849
rect 16373 2824 16817 2840
rect 16373 2822 16541 2824
rect 16737 2823 16817 2824
rect 16890 2823 17035 2848
rect 17177 2823 17222 2863
rect 17513 2903 17551 2905
rect 17513 2895 17556 2903
rect 17513 2877 17524 2895
rect 17542 2877 17556 2895
rect 17513 2850 17556 2877
rect 17700 2902 17738 2911
rect 17700 2882 17709 2902
rect 17729 2882 17738 2902
rect 17700 2874 17738 2882
rect 17804 2906 17889 2912
rect 17919 2911 17956 2912
rect 17804 2886 17812 2906
rect 17832 2886 17889 2906
rect 17804 2878 17889 2886
rect 17918 2902 17956 2911
rect 17918 2882 17927 2902
rect 17947 2882 17956 2902
rect 17804 2877 17840 2878
rect 17918 2874 17956 2882
rect 18022 2910 18166 2912
rect 18022 2906 18074 2910
rect 18022 2886 18030 2906
rect 18050 2890 18074 2906
rect 18094 2906 18166 2910
rect 18094 2890 18138 2906
rect 18050 2886 18138 2890
rect 18158 2886 18166 2906
rect 18022 2878 18166 2886
rect 18022 2877 18058 2878
rect 18130 2877 18166 2878
rect 18232 2911 18269 2912
rect 18232 2910 18270 2911
rect 18232 2902 18296 2910
rect 18232 2882 18241 2902
rect 18261 2888 18296 2902
rect 18316 2888 18319 2908
rect 18261 2883 18319 2888
rect 18261 2882 18296 2883
rect 16373 2644 16400 2822
rect 16440 2784 16504 2796
rect 16780 2792 16817 2823
rect 16998 2792 17035 2823
rect 17180 2816 17222 2823
rect 17514 2843 17556 2850
rect 17701 2843 17738 2874
rect 17919 2843 17956 2874
rect 18232 2870 18296 2882
rect 18336 2844 18363 3022
rect 16440 2783 16475 2784
rect 16417 2778 16475 2783
rect 16417 2758 16420 2778
rect 16440 2764 16475 2778
rect 16495 2764 16504 2784
rect 16440 2756 16504 2764
rect 16466 2755 16504 2756
rect 16467 2754 16504 2755
rect 16570 2788 16606 2789
rect 16678 2788 16714 2789
rect 16570 2780 16714 2788
rect 16570 2760 16578 2780
rect 16598 2776 16686 2780
rect 16598 2760 16642 2776
rect 16570 2756 16642 2760
rect 16662 2760 16686 2776
rect 16706 2760 16714 2780
rect 16662 2756 16714 2760
rect 16570 2754 16714 2756
rect 16780 2784 16818 2792
rect 16896 2788 16932 2789
rect 16780 2764 16789 2784
rect 16809 2764 16818 2784
rect 16780 2755 16818 2764
rect 16847 2780 16932 2788
rect 16847 2760 16904 2780
rect 16924 2760 16932 2780
rect 16780 2754 16817 2755
rect 16847 2754 16932 2760
rect 16998 2784 17036 2792
rect 16998 2764 17007 2784
rect 17027 2764 17036 2784
rect 16998 2755 17036 2764
rect 17180 2789 17223 2816
rect 17180 2771 17194 2789
rect 17212 2771 17223 2789
rect 17180 2763 17223 2771
rect 17185 2761 17223 2763
rect 17514 2803 17559 2843
rect 17701 2818 17846 2843
rect 17919 2842 17999 2843
rect 18195 2842 18363 2844
rect 17919 2826 18363 2842
rect 17703 2817 17846 2818
rect 17918 2816 18363 2826
rect 17514 2782 17561 2803
rect 17918 2782 17959 2816
rect 18195 2815 18363 2816
rect 18826 2820 18866 3044
rect 18992 3043 19160 3044
rect 19224 3076 19257 3409
rect 19224 3068 19261 3076
rect 19224 3049 19232 3068
rect 19253 3049 19261 3068
rect 19224 3043 19261 3049
rect 18826 2798 18834 2820
rect 18858 2798 18866 2820
rect 18826 2790 18866 2798
rect 16998 2754 17035 2755
rect 16459 2726 16549 2732
rect 16459 2706 16475 2726
rect 16495 2724 16549 2726
rect 16495 2706 16520 2724
rect 16459 2704 16520 2706
rect 16540 2704 16549 2724
rect 16459 2698 16549 2704
rect 16472 2644 16509 2645
rect 16568 2644 16605 2645
rect 16624 2644 16660 2754
rect 16847 2733 16878 2754
rect 17514 2752 17959 2782
rect 18997 2765 19062 2766
rect 17514 2749 17937 2752
rect 16843 2732 16878 2733
rect 16721 2722 16878 2732
rect 16721 2702 16738 2722
rect 16758 2702 16878 2722
rect 16721 2695 16878 2702
rect 16945 2725 17094 2733
rect 16945 2705 16956 2725
rect 16976 2705 17015 2725
rect 17035 2705 17094 2725
rect 16945 2698 17094 2705
rect 17514 2701 17561 2749
rect 16945 2697 16986 2698
rect 17182 2696 17219 2699
rect 16679 2644 16716 2645
rect 16372 2635 16510 2644
rect 15576 2596 16020 2622
rect 15576 2594 15744 2596
rect 15576 2416 15603 2594
rect 15643 2556 15707 2568
rect 15983 2564 16020 2596
rect 16046 2595 16237 2617
rect 16372 2615 16481 2635
rect 16501 2615 16510 2635
rect 16372 2608 16510 2615
rect 16568 2635 16716 2644
rect 16568 2615 16577 2635
rect 16597 2615 16687 2635
rect 16707 2615 16716 2635
rect 16372 2606 16468 2608
rect 16568 2605 16716 2615
rect 16775 2635 16812 2645
rect 16775 2615 16783 2635
rect 16803 2615 16812 2635
rect 16624 2604 16660 2605
rect 16201 2593 16237 2595
rect 16201 2564 16238 2593
rect 15643 2555 15678 2556
rect 15620 2550 15678 2555
rect 15620 2530 15623 2550
rect 15643 2536 15678 2550
rect 15698 2536 15707 2556
rect 15643 2530 15707 2536
rect 15620 2528 15707 2530
rect 15620 2524 15647 2528
rect 15669 2527 15707 2528
rect 15670 2526 15707 2527
rect 15773 2560 15809 2561
rect 15881 2560 15917 2561
rect 15773 2553 15917 2560
rect 15773 2552 15835 2553
rect 15773 2532 15781 2552
rect 15801 2535 15835 2552
rect 15854 2552 15917 2553
rect 15854 2535 15889 2552
rect 15801 2532 15889 2535
rect 15909 2532 15917 2552
rect 15773 2526 15917 2532
rect 15983 2556 16021 2564
rect 16099 2560 16135 2561
rect 15983 2536 15992 2556
rect 16012 2536 16021 2556
rect 15983 2527 16021 2536
rect 16050 2552 16135 2560
rect 16050 2532 16107 2552
rect 16127 2532 16135 2552
rect 15983 2526 16020 2527
rect 16050 2526 16135 2532
rect 16201 2556 16239 2564
rect 16201 2536 16210 2556
rect 16230 2536 16239 2556
rect 16472 2545 16509 2546
rect 16775 2545 16812 2615
rect 16847 2644 16878 2695
rect 17174 2690 17219 2696
rect 17174 2672 17192 2690
rect 17210 2672 17219 2690
rect 17514 2683 17524 2701
rect 17542 2683 17561 2701
rect 17514 2679 17561 2683
rect 18648 2740 18835 2764
rect 18866 2745 19259 2765
rect 19279 2745 19282 2765
rect 18866 2740 19282 2745
rect 17515 2674 17552 2679
rect 17174 2662 17219 2672
rect 18648 2669 18685 2740
rect 18866 2739 19207 2740
rect 18800 2679 18831 2680
rect 16897 2644 16934 2645
rect 16847 2635 16934 2644
rect 16847 2615 16905 2635
rect 16925 2615 16934 2635
rect 16847 2605 16934 2615
rect 16993 2635 17030 2645
rect 16993 2615 17001 2635
rect 17021 2615 17030 2635
rect 17174 2620 17217 2662
rect 18648 2649 18657 2669
rect 18677 2649 18685 2669
rect 18648 2639 18685 2649
rect 18744 2669 18831 2679
rect 18744 2649 18753 2669
rect 18773 2649 18831 2669
rect 18744 2640 18831 2649
rect 18744 2639 18781 2640
rect 17080 2618 17217 2620
rect 16847 2604 16878 2605
rect 16993 2545 17030 2615
rect 16471 2544 16812 2545
rect 16201 2527 16239 2536
rect 16396 2539 16812 2544
rect 16201 2526 16238 2527
rect 15662 2498 15752 2504
rect 15662 2478 15678 2498
rect 15698 2496 15752 2498
rect 15698 2478 15723 2496
rect 15662 2476 15723 2478
rect 15743 2476 15752 2496
rect 15662 2470 15752 2476
rect 15675 2416 15712 2417
rect 15771 2416 15808 2417
rect 15827 2416 15863 2526
rect 16050 2505 16081 2526
rect 16396 2519 16399 2539
rect 16419 2519 16812 2539
rect 16996 2529 17030 2545
rect 17074 2597 17217 2618
rect 17503 2612 17555 2614
rect 16772 2510 16812 2519
rect 17074 2510 17101 2597
rect 17174 2571 17217 2597
rect 17174 2553 17187 2571
rect 17205 2553 17217 2571
rect 17501 2608 17934 2612
rect 17501 2602 17940 2608
rect 17501 2584 17522 2602
rect 17540 2584 17940 2602
rect 18800 2589 18831 2640
rect 18866 2669 18903 2739
rect 19169 2738 19206 2739
rect 19018 2679 19054 2680
rect 18866 2649 18875 2669
rect 18895 2649 18903 2669
rect 18866 2639 18903 2649
rect 18962 2669 19110 2679
rect 19210 2676 19306 2678
rect 18962 2649 18971 2669
rect 18991 2649 19081 2669
rect 19101 2649 19110 2669
rect 18962 2640 19110 2649
rect 19168 2669 19306 2676
rect 19168 2649 19177 2669
rect 19197 2649 19306 2669
rect 19168 2640 19306 2649
rect 18962 2639 18999 2640
rect 18692 2586 18733 2587
rect 17501 2566 17940 2584
rect 17174 2542 17217 2553
rect 16046 2504 16081 2505
rect 15924 2494 16081 2504
rect 15924 2474 15941 2494
rect 15961 2474 16081 2494
rect 15924 2467 16081 2474
rect 16148 2497 16294 2505
rect 16148 2477 16159 2497
rect 16179 2477 16218 2497
rect 16238 2477 16294 2497
rect 16772 2493 17101 2510
rect 16772 2492 16812 2493
rect 16148 2470 16294 2477
rect 17169 2481 17209 2484
rect 17169 2475 17212 2481
rect 16794 2472 17212 2475
rect 16148 2469 16189 2470
rect 15882 2416 15919 2417
rect 15575 2407 15713 2416
rect 15575 2387 15684 2407
rect 15704 2387 15713 2407
rect 15575 2380 15713 2387
rect 15771 2407 15919 2416
rect 15771 2387 15780 2407
rect 15800 2387 15890 2407
rect 15910 2387 15919 2407
rect 15575 2378 15671 2380
rect 15771 2377 15919 2387
rect 15978 2407 16015 2417
rect 15978 2387 15986 2407
rect 16006 2387 16015 2407
rect 15827 2376 15863 2377
rect 15675 2317 15712 2318
rect 15978 2317 16015 2387
rect 16050 2416 16081 2467
rect 16794 2454 17185 2472
rect 17203 2454 17212 2472
rect 16794 2452 17212 2454
rect 16794 2444 16821 2452
rect 17062 2449 17212 2452
rect 16374 2438 16542 2439
rect 16793 2438 16821 2444
rect 16374 2422 16821 2438
rect 17169 2444 17212 2449
rect 16100 2416 16137 2417
rect 16050 2407 16137 2416
rect 16050 2387 16108 2407
rect 16128 2387 16137 2407
rect 16050 2377 16137 2387
rect 16196 2407 16233 2417
rect 16196 2387 16204 2407
rect 16224 2387 16233 2407
rect 16050 2376 16081 2377
rect 15674 2316 16015 2317
rect 16196 2316 16233 2387
rect 15599 2311 16015 2316
rect 15599 2291 15602 2311
rect 15622 2291 16015 2311
rect 16046 2292 16233 2316
rect 16374 2412 16818 2422
rect 16374 2410 16542 2412
rect 15474 2212 15516 2257
rect 16374 2232 16401 2410
rect 16441 2372 16505 2384
rect 16781 2380 16818 2412
rect 16844 2411 17035 2433
rect 16999 2409 17035 2411
rect 16999 2380 17036 2409
rect 17169 2388 17209 2444
rect 16441 2371 16476 2372
rect 16418 2366 16476 2371
rect 16418 2346 16421 2366
rect 16441 2352 16476 2366
rect 16496 2352 16505 2372
rect 16441 2344 16505 2352
rect 16467 2343 16505 2344
rect 16468 2342 16505 2343
rect 16571 2376 16607 2377
rect 16679 2376 16715 2377
rect 16571 2368 16715 2376
rect 16571 2348 16579 2368
rect 16599 2348 16634 2368
rect 16654 2348 16687 2368
rect 16707 2348 16715 2368
rect 16571 2342 16715 2348
rect 16781 2372 16819 2380
rect 16897 2376 16933 2377
rect 16781 2352 16790 2372
rect 16810 2352 16819 2372
rect 16781 2343 16819 2352
rect 16848 2368 16933 2376
rect 16848 2348 16905 2368
rect 16925 2348 16933 2368
rect 16781 2342 16818 2343
rect 16848 2342 16933 2348
rect 16999 2372 17037 2380
rect 16999 2352 17008 2372
rect 17028 2352 17037 2372
rect 17169 2370 17181 2388
rect 17199 2370 17209 2388
rect 17169 2360 17209 2370
rect 17503 2377 17555 2566
rect 17901 2541 17940 2566
rect 18584 2579 18733 2586
rect 18584 2559 18643 2579
rect 18663 2559 18702 2579
rect 18722 2559 18733 2579
rect 18584 2551 18733 2559
rect 18800 2582 18957 2589
rect 18800 2562 18920 2582
rect 18940 2562 18957 2582
rect 18800 2552 18957 2562
rect 18800 2551 18835 2552
rect 17685 2516 17872 2540
rect 17901 2521 18296 2541
rect 18316 2521 18319 2541
rect 18800 2530 18831 2551
rect 19018 2530 19054 2640
rect 19073 2639 19110 2640
rect 19169 2639 19206 2640
rect 19129 2580 19219 2586
rect 19129 2560 19138 2580
rect 19158 2578 19219 2580
rect 19158 2560 19183 2578
rect 19129 2558 19183 2560
rect 19203 2558 19219 2578
rect 19129 2552 19219 2558
rect 18643 2529 18680 2530
rect 17901 2516 18319 2521
rect 18642 2520 18680 2529
rect 17685 2445 17722 2516
rect 17901 2515 18244 2516
rect 17901 2512 17940 2515
rect 18206 2514 18243 2515
rect 17837 2455 17868 2456
rect 17685 2425 17694 2445
rect 17714 2425 17722 2445
rect 17685 2415 17722 2425
rect 17781 2445 17868 2455
rect 17781 2425 17790 2445
rect 17810 2425 17868 2445
rect 17781 2416 17868 2425
rect 17781 2415 17818 2416
rect 16999 2343 17037 2352
rect 17503 2359 17519 2377
rect 17537 2359 17555 2377
rect 17837 2365 17868 2416
rect 17903 2445 17940 2512
rect 18642 2500 18651 2520
rect 18671 2500 18680 2520
rect 18642 2492 18680 2500
rect 18746 2524 18831 2530
rect 18861 2529 18898 2530
rect 18746 2504 18754 2524
rect 18774 2504 18831 2524
rect 18746 2496 18831 2504
rect 18860 2520 18898 2529
rect 18860 2500 18869 2520
rect 18889 2500 18898 2520
rect 18746 2495 18782 2496
rect 18860 2492 18898 2500
rect 18964 2528 19108 2530
rect 18964 2524 19024 2528
rect 18964 2504 18972 2524
rect 18992 2506 19024 2524
rect 19047 2524 19108 2528
rect 19047 2506 19080 2524
rect 18992 2504 19080 2506
rect 19100 2504 19108 2524
rect 18964 2496 19108 2504
rect 18964 2495 19000 2496
rect 19072 2495 19108 2496
rect 19174 2529 19211 2530
rect 19174 2528 19212 2529
rect 19174 2520 19238 2528
rect 19174 2500 19183 2520
rect 19203 2506 19238 2520
rect 19258 2506 19261 2526
rect 19203 2501 19261 2506
rect 19203 2500 19238 2501
rect 18643 2463 18680 2492
rect 18644 2461 18680 2463
rect 18055 2455 18091 2456
rect 17903 2425 17912 2445
rect 17932 2425 17940 2445
rect 17903 2415 17940 2425
rect 17999 2445 18147 2455
rect 18247 2452 18343 2454
rect 17999 2425 18008 2445
rect 18028 2425 18118 2445
rect 18138 2425 18147 2445
rect 17999 2416 18147 2425
rect 18205 2445 18343 2452
rect 18205 2425 18214 2445
rect 18234 2425 18343 2445
rect 18644 2439 18835 2461
rect 18861 2460 18898 2492
rect 19174 2488 19238 2500
rect 18861 2459 19136 2460
rect 19278 2459 19305 2640
rect 18861 2434 19305 2459
rect 19441 2465 19480 4280
rect 19782 4267 19815 4600
rect 19879 4632 20047 4633
rect 20173 4632 20213 4856
rect 20676 4860 20844 4861
rect 21085 4860 21120 4877
rect 21477 4867 21524 4878
rect 20676 4834 21120 4860
rect 20676 4832 20844 4834
rect 21040 4833 21120 4834
rect 21275 4833 21342 4859
rect 21481 4833 21524 4867
rect 20676 4654 20703 4832
rect 20743 4794 20807 4806
rect 21083 4802 21120 4833
rect 21301 4802 21338 4833
rect 21483 4808 21524 4833
rect 21915 4892 21956 4917
rect 22101 4892 22138 4923
rect 22319 4892 22356 4923
rect 22632 4919 22696 4931
rect 22736 4893 22763 5071
rect 21915 4858 21958 4892
rect 22097 4866 22164 4892
rect 22319 4891 22399 4892
rect 22595 4891 22763 4893
rect 22319 4865 22763 4891
rect 21915 4847 21962 4858
rect 22319 4848 22354 4865
rect 22595 4864 22763 4865
rect 23226 4869 23266 5093
rect 23392 5092 23560 5093
rect 23624 5125 23657 5458
rect 23959 5445 23998 7260
rect 24134 7266 24578 7291
rect 24134 7085 24161 7266
rect 24303 7265 24578 7266
rect 24201 7225 24265 7237
rect 24541 7233 24578 7265
rect 24604 7264 24795 7286
rect 25096 7280 25205 7300
rect 25225 7280 25234 7300
rect 25096 7273 25234 7280
rect 25292 7300 25440 7309
rect 25292 7280 25301 7300
rect 25321 7280 25411 7300
rect 25431 7280 25440 7300
rect 25096 7271 25192 7273
rect 25292 7270 25440 7280
rect 25499 7300 25536 7310
rect 25499 7280 25507 7300
rect 25527 7280 25536 7300
rect 25348 7269 25384 7270
rect 24759 7262 24795 7264
rect 24759 7233 24796 7262
rect 24201 7224 24236 7225
rect 24178 7219 24236 7224
rect 24178 7199 24181 7219
rect 24201 7205 24236 7219
rect 24256 7205 24265 7225
rect 24201 7197 24265 7205
rect 24227 7196 24265 7197
rect 24228 7195 24265 7196
rect 24331 7229 24367 7230
rect 24439 7229 24475 7230
rect 24331 7221 24475 7229
rect 24331 7201 24339 7221
rect 24359 7219 24447 7221
rect 24359 7201 24392 7219
rect 24331 7197 24392 7201
rect 24415 7201 24447 7219
rect 24467 7201 24475 7221
rect 24415 7197 24475 7201
rect 24331 7195 24475 7197
rect 24541 7225 24579 7233
rect 24657 7229 24693 7230
rect 24541 7205 24550 7225
rect 24570 7205 24579 7225
rect 24541 7196 24579 7205
rect 24608 7221 24693 7229
rect 24608 7201 24665 7221
rect 24685 7201 24693 7221
rect 24541 7195 24578 7196
rect 24608 7195 24693 7201
rect 24759 7225 24797 7233
rect 24759 7205 24768 7225
rect 24788 7205 24797 7225
rect 25499 7213 25536 7280
rect 25571 7309 25602 7360
rect 25884 7348 25902 7366
rect 25920 7348 25936 7366
rect 25621 7309 25658 7310
rect 25571 7300 25658 7309
rect 25571 7280 25629 7300
rect 25649 7280 25658 7300
rect 25571 7270 25658 7280
rect 25717 7300 25754 7310
rect 25717 7280 25725 7300
rect 25745 7280 25754 7300
rect 25571 7269 25602 7270
rect 25196 7210 25233 7211
rect 25499 7210 25538 7213
rect 25195 7209 25538 7210
rect 25717 7209 25754 7280
rect 24759 7196 24797 7205
rect 25120 7204 25538 7209
rect 24759 7195 24796 7196
rect 24220 7167 24310 7173
rect 24220 7147 24236 7167
rect 24256 7165 24310 7167
rect 24256 7147 24281 7165
rect 24220 7145 24281 7147
rect 24301 7145 24310 7165
rect 24220 7139 24310 7145
rect 24233 7085 24270 7086
rect 24329 7085 24366 7086
rect 24385 7085 24421 7195
rect 24608 7174 24639 7195
rect 25120 7184 25123 7204
rect 25143 7184 25538 7204
rect 25567 7185 25754 7209
rect 24604 7173 24639 7174
rect 24482 7163 24639 7173
rect 24482 7143 24499 7163
rect 24519 7143 24639 7163
rect 24482 7136 24639 7143
rect 24706 7166 24855 7174
rect 24706 7146 24717 7166
rect 24737 7146 24776 7166
rect 24796 7146 24855 7166
rect 24706 7139 24855 7146
rect 25499 7159 25538 7184
rect 25884 7159 25936 7348
rect 26341 7375 26351 7393
rect 26369 7375 26381 7393
rect 26513 7391 26522 7411
rect 26542 7391 26551 7411
rect 26513 7383 26551 7391
rect 26617 7415 26702 7421
rect 26732 7420 26769 7421
rect 26617 7395 26625 7415
rect 26645 7395 26702 7415
rect 26617 7387 26702 7395
rect 26731 7411 26769 7420
rect 26731 7391 26740 7411
rect 26760 7391 26769 7411
rect 26617 7386 26653 7387
rect 26731 7383 26769 7391
rect 26835 7415 26979 7421
rect 26835 7395 26843 7415
rect 26863 7395 26896 7415
rect 26916 7395 26951 7415
rect 26971 7395 26979 7415
rect 26835 7387 26979 7395
rect 26835 7386 26871 7387
rect 26943 7386 26979 7387
rect 27045 7420 27082 7421
rect 27045 7419 27083 7420
rect 27045 7411 27109 7419
rect 27045 7391 27054 7411
rect 27074 7397 27109 7411
rect 27129 7397 27132 7417
rect 27074 7392 27132 7397
rect 27074 7391 27109 7392
rect 26341 7319 26381 7375
rect 26514 7354 26551 7383
rect 26515 7352 26551 7354
rect 26515 7330 26706 7352
rect 26732 7351 26769 7383
rect 27045 7379 27109 7391
rect 27149 7353 27176 7531
rect 28034 7506 28076 7551
rect 27008 7351 27176 7353
rect 26732 7341 27176 7351
rect 27317 7447 27504 7471
rect 27535 7452 27928 7472
rect 27948 7452 27951 7472
rect 27535 7447 27951 7452
rect 27317 7376 27354 7447
rect 27535 7446 27876 7447
rect 27469 7386 27500 7387
rect 27317 7356 27326 7376
rect 27346 7356 27354 7376
rect 27317 7346 27354 7356
rect 27413 7376 27500 7386
rect 27413 7356 27422 7376
rect 27442 7356 27500 7376
rect 27413 7347 27500 7356
rect 27413 7346 27450 7347
rect 26338 7314 26381 7319
rect 26729 7325 27176 7341
rect 26729 7319 26757 7325
rect 27008 7324 27176 7325
rect 26338 7311 26488 7314
rect 26729 7311 26756 7319
rect 26338 7309 26756 7311
rect 26338 7291 26347 7309
rect 26365 7291 26756 7309
rect 27469 7296 27500 7347
rect 27535 7376 27572 7446
rect 27838 7445 27875 7446
rect 27687 7386 27723 7387
rect 27535 7356 27544 7376
rect 27564 7356 27572 7376
rect 27535 7346 27572 7356
rect 27631 7376 27779 7386
rect 27879 7383 27975 7385
rect 27631 7356 27640 7376
rect 27660 7356 27750 7376
rect 27770 7356 27779 7376
rect 27631 7347 27779 7356
rect 27837 7376 27975 7383
rect 27837 7356 27846 7376
rect 27866 7356 27975 7376
rect 27837 7347 27975 7356
rect 27631 7346 27668 7347
rect 27361 7293 27402 7294
rect 26338 7288 26756 7291
rect 26338 7282 26381 7288
rect 26341 7279 26381 7282
rect 27256 7286 27402 7293
rect 26738 7270 26778 7271
rect 26449 7253 26778 7270
rect 27256 7266 27312 7286
rect 27332 7266 27371 7286
rect 27391 7266 27402 7286
rect 27256 7258 27402 7266
rect 27469 7289 27626 7296
rect 27469 7269 27589 7289
rect 27609 7269 27626 7289
rect 27469 7259 27626 7269
rect 27469 7258 27504 7259
rect 26333 7210 26376 7221
rect 26333 7192 26345 7210
rect 26363 7192 26376 7210
rect 26333 7166 26376 7192
rect 26449 7166 26476 7253
rect 26738 7244 26778 7253
rect 25499 7141 25938 7159
rect 24706 7138 24747 7139
rect 24440 7085 24477 7086
rect 24133 7076 24271 7085
rect 24133 7056 24242 7076
rect 24262 7056 24271 7076
rect 24133 7049 24271 7056
rect 24329 7076 24477 7085
rect 24329 7056 24338 7076
rect 24358 7056 24448 7076
rect 24468 7056 24477 7076
rect 24133 7047 24229 7049
rect 24329 7046 24477 7056
rect 24536 7076 24573 7086
rect 24536 7056 24544 7076
rect 24564 7056 24573 7076
rect 24385 7045 24421 7046
rect 24233 6986 24270 6987
rect 24536 6986 24573 7056
rect 24608 7085 24639 7136
rect 25499 7123 25899 7141
rect 25917 7123 25938 7141
rect 25499 7117 25938 7123
rect 25505 7113 25938 7117
rect 26333 7145 26476 7166
rect 26520 7218 26554 7234
rect 26738 7224 27131 7244
rect 27151 7224 27154 7244
rect 27469 7237 27500 7258
rect 27687 7237 27723 7347
rect 27742 7346 27779 7347
rect 27838 7346 27875 7347
rect 27798 7287 27888 7293
rect 27798 7267 27807 7287
rect 27827 7285 27888 7287
rect 27827 7267 27852 7285
rect 27798 7265 27852 7267
rect 27872 7265 27888 7285
rect 27798 7259 27888 7265
rect 27312 7236 27349 7237
rect 26738 7219 27154 7224
rect 27311 7227 27349 7236
rect 26738 7218 27079 7219
rect 26520 7148 26557 7218
rect 26672 7158 26703 7159
rect 26333 7143 26470 7145
rect 25884 7111 25936 7113
rect 26333 7101 26376 7143
rect 26520 7128 26529 7148
rect 26549 7128 26557 7148
rect 26520 7118 26557 7128
rect 26616 7148 26703 7158
rect 26616 7128 26625 7148
rect 26645 7128 26703 7148
rect 26616 7119 26703 7128
rect 26616 7118 26653 7119
rect 26331 7091 26376 7101
rect 24658 7085 24695 7086
rect 24608 7076 24695 7085
rect 24608 7056 24666 7076
rect 24686 7056 24695 7076
rect 24608 7046 24695 7056
rect 24754 7076 24791 7086
rect 24754 7056 24762 7076
rect 24782 7056 24791 7076
rect 26331 7073 26340 7091
rect 26358 7073 26376 7091
rect 26331 7067 26376 7073
rect 26672 7068 26703 7119
rect 26738 7148 26775 7218
rect 27041 7217 27078 7218
rect 27311 7207 27320 7227
rect 27340 7207 27349 7227
rect 27311 7199 27349 7207
rect 27415 7231 27500 7237
rect 27530 7236 27567 7237
rect 27415 7211 27423 7231
rect 27443 7211 27500 7231
rect 27415 7203 27500 7211
rect 27529 7227 27567 7236
rect 27529 7207 27538 7227
rect 27558 7207 27567 7227
rect 27415 7202 27451 7203
rect 27529 7199 27567 7207
rect 27633 7231 27777 7237
rect 27633 7211 27641 7231
rect 27661 7228 27749 7231
rect 27661 7211 27696 7228
rect 27633 7210 27696 7211
rect 27715 7211 27749 7228
rect 27769 7211 27777 7231
rect 27715 7210 27777 7211
rect 27633 7203 27777 7210
rect 27633 7202 27669 7203
rect 27741 7202 27777 7203
rect 27843 7236 27880 7237
rect 27843 7235 27881 7236
rect 27903 7235 27930 7239
rect 27843 7233 27930 7235
rect 27843 7227 27907 7233
rect 27843 7207 27852 7227
rect 27872 7213 27907 7227
rect 27927 7213 27930 7233
rect 27872 7208 27930 7213
rect 27872 7207 27907 7208
rect 27312 7170 27349 7199
rect 27313 7168 27349 7170
rect 26890 7158 26926 7159
rect 26738 7128 26747 7148
rect 26767 7128 26775 7148
rect 26738 7118 26775 7128
rect 26834 7148 26982 7158
rect 27082 7155 27178 7157
rect 26834 7128 26843 7148
rect 26863 7128 26953 7148
rect 26973 7128 26982 7148
rect 26834 7119 26982 7128
rect 27040 7148 27178 7155
rect 27040 7128 27049 7148
rect 27069 7128 27178 7148
rect 27313 7146 27504 7168
rect 27530 7167 27567 7199
rect 27843 7195 27907 7207
rect 27947 7169 27974 7347
rect 27806 7167 27974 7169
rect 27530 7141 27974 7167
rect 27040 7119 27178 7128
rect 26834 7118 26871 7119
rect 26331 7064 26368 7067
rect 26564 7065 26605 7066
rect 24608 7045 24639 7046
rect 24232 6985 24573 6986
rect 24754 6985 24791 7056
rect 26456 7058 26605 7065
rect 25887 7046 25924 7051
rect 24157 6980 24573 6985
rect 24157 6960 24160 6980
rect 24180 6960 24573 6980
rect 24604 6961 24791 6985
rect 25878 7042 25925 7046
rect 25878 7024 25897 7042
rect 25915 7024 25925 7042
rect 26456 7038 26515 7058
rect 26535 7038 26574 7058
rect 26594 7038 26605 7058
rect 26456 7030 26605 7038
rect 26672 7061 26829 7068
rect 26672 7041 26792 7061
rect 26812 7041 26829 7061
rect 26672 7031 26829 7041
rect 26672 7030 26707 7031
rect 25878 6976 25925 7024
rect 26672 7009 26703 7030
rect 26890 7009 26926 7119
rect 26945 7118 26982 7119
rect 27041 7118 27078 7119
rect 27001 7059 27091 7065
rect 27001 7039 27010 7059
rect 27030 7057 27091 7059
rect 27030 7039 27055 7057
rect 27001 7037 27055 7039
rect 27075 7037 27091 7057
rect 27001 7031 27091 7037
rect 26515 7008 26552 7009
rect 25502 6973 25925 6976
rect 24377 6959 24442 6960
rect 25480 6943 25925 6973
rect 26327 7000 26365 7002
rect 26327 6992 26370 7000
rect 26327 6974 26338 6992
rect 26356 6974 26370 6992
rect 26327 6947 26370 6974
rect 26514 6999 26552 7008
rect 26514 6979 26523 6999
rect 26543 6979 26552 6999
rect 26514 6971 26552 6979
rect 26618 7003 26703 7009
rect 26733 7008 26770 7009
rect 26618 6983 26626 7003
rect 26646 6983 26703 7003
rect 26618 6975 26703 6983
rect 26732 6999 26770 7008
rect 26732 6979 26741 6999
rect 26761 6979 26770 6999
rect 26618 6974 26654 6975
rect 26732 6971 26770 6979
rect 26836 7007 26980 7009
rect 26836 7003 26888 7007
rect 26836 6983 26844 7003
rect 26864 6987 26888 7003
rect 26908 7003 26980 7007
rect 26908 6987 26952 7003
rect 26864 6983 26952 6987
rect 26972 6983 26980 7003
rect 26836 6975 26980 6983
rect 26836 6974 26872 6975
rect 26944 6974 26980 6975
rect 27046 7008 27083 7009
rect 27046 7007 27084 7008
rect 27046 6999 27110 7007
rect 27046 6979 27055 6999
rect 27075 6985 27110 6999
rect 27130 6985 27133 7005
rect 27075 6980 27133 6985
rect 27075 6979 27110 6980
rect 24573 6927 24613 6935
rect 24573 6905 24581 6927
rect 24605 6905 24613 6927
rect 24178 6676 24215 6682
rect 24178 6657 24186 6676
rect 24207 6657 24215 6676
rect 24178 6649 24215 6657
rect 24182 6316 24215 6649
rect 24279 6681 24447 6682
rect 24573 6681 24613 6905
rect 25076 6909 25244 6910
rect 25480 6909 25521 6943
rect 25878 6922 25925 6943
rect 25076 6899 25521 6909
rect 25593 6907 25736 6908
rect 25076 6883 25520 6899
rect 25076 6881 25244 6883
rect 25440 6882 25520 6883
rect 25593 6882 25738 6907
rect 25880 6882 25925 6922
rect 25076 6703 25103 6881
rect 25143 6843 25207 6855
rect 25483 6851 25520 6882
rect 25701 6851 25738 6882
rect 25883 6875 25925 6882
rect 26328 6940 26370 6947
rect 26515 6940 26552 6971
rect 26733 6940 26770 6971
rect 27046 6967 27110 6979
rect 27150 6941 27177 7119
rect 26328 6900 26373 6940
rect 26515 6915 26660 6940
rect 26733 6939 26813 6940
rect 27009 6939 27177 6941
rect 26733 6923 27177 6939
rect 26517 6914 26660 6915
rect 26732 6913 27177 6923
rect 26328 6879 26375 6900
rect 26732 6879 26773 6913
rect 27009 6912 27177 6913
rect 27640 6917 27680 7141
rect 27806 7140 27974 7141
rect 28038 7173 28071 7506
rect 28676 7505 28703 7683
rect 28743 7645 28807 7657
rect 29083 7653 29120 7685
rect 29146 7684 29337 7706
rect 29472 7704 29581 7724
rect 29601 7704 29610 7724
rect 29472 7697 29610 7704
rect 29668 7724 29816 7733
rect 29668 7704 29677 7724
rect 29697 7704 29787 7724
rect 29807 7704 29816 7724
rect 29472 7695 29568 7697
rect 29668 7694 29816 7704
rect 29875 7724 29912 7734
rect 29875 7704 29883 7724
rect 29903 7704 29912 7724
rect 29724 7693 29760 7694
rect 29301 7682 29337 7684
rect 29301 7653 29338 7682
rect 28743 7644 28778 7645
rect 28720 7639 28778 7644
rect 28720 7619 28723 7639
rect 28743 7625 28778 7639
rect 28798 7625 28807 7645
rect 28743 7617 28807 7625
rect 28769 7616 28807 7617
rect 28770 7615 28807 7616
rect 28873 7649 28909 7650
rect 28981 7649 29017 7650
rect 28873 7641 29017 7649
rect 28873 7621 28881 7641
rect 28901 7640 28989 7641
rect 28901 7621 28936 7640
rect 28957 7621 28989 7640
rect 29009 7621 29017 7641
rect 28873 7615 29017 7621
rect 29083 7645 29121 7653
rect 29199 7649 29235 7650
rect 29083 7625 29092 7645
rect 29112 7625 29121 7645
rect 29083 7616 29121 7625
rect 29150 7641 29235 7649
rect 29150 7621 29207 7641
rect 29227 7621 29235 7641
rect 29083 7615 29120 7616
rect 29150 7615 29235 7621
rect 29301 7645 29339 7653
rect 29301 7625 29310 7645
rect 29330 7625 29339 7645
rect 29572 7634 29609 7635
rect 29875 7634 29912 7704
rect 29947 7733 29978 7784
rect 30274 7779 30319 7785
rect 30274 7761 30292 7779
rect 30310 7761 30319 7779
rect 31780 7779 31789 7799
rect 31809 7779 31817 7799
rect 31780 7769 31817 7779
rect 31876 7799 31963 7809
rect 31876 7779 31885 7799
rect 31905 7779 31963 7799
rect 31876 7770 31963 7779
rect 31876 7769 31913 7770
rect 30274 7751 30319 7761
rect 29997 7733 30034 7734
rect 29947 7724 30034 7733
rect 29947 7704 30005 7724
rect 30025 7704 30034 7724
rect 29947 7694 30034 7704
rect 30093 7724 30130 7734
rect 30093 7704 30101 7724
rect 30121 7704 30130 7724
rect 30274 7709 30317 7751
rect 30701 7740 30753 7742
rect 30180 7707 30317 7709
rect 29947 7693 29978 7694
rect 30093 7634 30130 7704
rect 29571 7633 29912 7634
rect 29301 7616 29339 7625
rect 29496 7628 29912 7633
rect 29301 7615 29338 7616
rect 28762 7587 28852 7593
rect 28762 7567 28778 7587
rect 28798 7585 28852 7587
rect 28798 7567 28823 7585
rect 28762 7565 28823 7567
rect 28843 7565 28852 7585
rect 28762 7559 28852 7565
rect 28775 7505 28812 7506
rect 28871 7505 28908 7506
rect 28927 7505 28963 7615
rect 29150 7594 29181 7615
rect 29496 7608 29499 7628
rect 29519 7608 29912 7628
rect 30096 7618 30130 7634
rect 30174 7686 30317 7707
rect 30699 7736 31132 7740
rect 30699 7730 31138 7736
rect 30699 7712 30720 7730
rect 30738 7712 31138 7730
rect 31932 7719 31963 7770
rect 31998 7799 32035 7869
rect 32301 7868 32338 7869
rect 32150 7809 32186 7810
rect 31998 7779 32007 7799
rect 32027 7779 32035 7799
rect 31998 7769 32035 7779
rect 32094 7799 32242 7809
rect 32342 7806 32438 7808
rect 32094 7779 32103 7799
rect 32123 7779 32213 7799
rect 32233 7779 32242 7799
rect 32094 7770 32242 7779
rect 32300 7799 32438 7806
rect 32300 7779 32309 7799
rect 32329 7779 32438 7799
rect 32300 7770 32438 7779
rect 32094 7769 32131 7770
rect 31824 7716 31865 7717
rect 30699 7694 31138 7712
rect 29872 7599 29912 7608
rect 30174 7599 30201 7686
rect 30274 7660 30317 7686
rect 30274 7642 30287 7660
rect 30305 7642 30317 7660
rect 30274 7631 30317 7642
rect 29146 7593 29181 7594
rect 29024 7583 29181 7593
rect 29024 7563 29041 7583
rect 29061 7563 29181 7583
rect 29024 7556 29181 7563
rect 29248 7586 29397 7594
rect 29248 7566 29259 7586
rect 29279 7566 29318 7586
rect 29338 7566 29397 7586
rect 29872 7582 30201 7599
rect 29872 7581 29912 7582
rect 29248 7559 29397 7566
rect 30269 7570 30309 7573
rect 30269 7564 30312 7570
rect 29894 7561 30312 7564
rect 29248 7558 29289 7559
rect 28982 7505 29019 7506
rect 28675 7496 28813 7505
rect 28538 7486 28574 7492
rect 28538 7468 28543 7486
rect 28565 7468 28574 7486
rect 28538 7464 28574 7468
rect 28675 7476 28784 7496
rect 28804 7476 28813 7496
rect 28675 7469 28813 7476
rect 28871 7496 29019 7505
rect 28871 7476 28880 7496
rect 28900 7476 28990 7496
rect 29010 7476 29019 7496
rect 28675 7467 28771 7469
rect 28871 7466 29019 7476
rect 29078 7496 29115 7506
rect 29078 7476 29086 7496
rect 29106 7476 29115 7496
rect 28927 7465 28963 7466
rect 28541 7305 28574 7464
rect 28775 7406 28812 7407
rect 29078 7406 29115 7476
rect 29150 7505 29181 7556
rect 29894 7543 30285 7561
rect 30303 7543 30312 7561
rect 29894 7541 30312 7543
rect 29894 7533 29921 7541
rect 30162 7538 30312 7541
rect 29474 7527 29642 7528
rect 29893 7527 29921 7533
rect 29474 7511 29921 7527
rect 30269 7533 30312 7538
rect 29200 7505 29237 7506
rect 29150 7496 29237 7505
rect 29150 7476 29208 7496
rect 29228 7476 29237 7496
rect 29150 7466 29237 7476
rect 29296 7496 29333 7506
rect 29296 7476 29304 7496
rect 29324 7476 29333 7496
rect 29150 7465 29181 7466
rect 28774 7405 29115 7406
rect 29296 7405 29333 7476
rect 28699 7400 29115 7405
rect 28699 7380 28702 7400
rect 28722 7380 29115 7400
rect 29146 7381 29333 7405
rect 29474 7501 29918 7511
rect 29474 7499 29642 7501
rect 29474 7321 29501 7499
rect 29541 7461 29605 7473
rect 29881 7469 29918 7501
rect 29944 7500 30135 7522
rect 30099 7498 30135 7500
rect 30099 7469 30136 7498
rect 30269 7477 30309 7533
rect 29541 7460 29576 7461
rect 29518 7455 29576 7460
rect 29518 7435 29521 7455
rect 29541 7441 29576 7455
rect 29596 7441 29605 7461
rect 29541 7433 29605 7441
rect 29567 7432 29605 7433
rect 29568 7431 29605 7432
rect 29671 7465 29707 7466
rect 29779 7465 29815 7466
rect 29671 7457 29815 7465
rect 29671 7437 29679 7457
rect 29699 7437 29734 7457
rect 29754 7437 29787 7457
rect 29807 7437 29815 7457
rect 29671 7431 29815 7437
rect 29881 7461 29919 7469
rect 29997 7465 30033 7466
rect 29881 7441 29890 7461
rect 29910 7441 29919 7461
rect 29881 7432 29919 7441
rect 29948 7457 30033 7465
rect 29948 7437 30005 7457
rect 30025 7437 30033 7457
rect 29881 7431 29918 7432
rect 29948 7431 30033 7437
rect 30099 7461 30137 7469
rect 30099 7441 30108 7461
rect 30128 7441 30137 7461
rect 30269 7459 30281 7477
rect 30299 7459 30309 7477
rect 30701 7505 30753 7694
rect 31099 7669 31138 7694
rect 31716 7709 31865 7716
rect 31716 7689 31775 7709
rect 31795 7689 31834 7709
rect 31854 7689 31865 7709
rect 31716 7681 31865 7689
rect 31932 7712 32089 7719
rect 31932 7692 32052 7712
rect 32072 7692 32089 7712
rect 31932 7682 32089 7692
rect 31932 7681 31967 7682
rect 30883 7644 31070 7668
rect 31099 7649 31494 7669
rect 31514 7649 31517 7669
rect 31932 7660 31963 7681
rect 32150 7660 32186 7770
rect 32205 7769 32242 7770
rect 32301 7769 32338 7770
rect 32261 7710 32351 7716
rect 32261 7690 32270 7710
rect 32290 7708 32351 7710
rect 32290 7690 32315 7708
rect 32261 7688 32315 7690
rect 32335 7688 32351 7708
rect 32261 7682 32351 7688
rect 31775 7659 31812 7660
rect 31099 7644 31517 7649
rect 31774 7650 31812 7659
rect 30883 7573 30920 7644
rect 31099 7643 31442 7644
rect 31099 7640 31138 7643
rect 31404 7642 31441 7643
rect 31035 7583 31066 7584
rect 30883 7553 30892 7573
rect 30912 7553 30920 7573
rect 30883 7543 30920 7553
rect 30979 7573 31066 7583
rect 30979 7553 30988 7573
rect 31008 7553 31066 7573
rect 30979 7544 31066 7553
rect 30979 7543 31016 7544
rect 30701 7487 30717 7505
rect 30735 7487 30753 7505
rect 31035 7493 31066 7544
rect 31101 7573 31138 7640
rect 31774 7630 31783 7650
rect 31803 7630 31812 7650
rect 31774 7622 31812 7630
rect 31878 7654 31963 7660
rect 31993 7659 32030 7660
rect 31878 7634 31886 7654
rect 31906 7634 31963 7654
rect 31878 7626 31963 7634
rect 31992 7650 32030 7659
rect 31992 7630 32001 7650
rect 32021 7630 32030 7650
rect 31878 7625 31914 7626
rect 31992 7622 32030 7630
rect 32096 7655 32240 7660
rect 32096 7654 32158 7655
rect 32096 7634 32104 7654
rect 32124 7636 32158 7654
rect 32179 7654 32240 7655
rect 32179 7636 32212 7654
rect 32124 7634 32212 7636
rect 32232 7634 32240 7654
rect 32096 7626 32240 7634
rect 32096 7625 32132 7626
rect 32204 7625 32240 7626
rect 32306 7659 32343 7660
rect 32306 7658 32344 7659
rect 32306 7650 32370 7658
rect 32306 7630 32315 7650
rect 32335 7636 32370 7650
rect 32390 7636 32393 7656
rect 32335 7631 32393 7636
rect 32335 7630 32370 7631
rect 31775 7593 31812 7622
rect 31776 7591 31812 7593
rect 31253 7583 31289 7584
rect 31101 7553 31110 7573
rect 31130 7553 31138 7573
rect 31101 7543 31138 7553
rect 31197 7573 31345 7583
rect 31445 7580 31541 7582
rect 31197 7553 31206 7573
rect 31226 7553 31316 7573
rect 31336 7553 31345 7573
rect 31197 7544 31345 7553
rect 31403 7573 31541 7580
rect 31403 7553 31412 7573
rect 31432 7553 31541 7573
rect 31776 7569 31967 7591
rect 31993 7590 32030 7622
rect 32306 7618 32370 7630
rect 32410 7592 32437 7770
rect 32269 7590 32437 7592
rect 31993 7576 32437 7590
rect 33040 7724 33208 7725
rect 33334 7724 33374 7948
rect 33837 7952 34005 7953
rect 34240 7952 34280 7985
rect 34636 7952 34683 7985
rect 33837 7951 34281 7952
rect 33837 7926 34282 7951
rect 33837 7924 34005 7926
rect 34201 7925 34282 7926
rect 34451 7925 34500 7951
rect 34636 7925 34685 7952
rect 33837 7746 33864 7924
rect 33904 7886 33968 7898
rect 34244 7894 34281 7925
rect 34462 7894 34499 7925
rect 34644 7900 34685 7925
rect 33904 7885 33939 7886
rect 33881 7880 33939 7885
rect 33881 7860 33884 7880
rect 33904 7866 33939 7880
rect 33959 7866 33968 7886
rect 33904 7858 33968 7866
rect 33930 7857 33968 7858
rect 33931 7856 33968 7857
rect 34034 7890 34070 7891
rect 34142 7890 34178 7891
rect 34034 7882 34178 7890
rect 34034 7862 34042 7882
rect 34062 7878 34150 7882
rect 34062 7862 34106 7878
rect 34034 7858 34106 7862
rect 34126 7862 34150 7878
rect 34170 7862 34178 7882
rect 34126 7858 34178 7862
rect 34034 7856 34178 7858
rect 34244 7886 34282 7894
rect 34360 7890 34396 7891
rect 34244 7866 34253 7886
rect 34273 7866 34282 7886
rect 34244 7857 34282 7866
rect 34311 7882 34396 7890
rect 34311 7862 34368 7882
rect 34388 7862 34396 7882
rect 34244 7856 34281 7857
rect 34311 7856 34396 7862
rect 34462 7886 34500 7894
rect 34462 7866 34471 7886
rect 34491 7866 34500 7886
rect 34462 7857 34500 7866
rect 34644 7891 34686 7900
rect 34644 7873 34658 7891
rect 34676 7873 34686 7891
rect 34644 7865 34686 7873
rect 34649 7863 34686 7865
rect 34462 7856 34499 7857
rect 33923 7828 34013 7834
rect 33923 7808 33939 7828
rect 33959 7826 34013 7828
rect 33959 7808 33984 7826
rect 33923 7806 33984 7808
rect 34004 7806 34013 7826
rect 33923 7800 34013 7806
rect 33936 7746 33973 7747
rect 34032 7746 34069 7747
rect 34088 7746 34124 7856
rect 34311 7835 34342 7856
rect 34307 7834 34342 7835
rect 34185 7824 34342 7834
rect 34185 7804 34202 7824
rect 34222 7804 34342 7824
rect 34185 7797 34342 7804
rect 34409 7827 34558 7835
rect 34409 7807 34420 7827
rect 34440 7807 34479 7827
rect 34499 7807 34558 7827
rect 34409 7800 34558 7807
rect 34409 7799 34450 7800
rect 34646 7798 34683 7801
rect 34143 7746 34180 7747
rect 33836 7737 33974 7746
rect 33040 7698 33484 7724
rect 33040 7696 33208 7698
rect 31993 7564 32440 7576
rect 32036 7562 32069 7564
rect 31403 7544 31541 7553
rect 31197 7543 31234 7544
rect 30927 7490 30968 7491
rect 30701 7469 30753 7487
rect 30819 7483 30968 7490
rect 30269 7449 30309 7459
rect 30819 7463 30878 7483
rect 30898 7463 30937 7483
rect 30957 7463 30968 7483
rect 30819 7455 30968 7463
rect 31035 7486 31192 7493
rect 31035 7466 31155 7486
rect 31175 7466 31192 7486
rect 31035 7456 31192 7466
rect 31035 7455 31070 7456
rect 30099 7432 30137 7441
rect 31035 7434 31066 7455
rect 31253 7434 31289 7544
rect 31308 7543 31345 7544
rect 31404 7543 31441 7544
rect 31364 7484 31454 7490
rect 31364 7464 31373 7484
rect 31393 7482 31454 7484
rect 31393 7464 31418 7482
rect 31364 7462 31418 7464
rect 31438 7462 31454 7482
rect 31364 7456 31454 7462
rect 30878 7433 30915 7434
rect 30099 7431 30136 7432
rect 29560 7403 29650 7409
rect 29560 7383 29576 7403
rect 29596 7401 29650 7403
rect 29596 7383 29621 7401
rect 29560 7381 29621 7383
rect 29641 7381 29650 7401
rect 29560 7375 29650 7381
rect 29573 7321 29610 7322
rect 29669 7321 29706 7322
rect 29725 7321 29761 7431
rect 29948 7410 29979 7431
rect 30877 7424 30915 7433
rect 29944 7409 29979 7410
rect 29822 7399 29979 7409
rect 29822 7379 29839 7399
rect 29859 7379 29979 7399
rect 29822 7372 29979 7379
rect 30046 7402 30195 7410
rect 30046 7382 30057 7402
rect 30077 7382 30116 7402
rect 30136 7382 30195 7402
rect 30705 7406 30745 7416
rect 30046 7375 30195 7382
rect 30261 7378 30313 7396
rect 30046 7374 30087 7375
rect 29780 7321 29817 7322
rect 29473 7312 29611 7321
rect 28540 7304 28577 7305
rect 28511 7303 28679 7304
rect 28805 7303 28845 7305
rect 28336 7294 28375 7300
rect 28336 7272 28344 7294
rect 28368 7272 28375 7294
rect 28038 7165 28075 7173
rect 28038 7146 28046 7165
rect 28067 7146 28075 7165
rect 28038 7140 28075 7146
rect 27640 6895 27648 6917
rect 27672 6895 27680 6917
rect 27640 6887 27680 6895
rect 25143 6842 25178 6843
rect 25120 6837 25178 6842
rect 25120 6817 25123 6837
rect 25143 6823 25178 6837
rect 25198 6823 25207 6843
rect 25143 6815 25207 6823
rect 25169 6814 25207 6815
rect 25170 6813 25207 6814
rect 25273 6847 25309 6848
rect 25381 6847 25417 6848
rect 25273 6839 25417 6847
rect 25273 6819 25281 6839
rect 25301 6835 25389 6839
rect 25301 6819 25345 6835
rect 25273 6815 25345 6819
rect 25365 6819 25389 6835
rect 25409 6819 25417 6839
rect 25365 6815 25417 6819
rect 25273 6813 25417 6815
rect 25483 6843 25521 6851
rect 25599 6847 25635 6848
rect 25483 6823 25492 6843
rect 25512 6823 25521 6843
rect 25483 6814 25521 6823
rect 25550 6839 25635 6847
rect 25550 6819 25607 6839
rect 25627 6819 25635 6839
rect 25483 6813 25520 6814
rect 25550 6813 25635 6819
rect 25701 6843 25739 6851
rect 25701 6823 25710 6843
rect 25730 6823 25739 6843
rect 25701 6814 25739 6823
rect 25883 6848 25926 6875
rect 25883 6830 25897 6848
rect 25915 6830 25926 6848
rect 25883 6822 25926 6830
rect 25888 6820 25926 6822
rect 26328 6849 26773 6879
rect 27811 6862 27876 6863
rect 26328 6846 26751 6849
rect 25701 6813 25738 6814
rect 25162 6785 25252 6791
rect 25162 6765 25178 6785
rect 25198 6783 25252 6785
rect 25198 6765 25223 6783
rect 25162 6763 25223 6765
rect 25243 6763 25252 6783
rect 25162 6757 25252 6763
rect 25175 6703 25212 6704
rect 25271 6703 25308 6704
rect 25327 6703 25363 6813
rect 25550 6792 25581 6813
rect 26328 6798 26375 6846
rect 25546 6791 25581 6792
rect 25424 6781 25581 6791
rect 25424 6761 25441 6781
rect 25461 6761 25581 6781
rect 25424 6754 25581 6761
rect 25648 6784 25797 6792
rect 25648 6764 25659 6784
rect 25679 6764 25718 6784
rect 25738 6764 25797 6784
rect 26328 6780 26338 6798
rect 26356 6780 26375 6798
rect 26328 6776 26375 6780
rect 27462 6837 27649 6861
rect 27680 6842 28073 6862
rect 28093 6842 28096 6862
rect 27680 6837 28096 6842
rect 26329 6771 26366 6776
rect 25648 6757 25797 6764
rect 27462 6766 27499 6837
rect 27680 6836 28021 6837
rect 27614 6776 27645 6777
rect 25648 6756 25689 6757
rect 25885 6755 25922 6758
rect 25382 6703 25419 6704
rect 25075 6694 25213 6703
rect 24279 6655 24723 6681
rect 24279 6653 24447 6655
rect 24279 6475 24306 6653
rect 24346 6615 24410 6627
rect 24686 6623 24723 6655
rect 24749 6654 24940 6676
rect 25075 6674 25184 6694
rect 25204 6674 25213 6694
rect 25075 6667 25213 6674
rect 25271 6694 25419 6703
rect 25271 6674 25280 6694
rect 25300 6674 25390 6694
rect 25410 6674 25419 6694
rect 25075 6665 25171 6667
rect 25271 6664 25419 6674
rect 25478 6694 25515 6704
rect 25478 6674 25486 6694
rect 25506 6674 25515 6694
rect 25327 6663 25363 6664
rect 24904 6652 24940 6654
rect 24904 6623 24941 6652
rect 24346 6614 24381 6615
rect 24323 6609 24381 6614
rect 24323 6589 24326 6609
rect 24346 6595 24381 6609
rect 24401 6595 24410 6615
rect 24346 6589 24410 6595
rect 24323 6587 24410 6589
rect 24323 6583 24350 6587
rect 24372 6586 24410 6587
rect 24373 6585 24410 6586
rect 24476 6619 24512 6620
rect 24584 6619 24620 6620
rect 24476 6612 24620 6619
rect 24476 6611 24538 6612
rect 24476 6591 24484 6611
rect 24504 6594 24538 6611
rect 24557 6611 24620 6612
rect 24557 6594 24592 6611
rect 24504 6591 24592 6594
rect 24612 6591 24620 6611
rect 24476 6585 24620 6591
rect 24686 6615 24724 6623
rect 24802 6619 24838 6620
rect 24686 6595 24695 6615
rect 24715 6595 24724 6615
rect 24686 6586 24724 6595
rect 24753 6611 24838 6619
rect 24753 6591 24810 6611
rect 24830 6591 24838 6611
rect 24686 6585 24723 6586
rect 24753 6585 24838 6591
rect 24904 6615 24942 6623
rect 24904 6595 24913 6615
rect 24933 6595 24942 6615
rect 25175 6604 25212 6605
rect 25478 6604 25515 6674
rect 25550 6703 25581 6754
rect 25877 6749 25922 6755
rect 25877 6731 25895 6749
rect 25913 6731 25922 6749
rect 27462 6746 27471 6766
rect 27491 6746 27499 6766
rect 27462 6736 27499 6746
rect 27558 6766 27645 6776
rect 27558 6746 27567 6766
rect 27587 6746 27645 6766
rect 27558 6737 27645 6746
rect 27558 6736 27595 6737
rect 25877 6721 25922 6731
rect 25600 6703 25637 6704
rect 25550 6694 25637 6703
rect 25550 6674 25608 6694
rect 25628 6674 25637 6694
rect 25550 6664 25637 6674
rect 25696 6694 25733 6704
rect 25696 6674 25704 6694
rect 25724 6674 25733 6694
rect 25877 6679 25920 6721
rect 26317 6709 26369 6711
rect 25783 6677 25920 6679
rect 25550 6663 25581 6664
rect 25696 6604 25733 6674
rect 25174 6603 25515 6604
rect 24904 6586 24942 6595
rect 25099 6598 25515 6603
rect 24904 6585 24941 6586
rect 24365 6557 24455 6563
rect 24365 6537 24381 6557
rect 24401 6555 24455 6557
rect 24401 6537 24426 6555
rect 24365 6535 24426 6537
rect 24446 6535 24455 6555
rect 24365 6529 24455 6535
rect 24378 6475 24415 6476
rect 24474 6475 24511 6476
rect 24530 6475 24566 6585
rect 24753 6564 24784 6585
rect 25099 6578 25102 6598
rect 25122 6578 25515 6598
rect 25699 6588 25733 6604
rect 25777 6656 25920 6677
rect 26315 6705 26748 6709
rect 26315 6699 26754 6705
rect 26315 6681 26336 6699
rect 26354 6681 26754 6699
rect 27614 6686 27645 6737
rect 27680 6766 27717 6836
rect 27983 6835 28020 6836
rect 27832 6776 27868 6777
rect 27680 6746 27689 6766
rect 27709 6746 27717 6766
rect 27680 6736 27717 6746
rect 27776 6766 27924 6776
rect 28024 6773 28120 6775
rect 27776 6746 27785 6766
rect 27805 6746 27895 6766
rect 27915 6746 27924 6766
rect 27776 6737 27924 6746
rect 27982 6766 28120 6773
rect 27982 6746 27991 6766
rect 28011 6746 28120 6766
rect 27982 6737 28120 6746
rect 27776 6736 27813 6737
rect 27506 6683 27547 6684
rect 26315 6663 26754 6681
rect 25475 6569 25515 6578
rect 25777 6569 25804 6656
rect 25877 6630 25920 6656
rect 25877 6612 25890 6630
rect 25908 6612 25920 6630
rect 25877 6601 25920 6612
rect 24749 6563 24784 6564
rect 24627 6553 24784 6563
rect 24627 6533 24644 6553
rect 24664 6533 24784 6553
rect 24627 6526 24784 6533
rect 24851 6556 24997 6564
rect 24851 6536 24862 6556
rect 24882 6536 24921 6556
rect 24941 6536 24997 6556
rect 25475 6552 25804 6569
rect 25475 6551 25515 6552
rect 24851 6529 24997 6536
rect 25872 6540 25912 6543
rect 25872 6534 25915 6540
rect 25497 6531 25915 6534
rect 24851 6528 24892 6529
rect 24585 6475 24622 6476
rect 24278 6466 24416 6475
rect 24278 6446 24387 6466
rect 24407 6446 24416 6466
rect 24278 6439 24416 6446
rect 24474 6466 24622 6475
rect 24474 6446 24483 6466
rect 24503 6446 24593 6466
rect 24613 6446 24622 6466
rect 24278 6437 24374 6439
rect 24474 6436 24622 6446
rect 24681 6466 24718 6476
rect 24681 6446 24689 6466
rect 24709 6446 24718 6466
rect 24530 6435 24566 6436
rect 24378 6376 24415 6377
rect 24681 6376 24718 6446
rect 24753 6475 24784 6526
rect 25497 6513 25888 6531
rect 25906 6513 25915 6531
rect 25497 6511 25915 6513
rect 25497 6503 25524 6511
rect 25765 6508 25915 6511
rect 25077 6497 25245 6498
rect 25496 6497 25524 6503
rect 25077 6481 25524 6497
rect 25872 6503 25915 6508
rect 24803 6475 24840 6476
rect 24753 6466 24840 6475
rect 24753 6446 24811 6466
rect 24831 6446 24840 6466
rect 24753 6436 24840 6446
rect 24899 6466 24936 6476
rect 24899 6446 24907 6466
rect 24927 6446 24936 6466
rect 24753 6435 24784 6436
rect 24377 6375 24718 6376
rect 24899 6375 24936 6446
rect 24302 6370 24718 6375
rect 24302 6350 24305 6370
rect 24325 6350 24718 6370
rect 24749 6351 24936 6375
rect 25077 6471 25521 6481
rect 25077 6469 25245 6471
rect 24177 6271 24219 6316
rect 25077 6291 25104 6469
rect 25144 6431 25208 6443
rect 25484 6439 25521 6471
rect 25547 6470 25738 6492
rect 25702 6468 25738 6470
rect 25702 6439 25739 6468
rect 25872 6447 25912 6503
rect 25144 6430 25179 6431
rect 25121 6425 25179 6430
rect 25121 6405 25124 6425
rect 25144 6411 25179 6425
rect 25199 6411 25208 6431
rect 25144 6403 25208 6411
rect 25170 6402 25208 6403
rect 25171 6401 25208 6402
rect 25274 6435 25310 6436
rect 25382 6435 25418 6436
rect 25274 6427 25418 6435
rect 25274 6407 25282 6427
rect 25302 6407 25337 6427
rect 25357 6407 25390 6427
rect 25410 6407 25418 6427
rect 25274 6401 25418 6407
rect 25484 6431 25522 6439
rect 25600 6435 25636 6436
rect 25484 6411 25493 6431
rect 25513 6411 25522 6431
rect 25484 6402 25522 6411
rect 25551 6427 25636 6435
rect 25551 6407 25608 6427
rect 25628 6407 25636 6427
rect 25484 6401 25521 6402
rect 25551 6401 25636 6407
rect 25702 6431 25740 6439
rect 25702 6411 25711 6431
rect 25731 6411 25740 6431
rect 25872 6429 25884 6447
rect 25902 6429 25912 6447
rect 26317 6474 26369 6663
rect 26715 6638 26754 6663
rect 27398 6676 27547 6683
rect 27398 6656 27457 6676
rect 27477 6656 27516 6676
rect 27536 6656 27547 6676
rect 27398 6648 27547 6656
rect 27614 6679 27771 6686
rect 27614 6659 27734 6679
rect 27754 6659 27771 6679
rect 27614 6649 27771 6659
rect 27614 6648 27649 6649
rect 26499 6613 26686 6637
rect 26715 6618 27110 6638
rect 27130 6618 27133 6638
rect 27614 6627 27645 6648
rect 27832 6627 27868 6737
rect 27887 6736 27924 6737
rect 27983 6736 28020 6737
rect 27943 6677 28033 6683
rect 27943 6657 27952 6677
rect 27972 6675 28033 6677
rect 27972 6657 27997 6675
rect 27943 6655 27997 6657
rect 28017 6655 28033 6675
rect 27943 6649 28033 6655
rect 27457 6626 27494 6627
rect 26715 6613 27133 6618
rect 27456 6617 27494 6626
rect 26499 6542 26536 6613
rect 26715 6612 27058 6613
rect 26715 6609 26754 6612
rect 27020 6611 27057 6612
rect 26651 6552 26682 6553
rect 26499 6522 26508 6542
rect 26528 6522 26536 6542
rect 26499 6512 26536 6522
rect 26595 6542 26682 6552
rect 26595 6522 26604 6542
rect 26624 6522 26682 6542
rect 26595 6513 26682 6522
rect 26595 6512 26632 6513
rect 26317 6456 26333 6474
rect 26351 6456 26369 6474
rect 26651 6462 26682 6513
rect 26717 6542 26754 6609
rect 27456 6597 27465 6617
rect 27485 6597 27494 6617
rect 27456 6589 27494 6597
rect 27560 6621 27645 6627
rect 27675 6626 27712 6627
rect 27560 6601 27568 6621
rect 27588 6601 27645 6621
rect 27560 6593 27645 6601
rect 27674 6617 27712 6626
rect 27674 6597 27683 6617
rect 27703 6597 27712 6617
rect 27560 6592 27596 6593
rect 27674 6589 27712 6597
rect 27778 6621 27922 6627
rect 27778 6601 27786 6621
rect 27806 6620 27894 6621
rect 27806 6602 27841 6620
rect 27859 6602 27894 6620
rect 27806 6601 27894 6602
rect 27914 6601 27922 6621
rect 27778 6593 27922 6601
rect 27778 6592 27814 6593
rect 27886 6592 27922 6593
rect 27988 6626 28025 6627
rect 27988 6625 28026 6626
rect 27988 6617 28052 6625
rect 27988 6597 27997 6617
rect 28017 6603 28052 6617
rect 28072 6603 28075 6623
rect 28017 6598 28075 6603
rect 28017 6597 28052 6598
rect 27457 6560 27494 6589
rect 27458 6558 27494 6560
rect 26869 6552 26905 6553
rect 26717 6522 26726 6542
rect 26746 6522 26754 6542
rect 26717 6512 26754 6522
rect 26813 6542 26961 6552
rect 27061 6549 27157 6551
rect 26813 6522 26822 6542
rect 26842 6522 26932 6542
rect 26952 6522 26961 6542
rect 26813 6513 26961 6522
rect 27019 6542 27157 6549
rect 27019 6522 27028 6542
rect 27048 6522 27157 6542
rect 27458 6536 27649 6558
rect 27675 6557 27712 6589
rect 27988 6585 28052 6597
rect 28092 6561 28119 6737
rect 28038 6559 28119 6561
rect 27951 6557 28119 6559
rect 27675 6531 28119 6557
rect 27785 6529 27825 6531
rect 27951 6530 28119 6531
rect 27019 6513 27157 6522
rect 28060 6528 28119 6530
rect 26813 6512 26850 6513
rect 26543 6459 26584 6460
rect 26317 6438 26369 6456
rect 26435 6452 26584 6459
rect 25872 6419 25912 6429
rect 26435 6432 26494 6452
rect 26514 6432 26553 6452
rect 26573 6432 26584 6452
rect 26435 6424 26584 6432
rect 26651 6455 26808 6462
rect 26651 6435 26771 6455
rect 26791 6435 26808 6455
rect 26651 6425 26808 6435
rect 26651 6424 26686 6425
rect 25702 6402 25740 6411
rect 26651 6403 26682 6424
rect 26869 6403 26905 6513
rect 26924 6512 26961 6513
rect 27020 6512 27057 6513
rect 26980 6453 27070 6459
rect 26980 6433 26989 6453
rect 27009 6451 27070 6453
rect 27009 6433 27034 6451
rect 26980 6431 27034 6433
rect 27054 6431 27070 6451
rect 26980 6425 27070 6431
rect 26494 6402 26531 6403
rect 25702 6401 25739 6402
rect 25163 6373 25253 6379
rect 25163 6353 25179 6373
rect 25199 6371 25253 6373
rect 25199 6353 25224 6371
rect 25163 6351 25224 6353
rect 25244 6351 25253 6371
rect 25163 6345 25253 6351
rect 25176 6291 25213 6292
rect 25272 6291 25309 6292
rect 25328 6291 25364 6401
rect 25551 6380 25582 6401
rect 26493 6393 26531 6402
rect 25547 6379 25582 6380
rect 25425 6369 25582 6379
rect 25425 6349 25442 6369
rect 25462 6349 25582 6369
rect 25425 6342 25582 6349
rect 25649 6372 25798 6380
rect 25649 6352 25660 6372
rect 25680 6352 25719 6372
rect 25739 6352 25798 6372
rect 26321 6375 26361 6385
rect 25649 6345 25798 6352
rect 25864 6348 25916 6366
rect 25649 6344 25690 6345
rect 25383 6291 25420 6292
rect 25076 6282 25214 6291
rect 24548 6271 24581 6273
rect 24177 6259 24624 6271
rect 24180 6245 24624 6259
rect 24180 6243 24348 6245
rect 24180 6065 24207 6243
rect 24247 6205 24311 6217
rect 24587 6213 24624 6245
rect 24650 6244 24841 6266
rect 25076 6262 25185 6282
rect 25205 6262 25214 6282
rect 25076 6255 25214 6262
rect 25272 6282 25420 6291
rect 25272 6262 25281 6282
rect 25301 6262 25391 6282
rect 25411 6262 25420 6282
rect 25076 6253 25172 6255
rect 25272 6252 25420 6262
rect 25479 6282 25516 6292
rect 25479 6262 25487 6282
rect 25507 6262 25516 6282
rect 25328 6251 25364 6252
rect 24805 6242 24841 6244
rect 24805 6213 24842 6242
rect 24247 6204 24282 6205
rect 24224 6199 24282 6204
rect 24224 6179 24227 6199
rect 24247 6185 24282 6199
rect 24302 6185 24311 6205
rect 24247 6177 24311 6185
rect 24273 6176 24311 6177
rect 24274 6175 24311 6176
rect 24377 6209 24413 6210
rect 24485 6209 24521 6210
rect 24377 6201 24521 6209
rect 24377 6181 24385 6201
rect 24405 6199 24493 6201
rect 24405 6181 24438 6199
rect 24377 6180 24438 6181
rect 24459 6181 24493 6199
rect 24513 6181 24521 6201
rect 24459 6180 24521 6181
rect 24377 6175 24521 6180
rect 24587 6205 24625 6213
rect 24703 6209 24739 6210
rect 24587 6185 24596 6205
rect 24616 6185 24625 6205
rect 24587 6176 24625 6185
rect 24654 6201 24739 6209
rect 24654 6181 24711 6201
rect 24731 6181 24739 6201
rect 24587 6175 24624 6176
rect 24654 6175 24739 6181
rect 24805 6205 24843 6213
rect 24805 6185 24814 6205
rect 24834 6185 24843 6205
rect 25479 6195 25516 6262
rect 25551 6291 25582 6342
rect 25864 6330 25882 6348
rect 25900 6330 25916 6348
rect 25601 6291 25638 6292
rect 25551 6282 25638 6291
rect 25551 6262 25609 6282
rect 25629 6262 25638 6282
rect 25551 6252 25638 6262
rect 25697 6282 25734 6292
rect 25697 6262 25705 6282
rect 25725 6262 25734 6282
rect 25551 6251 25582 6252
rect 25176 6192 25213 6193
rect 25479 6192 25518 6195
rect 25175 6191 25518 6192
rect 25697 6191 25734 6262
rect 24805 6176 24843 6185
rect 25100 6186 25518 6191
rect 24805 6175 24842 6176
rect 24266 6147 24356 6153
rect 24266 6127 24282 6147
rect 24302 6145 24356 6147
rect 24302 6127 24327 6145
rect 24266 6125 24327 6127
rect 24347 6125 24356 6145
rect 24266 6119 24356 6125
rect 24279 6065 24316 6066
rect 24375 6065 24412 6066
rect 24431 6065 24467 6175
rect 24654 6154 24685 6175
rect 25100 6166 25103 6186
rect 25123 6166 25518 6186
rect 25547 6167 25734 6191
rect 24650 6153 24685 6154
rect 24528 6143 24685 6153
rect 24528 6123 24545 6143
rect 24565 6123 24685 6143
rect 24528 6116 24685 6123
rect 24752 6146 24901 6154
rect 24752 6126 24763 6146
rect 24783 6126 24822 6146
rect 24842 6126 24901 6146
rect 24752 6119 24901 6126
rect 25479 6141 25518 6166
rect 25864 6141 25916 6330
rect 26321 6357 26331 6375
rect 26349 6357 26361 6375
rect 26493 6373 26502 6393
rect 26522 6373 26531 6393
rect 26493 6365 26531 6373
rect 26597 6397 26682 6403
rect 26712 6402 26749 6403
rect 26597 6377 26605 6397
rect 26625 6377 26682 6397
rect 26597 6369 26682 6377
rect 26711 6393 26749 6402
rect 26711 6373 26720 6393
rect 26740 6373 26749 6393
rect 26597 6368 26633 6369
rect 26711 6365 26749 6373
rect 26815 6397 26959 6403
rect 26815 6377 26823 6397
rect 26843 6377 26876 6397
rect 26896 6377 26931 6397
rect 26951 6377 26959 6397
rect 26815 6369 26959 6377
rect 26815 6368 26851 6369
rect 26923 6368 26959 6369
rect 27025 6402 27062 6403
rect 27025 6401 27063 6402
rect 27025 6393 27089 6401
rect 27025 6373 27034 6393
rect 27054 6379 27089 6393
rect 27109 6379 27112 6399
rect 27054 6374 27112 6379
rect 27054 6373 27089 6374
rect 26321 6301 26361 6357
rect 26494 6336 26531 6365
rect 26495 6334 26531 6336
rect 26495 6312 26686 6334
rect 26712 6333 26749 6365
rect 27025 6361 27089 6373
rect 27129 6335 27156 6513
rect 28060 6510 28089 6528
rect 26988 6333 27156 6335
rect 26712 6323 27156 6333
rect 27297 6429 27484 6453
rect 27515 6434 27908 6454
rect 27928 6434 27931 6454
rect 27515 6429 27931 6434
rect 27297 6358 27334 6429
rect 27515 6428 27856 6429
rect 27449 6368 27480 6369
rect 27297 6338 27306 6358
rect 27326 6338 27334 6358
rect 27297 6328 27334 6338
rect 27393 6358 27480 6368
rect 27393 6338 27402 6358
rect 27422 6338 27480 6358
rect 27393 6329 27480 6338
rect 27393 6328 27430 6329
rect 26318 6296 26361 6301
rect 26709 6307 27156 6323
rect 26709 6301 26737 6307
rect 26988 6306 27156 6307
rect 26318 6293 26468 6296
rect 26709 6293 26736 6301
rect 26318 6291 26736 6293
rect 26318 6273 26327 6291
rect 26345 6273 26736 6291
rect 27449 6278 27480 6329
rect 27515 6358 27552 6428
rect 27818 6427 27855 6428
rect 27667 6368 27703 6369
rect 27515 6338 27524 6358
rect 27544 6338 27552 6358
rect 27515 6328 27552 6338
rect 27611 6358 27759 6368
rect 27859 6365 27955 6367
rect 27611 6338 27620 6358
rect 27640 6338 27730 6358
rect 27750 6338 27759 6358
rect 27611 6329 27759 6338
rect 27817 6358 27955 6365
rect 27817 6338 27826 6358
rect 27846 6338 27955 6358
rect 27817 6329 27955 6338
rect 27611 6328 27648 6329
rect 27341 6275 27382 6276
rect 26318 6270 26736 6273
rect 26318 6264 26361 6270
rect 26321 6261 26361 6264
rect 27233 6268 27382 6275
rect 26718 6252 26758 6253
rect 26429 6235 26758 6252
rect 27233 6248 27292 6268
rect 27312 6248 27351 6268
rect 27371 6248 27382 6268
rect 27233 6240 27382 6248
rect 27449 6271 27606 6278
rect 27449 6251 27569 6271
rect 27589 6251 27606 6271
rect 27449 6241 27606 6251
rect 27449 6240 27484 6241
rect 26313 6192 26356 6203
rect 26313 6174 26325 6192
rect 26343 6174 26356 6192
rect 26313 6148 26356 6174
rect 26429 6148 26456 6235
rect 26718 6226 26758 6235
rect 25479 6123 25918 6141
rect 24752 6118 24793 6119
rect 24486 6065 24523 6066
rect 24179 6056 24317 6065
rect 24179 6036 24288 6056
rect 24308 6036 24317 6056
rect 24179 6029 24317 6036
rect 24375 6056 24523 6065
rect 24375 6036 24384 6056
rect 24404 6036 24494 6056
rect 24514 6036 24523 6056
rect 24179 6027 24275 6029
rect 24375 6026 24523 6036
rect 24582 6056 24619 6066
rect 24582 6036 24590 6056
rect 24610 6036 24619 6056
rect 24431 6025 24467 6026
rect 24279 5966 24316 5967
rect 24582 5966 24619 6036
rect 24654 6065 24685 6116
rect 25479 6105 25879 6123
rect 25897 6105 25918 6123
rect 25479 6099 25918 6105
rect 25485 6095 25918 6099
rect 26313 6127 26456 6148
rect 26500 6200 26534 6216
rect 26718 6206 27111 6226
rect 27131 6206 27134 6226
rect 27449 6219 27480 6240
rect 27667 6219 27703 6329
rect 27722 6328 27759 6329
rect 27818 6328 27855 6329
rect 27778 6269 27868 6275
rect 27778 6249 27787 6269
rect 27807 6267 27868 6269
rect 27807 6249 27832 6267
rect 27778 6247 27832 6249
rect 27852 6247 27868 6267
rect 27778 6241 27868 6247
rect 27292 6218 27329 6219
rect 26718 6201 27134 6206
rect 27291 6209 27329 6218
rect 26718 6200 27059 6201
rect 26500 6130 26537 6200
rect 26652 6140 26683 6141
rect 26313 6125 26450 6127
rect 25864 6093 25916 6095
rect 26313 6083 26356 6125
rect 26500 6110 26509 6130
rect 26529 6110 26537 6130
rect 26500 6100 26537 6110
rect 26596 6130 26683 6140
rect 26596 6110 26605 6130
rect 26625 6110 26683 6130
rect 26596 6101 26683 6110
rect 26596 6100 26633 6101
rect 26311 6073 26356 6083
rect 24704 6065 24741 6066
rect 24654 6056 24741 6065
rect 24654 6036 24712 6056
rect 24732 6036 24741 6056
rect 24654 6026 24741 6036
rect 24800 6056 24837 6066
rect 24800 6036 24808 6056
rect 24828 6036 24837 6056
rect 26311 6055 26320 6073
rect 26338 6055 26356 6073
rect 26311 6049 26356 6055
rect 26652 6050 26683 6101
rect 26718 6130 26755 6200
rect 27021 6199 27058 6200
rect 27291 6189 27300 6209
rect 27320 6189 27329 6209
rect 27291 6181 27329 6189
rect 27395 6213 27480 6219
rect 27510 6218 27547 6219
rect 27395 6193 27403 6213
rect 27423 6193 27480 6213
rect 27395 6185 27480 6193
rect 27509 6209 27547 6218
rect 27509 6189 27518 6209
rect 27538 6189 27547 6209
rect 27395 6184 27431 6185
rect 27509 6181 27547 6189
rect 27613 6213 27757 6219
rect 27613 6193 27621 6213
rect 27641 6194 27673 6213
rect 27694 6194 27729 6213
rect 27641 6193 27729 6194
rect 27749 6193 27757 6213
rect 27613 6185 27757 6193
rect 27613 6184 27649 6185
rect 27721 6184 27757 6185
rect 27823 6218 27860 6219
rect 27823 6217 27861 6218
rect 27823 6209 27887 6217
rect 27823 6189 27832 6209
rect 27852 6195 27887 6209
rect 27907 6195 27910 6215
rect 27852 6190 27910 6195
rect 27852 6189 27887 6190
rect 27292 6152 27329 6181
rect 27293 6150 27329 6152
rect 26870 6140 26906 6141
rect 26718 6110 26727 6130
rect 26747 6110 26755 6130
rect 26718 6100 26755 6110
rect 26814 6130 26962 6140
rect 27062 6137 27158 6139
rect 26814 6110 26823 6130
rect 26843 6110 26933 6130
rect 26953 6110 26962 6130
rect 26814 6101 26962 6110
rect 27020 6130 27158 6137
rect 27020 6110 27029 6130
rect 27049 6110 27158 6130
rect 27293 6128 27484 6150
rect 27510 6149 27547 6181
rect 27823 6177 27887 6189
rect 27927 6151 27954 6329
rect 27786 6149 27954 6151
rect 27510 6123 27954 6149
rect 27020 6101 27158 6110
rect 26814 6100 26851 6101
rect 26311 6046 26348 6049
rect 26544 6047 26585 6048
rect 24654 6025 24685 6026
rect 24278 5965 24619 5966
rect 24800 5965 24837 6036
rect 26436 6040 26585 6047
rect 25867 6028 25904 6033
rect 25858 6024 25905 6028
rect 25858 6006 25877 6024
rect 25895 6006 25905 6024
rect 26436 6020 26495 6040
rect 26515 6020 26554 6040
rect 26574 6020 26585 6040
rect 26436 6012 26585 6020
rect 26652 6043 26809 6050
rect 26652 6023 26772 6043
rect 26792 6023 26809 6043
rect 26652 6013 26809 6023
rect 26652 6012 26687 6013
rect 24203 5960 24619 5965
rect 24203 5940 24206 5960
rect 24226 5940 24619 5960
rect 24650 5941 24837 5965
rect 25462 5963 25502 5968
rect 25858 5963 25905 6006
rect 26652 5991 26683 6012
rect 26870 5991 26906 6101
rect 26925 6100 26962 6101
rect 27021 6100 27058 6101
rect 26981 6041 27071 6047
rect 26981 6021 26990 6041
rect 27010 6039 27071 6041
rect 27010 6021 27035 6039
rect 26981 6019 27035 6021
rect 27055 6019 27071 6039
rect 26981 6013 27071 6019
rect 26495 5990 26532 5991
rect 25462 5924 25905 5963
rect 26308 5982 26345 5984
rect 26308 5974 26350 5982
rect 26308 5956 26318 5974
rect 26336 5956 26350 5974
rect 26308 5947 26350 5956
rect 26494 5981 26532 5990
rect 26494 5961 26503 5981
rect 26523 5961 26532 5981
rect 26494 5953 26532 5961
rect 26598 5985 26683 5991
rect 26713 5990 26750 5991
rect 26598 5965 26606 5985
rect 26626 5965 26683 5985
rect 26598 5957 26683 5965
rect 26712 5981 26750 5990
rect 26712 5961 26721 5981
rect 26741 5961 26750 5981
rect 26598 5956 26634 5957
rect 26712 5953 26750 5961
rect 26816 5989 26960 5991
rect 26816 5985 26868 5989
rect 26816 5965 26824 5985
rect 26844 5969 26868 5985
rect 26888 5985 26960 5989
rect 26888 5969 26932 5985
rect 26844 5965 26932 5969
rect 26952 5965 26960 5985
rect 26816 5957 26960 5965
rect 26816 5956 26852 5957
rect 26924 5956 26960 5957
rect 27026 5990 27063 5991
rect 27026 5989 27064 5990
rect 27026 5981 27090 5989
rect 27026 5961 27035 5981
rect 27055 5967 27090 5981
rect 27110 5967 27113 5987
rect 27055 5962 27113 5967
rect 27055 5961 27090 5962
rect 24556 5909 24596 5917
rect 24556 5887 24564 5909
rect 24588 5887 24596 5909
rect 24262 5663 24430 5664
rect 24556 5663 24596 5887
rect 25059 5891 25227 5892
rect 25462 5891 25502 5924
rect 25858 5891 25905 5924
rect 26309 5922 26350 5947
rect 26495 5922 26532 5953
rect 26713 5922 26750 5953
rect 27026 5949 27090 5961
rect 27130 5923 27157 6101
rect 26309 5895 26358 5922
rect 26494 5896 26543 5922
rect 26712 5921 26793 5922
rect 26989 5921 27157 5923
rect 26712 5896 27157 5921
rect 26713 5895 27157 5896
rect 25059 5890 25503 5891
rect 25059 5865 25504 5890
rect 25059 5863 25227 5865
rect 25423 5864 25504 5865
rect 25673 5864 25722 5890
rect 25858 5864 25907 5891
rect 25059 5685 25086 5863
rect 25126 5825 25190 5837
rect 25466 5833 25503 5864
rect 25684 5833 25721 5864
rect 25866 5839 25907 5864
rect 26311 5862 26358 5895
rect 26714 5862 26754 5895
rect 26989 5894 27157 5895
rect 27620 5899 27660 6123
rect 27786 6122 27954 6123
rect 27620 5877 27628 5899
rect 27652 5877 27660 5899
rect 27620 5869 27660 5877
rect 25126 5824 25161 5825
rect 25103 5819 25161 5824
rect 25103 5799 25106 5819
rect 25126 5805 25161 5819
rect 25181 5805 25190 5825
rect 25126 5797 25190 5805
rect 25152 5796 25190 5797
rect 25153 5795 25190 5796
rect 25256 5829 25292 5830
rect 25364 5829 25400 5830
rect 25256 5821 25400 5829
rect 25256 5801 25264 5821
rect 25284 5817 25372 5821
rect 25284 5801 25328 5817
rect 25256 5797 25328 5801
rect 25348 5801 25372 5817
rect 25392 5801 25400 5821
rect 25348 5797 25400 5801
rect 25256 5795 25400 5797
rect 25466 5825 25504 5833
rect 25582 5829 25618 5830
rect 25466 5805 25475 5825
rect 25495 5805 25504 5825
rect 25466 5796 25504 5805
rect 25533 5821 25618 5829
rect 25533 5801 25590 5821
rect 25610 5801 25618 5821
rect 25466 5795 25503 5796
rect 25533 5795 25618 5801
rect 25684 5825 25722 5833
rect 25684 5805 25693 5825
rect 25713 5805 25722 5825
rect 25684 5796 25722 5805
rect 25866 5830 25908 5839
rect 25866 5812 25880 5830
rect 25898 5812 25908 5830
rect 25866 5804 25908 5812
rect 25871 5802 25908 5804
rect 26311 5823 26754 5862
rect 25684 5795 25721 5796
rect 25145 5767 25235 5773
rect 25145 5747 25161 5767
rect 25181 5765 25235 5767
rect 25181 5747 25206 5765
rect 25145 5745 25206 5747
rect 25226 5745 25235 5765
rect 25145 5739 25235 5745
rect 25158 5685 25195 5686
rect 25254 5685 25291 5686
rect 25310 5685 25346 5795
rect 25533 5774 25564 5795
rect 26311 5780 26358 5823
rect 26714 5818 26754 5823
rect 27379 5821 27566 5845
rect 27597 5826 27990 5846
rect 28010 5826 28013 5846
rect 27597 5821 28013 5826
rect 25529 5773 25564 5774
rect 25407 5763 25564 5773
rect 25407 5743 25424 5763
rect 25444 5743 25564 5763
rect 25407 5736 25564 5743
rect 25631 5766 25780 5774
rect 25631 5746 25642 5766
rect 25662 5746 25701 5766
rect 25721 5746 25780 5766
rect 26311 5762 26321 5780
rect 26339 5762 26358 5780
rect 26311 5758 26358 5762
rect 26312 5753 26349 5758
rect 25631 5739 25780 5746
rect 27379 5750 27416 5821
rect 27597 5820 27938 5821
rect 27531 5760 27562 5761
rect 25631 5738 25672 5739
rect 25868 5737 25905 5740
rect 25365 5685 25402 5686
rect 25058 5676 25196 5685
rect 24262 5637 24706 5663
rect 24262 5635 24430 5637
rect 24262 5457 24289 5635
rect 24329 5597 24393 5609
rect 24669 5605 24706 5637
rect 24732 5636 24923 5658
rect 25058 5656 25167 5676
rect 25187 5656 25196 5676
rect 25058 5649 25196 5656
rect 25254 5676 25402 5685
rect 25254 5656 25263 5676
rect 25283 5656 25373 5676
rect 25393 5656 25402 5676
rect 25058 5647 25154 5649
rect 25254 5646 25402 5656
rect 25461 5676 25498 5686
rect 25461 5656 25469 5676
rect 25489 5656 25498 5676
rect 25310 5645 25346 5646
rect 24887 5634 24923 5636
rect 24887 5605 24924 5634
rect 24329 5596 24364 5597
rect 24306 5591 24364 5596
rect 24306 5571 24309 5591
rect 24329 5577 24364 5591
rect 24384 5577 24393 5597
rect 24329 5569 24393 5577
rect 24355 5568 24393 5569
rect 24356 5567 24393 5568
rect 24459 5601 24495 5602
rect 24567 5601 24603 5602
rect 24459 5593 24603 5601
rect 24459 5573 24467 5593
rect 24487 5592 24575 5593
rect 24487 5573 24522 5592
rect 24543 5573 24575 5592
rect 24595 5573 24603 5593
rect 24459 5567 24603 5573
rect 24669 5597 24707 5605
rect 24785 5601 24821 5602
rect 24669 5577 24678 5597
rect 24698 5577 24707 5597
rect 24669 5568 24707 5577
rect 24736 5593 24821 5601
rect 24736 5573 24793 5593
rect 24813 5573 24821 5593
rect 24669 5567 24706 5568
rect 24736 5567 24821 5573
rect 24887 5597 24925 5605
rect 24887 5577 24896 5597
rect 24916 5577 24925 5597
rect 25158 5586 25195 5587
rect 25461 5586 25498 5656
rect 25533 5685 25564 5736
rect 25860 5731 25905 5737
rect 25860 5713 25878 5731
rect 25896 5713 25905 5731
rect 27379 5730 27388 5750
rect 27408 5730 27416 5750
rect 27379 5720 27416 5730
rect 27475 5750 27562 5760
rect 27475 5730 27484 5750
rect 27504 5730 27562 5750
rect 27475 5721 27562 5730
rect 27475 5720 27512 5721
rect 25860 5703 25905 5713
rect 25583 5685 25620 5686
rect 25533 5676 25620 5685
rect 25533 5656 25591 5676
rect 25611 5656 25620 5676
rect 25533 5646 25620 5656
rect 25679 5676 25716 5686
rect 25679 5656 25687 5676
rect 25707 5656 25716 5676
rect 25860 5661 25903 5703
rect 26300 5691 26352 5693
rect 25766 5659 25903 5661
rect 25533 5645 25564 5646
rect 25679 5586 25716 5656
rect 25157 5585 25498 5586
rect 24887 5568 24925 5577
rect 25082 5580 25498 5585
rect 24887 5567 24924 5568
rect 24348 5539 24438 5545
rect 24348 5519 24364 5539
rect 24384 5537 24438 5539
rect 24384 5519 24409 5537
rect 24348 5517 24409 5519
rect 24429 5517 24438 5537
rect 24348 5511 24438 5517
rect 24361 5457 24398 5458
rect 24457 5457 24494 5458
rect 24513 5457 24549 5567
rect 24736 5546 24767 5567
rect 25082 5560 25085 5580
rect 25105 5560 25498 5580
rect 25682 5570 25716 5586
rect 25760 5638 25903 5659
rect 26298 5687 26731 5691
rect 26298 5681 26737 5687
rect 26298 5663 26319 5681
rect 26337 5663 26737 5681
rect 27531 5670 27562 5721
rect 27597 5750 27634 5820
rect 27900 5819 27937 5820
rect 27749 5760 27785 5761
rect 27597 5730 27606 5750
rect 27626 5730 27634 5750
rect 27597 5720 27634 5730
rect 27693 5750 27841 5760
rect 27941 5757 28037 5759
rect 27693 5730 27702 5750
rect 27722 5730 27812 5750
rect 27832 5730 27841 5750
rect 27693 5721 27841 5730
rect 27899 5750 28037 5757
rect 27899 5730 27908 5750
rect 27928 5730 28037 5750
rect 27899 5721 28037 5730
rect 27693 5720 27730 5721
rect 27423 5667 27464 5668
rect 26298 5645 26737 5663
rect 25458 5551 25498 5560
rect 25760 5551 25787 5638
rect 25860 5612 25903 5638
rect 25860 5594 25873 5612
rect 25891 5594 25903 5612
rect 25860 5583 25903 5594
rect 24732 5545 24767 5546
rect 24610 5535 24767 5545
rect 24610 5515 24627 5535
rect 24647 5515 24767 5535
rect 24610 5508 24767 5515
rect 24834 5538 24983 5546
rect 24834 5518 24845 5538
rect 24865 5518 24904 5538
rect 24924 5518 24983 5538
rect 25458 5534 25787 5551
rect 25458 5533 25498 5534
rect 24834 5511 24983 5518
rect 25855 5522 25895 5525
rect 25855 5516 25898 5522
rect 25480 5513 25898 5516
rect 24834 5510 24875 5511
rect 24568 5457 24605 5458
rect 24261 5448 24399 5457
rect 23959 5273 23999 5445
rect 24261 5428 24370 5448
rect 24390 5428 24399 5448
rect 24261 5421 24399 5428
rect 24457 5448 24605 5457
rect 24457 5428 24466 5448
rect 24486 5428 24576 5448
rect 24596 5428 24605 5448
rect 24261 5419 24357 5421
rect 24457 5418 24605 5428
rect 24664 5448 24701 5458
rect 24664 5428 24672 5448
rect 24692 5428 24701 5448
rect 24513 5417 24549 5418
rect 24361 5358 24398 5359
rect 24664 5358 24701 5428
rect 24736 5457 24767 5508
rect 25480 5495 25871 5513
rect 25889 5495 25898 5513
rect 25480 5493 25898 5495
rect 25480 5485 25507 5493
rect 25748 5490 25898 5493
rect 25060 5479 25228 5480
rect 25479 5479 25507 5485
rect 25060 5463 25507 5479
rect 25855 5485 25898 5490
rect 24786 5457 24823 5458
rect 24736 5448 24823 5457
rect 24736 5428 24794 5448
rect 24814 5428 24823 5448
rect 24736 5418 24823 5428
rect 24882 5448 24919 5458
rect 24882 5428 24890 5448
rect 24910 5428 24919 5448
rect 24736 5417 24767 5418
rect 24360 5357 24701 5358
rect 24882 5357 24919 5428
rect 24285 5352 24701 5357
rect 24285 5332 24288 5352
rect 24308 5332 24701 5352
rect 24732 5333 24919 5357
rect 25060 5453 25504 5463
rect 25060 5451 25228 5453
rect 25060 5273 25087 5451
rect 25127 5413 25191 5425
rect 25467 5421 25504 5453
rect 25530 5452 25721 5474
rect 25685 5450 25721 5452
rect 25685 5421 25722 5450
rect 25855 5429 25895 5485
rect 25127 5412 25162 5413
rect 25104 5407 25162 5412
rect 25104 5387 25107 5407
rect 25127 5393 25162 5407
rect 25182 5393 25191 5413
rect 25127 5385 25191 5393
rect 25153 5384 25191 5385
rect 25154 5383 25191 5384
rect 25257 5417 25293 5418
rect 25365 5417 25401 5418
rect 25257 5409 25401 5417
rect 25257 5389 25265 5409
rect 25285 5389 25320 5409
rect 25340 5389 25373 5409
rect 25393 5389 25401 5409
rect 25257 5383 25401 5389
rect 25467 5413 25505 5421
rect 25583 5417 25619 5418
rect 25467 5393 25476 5413
rect 25496 5393 25505 5413
rect 25467 5384 25505 5393
rect 25534 5409 25619 5417
rect 25534 5389 25591 5409
rect 25611 5389 25619 5409
rect 25467 5383 25504 5384
rect 25534 5383 25619 5389
rect 25685 5413 25723 5421
rect 25685 5393 25694 5413
rect 25714 5393 25723 5413
rect 25855 5411 25867 5429
rect 25885 5411 25895 5429
rect 26300 5456 26352 5645
rect 26698 5620 26737 5645
rect 27315 5660 27464 5667
rect 27315 5640 27374 5660
rect 27394 5640 27433 5660
rect 27453 5640 27464 5660
rect 27315 5632 27464 5640
rect 27531 5663 27688 5670
rect 27531 5643 27651 5663
rect 27671 5643 27688 5663
rect 27531 5633 27688 5643
rect 27531 5632 27566 5633
rect 26482 5595 26669 5619
rect 26698 5600 27093 5620
rect 27113 5600 27116 5620
rect 27531 5611 27562 5632
rect 27749 5611 27785 5721
rect 27804 5720 27841 5721
rect 27900 5720 27937 5721
rect 27860 5661 27950 5667
rect 27860 5641 27869 5661
rect 27889 5659 27950 5661
rect 27889 5641 27914 5659
rect 27860 5639 27914 5641
rect 27934 5639 27950 5659
rect 27860 5633 27950 5639
rect 27374 5610 27411 5611
rect 26698 5595 27116 5600
rect 27373 5601 27411 5610
rect 26482 5524 26519 5595
rect 26698 5594 27041 5595
rect 26698 5591 26737 5594
rect 27003 5593 27040 5594
rect 26634 5534 26665 5535
rect 26482 5504 26491 5524
rect 26511 5504 26519 5524
rect 26482 5494 26519 5504
rect 26578 5524 26665 5534
rect 26578 5504 26587 5524
rect 26607 5504 26665 5524
rect 26578 5495 26665 5504
rect 26578 5494 26615 5495
rect 26300 5438 26316 5456
rect 26334 5438 26352 5456
rect 26634 5444 26665 5495
rect 26700 5524 26737 5591
rect 27373 5581 27382 5601
rect 27402 5581 27411 5601
rect 27373 5573 27411 5581
rect 27477 5605 27562 5611
rect 27592 5610 27629 5611
rect 27477 5585 27485 5605
rect 27505 5585 27562 5605
rect 27477 5577 27562 5585
rect 27591 5601 27629 5610
rect 27591 5581 27600 5601
rect 27620 5581 27629 5601
rect 27477 5576 27513 5577
rect 27591 5573 27629 5581
rect 27695 5605 27839 5611
rect 27695 5585 27703 5605
rect 27723 5600 27811 5605
rect 27723 5585 27759 5600
rect 27695 5583 27759 5585
rect 27778 5585 27811 5600
rect 27831 5585 27839 5605
rect 27778 5583 27839 5585
rect 27695 5577 27839 5583
rect 27695 5576 27731 5577
rect 27803 5576 27839 5577
rect 27905 5610 27942 5611
rect 27905 5609 27943 5610
rect 27905 5601 27969 5609
rect 27905 5581 27914 5601
rect 27934 5587 27969 5601
rect 27989 5587 27992 5607
rect 27934 5582 27992 5587
rect 27934 5581 27969 5582
rect 27374 5544 27411 5573
rect 27375 5542 27411 5544
rect 26852 5534 26888 5535
rect 26700 5504 26709 5524
rect 26729 5504 26737 5524
rect 26700 5494 26737 5504
rect 26796 5524 26944 5534
rect 27044 5531 27140 5533
rect 26796 5504 26805 5524
rect 26825 5504 26915 5524
rect 26935 5504 26944 5524
rect 26796 5495 26944 5504
rect 27002 5524 27140 5531
rect 27002 5504 27011 5524
rect 27031 5504 27140 5524
rect 27375 5520 27566 5542
rect 27592 5541 27629 5573
rect 27905 5569 27969 5581
rect 28009 5543 28036 5721
rect 27868 5541 28036 5543
rect 27592 5527 28036 5541
rect 28060 5564 28088 6510
rect 28060 5534 28105 5564
rect 27592 5515 28039 5527
rect 27635 5513 27668 5515
rect 27002 5495 27140 5504
rect 26796 5494 26833 5495
rect 26526 5441 26567 5442
rect 26300 5420 26352 5438
rect 26418 5434 26567 5441
rect 25855 5401 25895 5411
rect 26418 5414 26477 5434
rect 26497 5414 26536 5434
rect 26556 5414 26567 5434
rect 26418 5406 26567 5414
rect 26634 5437 26791 5444
rect 26634 5417 26754 5437
rect 26774 5417 26791 5437
rect 26634 5407 26791 5417
rect 26634 5406 26669 5407
rect 25685 5384 25723 5393
rect 26634 5385 26665 5406
rect 26852 5385 26888 5495
rect 26907 5494 26944 5495
rect 27003 5494 27040 5495
rect 26963 5435 27053 5441
rect 26963 5415 26972 5435
rect 26992 5433 27053 5435
rect 26992 5415 27017 5433
rect 26963 5413 27017 5415
rect 27037 5413 27053 5433
rect 26963 5407 27053 5413
rect 26477 5384 26514 5385
rect 25685 5383 25722 5384
rect 25146 5355 25236 5361
rect 25146 5335 25162 5355
rect 25182 5353 25236 5355
rect 25182 5335 25207 5353
rect 25146 5333 25207 5335
rect 25227 5333 25236 5353
rect 25146 5327 25236 5333
rect 25159 5273 25196 5274
rect 25255 5273 25292 5274
rect 25311 5273 25347 5383
rect 25534 5362 25565 5383
rect 26476 5375 26514 5384
rect 25530 5361 25565 5362
rect 25408 5351 25565 5361
rect 25408 5331 25425 5351
rect 25445 5331 25565 5351
rect 25408 5324 25565 5331
rect 25632 5354 25781 5362
rect 25632 5334 25643 5354
rect 25663 5334 25702 5354
rect 25722 5334 25781 5354
rect 26304 5357 26344 5367
rect 25632 5327 25781 5334
rect 25847 5330 25899 5348
rect 25632 5326 25673 5327
rect 25366 5273 25403 5274
rect 23960 5258 23999 5273
rect 25059 5264 25197 5273
rect 23960 5257 24126 5258
rect 24252 5257 24292 5259
rect 23960 5231 24402 5257
rect 23960 5229 24126 5231
rect 23624 5117 23661 5125
rect 23624 5098 23632 5117
rect 23653 5098 23661 5117
rect 23624 5092 23661 5098
rect 23960 5051 23985 5229
rect 24025 5191 24089 5203
rect 24365 5199 24402 5231
rect 24428 5230 24619 5252
rect 25059 5244 25168 5264
rect 25188 5244 25197 5264
rect 25059 5237 25197 5244
rect 25255 5264 25403 5273
rect 25255 5244 25264 5264
rect 25284 5244 25374 5264
rect 25394 5244 25403 5264
rect 25059 5235 25155 5237
rect 25255 5234 25403 5244
rect 25462 5264 25499 5274
rect 25462 5244 25470 5264
rect 25490 5244 25499 5264
rect 25311 5233 25347 5234
rect 24583 5228 24619 5230
rect 24583 5199 24620 5228
rect 24025 5190 24060 5191
rect 24002 5185 24060 5190
rect 24002 5165 24005 5185
rect 24025 5171 24060 5185
rect 24080 5171 24089 5191
rect 24025 5163 24089 5171
rect 24051 5162 24089 5163
rect 24052 5161 24089 5162
rect 24155 5195 24191 5196
rect 24263 5195 24299 5196
rect 24155 5190 24299 5195
rect 24155 5187 24217 5190
rect 24155 5167 24163 5187
rect 24183 5167 24217 5187
rect 24155 5164 24217 5167
rect 24243 5187 24299 5190
rect 24243 5167 24271 5187
rect 24291 5167 24299 5187
rect 24243 5164 24299 5167
rect 24155 5161 24299 5164
rect 24365 5191 24403 5199
rect 24481 5195 24517 5196
rect 24365 5171 24374 5191
rect 24394 5171 24403 5191
rect 24365 5162 24403 5171
rect 24432 5187 24517 5195
rect 24432 5167 24489 5187
rect 24509 5167 24517 5187
rect 24365 5161 24402 5162
rect 24432 5161 24517 5167
rect 24583 5191 24621 5199
rect 24583 5171 24592 5191
rect 24612 5171 24621 5191
rect 25462 5177 25499 5244
rect 25534 5273 25565 5324
rect 25847 5312 25865 5330
rect 25883 5312 25899 5330
rect 25584 5273 25621 5274
rect 25534 5264 25621 5273
rect 25534 5244 25592 5264
rect 25612 5244 25621 5264
rect 25534 5234 25621 5244
rect 25680 5264 25717 5274
rect 25680 5244 25688 5264
rect 25708 5244 25717 5264
rect 25534 5233 25565 5234
rect 25159 5174 25196 5175
rect 25462 5174 25501 5177
rect 25158 5173 25501 5174
rect 25680 5173 25717 5244
rect 24583 5162 24621 5171
rect 25083 5168 25501 5173
rect 24583 5161 24620 5162
rect 24044 5133 24134 5139
rect 24044 5113 24060 5133
rect 24080 5131 24134 5133
rect 24080 5113 24105 5131
rect 24044 5111 24105 5113
rect 24125 5111 24134 5131
rect 24044 5105 24134 5111
rect 24057 5051 24094 5052
rect 24153 5051 24190 5052
rect 24209 5051 24245 5161
rect 24432 5140 24463 5161
rect 25083 5148 25086 5168
rect 25106 5148 25501 5168
rect 25530 5149 25717 5173
rect 24428 5139 24463 5140
rect 24306 5129 24463 5139
rect 24306 5109 24323 5129
rect 24343 5109 24463 5129
rect 24306 5102 24463 5109
rect 24530 5132 24679 5140
rect 24530 5112 24541 5132
rect 24561 5112 24600 5132
rect 24620 5112 24679 5132
rect 24530 5105 24679 5112
rect 25462 5123 25501 5148
rect 25847 5123 25899 5312
rect 26304 5339 26314 5357
rect 26332 5339 26344 5357
rect 26476 5355 26485 5375
rect 26505 5355 26514 5375
rect 26476 5347 26514 5355
rect 26580 5379 26665 5385
rect 26695 5384 26732 5385
rect 26580 5359 26588 5379
rect 26608 5359 26665 5379
rect 26580 5351 26665 5359
rect 26694 5375 26732 5384
rect 26694 5355 26703 5375
rect 26723 5355 26732 5375
rect 26580 5350 26616 5351
rect 26694 5347 26732 5355
rect 26798 5379 26942 5385
rect 26798 5359 26806 5379
rect 26826 5359 26859 5379
rect 26879 5359 26914 5379
rect 26934 5359 26942 5379
rect 26798 5351 26942 5359
rect 26798 5350 26834 5351
rect 26906 5350 26942 5351
rect 27008 5384 27045 5385
rect 27008 5383 27046 5384
rect 27008 5375 27072 5383
rect 27008 5355 27017 5375
rect 27037 5361 27072 5375
rect 27092 5361 27095 5381
rect 27037 5356 27095 5361
rect 27037 5355 27072 5356
rect 26304 5283 26344 5339
rect 26477 5318 26514 5347
rect 26478 5316 26514 5318
rect 26478 5294 26669 5316
rect 26695 5315 26732 5347
rect 27008 5343 27072 5355
rect 27112 5317 27139 5495
rect 27997 5470 28039 5515
rect 28060 5516 28071 5534
rect 28093 5516 28105 5534
rect 28060 5510 28105 5516
rect 28061 5509 28105 5510
rect 26971 5315 27139 5317
rect 26695 5305 27139 5315
rect 27280 5411 27467 5435
rect 27498 5416 27891 5436
rect 27911 5416 27914 5436
rect 27498 5411 27914 5416
rect 27280 5340 27317 5411
rect 27498 5410 27839 5411
rect 27432 5350 27463 5351
rect 27280 5320 27289 5340
rect 27309 5320 27317 5340
rect 27280 5310 27317 5320
rect 27376 5340 27463 5350
rect 27376 5320 27385 5340
rect 27405 5320 27463 5340
rect 27376 5311 27463 5320
rect 27376 5310 27413 5311
rect 26301 5278 26344 5283
rect 26692 5289 27139 5305
rect 26692 5283 26720 5289
rect 26971 5288 27139 5289
rect 26301 5275 26451 5278
rect 26692 5275 26719 5283
rect 26301 5273 26719 5275
rect 26301 5255 26310 5273
rect 26328 5255 26719 5273
rect 27432 5260 27463 5311
rect 27498 5340 27535 5410
rect 27801 5409 27838 5410
rect 27650 5350 27686 5351
rect 27498 5320 27507 5340
rect 27527 5320 27535 5340
rect 27498 5310 27535 5320
rect 27594 5340 27742 5350
rect 27842 5347 27938 5349
rect 27594 5320 27603 5340
rect 27623 5320 27713 5340
rect 27733 5320 27742 5340
rect 27594 5311 27742 5320
rect 27800 5340 27938 5347
rect 27800 5320 27809 5340
rect 27829 5320 27938 5340
rect 27800 5311 27938 5320
rect 27594 5310 27631 5311
rect 27324 5257 27365 5258
rect 26301 5252 26719 5255
rect 26301 5246 26344 5252
rect 26304 5243 26344 5246
rect 27219 5250 27365 5257
rect 26701 5234 26741 5235
rect 26412 5217 26741 5234
rect 27219 5230 27275 5250
rect 27295 5230 27334 5250
rect 27354 5230 27365 5250
rect 27219 5222 27365 5230
rect 27432 5253 27589 5260
rect 27432 5233 27552 5253
rect 27572 5233 27589 5253
rect 27432 5223 27589 5233
rect 27432 5222 27467 5223
rect 26296 5174 26339 5185
rect 26296 5156 26308 5174
rect 26326 5156 26339 5174
rect 26296 5130 26339 5156
rect 26412 5130 26439 5217
rect 26701 5208 26741 5217
rect 25462 5105 25901 5123
rect 24530 5104 24571 5105
rect 24264 5051 24301 5052
rect 23960 5042 24095 5051
rect 23960 5022 24066 5042
rect 24086 5022 24095 5042
rect 23960 5015 24095 5022
rect 24153 5042 24301 5051
rect 24153 5022 24162 5042
rect 24182 5022 24272 5042
rect 24292 5022 24301 5042
rect 23960 5013 24053 5015
rect 24153 5012 24301 5022
rect 24360 5042 24397 5052
rect 24360 5022 24368 5042
rect 24388 5022 24397 5042
rect 24209 5011 24245 5012
rect 24057 4952 24094 4953
rect 24360 4952 24397 5022
rect 24432 5051 24463 5102
rect 25462 5087 25862 5105
rect 25880 5087 25901 5105
rect 25462 5081 25901 5087
rect 25468 5077 25901 5081
rect 26296 5109 26439 5130
rect 26483 5182 26517 5198
rect 26701 5188 27094 5208
rect 27114 5188 27117 5208
rect 27432 5201 27463 5222
rect 27650 5201 27686 5311
rect 27705 5310 27742 5311
rect 27801 5310 27838 5311
rect 27761 5251 27851 5257
rect 27761 5231 27770 5251
rect 27790 5249 27851 5251
rect 27790 5231 27815 5249
rect 27761 5229 27815 5231
rect 27835 5229 27851 5249
rect 27761 5223 27851 5229
rect 27275 5200 27312 5201
rect 26701 5183 27117 5188
rect 27274 5191 27312 5200
rect 26701 5182 27042 5183
rect 26483 5112 26520 5182
rect 26635 5122 26666 5123
rect 26296 5107 26433 5109
rect 25847 5075 25899 5077
rect 26296 5065 26339 5107
rect 26483 5092 26492 5112
rect 26512 5092 26520 5112
rect 26483 5082 26520 5092
rect 26579 5112 26666 5122
rect 26579 5092 26588 5112
rect 26608 5092 26666 5112
rect 26579 5083 26666 5092
rect 26579 5082 26616 5083
rect 26294 5055 26339 5065
rect 24482 5051 24519 5052
rect 24432 5042 24519 5051
rect 24432 5022 24490 5042
rect 24510 5022 24519 5042
rect 24432 5012 24519 5022
rect 24578 5042 24615 5052
rect 24578 5022 24586 5042
rect 24606 5022 24615 5042
rect 26294 5037 26303 5055
rect 26321 5037 26339 5055
rect 26294 5031 26339 5037
rect 26635 5032 26666 5083
rect 26701 5112 26738 5182
rect 27004 5181 27041 5182
rect 27274 5171 27283 5191
rect 27303 5171 27312 5191
rect 27274 5163 27312 5171
rect 27378 5195 27463 5201
rect 27493 5200 27530 5201
rect 27378 5175 27386 5195
rect 27406 5175 27463 5195
rect 27378 5167 27463 5175
rect 27492 5191 27530 5200
rect 27492 5171 27501 5191
rect 27521 5171 27530 5191
rect 27378 5166 27414 5167
rect 27492 5163 27530 5171
rect 27596 5195 27740 5201
rect 27596 5175 27604 5195
rect 27624 5192 27712 5195
rect 27624 5175 27659 5192
rect 27596 5174 27659 5175
rect 27678 5175 27712 5192
rect 27732 5175 27740 5195
rect 27678 5174 27740 5175
rect 27596 5167 27740 5174
rect 27596 5166 27632 5167
rect 27704 5166 27740 5167
rect 27806 5200 27843 5201
rect 27806 5199 27844 5200
rect 27866 5199 27893 5203
rect 27806 5197 27893 5199
rect 27806 5191 27870 5197
rect 27806 5171 27815 5191
rect 27835 5177 27870 5191
rect 27890 5177 27893 5197
rect 27835 5172 27893 5177
rect 27835 5171 27870 5172
rect 27275 5134 27312 5163
rect 27276 5132 27312 5134
rect 26853 5122 26889 5123
rect 26701 5092 26710 5112
rect 26730 5092 26738 5112
rect 26701 5082 26738 5092
rect 26797 5112 26945 5122
rect 27045 5119 27141 5121
rect 26797 5092 26806 5112
rect 26826 5092 26916 5112
rect 26936 5092 26945 5112
rect 26797 5083 26945 5092
rect 27003 5112 27141 5119
rect 27003 5092 27012 5112
rect 27032 5092 27141 5112
rect 27276 5110 27467 5132
rect 27493 5131 27530 5163
rect 27806 5159 27870 5171
rect 27910 5133 27937 5311
rect 27769 5131 27937 5133
rect 27493 5105 27937 5131
rect 27003 5083 27141 5092
rect 26797 5082 26834 5083
rect 26294 5028 26331 5031
rect 26527 5029 26568 5030
rect 24432 5011 24463 5012
rect 24056 4951 24397 4952
rect 24578 4951 24615 5022
rect 26419 5022 26568 5029
rect 25850 5010 25887 5015
rect 23981 4946 24397 4951
rect 23981 4926 23984 4946
rect 24004 4926 24397 4946
rect 24428 4927 24615 4951
rect 25841 5006 25888 5010
rect 25841 4988 25860 5006
rect 25878 4988 25888 5006
rect 26419 5002 26478 5022
rect 26498 5002 26537 5022
rect 26557 5002 26568 5022
rect 26419 4994 26568 5002
rect 26635 5025 26792 5032
rect 26635 5005 26755 5025
rect 26775 5005 26792 5025
rect 26635 4995 26792 5005
rect 26635 4994 26670 4995
rect 25449 4929 25487 4930
rect 25841 4929 25888 4988
rect 26635 4973 26666 4994
rect 26853 4973 26889 5083
rect 26908 5082 26945 5083
rect 27004 5082 27041 5083
rect 26964 5023 27054 5029
rect 26964 5003 26973 5023
rect 26993 5021 27054 5023
rect 26993 5003 27018 5021
rect 26964 5001 27018 5003
rect 27038 5001 27054 5021
rect 26964 4995 27054 5001
rect 26478 4972 26515 4973
rect 26291 4964 26328 4966
rect 26291 4956 26333 4964
rect 26291 4938 26301 4956
rect 26319 4938 26333 4956
rect 26291 4929 26333 4938
rect 26477 4963 26515 4972
rect 26477 4943 26486 4963
rect 26506 4943 26515 4963
rect 26477 4935 26515 4943
rect 26581 4967 26666 4973
rect 26696 4972 26733 4973
rect 26581 4947 26589 4967
rect 26609 4947 26666 4967
rect 26581 4939 26666 4947
rect 26695 4963 26733 4972
rect 26695 4943 26704 4963
rect 26724 4943 26733 4963
rect 26581 4938 26617 4939
rect 26695 4935 26733 4943
rect 26799 4971 26943 4973
rect 26799 4967 26851 4971
rect 26799 4947 26807 4967
rect 26827 4951 26851 4967
rect 26871 4967 26943 4971
rect 26871 4951 26915 4967
rect 26827 4947 26915 4951
rect 26935 4947 26943 4967
rect 26799 4939 26943 4947
rect 26799 4938 26835 4939
rect 26907 4938 26943 4939
rect 27009 4972 27046 4973
rect 27009 4971 27047 4972
rect 27009 4963 27073 4971
rect 27009 4943 27018 4963
rect 27038 4949 27073 4963
rect 27093 4949 27096 4969
rect 27038 4944 27096 4949
rect 27038 4943 27073 4944
rect 24201 4925 24266 4926
rect 22316 4847 22354 4848
rect 21915 4809 22354 4847
rect 23226 4847 23234 4869
rect 23258 4847 23266 4869
rect 23226 4839 23266 4847
rect 24537 4891 24577 4899
rect 24537 4869 24545 4891
rect 24569 4869 24577 4891
rect 25449 4891 25888 4929
rect 25449 4890 25487 4891
rect 23537 4812 23602 4813
rect 20743 4793 20778 4794
rect 20720 4788 20778 4793
rect 20720 4768 20723 4788
rect 20743 4774 20778 4788
rect 20798 4774 20807 4794
rect 20743 4766 20807 4774
rect 20769 4765 20807 4766
rect 20770 4764 20807 4765
rect 20873 4798 20909 4799
rect 20981 4798 21017 4799
rect 20873 4790 21017 4798
rect 20873 4770 20881 4790
rect 20901 4786 20989 4790
rect 20901 4770 20945 4786
rect 20873 4766 20945 4770
rect 20965 4770 20989 4786
rect 21009 4770 21017 4790
rect 20965 4766 21017 4770
rect 20873 4764 21017 4766
rect 21083 4794 21121 4802
rect 21199 4798 21235 4799
rect 21083 4774 21092 4794
rect 21112 4774 21121 4794
rect 21083 4765 21121 4774
rect 21150 4790 21235 4798
rect 21150 4770 21207 4790
rect 21227 4770 21235 4790
rect 21083 4764 21120 4765
rect 21150 4764 21235 4770
rect 21301 4794 21339 4802
rect 21301 4774 21310 4794
rect 21330 4774 21339 4794
rect 21301 4765 21339 4774
rect 21483 4799 21525 4808
rect 21483 4781 21497 4799
rect 21515 4781 21525 4799
rect 21483 4773 21525 4781
rect 21488 4771 21525 4773
rect 21301 4764 21338 4765
rect 20762 4736 20852 4742
rect 20762 4716 20778 4736
rect 20798 4734 20852 4736
rect 20798 4716 20823 4734
rect 20762 4714 20823 4716
rect 20843 4714 20852 4734
rect 20762 4708 20852 4714
rect 20775 4654 20812 4655
rect 20871 4654 20908 4655
rect 20927 4654 20963 4764
rect 21150 4743 21181 4764
rect 21915 4750 21962 4809
rect 22316 4808 22354 4809
rect 21146 4742 21181 4743
rect 21024 4732 21181 4742
rect 21024 4712 21041 4732
rect 21061 4712 21181 4732
rect 21024 4705 21181 4712
rect 21248 4735 21397 4743
rect 21248 4715 21259 4735
rect 21279 4715 21318 4735
rect 21338 4715 21397 4735
rect 21915 4732 21925 4750
rect 21943 4732 21962 4750
rect 21915 4728 21962 4732
rect 23188 4787 23375 4811
rect 23406 4792 23799 4812
rect 23819 4792 23822 4812
rect 23406 4787 23822 4792
rect 21916 4723 21953 4728
rect 21248 4708 21397 4715
rect 23188 4716 23225 4787
rect 23406 4786 23747 4787
rect 23340 4726 23371 4727
rect 21248 4707 21289 4708
rect 21485 4706 21522 4709
rect 20982 4654 21019 4655
rect 20675 4645 20813 4654
rect 19879 4606 20323 4632
rect 19879 4604 20047 4606
rect 19879 4426 19906 4604
rect 19946 4566 20010 4578
rect 20286 4574 20323 4606
rect 20349 4605 20540 4627
rect 20675 4625 20784 4645
rect 20804 4625 20813 4645
rect 20675 4618 20813 4625
rect 20871 4645 21019 4654
rect 20871 4625 20880 4645
rect 20900 4625 20990 4645
rect 21010 4625 21019 4645
rect 20675 4616 20771 4618
rect 20871 4615 21019 4625
rect 21078 4645 21115 4655
rect 21078 4625 21086 4645
rect 21106 4625 21115 4645
rect 20927 4614 20963 4615
rect 20504 4603 20540 4605
rect 20504 4574 20541 4603
rect 19946 4565 19981 4566
rect 19923 4560 19981 4565
rect 19923 4540 19926 4560
rect 19946 4546 19981 4560
rect 20001 4546 20010 4566
rect 19946 4540 20010 4546
rect 19923 4538 20010 4540
rect 19923 4534 19950 4538
rect 19972 4537 20010 4538
rect 19973 4536 20010 4537
rect 20076 4570 20112 4571
rect 20184 4570 20220 4571
rect 20076 4563 20220 4570
rect 20076 4562 20138 4563
rect 20076 4542 20084 4562
rect 20104 4545 20138 4562
rect 20157 4562 20220 4563
rect 20157 4545 20192 4562
rect 20104 4542 20192 4545
rect 20212 4542 20220 4562
rect 20076 4536 20220 4542
rect 20286 4566 20324 4574
rect 20402 4570 20438 4571
rect 20286 4546 20295 4566
rect 20315 4546 20324 4566
rect 20286 4537 20324 4546
rect 20353 4562 20438 4570
rect 20353 4542 20410 4562
rect 20430 4542 20438 4562
rect 20286 4536 20323 4537
rect 20353 4536 20438 4542
rect 20504 4566 20542 4574
rect 20504 4546 20513 4566
rect 20533 4546 20542 4566
rect 20775 4555 20812 4556
rect 21078 4555 21115 4625
rect 21150 4654 21181 4705
rect 21477 4700 21522 4706
rect 21477 4682 21495 4700
rect 21513 4682 21522 4700
rect 23188 4696 23197 4716
rect 23217 4696 23225 4716
rect 23188 4686 23225 4696
rect 23284 4716 23371 4726
rect 23284 4696 23293 4716
rect 23313 4696 23371 4716
rect 23284 4687 23371 4696
rect 23284 4686 23321 4687
rect 21477 4672 21522 4682
rect 21200 4654 21237 4655
rect 21150 4645 21237 4654
rect 21150 4625 21208 4645
rect 21228 4625 21237 4645
rect 21150 4615 21237 4625
rect 21296 4645 21333 4655
rect 21296 4625 21304 4645
rect 21324 4625 21333 4645
rect 21477 4630 21520 4672
rect 21904 4661 21956 4663
rect 21383 4628 21520 4630
rect 21150 4614 21181 4615
rect 21296 4555 21333 4625
rect 20774 4554 21115 4555
rect 20504 4537 20542 4546
rect 20699 4549 21115 4554
rect 20504 4536 20541 4537
rect 19965 4508 20055 4514
rect 19965 4488 19981 4508
rect 20001 4506 20055 4508
rect 20001 4488 20026 4506
rect 19965 4486 20026 4488
rect 20046 4486 20055 4506
rect 19965 4480 20055 4486
rect 19978 4426 20015 4427
rect 20074 4426 20111 4427
rect 20130 4426 20166 4536
rect 20353 4515 20384 4536
rect 20699 4529 20702 4549
rect 20722 4529 21115 4549
rect 21299 4539 21333 4555
rect 21377 4607 21520 4628
rect 21902 4657 22335 4661
rect 21902 4651 22341 4657
rect 21902 4633 21923 4651
rect 21941 4633 22341 4651
rect 23340 4636 23371 4687
rect 23406 4716 23443 4786
rect 23709 4785 23746 4786
rect 23558 4726 23594 4727
rect 23406 4696 23415 4716
rect 23435 4696 23443 4716
rect 23406 4686 23443 4696
rect 23502 4716 23650 4726
rect 23750 4723 23846 4725
rect 23502 4696 23511 4716
rect 23531 4696 23621 4716
rect 23641 4696 23650 4716
rect 23502 4687 23650 4696
rect 23708 4716 23846 4723
rect 23708 4696 23717 4716
rect 23737 4696 23846 4716
rect 23708 4687 23846 4696
rect 23502 4686 23539 4687
rect 23232 4633 23273 4634
rect 21902 4615 22341 4633
rect 21075 4520 21115 4529
rect 21377 4520 21404 4607
rect 21477 4581 21520 4607
rect 21477 4563 21490 4581
rect 21508 4563 21520 4581
rect 21477 4552 21520 4563
rect 20349 4514 20384 4515
rect 20227 4504 20384 4514
rect 20227 4484 20244 4504
rect 20264 4484 20384 4504
rect 20227 4477 20384 4484
rect 20451 4507 20597 4515
rect 20451 4487 20462 4507
rect 20482 4487 20521 4507
rect 20541 4487 20597 4507
rect 21075 4503 21404 4520
rect 21075 4502 21115 4503
rect 20451 4480 20597 4487
rect 21472 4491 21512 4494
rect 21472 4485 21515 4491
rect 21097 4482 21515 4485
rect 20451 4479 20492 4480
rect 20185 4426 20222 4427
rect 19878 4417 20016 4426
rect 19878 4397 19987 4417
rect 20007 4397 20016 4417
rect 19878 4390 20016 4397
rect 20074 4417 20222 4426
rect 20074 4397 20083 4417
rect 20103 4397 20193 4417
rect 20213 4397 20222 4417
rect 19878 4388 19974 4390
rect 20074 4387 20222 4397
rect 20281 4417 20318 4427
rect 20281 4397 20289 4417
rect 20309 4397 20318 4417
rect 20130 4386 20166 4387
rect 19978 4327 20015 4328
rect 20281 4327 20318 4397
rect 20353 4426 20384 4477
rect 21097 4464 21488 4482
rect 21506 4464 21515 4482
rect 21097 4462 21515 4464
rect 21097 4454 21124 4462
rect 21365 4459 21515 4462
rect 20677 4448 20845 4449
rect 21096 4448 21124 4454
rect 20677 4432 21124 4448
rect 21472 4454 21515 4459
rect 20403 4426 20440 4427
rect 20353 4417 20440 4426
rect 20353 4397 20411 4417
rect 20431 4397 20440 4417
rect 20353 4387 20440 4397
rect 20499 4417 20536 4427
rect 20499 4397 20507 4417
rect 20527 4397 20536 4417
rect 20353 4386 20384 4387
rect 19977 4326 20318 4327
rect 20499 4326 20536 4397
rect 19902 4321 20318 4326
rect 19902 4301 19905 4321
rect 19925 4301 20318 4321
rect 20349 4302 20536 4326
rect 20677 4422 21121 4432
rect 20677 4420 20845 4422
rect 19711 4227 19755 4228
rect 19711 4221 19756 4227
rect 19711 4203 19723 4221
rect 19745 4203 19756 4221
rect 19777 4222 19819 4267
rect 20677 4242 20704 4420
rect 20744 4382 20808 4394
rect 21084 4390 21121 4422
rect 21147 4421 21338 4443
rect 21302 4419 21338 4421
rect 21302 4390 21339 4419
rect 21472 4398 21512 4454
rect 20744 4381 20779 4382
rect 20721 4376 20779 4381
rect 20721 4356 20724 4376
rect 20744 4362 20779 4376
rect 20799 4362 20808 4382
rect 20744 4354 20808 4362
rect 20770 4353 20808 4354
rect 20771 4352 20808 4353
rect 20874 4386 20910 4387
rect 20982 4386 21018 4387
rect 20874 4378 21018 4386
rect 20874 4358 20882 4378
rect 20902 4358 20937 4378
rect 20957 4358 20990 4378
rect 21010 4358 21018 4378
rect 20874 4352 21018 4358
rect 21084 4382 21122 4390
rect 21200 4386 21236 4387
rect 21084 4362 21093 4382
rect 21113 4362 21122 4382
rect 21084 4353 21122 4362
rect 21151 4378 21236 4386
rect 21151 4358 21208 4378
rect 21228 4358 21236 4378
rect 21084 4352 21121 4353
rect 21151 4352 21236 4358
rect 21302 4382 21340 4390
rect 21302 4362 21311 4382
rect 21331 4362 21340 4382
rect 21472 4380 21484 4398
rect 21502 4380 21512 4398
rect 21904 4426 21956 4615
rect 22302 4590 22341 4615
rect 23124 4626 23273 4633
rect 23124 4606 23183 4626
rect 23203 4606 23242 4626
rect 23262 4606 23273 4626
rect 23124 4598 23273 4606
rect 23340 4629 23497 4636
rect 23340 4609 23460 4629
rect 23480 4609 23497 4629
rect 23340 4599 23497 4609
rect 23340 4598 23375 4599
rect 22086 4565 22273 4589
rect 22302 4570 22697 4590
rect 22717 4570 22720 4590
rect 23340 4577 23371 4598
rect 23558 4577 23594 4687
rect 23613 4686 23650 4687
rect 23709 4686 23746 4687
rect 23669 4627 23759 4633
rect 23669 4607 23678 4627
rect 23698 4625 23759 4627
rect 23698 4607 23723 4625
rect 23669 4605 23723 4607
rect 23743 4605 23759 4625
rect 23669 4599 23759 4605
rect 23183 4576 23220 4577
rect 22302 4565 22720 4570
rect 23182 4567 23220 4576
rect 22086 4494 22123 4565
rect 22302 4564 22645 4565
rect 22302 4561 22341 4564
rect 22607 4563 22644 4564
rect 22238 4504 22269 4505
rect 22086 4474 22095 4494
rect 22115 4474 22123 4494
rect 22086 4464 22123 4474
rect 22182 4494 22269 4504
rect 22182 4474 22191 4494
rect 22211 4474 22269 4494
rect 22182 4465 22269 4474
rect 22182 4464 22219 4465
rect 21904 4408 21920 4426
rect 21938 4408 21956 4426
rect 22238 4414 22269 4465
rect 22304 4494 22341 4561
rect 23182 4547 23191 4567
rect 23211 4547 23220 4567
rect 23182 4539 23220 4547
rect 23286 4571 23371 4577
rect 23401 4576 23438 4577
rect 23286 4551 23294 4571
rect 23314 4551 23371 4571
rect 23286 4543 23371 4551
rect 23400 4567 23438 4576
rect 23400 4547 23409 4567
rect 23429 4547 23438 4567
rect 23286 4542 23322 4543
rect 23400 4539 23438 4547
rect 23504 4571 23648 4577
rect 23504 4551 23512 4571
rect 23532 4565 23620 4571
rect 23532 4551 23561 4565
rect 23504 4543 23561 4551
rect 23504 4542 23540 4543
rect 23584 4551 23620 4565
rect 23640 4551 23648 4571
rect 23584 4543 23648 4551
rect 23612 4542 23648 4543
rect 23714 4576 23751 4577
rect 23714 4575 23752 4576
rect 23714 4567 23778 4575
rect 23714 4547 23723 4567
rect 23743 4553 23778 4567
rect 23798 4553 23801 4573
rect 23743 4548 23801 4553
rect 23743 4547 23778 4548
rect 23183 4510 23220 4539
rect 23184 4508 23220 4510
rect 22456 4504 22492 4505
rect 22304 4474 22313 4494
rect 22333 4474 22341 4494
rect 22304 4464 22341 4474
rect 22400 4494 22548 4504
rect 22648 4501 22744 4503
rect 22400 4474 22409 4494
rect 22429 4474 22519 4494
rect 22539 4474 22548 4494
rect 22400 4465 22548 4474
rect 22606 4494 22744 4501
rect 22606 4474 22615 4494
rect 22635 4474 22744 4494
rect 23184 4486 23375 4508
rect 23401 4507 23438 4539
rect 23714 4535 23778 4547
rect 23818 4509 23845 4687
rect 24142 4640 24179 4646
rect 24142 4621 24150 4640
rect 24171 4621 24179 4640
rect 24142 4613 24179 4621
rect 23677 4507 23845 4509
rect 23401 4481 23845 4507
rect 23511 4479 23551 4481
rect 23677 4480 23845 4481
rect 22606 4465 22744 4474
rect 23804 4475 23845 4480
rect 22400 4464 22437 4465
rect 22130 4411 22171 4412
rect 21904 4390 21956 4408
rect 22022 4404 22171 4411
rect 21472 4370 21512 4380
rect 22022 4384 22081 4404
rect 22101 4384 22140 4404
rect 22160 4384 22171 4404
rect 22022 4376 22171 4384
rect 22238 4407 22395 4414
rect 22238 4387 22358 4407
rect 22378 4387 22395 4407
rect 22238 4377 22395 4387
rect 22238 4376 22273 4377
rect 21302 4353 21340 4362
rect 22238 4355 22269 4376
rect 22456 4355 22492 4465
rect 22511 4464 22548 4465
rect 22607 4464 22644 4465
rect 22567 4405 22657 4411
rect 22567 4385 22576 4405
rect 22596 4403 22657 4405
rect 22596 4385 22621 4403
rect 22567 4383 22621 4385
rect 22641 4383 22657 4403
rect 22567 4377 22657 4383
rect 22081 4354 22118 4355
rect 21302 4352 21339 4353
rect 20763 4324 20853 4330
rect 20763 4304 20779 4324
rect 20799 4322 20853 4324
rect 20799 4304 20824 4322
rect 20763 4302 20824 4304
rect 20844 4302 20853 4322
rect 20763 4296 20853 4302
rect 20776 4242 20813 4243
rect 20872 4242 20909 4243
rect 20928 4242 20964 4352
rect 21151 4331 21182 4352
rect 22080 4345 22118 4354
rect 21147 4330 21182 4331
rect 21025 4320 21182 4330
rect 21025 4300 21042 4320
rect 21062 4300 21182 4320
rect 21025 4293 21182 4300
rect 21249 4323 21398 4331
rect 21249 4303 21260 4323
rect 21280 4303 21319 4323
rect 21339 4303 21398 4323
rect 21908 4327 21948 4337
rect 21249 4296 21398 4303
rect 21464 4299 21516 4317
rect 21249 4295 21290 4296
rect 20983 4242 21020 4243
rect 20676 4233 20814 4242
rect 20148 4222 20181 4224
rect 19777 4210 20224 4222
rect 19711 4173 19756 4203
rect 19728 3227 19756 4173
rect 19780 4196 20224 4210
rect 19780 4194 19948 4196
rect 19780 4016 19807 4194
rect 19847 4156 19911 4168
rect 20187 4164 20224 4196
rect 20250 4195 20441 4217
rect 20676 4213 20785 4233
rect 20805 4213 20814 4233
rect 20676 4206 20814 4213
rect 20872 4233 21020 4242
rect 20872 4213 20881 4233
rect 20901 4213 20991 4233
rect 21011 4213 21020 4233
rect 20676 4204 20772 4206
rect 20872 4203 21020 4213
rect 21079 4233 21116 4243
rect 21079 4213 21087 4233
rect 21107 4213 21116 4233
rect 20928 4202 20964 4203
rect 20405 4193 20441 4195
rect 20405 4164 20442 4193
rect 19847 4155 19882 4156
rect 19824 4150 19882 4155
rect 19824 4130 19827 4150
rect 19847 4136 19882 4150
rect 19902 4136 19911 4156
rect 19847 4128 19911 4136
rect 19873 4127 19911 4128
rect 19874 4126 19911 4127
rect 19977 4160 20013 4161
rect 20085 4160 20121 4161
rect 19977 4154 20121 4160
rect 19977 4152 20038 4154
rect 19977 4132 19985 4152
rect 20005 4137 20038 4152
rect 20057 4152 20121 4154
rect 20057 4137 20093 4152
rect 20005 4132 20093 4137
rect 20113 4132 20121 4152
rect 19977 4126 20121 4132
rect 20187 4156 20225 4164
rect 20303 4160 20339 4161
rect 20187 4136 20196 4156
rect 20216 4136 20225 4156
rect 20187 4127 20225 4136
rect 20254 4152 20339 4160
rect 20254 4132 20311 4152
rect 20331 4132 20339 4152
rect 20187 4126 20224 4127
rect 20254 4126 20339 4132
rect 20405 4156 20443 4164
rect 20405 4136 20414 4156
rect 20434 4136 20443 4156
rect 21079 4146 21116 4213
rect 21151 4242 21182 4293
rect 21464 4281 21482 4299
rect 21500 4281 21516 4299
rect 21201 4242 21238 4243
rect 21151 4233 21238 4242
rect 21151 4213 21209 4233
rect 21229 4213 21238 4233
rect 21151 4203 21238 4213
rect 21297 4233 21334 4243
rect 21297 4213 21305 4233
rect 21325 4213 21334 4233
rect 21151 4202 21182 4203
rect 20776 4143 20813 4144
rect 21079 4143 21118 4146
rect 20775 4142 21118 4143
rect 21297 4142 21334 4213
rect 20405 4127 20443 4136
rect 20700 4137 21118 4142
rect 20405 4126 20442 4127
rect 19866 4098 19956 4104
rect 19866 4078 19882 4098
rect 19902 4096 19956 4098
rect 19902 4078 19927 4096
rect 19866 4076 19927 4078
rect 19947 4076 19956 4096
rect 19866 4070 19956 4076
rect 19879 4016 19916 4017
rect 19975 4016 20012 4017
rect 20031 4016 20067 4126
rect 20254 4105 20285 4126
rect 20700 4117 20703 4137
rect 20723 4117 21118 4137
rect 21147 4118 21334 4142
rect 20250 4104 20285 4105
rect 20128 4094 20285 4104
rect 20128 4074 20145 4094
rect 20165 4074 20285 4094
rect 20128 4067 20285 4074
rect 20352 4097 20501 4105
rect 20352 4077 20363 4097
rect 20383 4077 20422 4097
rect 20442 4077 20501 4097
rect 20352 4070 20501 4077
rect 21079 4092 21118 4117
rect 21464 4092 21516 4281
rect 21908 4309 21918 4327
rect 21936 4309 21948 4327
rect 22080 4325 22089 4345
rect 22109 4325 22118 4345
rect 22080 4317 22118 4325
rect 22184 4349 22269 4355
rect 22299 4354 22336 4355
rect 22184 4329 22192 4349
rect 22212 4329 22269 4349
rect 22184 4321 22269 4329
rect 22298 4345 22336 4354
rect 22298 4325 22307 4345
rect 22327 4325 22336 4345
rect 22184 4320 22220 4321
rect 22298 4317 22336 4325
rect 22402 4349 22546 4355
rect 22402 4329 22410 4349
rect 22430 4329 22463 4349
rect 22483 4329 22518 4349
rect 22538 4329 22546 4349
rect 22402 4321 22546 4329
rect 22402 4320 22438 4321
rect 22510 4320 22546 4321
rect 22612 4354 22649 4355
rect 22612 4353 22650 4354
rect 22612 4345 22676 4353
rect 22612 4325 22621 4345
rect 22641 4331 22676 4345
rect 22696 4331 22699 4351
rect 22641 4326 22699 4331
rect 22641 4325 22676 4326
rect 21908 4253 21948 4309
rect 22081 4288 22118 4317
rect 22082 4286 22118 4288
rect 22082 4264 22273 4286
rect 22299 4285 22336 4317
rect 22612 4313 22676 4325
rect 22716 4287 22743 4465
rect 22575 4285 22743 4287
rect 22299 4275 22743 4285
rect 22884 4381 23071 4405
rect 23102 4386 23495 4406
rect 23515 4386 23518 4406
rect 23102 4381 23518 4386
rect 22884 4310 22921 4381
rect 23102 4380 23443 4381
rect 23036 4320 23067 4321
rect 22884 4290 22893 4310
rect 22913 4290 22921 4310
rect 22884 4280 22921 4290
rect 22980 4310 23067 4320
rect 22980 4290 22989 4310
rect 23009 4290 23067 4310
rect 22980 4281 23067 4290
rect 22980 4280 23017 4281
rect 21905 4248 21948 4253
rect 22296 4259 22743 4275
rect 22296 4253 22324 4259
rect 22575 4258 22743 4259
rect 21905 4245 22055 4248
rect 22296 4245 22323 4253
rect 21905 4243 22323 4245
rect 21905 4225 21914 4243
rect 21932 4225 22323 4243
rect 23036 4230 23067 4281
rect 23102 4310 23139 4380
rect 23405 4379 23442 4380
rect 23254 4320 23290 4321
rect 23102 4290 23111 4310
rect 23131 4290 23139 4310
rect 23102 4280 23139 4290
rect 23198 4310 23346 4320
rect 23446 4317 23542 4319
rect 23198 4290 23207 4310
rect 23227 4290 23317 4310
rect 23337 4290 23346 4310
rect 23198 4281 23346 4290
rect 23404 4310 23542 4317
rect 23404 4290 23413 4310
rect 23433 4290 23542 4310
rect 23804 4293 23844 4475
rect 23404 4281 23542 4290
rect 23198 4280 23235 4281
rect 22928 4227 22969 4228
rect 21905 4222 22323 4225
rect 21905 4216 21948 4222
rect 21908 4213 21948 4216
rect 22820 4220 22969 4227
rect 22305 4204 22345 4205
rect 22016 4187 22345 4204
rect 22820 4200 22879 4220
rect 22899 4200 22938 4220
rect 22958 4200 22969 4220
rect 22820 4192 22969 4200
rect 23036 4223 23193 4230
rect 23036 4203 23156 4223
rect 23176 4203 23193 4223
rect 23036 4193 23193 4203
rect 23036 4192 23071 4193
rect 21900 4144 21943 4155
rect 21900 4126 21912 4144
rect 21930 4126 21943 4144
rect 21900 4100 21943 4126
rect 22016 4100 22043 4187
rect 22305 4178 22345 4187
rect 21079 4074 21518 4092
rect 20352 4069 20393 4070
rect 20086 4016 20123 4017
rect 19779 4007 19917 4016
rect 19779 3987 19888 4007
rect 19908 3987 19917 4007
rect 19779 3980 19917 3987
rect 19975 4007 20123 4016
rect 19975 3987 19984 4007
rect 20004 3987 20094 4007
rect 20114 3987 20123 4007
rect 19779 3978 19875 3980
rect 19975 3977 20123 3987
rect 20182 4007 20219 4017
rect 20182 3987 20190 4007
rect 20210 3987 20219 4007
rect 20031 3976 20067 3977
rect 19879 3917 19916 3918
rect 20182 3917 20219 3987
rect 20254 4016 20285 4067
rect 21079 4056 21479 4074
rect 21497 4056 21518 4074
rect 21079 4050 21518 4056
rect 21085 4046 21518 4050
rect 21900 4079 22043 4100
rect 22087 4152 22121 4168
rect 22305 4158 22698 4178
rect 22718 4158 22721 4178
rect 23036 4171 23067 4192
rect 23254 4171 23290 4281
rect 23309 4280 23346 4281
rect 23405 4280 23442 4281
rect 23365 4221 23455 4227
rect 23365 4201 23374 4221
rect 23394 4219 23455 4221
rect 23394 4201 23419 4219
rect 23365 4199 23419 4201
rect 23439 4199 23455 4219
rect 23365 4193 23455 4199
rect 22879 4170 22916 4171
rect 22305 4153 22721 4158
rect 22878 4161 22916 4170
rect 22305 4152 22646 4153
rect 22087 4082 22124 4152
rect 22239 4092 22270 4093
rect 21900 4077 22037 4079
rect 21464 4044 21516 4046
rect 21900 4035 21943 4077
rect 22087 4062 22096 4082
rect 22116 4062 22124 4082
rect 22087 4052 22124 4062
rect 22183 4082 22270 4092
rect 22183 4062 22192 4082
rect 22212 4062 22270 4082
rect 22183 4053 22270 4062
rect 22183 4052 22220 4053
rect 21898 4025 21943 4035
rect 20304 4016 20341 4017
rect 20254 4007 20341 4016
rect 20254 3987 20312 4007
rect 20332 3987 20341 4007
rect 20254 3977 20341 3987
rect 20400 4007 20437 4017
rect 20400 3987 20408 4007
rect 20428 3987 20437 4007
rect 21898 4007 21907 4025
rect 21925 4007 21943 4025
rect 21898 4001 21943 4007
rect 22239 4002 22270 4053
rect 22305 4082 22342 4152
rect 22608 4151 22645 4152
rect 22878 4141 22887 4161
rect 22907 4141 22916 4161
rect 22878 4133 22916 4141
rect 22982 4165 23067 4171
rect 23097 4170 23134 4171
rect 22982 4145 22990 4165
rect 23010 4145 23067 4165
rect 22982 4137 23067 4145
rect 23096 4161 23134 4170
rect 23096 4141 23105 4161
rect 23125 4141 23134 4161
rect 22982 4136 23018 4137
rect 23096 4133 23134 4141
rect 23200 4165 23344 4171
rect 23200 4145 23208 4165
rect 23228 4146 23260 4165
rect 23281 4146 23316 4165
rect 23228 4145 23316 4146
rect 23336 4145 23344 4165
rect 23200 4137 23344 4145
rect 23200 4136 23236 4137
rect 23308 4136 23344 4137
rect 23410 4170 23447 4171
rect 23410 4169 23448 4170
rect 23410 4161 23474 4169
rect 23410 4141 23419 4161
rect 23439 4147 23474 4161
rect 23494 4147 23497 4167
rect 23439 4142 23497 4147
rect 23439 4141 23474 4142
rect 22879 4104 22916 4133
rect 22880 4102 22916 4104
rect 22457 4092 22493 4093
rect 22305 4062 22314 4082
rect 22334 4062 22342 4082
rect 22305 4052 22342 4062
rect 22401 4082 22549 4092
rect 22649 4089 22745 4091
rect 22401 4062 22410 4082
rect 22430 4062 22520 4082
rect 22540 4062 22549 4082
rect 22401 4053 22549 4062
rect 22607 4082 22745 4089
rect 22607 4062 22616 4082
rect 22636 4062 22745 4082
rect 22880 4080 23071 4102
rect 23097 4101 23134 4133
rect 23410 4129 23474 4141
rect 23514 4103 23541 4281
rect 23373 4101 23541 4103
rect 23097 4075 23541 4101
rect 22607 4053 22745 4062
rect 22401 4052 22438 4053
rect 21898 3998 21935 4001
rect 22131 3999 22172 4000
rect 20254 3976 20285 3977
rect 19878 3916 20219 3917
rect 20400 3916 20437 3987
rect 22023 3992 22172 3999
rect 21467 3979 21504 3984
rect 21458 3975 21505 3979
rect 21458 3957 21477 3975
rect 21495 3957 21505 3975
rect 22023 3972 22082 3992
rect 22102 3972 22141 3992
rect 22161 3972 22172 3992
rect 22023 3964 22172 3972
rect 22239 3995 22396 4002
rect 22239 3975 22359 3995
rect 22379 3975 22396 3995
rect 22239 3965 22396 3975
rect 22239 3964 22274 3965
rect 19803 3911 20219 3916
rect 19803 3891 19806 3911
rect 19826 3891 20219 3911
rect 20250 3892 20437 3916
rect 21062 3914 21102 3919
rect 21458 3914 21505 3957
rect 22239 3943 22270 3964
rect 22457 3943 22493 4053
rect 22512 4052 22549 4053
rect 22608 4052 22645 4053
rect 22568 3993 22658 3999
rect 22568 3973 22577 3993
rect 22597 3991 22658 3993
rect 22597 3973 22622 3991
rect 22568 3971 22622 3973
rect 22642 3971 22658 3991
rect 22568 3965 22658 3971
rect 22082 3942 22119 3943
rect 21062 3875 21505 3914
rect 21895 3934 21932 3936
rect 21895 3926 21937 3934
rect 21895 3908 21905 3926
rect 21923 3908 21937 3926
rect 21895 3899 21937 3908
rect 22081 3933 22119 3942
rect 22081 3913 22090 3933
rect 22110 3913 22119 3933
rect 22081 3905 22119 3913
rect 22185 3937 22270 3943
rect 22300 3942 22337 3943
rect 22185 3917 22193 3937
rect 22213 3917 22270 3937
rect 22185 3909 22270 3917
rect 22299 3933 22337 3942
rect 22299 3913 22308 3933
rect 22328 3913 22337 3933
rect 22185 3908 22221 3909
rect 22299 3905 22337 3913
rect 22403 3941 22547 3943
rect 22403 3937 22455 3941
rect 22403 3917 22411 3937
rect 22431 3921 22455 3937
rect 22475 3937 22547 3941
rect 22475 3921 22519 3937
rect 22431 3917 22519 3921
rect 22539 3917 22547 3937
rect 22403 3909 22547 3917
rect 22403 3908 22439 3909
rect 22511 3908 22547 3909
rect 22613 3942 22650 3943
rect 22613 3941 22651 3942
rect 22613 3933 22677 3941
rect 22613 3913 22622 3933
rect 22642 3919 22677 3933
rect 22697 3919 22700 3939
rect 22642 3914 22700 3919
rect 22642 3913 22677 3914
rect 20156 3860 20196 3868
rect 20156 3838 20164 3860
rect 20188 3838 20196 3860
rect 19862 3614 20030 3615
rect 20156 3614 20196 3838
rect 20659 3842 20827 3843
rect 21062 3842 21102 3875
rect 21458 3842 21505 3875
rect 21896 3874 21937 3899
rect 22082 3874 22119 3905
rect 22300 3874 22337 3905
rect 22613 3901 22677 3913
rect 22717 3875 22744 4053
rect 21896 3847 21945 3874
rect 22081 3848 22130 3874
rect 22299 3873 22380 3874
rect 22576 3873 22744 3875
rect 22299 3848 22744 3873
rect 22300 3847 22744 3848
rect 20659 3841 21103 3842
rect 20659 3816 21104 3841
rect 20659 3814 20827 3816
rect 21023 3815 21104 3816
rect 21273 3815 21322 3841
rect 21458 3815 21507 3842
rect 20659 3636 20686 3814
rect 20726 3776 20790 3788
rect 21066 3784 21103 3815
rect 21284 3784 21321 3815
rect 21466 3790 21507 3815
rect 21898 3814 21945 3847
rect 22301 3814 22341 3847
rect 22576 3846 22744 3847
rect 23207 3851 23247 4075
rect 23373 4074 23541 4075
rect 23207 3829 23215 3851
rect 23239 3829 23247 3851
rect 23207 3821 23247 3829
rect 20726 3775 20761 3776
rect 20703 3770 20761 3775
rect 20703 3750 20706 3770
rect 20726 3756 20761 3770
rect 20781 3756 20790 3776
rect 20726 3748 20790 3756
rect 20752 3747 20790 3748
rect 20753 3746 20790 3747
rect 20856 3780 20892 3781
rect 20964 3780 21000 3781
rect 20856 3772 21000 3780
rect 20856 3752 20864 3772
rect 20884 3768 20972 3772
rect 20884 3752 20928 3768
rect 20856 3748 20928 3752
rect 20948 3752 20972 3768
rect 20992 3752 21000 3772
rect 20948 3748 21000 3752
rect 20856 3746 21000 3748
rect 21066 3776 21104 3784
rect 21182 3780 21218 3781
rect 21066 3756 21075 3776
rect 21095 3756 21104 3776
rect 21066 3747 21104 3756
rect 21133 3772 21218 3780
rect 21133 3752 21190 3772
rect 21210 3752 21218 3772
rect 21066 3746 21103 3747
rect 21133 3746 21218 3752
rect 21284 3776 21322 3784
rect 21284 3756 21293 3776
rect 21313 3756 21322 3776
rect 21284 3747 21322 3756
rect 21466 3781 21508 3790
rect 21466 3763 21480 3781
rect 21498 3763 21508 3781
rect 21466 3755 21508 3763
rect 21471 3753 21508 3755
rect 21898 3775 22341 3814
rect 21284 3746 21321 3747
rect 20745 3718 20835 3724
rect 20745 3698 20761 3718
rect 20781 3716 20835 3718
rect 20781 3698 20806 3716
rect 20745 3696 20806 3698
rect 20826 3696 20835 3716
rect 20745 3690 20835 3696
rect 20758 3636 20795 3637
rect 20854 3636 20891 3637
rect 20910 3636 20946 3746
rect 21133 3725 21164 3746
rect 21898 3732 21945 3775
rect 22301 3770 22341 3775
rect 22966 3773 23153 3797
rect 23184 3778 23577 3798
rect 23597 3778 23600 3798
rect 23184 3773 23600 3778
rect 21129 3724 21164 3725
rect 21007 3714 21164 3724
rect 21007 3694 21024 3714
rect 21044 3694 21164 3714
rect 21007 3687 21164 3694
rect 21231 3717 21380 3725
rect 21231 3697 21242 3717
rect 21262 3697 21301 3717
rect 21321 3697 21380 3717
rect 21898 3714 21908 3732
rect 21926 3714 21945 3732
rect 21898 3710 21945 3714
rect 21899 3705 21936 3710
rect 21231 3690 21380 3697
rect 22966 3702 23003 3773
rect 23184 3772 23525 3773
rect 23118 3712 23149 3713
rect 21231 3689 21272 3690
rect 21468 3688 21505 3691
rect 20965 3636 21002 3637
rect 20658 3627 20796 3636
rect 19862 3588 20306 3614
rect 19862 3586 20030 3588
rect 19862 3408 19889 3586
rect 19929 3548 19993 3560
rect 20269 3556 20306 3588
rect 20332 3587 20523 3609
rect 20658 3607 20767 3627
rect 20787 3607 20796 3627
rect 20658 3600 20796 3607
rect 20854 3627 21002 3636
rect 20854 3607 20863 3627
rect 20883 3607 20973 3627
rect 20993 3607 21002 3627
rect 20658 3598 20754 3600
rect 20854 3597 21002 3607
rect 21061 3627 21098 3637
rect 21061 3607 21069 3627
rect 21089 3607 21098 3627
rect 20910 3596 20946 3597
rect 20487 3585 20523 3587
rect 20487 3556 20524 3585
rect 19929 3547 19964 3548
rect 19906 3542 19964 3547
rect 19906 3522 19909 3542
rect 19929 3528 19964 3542
rect 19984 3528 19993 3548
rect 19929 3520 19993 3528
rect 19955 3519 19993 3520
rect 19956 3518 19993 3519
rect 20059 3552 20095 3553
rect 20167 3552 20203 3553
rect 20059 3544 20203 3552
rect 20059 3524 20067 3544
rect 20087 3543 20175 3544
rect 20087 3524 20122 3543
rect 20143 3524 20175 3543
rect 20195 3524 20203 3544
rect 20059 3518 20203 3524
rect 20269 3548 20307 3556
rect 20385 3552 20421 3553
rect 20269 3528 20278 3548
rect 20298 3528 20307 3548
rect 20269 3519 20307 3528
rect 20336 3544 20421 3552
rect 20336 3524 20393 3544
rect 20413 3524 20421 3544
rect 20269 3518 20306 3519
rect 20336 3518 20421 3524
rect 20487 3548 20525 3556
rect 20487 3528 20496 3548
rect 20516 3528 20525 3548
rect 20758 3537 20795 3538
rect 21061 3537 21098 3607
rect 21133 3636 21164 3687
rect 21460 3682 21505 3688
rect 21460 3664 21478 3682
rect 21496 3664 21505 3682
rect 22966 3682 22975 3702
rect 22995 3682 23003 3702
rect 22966 3672 23003 3682
rect 23062 3702 23149 3712
rect 23062 3682 23071 3702
rect 23091 3682 23149 3702
rect 23062 3673 23149 3682
rect 23062 3672 23099 3673
rect 21460 3654 21505 3664
rect 21183 3636 21220 3637
rect 21133 3627 21220 3636
rect 21133 3607 21191 3627
rect 21211 3607 21220 3627
rect 21133 3597 21220 3607
rect 21279 3627 21316 3637
rect 21279 3607 21287 3627
rect 21307 3607 21316 3627
rect 21460 3612 21503 3654
rect 21887 3643 21939 3645
rect 21366 3610 21503 3612
rect 21133 3596 21164 3597
rect 21279 3537 21316 3607
rect 20757 3536 21098 3537
rect 20487 3519 20525 3528
rect 20682 3531 21098 3536
rect 20487 3518 20524 3519
rect 19948 3490 20038 3496
rect 19948 3470 19964 3490
rect 19984 3488 20038 3490
rect 19984 3470 20009 3488
rect 19948 3468 20009 3470
rect 20029 3468 20038 3488
rect 19948 3462 20038 3468
rect 19961 3408 19998 3409
rect 20057 3408 20094 3409
rect 20113 3408 20149 3518
rect 20336 3497 20367 3518
rect 20682 3511 20685 3531
rect 20705 3511 21098 3531
rect 21282 3521 21316 3537
rect 21360 3589 21503 3610
rect 21885 3639 22318 3643
rect 21885 3633 22324 3639
rect 21885 3615 21906 3633
rect 21924 3615 22324 3633
rect 23118 3622 23149 3673
rect 23184 3702 23221 3772
rect 23487 3771 23524 3772
rect 23336 3712 23372 3713
rect 23184 3682 23193 3702
rect 23213 3682 23221 3702
rect 23184 3672 23221 3682
rect 23280 3702 23428 3712
rect 23528 3709 23624 3711
rect 23280 3682 23289 3702
rect 23309 3682 23399 3702
rect 23419 3682 23428 3702
rect 23280 3673 23428 3682
rect 23486 3702 23624 3709
rect 23486 3682 23495 3702
rect 23515 3682 23624 3702
rect 23486 3673 23624 3682
rect 23280 3672 23317 3673
rect 23010 3619 23051 3620
rect 21885 3597 22324 3615
rect 21058 3502 21098 3511
rect 21360 3502 21387 3589
rect 21460 3563 21503 3589
rect 21460 3545 21473 3563
rect 21491 3545 21503 3563
rect 21460 3534 21503 3545
rect 20332 3496 20367 3497
rect 20210 3486 20367 3496
rect 20210 3466 20227 3486
rect 20247 3466 20367 3486
rect 20210 3459 20367 3466
rect 20434 3489 20583 3497
rect 20434 3469 20445 3489
rect 20465 3469 20504 3489
rect 20524 3469 20583 3489
rect 21058 3485 21387 3502
rect 21058 3484 21098 3485
rect 20434 3462 20583 3469
rect 21455 3473 21495 3476
rect 21455 3467 21498 3473
rect 21080 3464 21498 3467
rect 20434 3461 20475 3462
rect 20168 3408 20205 3409
rect 19861 3399 19999 3408
rect 19861 3379 19970 3399
rect 19990 3379 19999 3399
rect 19861 3372 19999 3379
rect 20057 3399 20205 3408
rect 20057 3379 20066 3399
rect 20086 3379 20176 3399
rect 20196 3379 20205 3399
rect 19861 3370 19957 3372
rect 20057 3369 20205 3379
rect 20264 3399 20301 3409
rect 20264 3379 20272 3399
rect 20292 3379 20301 3399
rect 20113 3368 20149 3369
rect 19961 3309 19998 3310
rect 20264 3309 20301 3379
rect 20336 3408 20367 3459
rect 21080 3446 21471 3464
rect 21489 3446 21498 3464
rect 21080 3444 21498 3446
rect 21080 3436 21107 3444
rect 21348 3441 21498 3444
rect 20660 3430 20828 3431
rect 21079 3430 21107 3436
rect 20660 3414 21107 3430
rect 21455 3436 21498 3441
rect 20386 3408 20423 3409
rect 20336 3399 20423 3408
rect 20336 3379 20394 3399
rect 20414 3379 20423 3399
rect 20336 3369 20423 3379
rect 20482 3399 20519 3409
rect 20482 3379 20490 3399
rect 20510 3379 20519 3399
rect 20336 3368 20367 3369
rect 19960 3308 20301 3309
rect 20482 3308 20519 3379
rect 19885 3303 20301 3308
rect 19885 3283 19888 3303
rect 19908 3283 20301 3303
rect 20332 3284 20519 3308
rect 20660 3404 21104 3414
rect 20660 3402 20828 3404
rect 19727 3209 19756 3227
rect 20660 3224 20687 3402
rect 20727 3364 20791 3376
rect 21067 3372 21104 3404
rect 21130 3403 21321 3425
rect 21285 3401 21321 3403
rect 21285 3372 21322 3401
rect 21455 3380 21495 3436
rect 20727 3363 20762 3364
rect 20704 3358 20762 3363
rect 20704 3338 20707 3358
rect 20727 3344 20762 3358
rect 20782 3344 20791 3364
rect 20727 3336 20791 3344
rect 20753 3335 20791 3336
rect 20754 3334 20791 3335
rect 20857 3368 20893 3369
rect 20965 3368 21001 3369
rect 20857 3360 21001 3368
rect 20857 3340 20865 3360
rect 20885 3340 20920 3360
rect 20940 3340 20973 3360
rect 20993 3340 21001 3360
rect 20857 3334 21001 3340
rect 21067 3364 21105 3372
rect 21183 3368 21219 3369
rect 21067 3344 21076 3364
rect 21096 3344 21105 3364
rect 21067 3335 21105 3344
rect 21134 3360 21219 3368
rect 21134 3340 21191 3360
rect 21211 3340 21219 3360
rect 21067 3334 21104 3335
rect 21134 3334 21219 3340
rect 21285 3364 21323 3372
rect 21285 3344 21294 3364
rect 21314 3344 21323 3364
rect 21455 3362 21467 3380
rect 21485 3362 21495 3380
rect 21887 3408 21939 3597
rect 22285 3572 22324 3597
rect 22902 3612 23051 3619
rect 22902 3592 22961 3612
rect 22981 3592 23020 3612
rect 23040 3592 23051 3612
rect 22902 3584 23051 3592
rect 23118 3615 23275 3622
rect 23118 3595 23238 3615
rect 23258 3595 23275 3615
rect 23118 3585 23275 3595
rect 23118 3584 23153 3585
rect 22069 3547 22256 3571
rect 22285 3552 22680 3572
rect 22700 3552 22703 3572
rect 23118 3563 23149 3584
rect 23336 3563 23372 3673
rect 23391 3672 23428 3673
rect 23487 3672 23524 3673
rect 23447 3613 23537 3619
rect 23447 3593 23456 3613
rect 23476 3611 23537 3613
rect 23476 3593 23501 3611
rect 23447 3591 23501 3593
rect 23521 3591 23537 3611
rect 23447 3585 23537 3591
rect 22961 3562 22998 3563
rect 22285 3547 22703 3552
rect 22960 3553 22998 3562
rect 22069 3476 22106 3547
rect 22285 3546 22628 3547
rect 22285 3543 22324 3546
rect 22590 3545 22627 3546
rect 22221 3486 22252 3487
rect 22069 3456 22078 3476
rect 22098 3456 22106 3476
rect 22069 3446 22106 3456
rect 22165 3476 22252 3486
rect 22165 3456 22174 3476
rect 22194 3456 22252 3476
rect 22165 3447 22252 3456
rect 22165 3446 22202 3447
rect 21887 3390 21903 3408
rect 21921 3390 21939 3408
rect 22221 3396 22252 3447
rect 22287 3476 22324 3543
rect 22960 3533 22969 3553
rect 22989 3533 22998 3553
rect 22960 3525 22998 3533
rect 23064 3557 23149 3563
rect 23179 3562 23216 3563
rect 23064 3537 23072 3557
rect 23092 3537 23149 3557
rect 23064 3529 23149 3537
rect 23178 3553 23216 3562
rect 23178 3533 23187 3553
rect 23207 3533 23216 3553
rect 23064 3528 23100 3529
rect 23178 3525 23216 3533
rect 23282 3558 23426 3563
rect 23282 3557 23344 3558
rect 23282 3537 23290 3557
rect 23310 3539 23344 3557
rect 23365 3557 23426 3558
rect 23365 3539 23398 3557
rect 23310 3537 23398 3539
rect 23418 3537 23426 3557
rect 23282 3529 23426 3537
rect 23282 3528 23318 3529
rect 23390 3528 23426 3529
rect 23492 3562 23529 3563
rect 23492 3561 23530 3562
rect 23492 3553 23556 3561
rect 23492 3533 23501 3553
rect 23521 3539 23556 3553
rect 23576 3539 23579 3559
rect 23521 3534 23579 3539
rect 23521 3533 23556 3534
rect 22961 3496 22998 3525
rect 22962 3494 22998 3496
rect 22439 3486 22475 3487
rect 22287 3456 22296 3476
rect 22316 3456 22324 3476
rect 22287 3446 22324 3456
rect 22383 3476 22531 3486
rect 22631 3483 22727 3485
rect 22383 3456 22392 3476
rect 22412 3456 22502 3476
rect 22522 3456 22531 3476
rect 22383 3447 22531 3456
rect 22589 3476 22727 3483
rect 22589 3456 22598 3476
rect 22618 3456 22727 3476
rect 22962 3472 23153 3494
rect 23179 3493 23216 3525
rect 23492 3521 23556 3533
rect 23596 3495 23623 3673
rect 23455 3493 23623 3495
rect 23179 3479 23623 3493
rect 23179 3467 23626 3479
rect 23222 3465 23255 3467
rect 22589 3447 22727 3456
rect 22383 3446 22420 3447
rect 22113 3393 22154 3394
rect 21887 3372 21939 3390
rect 22005 3386 22154 3393
rect 21455 3352 21495 3362
rect 22005 3366 22064 3386
rect 22084 3366 22123 3386
rect 22143 3366 22154 3386
rect 22005 3358 22154 3366
rect 22221 3389 22378 3396
rect 22221 3369 22341 3389
rect 22361 3369 22378 3389
rect 22221 3359 22378 3369
rect 22221 3358 22256 3359
rect 21285 3335 21323 3344
rect 22221 3337 22252 3358
rect 22439 3337 22475 3447
rect 22494 3446 22531 3447
rect 22590 3446 22627 3447
rect 22550 3387 22640 3393
rect 22550 3367 22559 3387
rect 22579 3385 22640 3387
rect 22579 3367 22604 3385
rect 22550 3365 22604 3367
rect 22624 3365 22640 3385
rect 22550 3359 22640 3365
rect 22064 3336 22101 3337
rect 21285 3334 21322 3335
rect 20746 3306 20836 3312
rect 20746 3286 20762 3306
rect 20782 3304 20836 3306
rect 20782 3286 20807 3304
rect 20746 3284 20807 3286
rect 20827 3284 20836 3304
rect 20746 3278 20836 3284
rect 20759 3224 20796 3225
rect 20855 3224 20892 3225
rect 20911 3224 20947 3334
rect 21134 3313 21165 3334
rect 22063 3327 22101 3336
rect 21130 3312 21165 3313
rect 21008 3302 21165 3312
rect 21008 3282 21025 3302
rect 21045 3282 21165 3302
rect 21008 3275 21165 3282
rect 21232 3305 21381 3313
rect 21232 3285 21243 3305
rect 21263 3285 21302 3305
rect 21322 3285 21381 3305
rect 21891 3309 21931 3319
rect 21232 3278 21381 3285
rect 21447 3281 21499 3299
rect 21232 3277 21273 3278
rect 20966 3224 21003 3225
rect 19697 3207 19756 3209
rect 20659 3215 20797 3224
rect 19697 3206 19865 3207
rect 19991 3206 20031 3208
rect 19697 3180 20141 3206
rect 19697 3178 19865 3180
rect 19697 3176 19778 3178
rect 19697 3000 19724 3176
rect 19764 3140 19828 3152
rect 20104 3148 20141 3180
rect 20167 3179 20358 3201
rect 20659 3195 20768 3215
rect 20788 3195 20797 3215
rect 20659 3188 20797 3195
rect 20855 3215 21003 3224
rect 20855 3195 20864 3215
rect 20884 3195 20974 3215
rect 20994 3195 21003 3215
rect 20659 3186 20755 3188
rect 20855 3185 21003 3195
rect 21062 3215 21099 3225
rect 21062 3195 21070 3215
rect 21090 3195 21099 3215
rect 20911 3184 20947 3185
rect 20322 3177 20358 3179
rect 20322 3148 20359 3177
rect 19764 3139 19799 3140
rect 19741 3134 19799 3139
rect 19741 3114 19744 3134
rect 19764 3120 19799 3134
rect 19819 3120 19828 3140
rect 19764 3112 19828 3120
rect 19790 3111 19828 3112
rect 19791 3110 19828 3111
rect 19894 3144 19930 3145
rect 20002 3144 20038 3145
rect 19894 3136 20038 3144
rect 19894 3116 19902 3136
rect 19922 3135 20010 3136
rect 19922 3117 19957 3135
rect 19975 3117 20010 3135
rect 19922 3116 20010 3117
rect 20030 3116 20038 3136
rect 19894 3110 20038 3116
rect 20104 3140 20142 3148
rect 20220 3144 20256 3145
rect 20104 3120 20113 3140
rect 20133 3120 20142 3140
rect 20104 3111 20142 3120
rect 20171 3136 20256 3144
rect 20171 3116 20228 3136
rect 20248 3116 20256 3136
rect 20104 3110 20141 3111
rect 20171 3110 20256 3116
rect 20322 3140 20360 3148
rect 20322 3120 20331 3140
rect 20351 3120 20360 3140
rect 21062 3128 21099 3195
rect 21134 3224 21165 3275
rect 21447 3263 21465 3281
rect 21483 3263 21499 3281
rect 21184 3224 21221 3225
rect 21134 3215 21221 3224
rect 21134 3195 21192 3215
rect 21212 3195 21221 3215
rect 21134 3185 21221 3195
rect 21280 3215 21317 3225
rect 21280 3195 21288 3215
rect 21308 3195 21317 3215
rect 21134 3184 21165 3185
rect 20759 3125 20796 3126
rect 21062 3125 21101 3128
rect 20758 3124 21101 3125
rect 21280 3124 21317 3195
rect 20322 3111 20360 3120
rect 20683 3119 21101 3124
rect 20322 3110 20359 3111
rect 19783 3082 19873 3088
rect 19783 3062 19799 3082
rect 19819 3080 19873 3082
rect 19819 3062 19844 3080
rect 19783 3060 19844 3062
rect 19864 3060 19873 3080
rect 19783 3054 19873 3060
rect 19796 3000 19833 3001
rect 19892 3000 19929 3001
rect 19948 3000 19984 3110
rect 20171 3089 20202 3110
rect 20683 3099 20686 3119
rect 20706 3099 21101 3119
rect 21130 3100 21317 3124
rect 20167 3088 20202 3089
rect 20045 3078 20202 3088
rect 20045 3058 20062 3078
rect 20082 3058 20202 3078
rect 20045 3051 20202 3058
rect 20269 3081 20418 3089
rect 20269 3061 20280 3081
rect 20300 3061 20339 3081
rect 20359 3061 20418 3081
rect 20269 3054 20418 3061
rect 21062 3074 21101 3099
rect 21447 3074 21499 3263
rect 21891 3291 21901 3309
rect 21919 3291 21931 3309
rect 22063 3307 22072 3327
rect 22092 3307 22101 3327
rect 22063 3299 22101 3307
rect 22167 3331 22252 3337
rect 22282 3336 22319 3337
rect 22167 3311 22175 3331
rect 22195 3311 22252 3331
rect 22167 3303 22252 3311
rect 22281 3327 22319 3336
rect 22281 3307 22290 3327
rect 22310 3307 22319 3327
rect 22167 3302 22203 3303
rect 22281 3299 22319 3307
rect 22385 3331 22529 3337
rect 22385 3311 22393 3331
rect 22413 3311 22446 3331
rect 22466 3311 22501 3331
rect 22521 3311 22529 3331
rect 22385 3303 22529 3311
rect 22385 3302 22421 3303
rect 22493 3302 22529 3303
rect 22595 3336 22632 3337
rect 22595 3335 22633 3336
rect 22595 3327 22659 3335
rect 22595 3307 22604 3327
rect 22624 3313 22659 3327
rect 22679 3313 22682 3333
rect 22624 3308 22682 3313
rect 22624 3307 22659 3308
rect 21891 3235 21931 3291
rect 22064 3270 22101 3299
rect 22065 3268 22101 3270
rect 22065 3246 22256 3268
rect 22282 3267 22319 3299
rect 22595 3295 22659 3307
rect 22699 3269 22726 3447
rect 23584 3422 23626 3467
rect 22558 3267 22726 3269
rect 22282 3257 22726 3267
rect 22867 3363 23054 3387
rect 23085 3368 23478 3388
rect 23498 3368 23501 3388
rect 23085 3363 23501 3368
rect 22867 3292 22904 3363
rect 23085 3362 23426 3363
rect 23019 3302 23050 3303
rect 22867 3272 22876 3292
rect 22896 3272 22904 3292
rect 22867 3262 22904 3272
rect 22963 3292 23050 3302
rect 22963 3272 22972 3292
rect 22992 3272 23050 3292
rect 22963 3263 23050 3272
rect 22963 3262 23000 3263
rect 21888 3230 21931 3235
rect 22279 3241 22726 3257
rect 22279 3235 22307 3241
rect 22558 3240 22726 3241
rect 21888 3227 22038 3230
rect 22279 3227 22306 3235
rect 21888 3225 22306 3227
rect 21888 3207 21897 3225
rect 21915 3207 22306 3225
rect 23019 3212 23050 3263
rect 23085 3292 23122 3362
rect 23388 3361 23425 3362
rect 23237 3302 23273 3303
rect 23085 3272 23094 3292
rect 23114 3272 23122 3292
rect 23085 3262 23122 3272
rect 23181 3292 23329 3302
rect 23429 3299 23525 3301
rect 23181 3272 23190 3292
rect 23210 3272 23300 3292
rect 23320 3272 23329 3292
rect 23181 3263 23329 3272
rect 23387 3292 23525 3299
rect 23387 3272 23396 3292
rect 23416 3272 23525 3292
rect 23387 3263 23525 3272
rect 23181 3262 23218 3263
rect 22911 3209 22952 3210
rect 21888 3204 22306 3207
rect 21888 3198 21931 3204
rect 21891 3195 21931 3198
rect 22806 3202 22952 3209
rect 22288 3186 22328 3187
rect 21999 3169 22328 3186
rect 22806 3182 22862 3202
rect 22882 3182 22921 3202
rect 22941 3182 22952 3202
rect 22806 3174 22952 3182
rect 23019 3205 23176 3212
rect 23019 3185 23139 3205
rect 23159 3185 23176 3205
rect 23019 3175 23176 3185
rect 23019 3174 23054 3175
rect 21883 3126 21926 3137
rect 21883 3108 21895 3126
rect 21913 3108 21926 3126
rect 21883 3082 21926 3108
rect 21999 3082 22026 3169
rect 22288 3160 22328 3169
rect 21062 3056 21501 3074
rect 20269 3053 20310 3054
rect 20003 3000 20040 3001
rect 19696 2991 19834 3000
rect 19696 2971 19805 2991
rect 19825 2971 19834 2991
rect 19696 2964 19834 2971
rect 19892 2991 20040 3000
rect 19892 2971 19901 2991
rect 19921 2971 20011 2991
rect 20031 2971 20040 2991
rect 19696 2962 19792 2964
rect 19892 2961 20040 2971
rect 20099 2991 20136 3001
rect 20099 2971 20107 2991
rect 20127 2971 20136 2991
rect 19948 2960 19984 2961
rect 19796 2901 19833 2902
rect 20099 2901 20136 2971
rect 20171 3000 20202 3051
rect 21062 3038 21462 3056
rect 21480 3038 21501 3056
rect 21062 3032 21501 3038
rect 21068 3028 21501 3032
rect 21883 3061 22026 3082
rect 22070 3134 22104 3150
rect 22288 3140 22681 3160
rect 22701 3140 22704 3160
rect 23019 3153 23050 3174
rect 23237 3153 23273 3263
rect 23292 3262 23329 3263
rect 23388 3262 23425 3263
rect 23348 3203 23438 3209
rect 23348 3183 23357 3203
rect 23377 3201 23438 3203
rect 23377 3183 23402 3201
rect 23348 3181 23402 3183
rect 23422 3181 23438 3201
rect 23348 3175 23438 3181
rect 22862 3152 22899 3153
rect 22288 3135 22704 3140
rect 22861 3143 22899 3152
rect 22288 3134 22629 3135
rect 22070 3064 22107 3134
rect 22222 3074 22253 3075
rect 21883 3059 22020 3061
rect 21447 3026 21499 3028
rect 21883 3017 21926 3059
rect 22070 3044 22079 3064
rect 22099 3044 22107 3064
rect 22070 3034 22107 3044
rect 22166 3064 22253 3074
rect 22166 3044 22175 3064
rect 22195 3044 22253 3064
rect 22166 3035 22253 3044
rect 22166 3034 22203 3035
rect 21881 3007 21926 3017
rect 20221 3000 20258 3001
rect 20171 2991 20258 3000
rect 20171 2971 20229 2991
rect 20249 2971 20258 2991
rect 20171 2961 20258 2971
rect 20317 2991 20354 3001
rect 20317 2971 20325 2991
rect 20345 2971 20354 2991
rect 21881 2989 21890 3007
rect 21908 2989 21926 3007
rect 21881 2983 21926 2989
rect 22222 2984 22253 3035
rect 22288 3064 22325 3134
rect 22591 3133 22628 3134
rect 22861 3123 22870 3143
rect 22890 3123 22899 3143
rect 22861 3115 22899 3123
rect 22965 3147 23050 3153
rect 23080 3152 23117 3153
rect 22965 3127 22973 3147
rect 22993 3127 23050 3147
rect 22965 3119 23050 3127
rect 23079 3143 23117 3152
rect 23079 3123 23088 3143
rect 23108 3123 23117 3143
rect 22965 3118 23001 3119
rect 23079 3115 23117 3123
rect 23183 3147 23327 3153
rect 23183 3127 23191 3147
rect 23211 3144 23299 3147
rect 23211 3127 23246 3144
rect 23183 3126 23246 3127
rect 23265 3127 23299 3144
rect 23319 3127 23327 3147
rect 23265 3126 23327 3127
rect 23183 3119 23327 3126
rect 23183 3118 23219 3119
rect 23291 3118 23327 3119
rect 23393 3152 23430 3153
rect 23393 3151 23431 3152
rect 23453 3151 23480 3155
rect 23393 3149 23480 3151
rect 23393 3143 23457 3149
rect 23393 3123 23402 3143
rect 23422 3129 23457 3143
rect 23477 3129 23480 3149
rect 23422 3124 23480 3129
rect 23422 3123 23457 3124
rect 22862 3086 22899 3115
rect 22863 3084 22899 3086
rect 22440 3074 22476 3075
rect 22288 3044 22297 3064
rect 22317 3044 22325 3064
rect 22288 3034 22325 3044
rect 22384 3064 22532 3074
rect 22632 3071 22728 3073
rect 22384 3044 22393 3064
rect 22413 3044 22503 3064
rect 22523 3044 22532 3064
rect 22384 3035 22532 3044
rect 22590 3064 22728 3071
rect 22590 3044 22599 3064
rect 22619 3044 22728 3064
rect 22863 3062 23054 3084
rect 23080 3083 23117 3115
rect 23393 3111 23457 3123
rect 23497 3085 23524 3263
rect 23356 3083 23524 3085
rect 23080 3057 23524 3083
rect 22590 3035 22728 3044
rect 22384 3034 22421 3035
rect 21881 2980 21918 2983
rect 22114 2981 22155 2982
rect 20171 2960 20202 2961
rect 19795 2900 20136 2901
rect 20317 2900 20354 2971
rect 22006 2974 22155 2981
rect 21450 2961 21487 2966
rect 19720 2895 20136 2900
rect 19720 2875 19723 2895
rect 19743 2875 20136 2895
rect 20167 2876 20354 2900
rect 21441 2957 21488 2961
rect 21441 2939 21460 2957
rect 21478 2939 21488 2957
rect 22006 2954 22065 2974
rect 22085 2954 22124 2974
rect 22144 2954 22155 2974
rect 22006 2946 22155 2954
rect 22222 2977 22379 2984
rect 22222 2957 22342 2977
rect 22362 2957 22379 2977
rect 22222 2947 22379 2957
rect 22222 2946 22257 2947
rect 21441 2891 21488 2939
rect 22222 2925 22253 2946
rect 22440 2925 22476 3035
rect 22495 3034 22532 3035
rect 22591 3034 22628 3035
rect 22551 2975 22641 2981
rect 22551 2955 22560 2975
rect 22580 2973 22641 2975
rect 22580 2955 22605 2973
rect 22551 2953 22605 2955
rect 22625 2953 22641 2973
rect 22551 2947 22641 2953
rect 22065 2924 22102 2925
rect 21065 2888 21488 2891
rect 19940 2874 20005 2875
rect 21043 2858 21488 2888
rect 21877 2916 21915 2918
rect 21877 2908 21920 2916
rect 21877 2890 21888 2908
rect 21906 2890 21920 2908
rect 21877 2863 21920 2890
rect 22064 2915 22102 2924
rect 22064 2895 22073 2915
rect 22093 2895 22102 2915
rect 22064 2887 22102 2895
rect 22168 2919 22253 2925
rect 22283 2924 22320 2925
rect 22168 2899 22176 2919
rect 22196 2899 22253 2919
rect 22168 2891 22253 2899
rect 22282 2915 22320 2924
rect 22282 2895 22291 2915
rect 22311 2895 22320 2915
rect 22168 2890 22204 2891
rect 22282 2887 22320 2895
rect 22386 2923 22530 2925
rect 22386 2919 22438 2923
rect 22386 2899 22394 2919
rect 22414 2903 22438 2919
rect 22458 2919 22530 2923
rect 22458 2903 22502 2919
rect 22414 2899 22502 2903
rect 22522 2899 22530 2919
rect 22386 2891 22530 2899
rect 22386 2890 22422 2891
rect 22494 2890 22530 2891
rect 22596 2924 22633 2925
rect 22596 2923 22634 2924
rect 22596 2915 22660 2923
rect 22596 2895 22605 2915
rect 22625 2901 22660 2915
rect 22680 2901 22683 2921
rect 22625 2896 22683 2901
rect 22625 2895 22660 2896
rect 20136 2842 20176 2850
rect 20136 2820 20144 2842
rect 20168 2820 20176 2842
rect 19741 2591 19778 2597
rect 19741 2572 19749 2591
rect 19770 2572 19778 2591
rect 19741 2564 19778 2572
rect 19441 2443 19448 2465
rect 19472 2443 19480 2465
rect 19441 2437 19480 2443
rect 18971 2432 19011 2434
rect 19137 2433 19305 2434
rect 19239 2432 19276 2433
rect 18205 2416 18343 2425
rect 17999 2415 18036 2416
rect 17729 2362 17770 2363
rect 16999 2342 17036 2343
rect 16460 2314 16550 2320
rect 16460 2294 16476 2314
rect 16496 2312 16550 2314
rect 16496 2294 16521 2312
rect 16460 2292 16521 2294
rect 16541 2292 16550 2312
rect 16460 2286 16550 2292
rect 16473 2232 16510 2233
rect 16569 2232 16606 2233
rect 16625 2232 16661 2342
rect 16848 2321 16879 2342
rect 17503 2341 17555 2359
rect 17621 2355 17770 2362
rect 17621 2335 17680 2355
rect 17700 2335 17739 2355
rect 17759 2335 17770 2355
rect 17621 2327 17770 2335
rect 17837 2358 17994 2365
rect 17837 2338 17957 2358
rect 17977 2338 17994 2358
rect 17837 2328 17994 2338
rect 17837 2327 17872 2328
rect 16844 2320 16879 2321
rect 16722 2310 16879 2320
rect 16722 2290 16739 2310
rect 16759 2290 16879 2310
rect 16722 2283 16879 2290
rect 16946 2313 17095 2321
rect 16946 2293 16957 2313
rect 16977 2293 17016 2313
rect 17036 2293 17095 2313
rect 16946 2286 17095 2293
rect 17161 2289 17213 2307
rect 17837 2306 17868 2327
rect 18055 2306 18091 2416
rect 18110 2415 18147 2416
rect 18206 2415 18243 2416
rect 18166 2356 18256 2362
rect 18166 2336 18175 2356
rect 18195 2354 18256 2356
rect 18195 2336 18220 2354
rect 18166 2334 18220 2336
rect 18240 2334 18256 2354
rect 18166 2328 18256 2334
rect 17680 2305 17717 2306
rect 16946 2285 16987 2286
rect 16680 2232 16717 2233
rect 16373 2223 16511 2232
rect 15845 2212 15878 2214
rect 15474 2200 15921 2212
rect 14706 2078 14874 2080
rect 14430 2052 14874 2078
rect 13940 2030 14078 2039
rect 13734 2029 13771 2030
rect 13231 1975 13268 1978
rect 13464 1976 13505 1977
rect 11587 1953 11618 1954
rect 11211 1893 11552 1894
rect 11733 1893 11770 1964
rect 13356 1969 13505 1976
rect 12800 1956 12837 1961
rect 12791 1952 12838 1956
rect 12791 1934 12810 1952
rect 12828 1934 12838 1952
rect 13356 1949 13415 1969
rect 13435 1949 13474 1969
rect 13494 1949 13505 1969
rect 13356 1941 13505 1949
rect 13572 1972 13729 1979
rect 13572 1952 13692 1972
rect 13712 1952 13729 1972
rect 13572 1942 13729 1952
rect 13572 1941 13607 1942
rect 11136 1888 11552 1893
rect 11136 1868 11139 1888
rect 11159 1868 11552 1888
rect 11583 1869 11770 1893
rect 12395 1891 12435 1896
rect 12791 1891 12838 1934
rect 13572 1920 13603 1941
rect 13790 1920 13826 2030
rect 13845 2029 13882 2030
rect 13941 2029 13978 2030
rect 13901 1970 13991 1976
rect 13901 1950 13910 1970
rect 13930 1968 13991 1970
rect 13930 1950 13955 1968
rect 13901 1948 13955 1950
rect 13975 1948 13991 1968
rect 13901 1942 13991 1948
rect 13415 1919 13452 1920
rect 12395 1852 12838 1891
rect 13228 1911 13265 1913
rect 13228 1903 13270 1911
rect 13228 1885 13238 1903
rect 13256 1885 13270 1903
rect 13228 1876 13270 1885
rect 13414 1910 13452 1919
rect 13414 1890 13423 1910
rect 13443 1890 13452 1910
rect 13414 1882 13452 1890
rect 13518 1914 13603 1920
rect 13633 1919 13670 1920
rect 13518 1894 13526 1914
rect 13546 1894 13603 1914
rect 13518 1886 13603 1894
rect 13632 1910 13670 1919
rect 13632 1890 13641 1910
rect 13661 1890 13670 1910
rect 13518 1885 13554 1886
rect 13632 1882 13670 1890
rect 13736 1918 13880 1920
rect 13736 1914 13788 1918
rect 13736 1894 13744 1914
rect 13764 1898 13788 1914
rect 13808 1914 13880 1918
rect 13808 1898 13852 1914
rect 13764 1894 13852 1898
rect 13872 1894 13880 1914
rect 13736 1886 13880 1894
rect 13736 1885 13772 1886
rect 13844 1885 13880 1886
rect 13946 1919 13983 1920
rect 13946 1918 13984 1919
rect 13946 1910 14010 1918
rect 13946 1890 13955 1910
rect 13975 1896 14010 1910
rect 14030 1896 14033 1916
rect 13975 1891 14033 1896
rect 13975 1890 14010 1891
rect 10176 1793 10184 1815
rect 10208 1793 10216 1815
rect 10176 1785 10216 1793
rect 11489 1837 11529 1845
rect 11489 1815 11497 1837
rect 11521 1815 11529 1837
rect 7682 1740 7717 1741
rect 7659 1735 7717 1740
rect 7659 1715 7662 1735
rect 7682 1721 7717 1735
rect 7737 1721 7746 1741
rect 7682 1713 7746 1721
rect 7708 1712 7746 1713
rect 7709 1711 7746 1712
rect 7812 1745 7848 1746
rect 7920 1745 7956 1746
rect 7812 1737 7956 1745
rect 7812 1717 7820 1737
rect 7840 1733 7928 1737
rect 7840 1717 7884 1733
rect 7812 1713 7884 1717
rect 7904 1717 7928 1733
rect 7948 1717 7956 1737
rect 7904 1713 7956 1717
rect 7812 1711 7956 1713
rect 8022 1741 8060 1749
rect 8138 1745 8174 1746
rect 8022 1721 8031 1741
rect 8051 1721 8060 1741
rect 8022 1712 8060 1721
rect 8089 1737 8174 1745
rect 8089 1717 8146 1737
rect 8166 1717 8174 1737
rect 8022 1711 8059 1712
rect 8089 1711 8174 1717
rect 8240 1741 8278 1749
rect 8240 1721 8249 1741
rect 8269 1721 8278 1741
rect 8240 1712 8278 1721
rect 8422 1746 8464 1755
rect 8422 1728 8436 1746
rect 8454 1728 8464 1746
rect 8422 1720 8464 1728
rect 8427 1718 8464 1720
rect 8867 1739 9310 1778
rect 8240 1711 8277 1712
rect 7701 1683 7791 1689
rect 7701 1663 7717 1683
rect 7737 1681 7791 1683
rect 7737 1663 7762 1681
rect 7701 1661 7762 1663
rect 7782 1661 7791 1681
rect 7701 1655 7791 1661
rect 7714 1601 7751 1602
rect 7810 1601 7847 1602
rect 7866 1601 7902 1711
rect 8089 1690 8120 1711
rect 8867 1696 8914 1739
rect 9270 1734 9310 1739
rect 9935 1737 10122 1761
rect 10153 1742 10546 1762
rect 10566 1742 10569 1762
rect 10153 1737 10569 1742
rect 8085 1689 8120 1690
rect 7963 1679 8120 1689
rect 7963 1659 7980 1679
rect 8000 1659 8120 1679
rect 7963 1652 8120 1659
rect 8187 1682 8336 1690
rect 8187 1662 8198 1682
rect 8218 1662 8257 1682
rect 8277 1662 8336 1682
rect 8867 1678 8877 1696
rect 8895 1678 8914 1696
rect 8867 1674 8914 1678
rect 8868 1669 8905 1674
rect 8187 1655 8336 1662
rect 9935 1666 9972 1737
rect 10153 1736 10494 1737
rect 10087 1676 10118 1677
rect 8187 1654 8228 1655
rect 8424 1653 8461 1656
rect 7921 1601 7958 1602
rect 7614 1592 7752 1601
rect 6818 1553 7262 1579
rect 6818 1551 6986 1553
rect 5771 1419 6218 1431
rect 5814 1417 5847 1419
rect 5181 1399 5319 1408
rect 4975 1398 5012 1399
rect 4705 1345 4746 1346
rect 4479 1324 4531 1342
rect 4597 1338 4746 1345
rect 4047 1304 4087 1314
rect 4597 1318 4656 1338
rect 4676 1318 4715 1338
rect 4735 1318 4746 1338
rect 4597 1310 4746 1318
rect 4813 1341 4970 1348
rect 4813 1321 4933 1341
rect 4953 1321 4970 1341
rect 4813 1311 4970 1321
rect 4813 1310 4848 1311
rect 3877 1287 3915 1296
rect 4813 1289 4844 1310
rect 5031 1289 5067 1399
rect 5086 1398 5123 1399
rect 5182 1398 5219 1399
rect 5142 1339 5232 1345
rect 5142 1319 5151 1339
rect 5171 1337 5232 1339
rect 5171 1319 5196 1337
rect 5142 1317 5196 1319
rect 5216 1317 5232 1337
rect 5142 1311 5232 1317
rect 4656 1288 4693 1289
rect 3877 1286 3914 1287
rect 3338 1258 3428 1264
rect 3338 1238 3354 1258
rect 3374 1256 3428 1258
rect 3374 1238 3399 1256
rect 3338 1236 3399 1238
rect 3419 1236 3428 1256
rect 3338 1230 3428 1236
rect 3351 1176 3388 1177
rect 3447 1176 3484 1177
rect 3503 1176 3539 1286
rect 3726 1265 3757 1286
rect 4655 1279 4693 1288
rect 3722 1264 3757 1265
rect 3600 1254 3757 1264
rect 3600 1234 3617 1254
rect 3637 1234 3757 1254
rect 3600 1227 3757 1234
rect 3824 1257 3973 1265
rect 3824 1237 3835 1257
rect 3855 1237 3894 1257
rect 3914 1237 3973 1257
rect 4483 1261 4523 1271
rect 3824 1230 3973 1237
rect 4039 1233 4091 1251
rect 3824 1229 3865 1230
rect 3558 1176 3595 1177
rect 3251 1167 3389 1176
rect 3251 1147 3360 1167
rect 3380 1147 3389 1167
rect 3251 1140 3389 1147
rect 3447 1167 3595 1176
rect 3447 1147 3456 1167
rect 3476 1147 3566 1167
rect 3586 1147 3595 1167
rect 3251 1138 3347 1140
rect 3447 1137 3595 1147
rect 3654 1167 3691 1177
rect 3654 1147 3662 1167
rect 3682 1147 3691 1167
rect 3503 1136 3539 1137
rect 3654 1080 3691 1147
rect 3726 1176 3757 1227
rect 4039 1215 4057 1233
rect 4075 1215 4091 1233
rect 3776 1176 3813 1177
rect 3726 1167 3813 1176
rect 3726 1147 3784 1167
rect 3804 1147 3813 1167
rect 3726 1137 3813 1147
rect 3872 1167 3909 1177
rect 3872 1147 3880 1167
rect 3900 1147 3909 1167
rect 3726 1136 3757 1137
rect 3351 1077 3388 1078
rect 3654 1077 3693 1080
rect 3350 1076 3693 1077
rect 3872 1076 3909 1147
rect 3275 1071 3693 1076
rect 3275 1051 3278 1071
rect 3298 1051 3693 1071
rect 3722 1052 3909 1076
rect 1816 1020 1853 1028
rect 1816 1001 1824 1020
rect 1845 1001 1853 1020
rect 1816 995 1853 1001
rect 3654 1026 3693 1051
rect 4039 1026 4091 1215
rect 4483 1243 4493 1261
rect 4511 1243 4523 1261
rect 4655 1259 4664 1279
rect 4684 1259 4693 1279
rect 4655 1251 4693 1259
rect 4759 1283 4844 1289
rect 4874 1288 4911 1289
rect 4759 1263 4767 1283
rect 4787 1263 4844 1283
rect 4759 1255 4844 1263
rect 4873 1279 4911 1288
rect 4873 1259 4882 1279
rect 4902 1259 4911 1279
rect 4759 1254 4795 1255
rect 4873 1251 4911 1259
rect 4977 1283 5121 1289
rect 4977 1263 4985 1283
rect 5005 1263 5038 1283
rect 5058 1263 5093 1283
rect 5113 1263 5121 1283
rect 4977 1255 5121 1263
rect 4977 1254 5013 1255
rect 5085 1254 5121 1255
rect 5187 1288 5224 1289
rect 5187 1287 5225 1288
rect 5187 1279 5251 1287
rect 5187 1259 5196 1279
rect 5216 1265 5251 1279
rect 5271 1265 5274 1285
rect 5216 1260 5274 1265
rect 5216 1259 5251 1260
rect 4483 1187 4523 1243
rect 4656 1222 4693 1251
rect 4657 1220 4693 1222
rect 4657 1198 4848 1220
rect 4874 1219 4911 1251
rect 5187 1247 5251 1259
rect 5291 1221 5318 1399
rect 6176 1374 6218 1419
rect 5150 1219 5318 1221
rect 4874 1209 5318 1219
rect 5459 1315 5646 1339
rect 5677 1320 6070 1340
rect 6090 1320 6093 1340
rect 5677 1315 6093 1320
rect 5459 1244 5496 1315
rect 5677 1314 6018 1315
rect 5611 1254 5642 1255
rect 5459 1224 5468 1244
rect 5488 1224 5496 1244
rect 5459 1214 5496 1224
rect 5555 1244 5642 1254
rect 5555 1224 5564 1244
rect 5584 1224 5642 1244
rect 5555 1215 5642 1224
rect 5555 1214 5592 1215
rect 4480 1182 4523 1187
rect 4871 1193 5318 1209
rect 4871 1187 4899 1193
rect 5150 1192 5318 1193
rect 4480 1179 4630 1182
rect 4871 1179 4898 1187
rect 4480 1177 4898 1179
rect 4480 1159 4489 1177
rect 4507 1159 4898 1177
rect 5611 1164 5642 1215
rect 5677 1244 5714 1314
rect 5980 1313 6017 1314
rect 5829 1254 5865 1255
rect 5677 1224 5686 1244
rect 5706 1224 5714 1244
rect 5677 1214 5714 1224
rect 5773 1244 5921 1254
rect 6021 1251 6117 1253
rect 5773 1224 5782 1244
rect 5802 1224 5892 1244
rect 5912 1224 5921 1244
rect 5773 1215 5921 1224
rect 5979 1244 6117 1251
rect 5979 1224 5988 1244
rect 6008 1224 6117 1244
rect 5979 1215 6117 1224
rect 5773 1214 5810 1215
rect 5503 1161 5544 1162
rect 4480 1156 4898 1159
rect 4480 1150 4523 1156
rect 4483 1147 4523 1150
rect 5398 1154 5544 1161
rect 4880 1138 4920 1139
rect 4591 1121 4920 1138
rect 5398 1134 5454 1154
rect 5474 1134 5513 1154
rect 5533 1134 5544 1154
rect 5398 1126 5544 1134
rect 5611 1157 5768 1164
rect 5611 1137 5731 1157
rect 5751 1137 5768 1157
rect 5611 1127 5768 1137
rect 5611 1126 5646 1127
rect 4475 1078 4518 1089
rect 4475 1060 4487 1078
rect 4505 1060 4518 1078
rect 4475 1034 4518 1060
rect 4591 1034 4618 1121
rect 4880 1112 4920 1121
rect 3654 1008 4093 1026
rect 3654 990 4054 1008
rect 4072 990 4093 1008
rect 3654 984 4093 990
rect 3660 980 4093 984
rect 4475 1013 4618 1034
rect 4662 1086 4696 1102
rect 4880 1092 5273 1112
rect 5293 1092 5296 1112
rect 5611 1105 5642 1126
rect 5829 1105 5865 1215
rect 5884 1214 5921 1215
rect 5980 1214 6017 1215
rect 5940 1155 6030 1161
rect 5940 1135 5949 1155
rect 5969 1153 6030 1155
rect 5969 1135 5994 1153
rect 5940 1133 5994 1135
rect 6014 1133 6030 1153
rect 5940 1127 6030 1133
rect 5454 1104 5491 1105
rect 4880 1087 5296 1092
rect 5453 1095 5491 1104
rect 4880 1086 5221 1087
rect 4662 1016 4699 1086
rect 4814 1026 4845 1027
rect 4475 1011 4612 1013
rect 4039 978 4091 980
rect 4475 969 4518 1011
rect 4662 996 4671 1016
rect 4691 996 4699 1016
rect 4662 986 4699 996
rect 4758 1016 4845 1026
rect 4758 996 4767 1016
rect 4787 996 4845 1016
rect 4758 987 4845 996
rect 4758 986 4795 987
rect 4473 959 4518 969
rect 4473 941 4482 959
rect 4500 941 4518 959
rect 4473 935 4518 941
rect 4814 936 4845 987
rect 4880 1016 4917 1086
rect 5183 1085 5220 1086
rect 5453 1075 5462 1095
rect 5482 1075 5491 1095
rect 5453 1067 5491 1075
rect 5557 1099 5642 1105
rect 5672 1104 5709 1105
rect 5557 1079 5565 1099
rect 5585 1079 5642 1099
rect 5557 1071 5642 1079
rect 5671 1095 5709 1104
rect 5671 1075 5680 1095
rect 5700 1075 5709 1095
rect 5557 1070 5593 1071
rect 5671 1067 5709 1075
rect 5775 1099 5919 1105
rect 5775 1079 5783 1099
rect 5803 1096 5891 1099
rect 5803 1079 5838 1096
rect 5775 1078 5838 1079
rect 5857 1079 5891 1096
rect 5911 1079 5919 1099
rect 5857 1078 5919 1079
rect 5775 1071 5919 1078
rect 5775 1070 5811 1071
rect 5883 1070 5919 1071
rect 5985 1104 6022 1105
rect 5985 1103 6023 1104
rect 6045 1103 6072 1107
rect 5985 1101 6072 1103
rect 5985 1095 6049 1101
rect 5985 1075 5994 1095
rect 6014 1081 6049 1095
rect 6069 1081 6072 1101
rect 6014 1076 6072 1081
rect 6014 1075 6049 1076
rect 5454 1038 5491 1067
rect 5455 1036 5491 1038
rect 5032 1026 5068 1027
rect 4880 996 4889 1016
rect 4909 996 4917 1016
rect 4880 986 4917 996
rect 4976 1016 5124 1026
rect 5224 1023 5320 1025
rect 4976 996 4985 1016
rect 5005 996 5095 1016
rect 5115 996 5124 1016
rect 4976 987 5124 996
rect 5182 1016 5320 1023
rect 5182 996 5191 1016
rect 5211 996 5320 1016
rect 5455 1014 5646 1036
rect 5672 1035 5709 1067
rect 5985 1063 6049 1075
rect 6089 1037 6116 1215
rect 5948 1035 6116 1037
rect 5672 1009 6116 1035
rect 5182 987 5320 996
rect 4976 986 5013 987
rect 4473 932 4510 935
rect 4706 933 4747 934
rect 4598 926 4747 933
rect 4042 913 4079 918
rect 4033 909 4080 913
rect 4033 891 4052 909
rect 4070 891 4080 909
rect 4598 906 4657 926
rect 4677 906 4716 926
rect 4736 906 4747 926
rect 4598 898 4747 906
rect 4814 929 4971 936
rect 4814 909 4934 929
rect 4954 909 4971 929
rect 4814 899 4971 909
rect 4814 898 4849 899
rect 4033 828 4080 891
rect 4814 877 4845 898
rect 5032 877 5068 987
rect 5087 986 5124 987
rect 5183 986 5220 987
rect 5143 927 5233 933
rect 5143 907 5152 927
rect 5172 925 5233 927
rect 5172 907 5197 925
rect 5143 905 5197 907
rect 5217 905 5233 925
rect 5143 899 5233 905
rect 4657 876 4694 877
rect 4470 868 4507 870
rect 4470 860 4512 868
rect 4470 842 4480 860
rect 4498 842 4512 860
rect 4470 833 4512 842
rect 4656 867 4694 876
rect 4656 847 4665 867
rect 4685 847 4694 867
rect 4656 839 4694 847
rect 4760 871 4845 877
rect 4875 876 4912 877
rect 4760 851 4768 871
rect 4788 851 4845 871
rect 4760 843 4845 851
rect 4874 867 4912 876
rect 4874 847 4883 867
rect 4903 847 4912 867
rect 4760 842 4796 843
rect 4874 839 4912 847
rect 4978 875 5122 877
rect 4978 871 5030 875
rect 4978 851 4986 871
rect 5006 855 5030 871
rect 5050 871 5122 875
rect 5050 855 5094 871
rect 5006 851 5094 855
rect 5114 851 5122 871
rect 4978 843 5122 851
rect 4978 842 5014 843
rect 5086 842 5122 843
rect 5188 876 5225 877
rect 5188 875 5226 876
rect 5188 867 5252 875
rect 5188 847 5197 867
rect 5217 853 5252 867
rect 5272 853 5275 873
rect 5217 848 5275 853
rect 5217 847 5252 848
rect 4033 813 4083 828
rect 4033 788 4047 813
rect 4079 788 4083 813
rect 4471 808 4512 833
rect 4657 808 4694 839
rect 4875 817 4912 839
rect 5188 835 5252 847
rect 4870 808 4912 817
rect 5292 809 5319 987
rect 4471 796 4516 808
rect 4033 775 4080 788
rect 1418 750 1426 772
rect 1450 750 1458 772
rect 1418 742 1458 750
rect 4467 738 4516 796
rect 4657 782 4719 808
rect 4870 807 4955 808
rect 5151 807 5319 809
rect 4870 781 5319 807
rect 4870 738 4909 781
rect 5151 780 5319 781
rect 5782 785 5822 1009
rect 5948 1008 6116 1009
rect 6180 1041 6213 1374
rect 6818 1373 6845 1551
rect 6885 1513 6949 1525
rect 7225 1521 7262 1553
rect 7288 1552 7479 1574
rect 7614 1572 7723 1592
rect 7743 1572 7752 1592
rect 7614 1565 7752 1572
rect 7810 1592 7958 1601
rect 7810 1572 7819 1592
rect 7839 1572 7929 1592
rect 7949 1572 7958 1592
rect 7614 1563 7710 1565
rect 7810 1562 7958 1572
rect 8017 1592 8054 1602
rect 8017 1572 8025 1592
rect 8045 1572 8054 1592
rect 7866 1561 7902 1562
rect 7443 1550 7479 1552
rect 7443 1521 7480 1550
rect 6885 1512 6920 1513
rect 6862 1507 6920 1512
rect 6862 1487 6865 1507
rect 6885 1493 6920 1507
rect 6940 1493 6949 1513
rect 6885 1485 6949 1493
rect 6911 1484 6949 1485
rect 6912 1483 6949 1484
rect 7015 1517 7051 1518
rect 7123 1517 7159 1518
rect 7015 1509 7159 1517
rect 7015 1489 7023 1509
rect 7043 1508 7131 1509
rect 7043 1489 7078 1508
rect 7099 1489 7131 1508
rect 7151 1489 7159 1509
rect 7015 1483 7159 1489
rect 7225 1513 7263 1521
rect 7341 1517 7377 1518
rect 7225 1493 7234 1513
rect 7254 1493 7263 1513
rect 7225 1484 7263 1493
rect 7292 1509 7377 1517
rect 7292 1489 7349 1509
rect 7369 1489 7377 1509
rect 7225 1483 7262 1484
rect 7292 1483 7377 1489
rect 7443 1513 7481 1521
rect 7443 1493 7452 1513
rect 7472 1493 7481 1513
rect 7714 1502 7751 1503
rect 8017 1502 8054 1572
rect 8089 1601 8120 1652
rect 8416 1647 8461 1653
rect 8416 1629 8434 1647
rect 8452 1629 8461 1647
rect 9935 1646 9944 1666
rect 9964 1646 9972 1666
rect 9935 1636 9972 1646
rect 10031 1666 10118 1676
rect 10031 1646 10040 1666
rect 10060 1646 10118 1666
rect 10031 1637 10118 1646
rect 10031 1636 10068 1637
rect 8416 1619 8461 1629
rect 8139 1601 8176 1602
rect 8089 1592 8176 1601
rect 8089 1572 8147 1592
rect 8167 1572 8176 1592
rect 8089 1562 8176 1572
rect 8235 1592 8272 1602
rect 8235 1572 8243 1592
rect 8263 1572 8272 1592
rect 8416 1577 8459 1619
rect 8856 1607 8908 1609
rect 8322 1575 8459 1577
rect 8089 1561 8120 1562
rect 8235 1502 8272 1572
rect 7713 1501 8054 1502
rect 7443 1484 7481 1493
rect 7638 1496 8054 1501
rect 7443 1483 7480 1484
rect 6904 1455 6994 1461
rect 6904 1435 6920 1455
rect 6940 1453 6994 1455
rect 6940 1435 6965 1453
rect 6904 1433 6965 1435
rect 6985 1433 6994 1453
rect 6904 1427 6994 1433
rect 6917 1373 6954 1374
rect 7013 1373 7050 1374
rect 7069 1373 7105 1483
rect 7292 1462 7323 1483
rect 7638 1476 7641 1496
rect 7661 1476 8054 1496
rect 8238 1486 8272 1502
rect 8316 1554 8459 1575
rect 8854 1603 9287 1607
rect 8854 1597 9293 1603
rect 8854 1579 8875 1597
rect 8893 1579 9293 1597
rect 10087 1586 10118 1637
rect 10153 1666 10190 1736
rect 10456 1735 10493 1736
rect 10305 1676 10341 1677
rect 10153 1646 10162 1666
rect 10182 1646 10190 1666
rect 10153 1636 10190 1646
rect 10249 1666 10397 1676
rect 10497 1673 10593 1675
rect 10249 1646 10258 1666
rect 10278 1646 10368 1666
rect 10388 1646 10397 1666
rect 10249 1637 10397 1646
rect 10455 1666 10593 1673
rect 10455 1646 10464 1666
rect 10484 1646 10593 1666
rect 10455 1637 10593 1646
rect 10249 1636 10286 1637
rect 9979 1583 10020 1584
rect 8854 1561 9293 1579
rect 8014 1467 8054 1476
rect 8316 1467 8343 1554
rect 8416 1528 8459 1554
rect 8416 1510 8429 1528
rect 8447 1510 8459 1528
rect 8416 1499 8459 1510
rect 7288 1461 7323 1462
rect 7166 1451 7323 1461
rect 7166 1431 7183 1451
rect 7203 1431 7323 1451
rect 7166 1424 7323 1431
rect 7390 1454 7539 1462
rect 7390 1434 7401 1454
rect 7421 1434 7460 1454
rect 7480 1434 7539 1454
rect 8014 1450 8343 1467
rect 8014 1449 8054 1450
rect 7390 1427 7539 1434
rect 8411 1438 8451 1441
rect 8411 1432 8454 1438
rect 8036 1429 8454 1432
rect 7390 1426 7431 1427
rect 7124 1373 7161 1374
rect 6817 1364 6955 1373
rect 6817 1344 6926 1364
rect 6946 1344 6955 1364
rect 6817 1337 6955 1344
rect 7013 1364 7161 1373
rect 7013 1344 7022 1364
rect 7042 1344 7132 1364
rect 7152 1344 7161 1364
rect 6817 1335 6913 1337
rect 7013 1334 7161 1344
rect 7220 1364 7257 1374
rect 7220 1344 7228 1364
rect 7248 1344 7257 1364
rect 7069 1333 7105 1334
rect 6917 1274 6954 1275
rect 7220 1274 7257 1344
rect 7292 1373 7323 1424
rect 8036 1411 8427 1429
rect 8445 1411 8454 1429
rect 8036 1409 8454 1411
rect 8036 1401 8063 1409
rect 8304 1406 8454 1409
rect 7616 1395 7784 1396
rect 8035 1395 8063 1401
rect 7616 1379 8063 1395
rect 8411 1401 8454 1406
rect 7342 1373 7379 1374
rect 7292 1364 7379 1373
rect 7292 1344 7350 1364
rect 7370 1344 7379 1364
rect 7292 1334 7379 1344
rect 7438 1364 7475 1374
rect 7438 1344 7446 1364
rect 7466 1344 7475 1364
rect 7292 1333 7323 1334
rect 6916 1273 7257 1274
rect 7438 1273 7475 1344
rect 6841 1268 7257 1273
rect 6841 1248 6844 1268
rect 6864 1248 7257 1268
rect 7288 1249 7475 1273
rect 7616 1369 8060 1379
rect 7616 1367 7784 1369
rect 7616 1189 7643 1367
rect 7683 1329 7747 1341
rect 8023 1337 8060 1369
rect 8086 1368 8277 1390
rect 8241 1366 8277 1368
rect 8241 1337 8278 1366
rect 8411 1345 8451 1401
rect 7683 1328 7718 1329
rect 7660 1323 7718 1328
rect 7660 1303 7663 1323
rect 7683 1309 7718 1323
rect 7738 1309 7747 1329
rect 7683 1301 7747 1309
rect 7709 1300 7747 1301
rect 7710 1299 7747 1300
rect 7813 1333 7849 1334
rect 7921 1333 7957 1334
rect 7813 1325 7957 1333
rect 7813 1305 7821 1325
rect 7841 1305 7876 1325
rect 7896 1305 7929 1325
rect 7949 1305 7957 1325
rect 7813 1299 7957 1305
rect 8023 1329 8061 1337
rect 8139 1333 8175 1334
rect 8023 1309 8032 1329
rect 8052 1309 8061 1329
rect 8023 1300 8061 1309
rect 8090 1325 8175 1333
rect 8090 1305 8147 1325
rect 8167 1305 8175 1325
rect 8023 1299 8060 1300
rect 8090 1299 8175 1305
rect 8241 1329 8279 1337
rect 8241 1309 8250 1329
rect 8270 1309 8279 1329
rect 8411 1327 8423 1345
rect 8441 1327 8451 1345
rect 8856 1372 8908 1561
rect 9254 1536 9293 1561
rect 9871 1576 10020 1583
rect 9871 1556 9930 1576
rect 9950 1556 9989 1576
rect 10009 1556 10020 1576
rect 9871 1548 10020 1556
rect 10087 1579 10244 1586
rect 10087 1559 10207 1579
rect 10227 1559 10244 1579
rect 10087 1549 10244 1559
rect 10087 1548 10122 1549
rect 9038 1511 9225 1535
rect 9254 1516 9649 1536
rect 9669 1516 9672 1536
rect 10087 1527 10118 1548
rect 10305 1527 10341 1637
rect 10360 1636 10397 1637
rect 10456 1636 10493 1637
rect 10416 1577 10506 1583
rect 10416 1557 10425 1577
rect 10445 1575 10506 1577
rect 10445 1557 10470 1575
rect 10416 1555 10470 1557
rect 10490 1555 10506 1575
rect 10416 1549 10506 1555
rect 9930 1526 9967 1527
rect 9254 1511 9672 1516
rect 9929 1517 9967 1526
rect 9038 1440 9075 1511
rect 9254 1510 9597 1511
rect 9254 1507 9293 1510
rect 9559 1509 9596 1510
rect 9190 1450 9221 1451
rect 9038 1420 9047 1440
rect 9067 1420 9075 1440
rect 9038 1410 9075 1420
rect 9134 1440 9221 1450
rect 9134 1420 9143 1440
rect 9163 1420 9221 1440
rect 9134 1411 9221 1420
rect 9134 1410 9171 1411
rect 8856 1354 8872 1372
rect 8890 1354 8908 1372
rect 9190 1360 9221 1411
rect 9256 1440 9293 1507
rect 9929 1497 9938 1517
rect 9958 1497 9967 1517
rect 9929 1489 9967 1497
rect 10033 1521 10118 1527
rect 10148 1526 10185 1527
rect 10033 1501 10041 1521
rect 10061 1501 10118 1521
rect 10033 1493 10118 1501
rect 10147 1517 10185 1526
rect 10147 1497 10156 1517
rect 10176 1497 10185 1517
rect 10033 1492 10069 1493
rect 10147 1489 10185 1497
rect 10251 1521 10395 1527
rect 10251 1501 10259 1521
rect 10279 1516 10367 1521
rect 10279 1501 10315 1516
rect 10251 1499 10315 1501
rect 10334 1501 10367 1516
rect 10387 1501 10395 1521
rect 10334 1499 10395 1501
rect 10251 1493 10395 1499
rect 10251 1492 10287 1493
rect 10359 1492 10395 1493
rect 10461 1526 10498 1527
rect 10461 1525 10499 1526
rect 10461 1517 10525 1525
rect 10461 1497 10470 1517
rect 10490 1503 10525 1517
rect 10545 1503 10548 1523
rect 10490 1498 10548 1503
rect 10490 1497 10525 1498
rect 9930 1460 9967 1489
rect 9931 1458 9967 1460
rect 9408 1450 9444 1451
rect 9256 1420 9265 1440
rect 9285 1420 9293 1440
rect 9256 1410 9293 1420
rect 9352 1440 9500 1450
rect 9600 1447 9696 1449
rect 9352 1420 9361 1440
rect 9381 1420 9471 1440
rect 9491 1420 9500 1440
rect 9352 1411 9500 1420
rect 9558 1440 9696 1447
rect 9558 1420 9567 1440
rect 9587 1420 9696 1440
rect 9931 1436 10122 1458
rect 10148 1457 10185 1489
rect 10461 1485 10525 1497
rect 10565 1459 10592 1637
rect 10424 1457 10592 1459
rect 10148 1443 10592 1457
rect 11195 1591 11363 1592
rect 11489 1591 11529 1815
rect 11992 1819 12160 1820
rect 12395 1819 12435 1852
rect 12791 1819 12838 1852
rect 13229 1851 13270 1876
rect 13415 1851 13452 1882
rect 13633 1851 13670 1882
rect 13946 1878 14010 1890
rect 14050 1852 14077 2030
rect 13229 1824 13278 1851
rect 13414 1825 13463 1851
rect 13632 1850 13713 1851
rect 13909 1850 14077 1852
rect 13632 1825 14077 1850
rect 13633 1824 14077 1825
rect 11992 1818 12436 1819
rect 11992 1793 12437 1818
rect 11992 1791 12160 1793
rect 12356 1792 12437 1793
rect 12606 1792 12655 1818
rect 12791 1792 12840 1819
rect 11992 1613 12019 1791
rect 12059 1753 12123 1765
rect 12399 1761 12436 1792
rect 12617 1761 12654 1792
rect 12799 1767 12840 1792
rect 13231 1791 13278 1824
rect 13634 1791 13674 1824
rect 13909 1823 14077 1824
rect 14540 1828 14580 2052
rect 14706 2051 14874 2052
rect 15477 2186 15921 2200
rect 15477 2184 15645 2186
rect 15477 2006 15504 2184
rect 15544 2146 15608 2158
rect 15884 2154 15921 2186
rect 15947 2185 16138 2207
rect 16373 2203 16482 2223
rect 16502 2203 16511 2223
rect 16373 2196 16511 2203
rect 16569 2223 16717 2232
rect 16569 2203 16578 2223
rect 16598 2203 16688 2223
rect 16708 2203 16717 2223
rect 16373 2194 16469 2196
rect 16569 2193 16717 2203
rect 16776 2223 16813 2233
rect 16776 2203 16784 2223
rect 16804 2203 16813 2223
rect 16625 2192 16661 2193
rect 16102 2183 16138 2185
rect 16102 2154 16139 2183
rect 15544 2145 15579 2146
rect 15521 2140 15579 2145
rect 15521 2120 15524 2140
rect 15544 2126 15579 2140
rect 15599 2126 15608 2146
rect 15544 2118 15608 2126
rect 15570 2117 15608 2118
rect 15571 2116 15608 2117
rect 15674 2150 15710 2151
rect 15782 2150 15818 2151
rect 15674 2142 15818 2150
rect 15674 2122 15682 2142
rect 15702 2140 15790 2142
rect 15702 2122 15735 2140
rect 15674 2121 15735 2122
rect 15756 2122 15790 2140
rect 15810 2122 15818 2142
rect 15756 2121 15818 2122
rect 15674 2116 15818 2121
rect 15884 2146 15922 2154
rect 16000 2150 16036 2151
rect 15884 2126 15893 2146
rect 15913 2126 15922 2146
rect 15884 2117 15922 2126
rect 15951 2142 16036 2150
rect 15951 2122 16008 2142
rect 16028 2122 16036 2142
rect 15884 2116 15921 2117
rect 15951 2116 16036 2122
rect 16102 2146 16140 2154
rect 16102 2126 16111 2146
rect 16131 2126 16140 2146
rect 16776 2136 16813 2203
rect 16848 2232 16879 2283
rect 17161 2271 17179 2289
rect 17197 2271 17213 2289
rect 17679 2296 17717 2305
rect 16898 2232 16935 2233
rect 16848 2223 16935 2232
rect 16848 2203 16906 2223
rect 16926 2203 16935 2223
rect 16848 2193 16935 2203
rect 16994 2223 17031 2233
rect 16994 2203 17002 2223
rect 17022 2203 17031 2223
rect 16848 2192 16879 2193
rect 16473 2133 16510 2134
rect 16776 2133 16815 2136
rect 16472 2132 16815 2133
rect 16994 2132 17031 2203
rect 16102 2117 16140 2126
rect 16397 2127 16815 2132
rect 16102 2116 16139 2117
rect 15563 2088 15653 2094
rect 15563 2068 15579 2088
rect 15599 2086 15653 2088
rect 15599 2068 15624 2086
rect 15563 2066 15624 2068
rect 15644 2066 15653 2086
rect 15563 2060 15653 2066
rect 15576 2006 15613 2007
rect 15672 2006 15709 2007
rect 15728 2006 15764 2116
rect 15951 2095 15982 2116
rect 16397 2107 16400 2127
rect 16420 2107 16815 2127
rect 16844 2108 17031 2132
rect 15947 2094 15982 2095
rect 15825 2084 15982 2094
rect 15825 2064 15842 2084
rect 15862 2064 15982 2084
rect 15825 2057 15982 2064
rect 16049 2087 16198 2095
rect 16049 2067 16060 2087
rect 16080 2067 16119 2087
rect 16139 2067 16198 2087
rect 16049 2060 16198 2067
rect 16776 2082 16815 2107
rect 17161 2082 17213 2271
rect 17507 2278 17547 2288
rect 17507 2260 17517 2278
rect 17535 2260 17547 2278
rect 17679 2276 17688 2296
rect 17708 2276 17717 2296
rect 17679 2268 17717 2276
rect 17783 2300 17868 2306
rect 17898 2305 17935 2306
rect 17783 2280 17791 2300
rect 17811 2280 17868 2300
rect 17783 2272 17868 2280
rect 17897 2296 17935 2305
rect 17897 2276 17906 2296
rect 17926 2276 17935 2296
rect 17783 2271 17819 2272
rect 17897 2268 17935 2276
rect 18001 2300 18145 2306
rect 18001 2280 18009 2300
rect 18029 2280 18062 2300
rect 18082 2280 18117 2300
rect 18137 2280 18145 2300
rect 18001 2272 18145 2280
rect 18001 2271 18037 2272
rect 18109 2271 18145 2272
rect 18211 2305 18248 2306
rect 18211 2304 18249 2305
rect 18211 2296 18275 2304
rect 18211 2276 18220 2296
rect 18240 2282 18275 2296
rect 18295 2282 18298 2302
rect 18240 2277 18298 2282
rect 18240 2276 18275 2277
rect 17507 2204 17547 2260
rect 17680 2239 17717 2268
rect 17681 2237 17717 2239
rect 17681 2215 17872 2237
rect 17898 2236 17935 2268
rect 18211 2264 18275 2276
rect 18315 2238 18342 2416
rect 18174 2236 18342 2238
rect 17898 2226 18342 2236
rect 18483 2332 18670 2356
rect 18701 2337 19094 2357
rect 19114 2337 19117 2357
rect 18701 2332 19117 2337
rect 18483 2261 18520 2332
rect 18701 2331 19042 2332
rect 18635 2271 18666 2272
rect 18483 2241 18492 2261
rect 18512 2241 18520 2261
rect 18483 2231 18520 2241
rect 18579 2261 18666 2271
rect 18579 2241 18588 2261
rect 18608 2241 18666 2261
rect 18579 2232 18666 2241
rect 18579 2231 18616 2232
rect 17504 2199 17547 2204
rect 17895 2210 18342 2226
rect 17895 2204 17923 2210
rect 18174 2209 18342 2210
rect 17504 2196 17654 2199
rect 17895 2196 17922 2204
rect 17504 2194 17922 2196
rect 17504 2176 17513 2194
rect 17531 2176 17922 2194
rect 18635 2181 18666 2232
rect 18701 2261 18738 2331
rect 19004 2330 19041 2331
rect 19242 2273 19275 2432
rect 18853 2271 18889 2272
rect 18701 2241 18710 2261
rect 18730 2241 18738 2261
rect 18701 2231 18738 2241
rect 18797 2261 18945 2271
rect 19045 2268 19141 2270
rect 18797 2241 18806 2261
rect 18826 2241 18916 2261
rect 18936 2241 18945 2261
rect 18797 2232 18945 2241
rect 19003 2261 19141 2268
rect 19003 2241 19012 2261
rect 19032 2241 19141 2261
rect 19242 2269 19278 2273
rect 19242 2251 19251 2269
rect 19273 2251 19278 2269
rect 19242 2245 19278 2251
rect 19003 2232 19141 2241
rect 18797 2231 18834 2232
rect 18527 2178 18568 2179
rect 17504 2173 17922 2176
rect 17504 2167 17547 2173
rect 17507 2164 17547 2167
rect 18419 2171 18568 2178
rect 17904 2155 17944 2156
rect 17615 2138 17944 2155
rect 18419 2151 18478 2171
rect 18498 2151 18537 2171
rect 18557 2151 18568 2171
rect 18419 2143 18568 2151
rect 18635 2174 18792 2181
rect 18635 2154 18755 2174
rect 18775 2154 18792 2174
rect 18635 2144 18792 2154
rect 18635 2143 18670 2144
rect 17499 2095 17542 2106
rect 16776 2064 17215 2082
rect 16049 2059 16090 2060
rect 15783 2006 15820 2007
rect 15476 1997 15614 2006
rect 15476 1977 15585 1997
rect 15605 1977 15614 1997
rect 15476 1970 15614 1977
rect 15672 1997 15820 2006
rect 15672 1977 15681 1997
rect 15701 1977 15791 1997
rect 15811 1977 15820 1997
rect 15476 1968 15572 1970
rect 15672 1967 15820 1977
rect 15879 1997 15916 2007
rect 15879 1977 15887 1997
rect 15907 1977 15916 1997
rect 15728 1966 15764 1967
rect 15576 1907 15613 1908
rect 15879 1907 15916 1977
rect 15951 2006 15982 2057
rect 16776 2046 17176 2064
rect 17194 2046 17215 2064
rect 16776 2040 17215 2046
rect 16782 2036 17215 2040
rect 17499 2077 17511 2095
rect 17529 2077 17542 2095
rect 17499 2051 17542 2077
rect 17615 2051 17642 2138
rect 17904 2129 17944 2138
rect 17161 2034 17213 2036
rect 17499 2030 17642 2051
rect 17686 2103 17720 2119
rect 17904 2109 18297 2129
rect 18317 2109 18320 2129
rect 18635 2122 18666 2143
rect 18853 2122 18889 2232
rect 18908 2231 18945 2232
rect 19004 2231 19041 2232
rect 18964 2172 19054 2178
rect 18964 2152 18973 2172
rect 18993 2170 19054 2172
rect 18993 2152 19018 2170
rect 18964 2150 19018 2152
rect 19038 2150 19054 2170
rect 18964 2144 19054 2150
rect 18478 2121 18515 2122
rect 17904 2104 18320 2109
rect 18477 2112 18515 2121
rect 17904 2103 18245 2104
rect 17686 2033 17723 2103
rect 17838 2043 17869 2044
rect 17499 2028 17636 2030
rect 16001 2006 16038 2007
rect 15951 1997 16038 2006
rect 15951 1977 16009 1997
rect 16029 1977 16038 1997
rect 15951 1967 16038 1977
rect 16097 1997 16134 2007
rect 16097 1977 16105 1997
rect 16125 1977 16134 1997
rect 17499 1986 17542 2028
rect 17686 2013 17695 2033
rect 17715 2013 17723 2033
rect 17686 2003 17723 2013
rect 17782 2033 17869 2043
rect 17782 2013 17791 2033
rect 17811 2013 17869 2033
rect 17782 2004 17869 2013
rect 17782 2003 17819 2004
rect 15951 1966 15982 1967
rect 15575 1906 15916 1907
rect 16097 1906 16134 1977
rect 17497 1976 17542 1986
rect 17164 1969 17201 1974
rect 17155 1965 17202 1969
rect 17155 1947 17174 1965
rect 17192 1947 17202 1965
rect 17497 1958 17506 1976
rect 17524 1958 17542 1976
rect 17497 1952 17542 1958
rect 17838 1953 17869 2004
rect 17904 2033 17941 2103
rect 18207 2102 18244 2103
rect 18477 2092 18486 2112
rect 18506 2092 18515 2112
rect 18477 2084 18515 2092
rect 18581 2116 18666 2122
rect 18696 2121 18733 2122
rect 18581 2096 18589 2116
rect 18609 2096 18666 2116
rect 18581 2088 18666 2096
rect 18695 2112 18733 2121
rect 18695 2092 18704 2112
rect 18724 2092 18733 2112
rect 18581 2087 18617 2088
rect 18695 2084 18733 2092
rect 18799 2116 18943 2122
rect 18799 2096 18807 2116
rect 18827 2097 18859 2116
rect 18880 2097 18915 2116
rect 18827 2096 18915 2097
rect 18935 2096 18943 2116
rect 18799 2088 18943 2096
rect 18799 2087 18835 2088
rect 18907 2087 18943 2088
rect 19009 2121 19046 2122
rect 19009 2120 19047 2121
rect 19009 2112 19073 2120
rect 19009 2092 19018 2112
rect 19038 2098 19073 2112
rect 19093 2098 19096 2118
rect 19038 2093 19096 2098
rect 19038 2092 19073 2093
rect 18478 2055 18515 2084
rect 18479 2053 18515 2055
rect 18056 2043 18092 2044
rect 17904 2013 17913 2033
rect 17933 2013 17941 2033
rect 17904 2003 17941 2013
rect 18000 2033 18148 2043
rect 18248 2040 18344 2042
rect 18000 2013 18009 2033
rect 18029 2013 18119 2033
rect 18139 2013 18148 2033
rect 18000 2004 18148 2013
rect 18206 2033 18344 2040
rect 18206 2013 18215 2033
rect 18235 2013 18344 2033
rect 18479 2031 18670 2053
rect 18696 2052 18733 2084
rect 19009 2080 19073 2092
rect 19113 2054 19140 2232
rect 19745 2231 19778 2564
rect 19842 2596 20010 2597
rect 20136 2596 20176 2820
rect 20639 2824 20807 2825
rect 21043 2824 21084 2858
rect 21441 2837 21488 2858
rect 20639 2814 21084 2824
rect 21156 2822 21299 2823
rect 20639 2798 21083 2814
rect 20639 2796 20807 2798
rect 21003 2797 21083 2798
rect 21156 2797 21301 2822
rect 21443 2797 21488 2837
rect 20639 2618 20666 2796
rect 20706 2758 20770 2770
rect 21046 2766 21083 2797
rect 21264 2766 21301 2797
rect 21446 2790 21488 2797
rect 21878 2856 21920 2863
rect 22065 2856 22102 2887
rect 22283 2856 22320 2887
rect 22596 2883 22660 2895
rect 22700 2857 22727 3035
rect 21878 2816 21923 2856
rect 22065 2831 22210 2856
rect 22283 2855 22363 2856
rect 22559 2855 22727 2857
rect 22283 2839 22727 2855
rect 22067 2830 22210 2831
rect 22282 2829 22727 2839
rect 21878 2795 21925 2816
rect 22282 2795 22323 2829
rect 22559 2828 22727 2829
rect 23190 2833 23230 3057
rect 23356 3056 23524 3057
rect 23588 3089 23621 3422
rect 23588 3081 23625 3089
rect 23588 3062 23596 3081
rect 23617 3062 23625 3081
rect 23588 3056 23625 3062
rect 23190 2811 23198 2833
rect 23222 2811 23230 2833
rect 23190 2803 23230 2811
rect 20706 2757 20741 2758
rect 20683 2752 20741 2757
rect 20683 2732 20686 2752
rect 20706 2738 20741 2752
rect 20761 2738 20770 2758
rect 20706 2730 20770 2738
rect 20732 2729 20770 2730
rect 20733 2728 20770 2729
rect 20836 2762 20872 2763
rect 20944 2762 20980 2763
rect 20836 2754 20980 2762
rect 20836 2734 20844 2754
rect 20864 2750 20952 2754
rect 20864 2734 20908 2750
rect 20836 2730 20908 2734
rect 20928 2734 20952 2750
rect 20972 2734 20980 2754
rect 20928 2730 20980 2734
rect 20836 2728 20980 2730
rect 21046 2758 21084 2766
rect 21162 2762 21198 2763
rect 21046 2738 21055 2758
rect 21075 2738 21084 2758
rect 21046 2729 21084 2738
rect 21113 2754 21198 2762
rect 21113 2734 21170 2754
rect 21190 2734 21198 2754
rect 21046 2728 21083 2729
rect 21113 2728 21198 2734
rect 21264 2758 21302 2766
rect 21264 2738 21273 2758
rect 21293 2738 21302 2758
rect 21264 2729 21302 2738
rect 21446 2763 21489 2790
rect 21446 2745 21460 2763
rect 21478 2745 21489 2763
rect 21446 2737 21489 2745
rect 21451 2735 21489 2737
rect 21878 2765 22323 2795
rect 23361 2778 23426 2779
rect 21878 2762 22301 2765
rect 21264 2728 21301 2729
rect 20725 2700 20815 2706
rect 20725 2680 20741 2700
rect 20761 2698 20815 2700
rect 20761 2680 20786 2698
rect 20725 2678 20786 2680
rect 20806 2678 20815 2698
rect 20725 2672 20815 2678
rect 20738 2618 20775 2619
rect 20834 2618 20871 2619
rect 20890 2618 20926 2728
rect 21113 2707 21144 2728
rect 21878 2714 21925 2762
rect 21109 2706 21144 2707
rect 20987 2696 21144 2706
rect 20987 2676 21004 2696
rect 21024 2676 21144 2696
rect 20987 2669 21144 2676
rect 21211 2699 21360 2707
rect 21211 2679 21222 2699
rect 21242 2679 21281 2699
rect 21301 2679 21360 2699
rect 21878 2696 21888 2714
rect 21906 2696 21925 2714
rect 21878 2692 21925 2696
rect 23012 2753 23199 2777
rect 23230 2758 23623 2778
rect 23643 2758 23646 2778
rect 23230 2753 23646 2758
rect 21879 2687 21916 2692
rect 21211 2672 21360 2679
rect 23012 2682 23049 2753
rect 23230 2752 23571 2753
rect 23164 2692 23195 2693
rect 21211 2671 21252 2672
rect 21448 2670 21485 2673
rect 20945 2618 20982 2619
rect 20638 2609 20776 2618
rect 19842 2570 20286 2596
rect 19842 2568 20010 2570
rect 19842 2390 19869 2568
rect 19909 2530 19973 2542
rect 20249 2538 20286 2570
rect 20312 2569 20503 2591
rect 20638 2589 20747 2609
rect 20767 2589 20776 2609
rect 20638 2582 20776 2589
rect 20834 2609 20982 2618
rect 20834 2589 20843 2609
rect 20863 2589 20953 2609
rect 20973 2589 20982 2609
rect 20638 2580 20734 2582
rect 20834 2579 20982 2589
rect 21041 2609 21078 2619
rect 21041 2589 21049 2609
rect 21069 2589 21078 2609
rect 20890 2578 20926 2579
rect 20467 2567 20503 2569
rect 20467 2538 20504 2567
rect 19909 2529 19944 2530
rect 19886 2524 19944 2529
rect 19886 2504 19889 2524
rect 19909 2510 19944 2524
rect 19964 2510 19973 2530
rect 19909 2504 19973 2510
rect 19886 2502 19973 2504
rect 19886 2498 19913 2502
rect 19935 2501 19973 2502
rect 19936 2500 19973 2501
rect 20039 2534 20075 2535
rect 20147 2534 20183 2535
rect 20039 2527 20183 2534
rect 20039 2526 20101 2527
rect 20039 2506 20047 2526
rect 20067 2509 20101 2526
rect 20120 2526 20183 2527
rect 20120 2509 20155 2526
rect 20067 2506 20155 2509
rect 20175 2506 20183 2526
rect 20039 2500 20183 2506
rect 20249 2530 20287 2538
rect 20365 2534 20401 2535
rect 20249 2510 20258 2530
rect 20278 2510 20287 2530
rect 20249 2501 20287 2510
rect 20316 2526 20401 2534
rect 20316 2506 20373 2526
rect 20393 2506 20401 2526
rect 20249 2500 20286 2501
rect 20316 2500 20401 2506
rect 20467 2530 20505 2538
rect 20467 2510 20476 2530
rect 20496 2510 20505 2530
rect 20738 2519 20775 2520
rect 21041 2519 21078 2589
rect 21113 2618 21144 2669
rect 21440 2664 21485 2670
rect 21440 2646 21458 2664
rect 21476 2646 21485 2664
rect 23012 2662 23021 2682
rect 23041 2662 23049 2682
rect 23012 2652 23049 2662
rect 23108 2682 23195 2692
rect 23108 2662 23117 2682
rect 23137 2662 23195 2682
rect 23108 2653 23195 2662
rect 23108 2652 23145 2653
rect 21440 2636 21485 2646
rect 21163 2618 21200 2619
rect 21113 2609 21200 2618
rect 21113 2589 21171 2609
rect 21191 2589 21200 2609
rect 21113 2579 21200 2589
rect 21259 2609 21296 2619
rect 21259 2589 21267 2609
rect 21287 2589 21296 2609
rect 21440 2594 21483 2636
rect 21867 2625 21919 2627
rect 21346 2592 21483 2594
rect 21113 2578 21144 2579
rect 21259 2519 21296 2589
rect 20737 2518 21078 2519
rect 20467 2501 20505 2510
rect 20662 2513 21078 2518
rect 20467 2500 20504 2501
rect 19928 2472 20018 2478
rect 19928 2452 19944 2472
rect 19964 2470 20018 2472
rect 19964 2452 19989 2470
rect 19928 2450 19989 2452
rect 20009 2450 20018 2470
rect 19928 2444 20018 2450
rect 19941 2390 19978 2391
rect 20037 2390 20074 2391
rect 20093 2390 20129 2500
rect 20316 2479 20347 2500
rect 20662 2493 20665 2513
rect 20685 2493 21078 2513
rect 21262 2503 21296 2519
rect 21340 2571 21483 2592
rect 21865 2621 22298 2625
rect 21865 2615 22304 2621
rect 21865 2597 21886 2615
rect 21904 2597 22304 2615
rect 23164 2602 23195 2653
rect 23230 2682 23267 2752
rect 23533 2751 23570 2752
rect 23382 2692 23418 2693
rect 23230 2662 23239 2682
rect 23259 2662 23267 2682
rect 23230 2652 23267 2662
rect 23326 2682 23474 2692
rect 23574 2689 23670 2691
rect 23326 2662 23335 2682
rect 23355 2662 23445 2682
rect 23465 2662 23474 2682
rect 23326 2653 23474 2662
rect 23532 2682 23670 2689
rect 23532 2662 23541 2682
rect 23561 2662 23670 2682
rect 23532 2653 23670 2662
rect 23326 2652 23363 2653
rect 23056 2599 23097 2600
rect 21865 2579 22304 2597
rect 21038 2484 21078 2493
rect 21340 2484 21367 2571
rect 21440 2545 21483 2571
rect 21440 2527 21453 2545
rect 21471 2527 21483 2545
rect 21440 2516 21483 2527
rect 20312 2478 20347 2479
rect 20190 2468 20347 2478
rect 20190 2448 20207 2468
rect 20227 2448 20347 2468
rect 20190 2441 20347 2448
rect 20414 2471 20560 2479
rect 20414 2451 20425 2471
rect 20445 2451 20484 2471
rect 20504 2451 20560 2471
rect 21038 2467 21367 2484
rect 21038 2466 21078 2467
rect 20414 2444 20560 2451
rect 21435 2455 21475 2458
rect 21435 2449 21478 2455
rect 21060 2446 21478 2449
rect 20414 2443 20455 2444
rect 20148 2390 20185 2391
rect 19841 2381 19979 2390
rect 19841 2361 19950 2381
rect 19970 2361 19979 2381
rect 19841 2354 19979 2361
rect 20037 2381 20185 2390
rect 20037 2361 20046 2381
rect 20066 2361 20156 2381
rect 20176 2361 20185 2381
rect 19841 2352 19937 2354
rect 20037 2351 20185 2361
rect 20244 2381 20281 2391
rect 20244 2361 20252 2381
rect 20272 2361 20281 2381
rect 20093 2350 20129 2351
rect 19941 2291 19978 2292
rect 20244 2291 20281 2361
rect 20316 2390 20347 2441
rect 21060 2428 21451 2446
rect 21469 2428 21478 2446
rect 21060 2426 21478 2428
rect 21060 2418 21087 2426
rect 21328 2423 21478 2426
rect 20640 2412 20808 2413
rect 21059 2412 21087 2418
rect 20640 2396 21087 2412
rect 21435 2418 21478 2423
rect 20366 2390 20403 2391
rect 20316 2381 20403 2390
rect 20316 2361 20374 2381
rect 20394 2361 20403 2381
rect 20316 2351 20403 2361
rect 20462 2381 20499 2391
rect 20462 2361 20470 2381
rect 20490 2361 20499 2381
rect 20316 2350 20347 2351
rect 19940 2290 20281 2291
rect 20462 2290 20499 2361
rect 19865 2285 20281 2290
rect 19865 2265 19868 2285
rect 19888 2265 20281 2285
rect 20312 2266 20499 2290
rect 20640 2386 21084 2396
rect 20640 2384 20808 2386
rect 19740 2186 19782 2231
rect 20640 2206 20667 2384
rect 20707 2346 20771 2358
rect 21047 2354 21084 2386
rect 21110 2385 21301 2407
rect 21265 2383 21301 2385
rect 21265 2354 21302 2383
rect 21435 2362 21475 2418
rect 20707 2345 20742 2346
rect 20684 2340 20742 2345
rect 20684 2320 20687 2340
rect 20707 2326 20742 2340
rect 20762 2326 20771 2346
rect 20707 2318 20771 2326
rect 20733 2317 20771 2318
rect 20734 2316 20771 2317
rect 20837 2350 20873 2351
rect 20945 2350 20981 2351
rect 20837 2342 20981 2350
rect 20837 2322 20845 2342
rect 20865 2322 20900 2342
rect 20920 2322 20953 2342
rect 20973 2322 20981 2342
rect 20837 2316 20981 2322
rect 21047 2346 21085 2354
rect 21163 2350 21199 2351
rect 21047 2326 21056 2346
rect 21076 2326 21085 2346
rect 21047 2317 21085 2326
rect 21114 2342 21199 2350
rect 21114 2322 21171 2342
rect 21191 2322 21199 2342
rect 21047 2316 21084 2317
rect 21114 2316 21199 2322
rect 21265 2346 21303 2354
rect 21265 2326 21274 2346
rect 21294 2326 21303 2346
rect 21435 2344 21447 2362
rect 21465 2344 21475 2362
rect 21867 2390 21919 2579
rect 22265 2554 22304 2579
rect 22948 2592 23097 2599
rect 22948 2572 23007 2592
rect 23027 2572 23066 2592
rect 23086 2572 23097 2592
rect 22948 2564 23097 2572
rect 23164 2595 23321 2602
rect 23164 2575 23284 2595
rect 23304 2575 23321 2595
rect 23164 2565 23321 2575
rect 23164 2564 23199 2565
rect 22049 2529 22236 2553
rect 22265 2534 22660 2554
rect 22680 2534 22683 2554
rect 23164 2543 23195 2564
rect 23382 2543 23418 2653
rect 23437 2652 23474 2653
rect 23533 2652 23570 2653
rect 23493 2593 23583 2599
rect 23493 2573 23502 2593
rect 23522 2591 23583 2593
rect 23522 2573 23547 2591
rect 23493 2571 23547 2573
rect 23567 2571 23583 2591
rect 23493 2565 23583 2571
rect 23007 2542 23044 2543
rect 22265 2529 22683 2534
rect 23006 2533 23044 2542
rect 22049 2458 22086 2529
rect 22265 2528 22608 2529
rect 22265 2525 22304 2528
rect 22570 2527 22607 2528
rect 22201 2468 22232 2469
rect 22049 2438 22058 2458
rect 22078 2438 22086 2458
rect 22049 2428 22086 2438
rect 22145 2458 22232 2468
rect 22145 2438 22154 2458
rect 22174 2438 22232 2458
rect 22145 2429 22232 2438
rect 22145 2428 22182 2429
rect 21867 2372 21883 2390
rect 21901 2372 21919 2390
rect 22201 2378 22232 2429
rect 22267 2458 22304 2525
rect 23006 2513 23015 2533
rect 23035 2513 23044 2533
rect 23006 2505 23044 2513
rect 23110 2537 23195 2543
rect 23225 2542 23262 2543
rect 23110 2517 23118 2537
rect 23138 2517 23195 2537
rect 23110 2509 23195 2517
rect 23224 2533 23262 2542
rect 23224 2513 23233 2533
rect 23253 2513 23262 2533
rect 23110 2508 23146 2509
rect 23224 2505 23262 2513
rect 23328 2541 23472 2543
rect 23328 2537 23388 2541
rect 23328 2517 23336 2537
rect 23356 2519 23388 2537
rect 23411 2537 23472 2541
rect 23411 2519 23444 2537
rect 23356 2517 23444 2519
rect 23464 2517 23472 2537
rect 23328 2509 23472 2517
rect 23328 2508 23364 2509
rect 23436 2508 23472 2509
rect 23538 2542 23575 2543
rect 23538 2541 23576 2542
rect 23538 2533 23602 2541
rect 23538 2513 23547 2533
rect 23567 2519 23602 2533
rect 23622 2519 23625 2539
rect 23567 2514 23625 2519
rect 23567 2513 23602 2514
rect 23007 2476 23044 2505
rect 23008 2474 23044 2476
rect 22419 2468 22455 2469
rect 22267 2438 22276 2458
rect 22296 2438 22304 2458
rect 22267 2428 22304 2438
rect 22363 2458 22511 2468
rect 22611 2465 22707 2467
rect 22363 2438 22372 2458
rect 22392 2438 22482 2458
rect 22502 2438 22511 2458
rect 22363 2429 22511 2438
rect 22569 2458 22707 2465
rect 22569 2438 22578 2458
rect 22598 2438 22707 2458
rect 23008 2452 23199 2474
rect 23225 2473 23262 2505
rect 23538 2501 23602 2513
rect 23225 2472 23500 2473
rect 23642 2472 23669 2653
rect 23225 2447 23669 2472
rect 23805 2478 23844 4293
rect 24146 4280 24179 4613
rect 24243 4645 24411 4646
rect 24537 4645 24577 4869
rect 25040 4873 25208 4874
rect 25449 4873 25484 4890
rect 25841 4880 25888 4891
rect 25040 4847 25484 4873
rect 25040 4845 25208 4847
rect 25404 4846 25484 4847
rect 25639 4846 25706 4872
rect 25845 4846 25888 4880
rect 25040 4667 25067 4845
rect 25107 4807 25171 4819
rect 25447 4815 25484 4846
rect 25665 4815 25702 4846
rect 25847 4821 25888 4846
rect 26292 4904 26333 4929
rect 26478 4904 26515 4935
rect 26696 4904 26733 4935
rect 27009 4931 27073 4943
rect 27113 4905 27140 5083
rect 26292 4870 26335 4904
rect 26474 4878 26541 4904
rect 26696 4903 26776 4904
rect 26972 4903 27140 4905
rect 26696 4877 27140 4903
rect 26292 4859 26339 4870
rect 26696 4860 26731 4877
rect 26972 4876 27140 4877
rect 27603 4881 27643 5105
rect 27769 5104 27937 5105
rect 28001 5137 28034 5470
rect 28336 5457 28375 7272
rect 28511 7278 28955 7303
rect 28511 7097 28538 7278
rect 28680 7277 28955 7278
rect 28578 7237 28642 7249
rect 28918 7245 28955 7277
rect 28981 7276 29172 7298
rect 29473 7292 29582 7312
rect 29602 7292 29611 7312
rect 29473 7285 29611 7292
rect 29669 7312 29817 7321
rect 29669 7292 29678 7312
rect 29698 7292 29788 7312
rect 29808 7292 29817 7312
rect 29473 7283 29569 7285
rect 29669 7282 29817 7292
rect 29876 7312 29913 7322
rect 29876 7292 29884 7312
rect 29904 7292 29913 7312
rect 29725 7281 29761 7282
rect 29136 7274 29172 7276
rect 29136 7245 29173 7274
rect 28578 7236 28613 7237
rect 28555 7231 28613 7236
rect 28555 7211 28558 7231
rect 28578 7217 28613 7231
rect 28633 7217 28642 7237
rect 28578 7209 28642 7217
rect 28604 7208 28642 7209
rect 28605 7207 28642 7208
rect 28708 7241 28744 7242
rect 28816 7241 28852 7242
rect 28708 7233 28852 7241
rect 28708 7213 28716 7233
rect 28736 7231 28824 7233
rect 28736 7213 28769 7231
rect 28708 7209 28769 7213
rect 28792 7213 28824 7231
rect 28844 7213 28852 7233
rect 28792 7209 28852 7213
rect 28708 7207 28852 7209
rect 28918 7237 28956 7245
rect 29034 7241 29070 7242
rect 28918 7217 28927 7237
rect 28947 7217 28956 7237
rect 28918 7208 28956 7217
rect 28985 7233 29070 7241
rect 28985 7213 29042 7233
rect 29062 7213 29070 7233
rect 28918 7207 28955 7208
rect 28985 7207 29070 7213
rect 29136 7237 29174 7245
rect 29136 7217 29145 7237
rect 29165 7217 29174 7237
rect 29876 7225 29913 7292
rect 29948 7321 29979 7372
rect 30261 7360 30279 7378
rect 30297 7360 30313 7378
rect 29998 7321 30035 7322
rect 29948 7312 30035 7321
rect 29948 7292 30006 7312
rect 30026 7292 30035 7312
rect 29948 7282 30035 7292
rect 30094 7312 30131 7322
rect 30094 7292 30102 7312
rect 30122 7292 30131 7312
rect 29948 7281 29979 7282
rect 29573 7222 29610 7223
rect 29876 7222 29915 7225
rect 29572 7221 29915 7222
rect 30094 7221 30131 7292
rect 29136 7208 29174 7217
rect 29497 7216 29915 7221
rect 29136 7207 29173 7208
rect 28597 7179 28687 7185
rect 28597 7159 28613 7179
rect 28633 7177 28687 7179
rect 28633 7159 28658 7177
rect 28597 7157 28658 7159
rect 28678 7157 28687 7177
rect 28597 7151 28687 7157
rect 28610 7097 28647 7098
rect 28706 7097 28743 7098
rect 28762 7097 28798 7207
rect 28985 7186 29016 7207
rect 29497 7196 29500 7216
rect 29520 7196 29915 7216
rect 29944 7197 30131 7221
rect 28981 7185 29016 7186
rect 28859 7175 29016 7185
rect 28859 7155 28876 7175
rect 28896 7155 29016 7175
rect 28859 7148 29016 7155
rect 29083 7178 29232 7186
rect 29083 7158 29094 7178
rect 29114 7158 29153 7178
rect 29173 7158 29232 7178
rect 29083 7151 29232 7158
rect 29876 7171 29915 7196
rect 30261 7171 30313 7360
rect 30705 7388 30715 7406
rect 30733 7388 30745 7406
rect 30877 7404 30886 7424
rect 30906 7404 30915 7424
rect 30877 7396 30915 7404
rect 30981 7428 31066 7434
rect 31096 7433 31133 7434
rect 30981 7408 30989 7428
rect 31009 7408 31066 7428
rect 30981 7400 31066 7408
rect 31095 7424 31133 7433
rect 31095 7404 31104 7424
rect 31124 7404 31133 7424
rect 30981 7399 31017 7400
rect 31095 7396 31133 7404
rect 31199 7428 31343 7434
rect 31199 7408 31207 7428
rect 31227 7408 31260 7428
rect 31280 7408 31315 7428
rect 31335 7408 31343 7428
rect 31199 7400 31343 7408
rect 31199 7399 31235 7400
rect 31307 7399 31343 7400
rect 31409 7433 31446 7434
rect 31409 7432 31447 7433
rect 31409 7424 31473 7432
rect 31409 7404 31418 7424
rect 31438 7410 31473 7424
rect 31493 7410 31496 7430
rect 31438 7405 31496 7410
rect 31438 7404 31473 7405
rect 30705 7332 30745 7388
rect 30878 7367 30915 7396
rect 30879 7365 30915 7367
rect 30879 7343 31070 7365
rect 31096 7364 31133 7396
rect 31409 7392 31473 7404
rect 31513 7366 31540 7544
rect 32398 7519 32440 7564
rect 31372 7364 31540 7366
rect 31096 7354 31540 7364
rect 31681 7460 31868 7484
rect 31899 7465 32292 7485
rect 32312 7465 32315 7485
rect 31899 7460 32315 7465
rect 31681 7389 31718 7460
rect 31899 7459 32240 7460
rect 31833 7399 31864 7400
rect 31681 7369 31690 7389
rect 31710 7369 31718 7389
rect 31681 7359 31718 7369
rect 31777 7389 31864 7399
rect 31777 7369 31786 7389
rect 31806 7369 31864 7389
rect 31777 7360 31864 7369
rect 31777 7359 31814 7360
rect 30702 7327 30745 7332
rect 31093 7338 31540 7354
rect 31093 7332 31121 7338
rect 31372 7337 31540 7338
rect 30702 7324 30852 7327
rect 31093 7324 31120 7332
rect 30702 7322 31120 7324
rect 30702 7304 30711 7322
rect 30729 7304 31120 7322
rect 31833 7309 31864 7360
rect 31899 7389 31936 7459
rect 32202 7458 32239 7459
rect 32051 7399 32087 7400
rect 31899 7369 31908 7389
rect 31928 7369 31936 7389
rect 31899 7359 31936 7369
rect 31995 7389 32143 7399
rect 32243 7396 32339 7398
rect 31995 7369 32004 7389
rect 32024 7369 32114 7389
rect 32134 7369 32143 7389
rect 31995 7360 32143 7369
rect 32201 7389 32339 7396
rect 32201 7369 32210 7389
rect 32230 7369 32339 7389
rect 32201 7360 32339 7369
rect 31995 7359 32032 7360
rect 31725 7306 31766 7307
rect 30702 7301 31120 7304
rect 30702 7295 30745 7301
rect 30705 7292 30745 7295
rect 31620 7299 31766 7306
rect 31102 7283 31142 7284
rect 30813 7266 31142 7283
rect 31620 7279 31676 7299
rect 31696 7279 31735 7299
rect 31755 7279 31766 7299
rect 31620 7271 31766 7279
rect 31833 7302 31990 7309
rect 31833 7282 31953 7302
rect 31973 7282 31990 7302
rect 31833 7272 31990 7282
rect 31833 7271 31868 7272
rect 30697 7223 30740 7234
rect 30697 7205 30709 7223
rect 30727 7205 30740 7223
rect 30697 7179 30740 7205
rect 30813 7179 30840 7266
rect 31102 7257 31142 7266
rect 29876 7153 30315 7171
rect 29083 7150 29124 7151
rect 28817 7097 28854 7098
rect 28510 7088 28648 7097
rect 28510 7068 28619 7088
rect 28639 7068 28648 7088
rect 28510 7061 28648 7068
rect 28706 7088 28854 7097
rect 28706 7068 28715 7088
rect 28735 7068 28825 7088
rect 28845 7068 28854 7088
rect 28510 7059 28606 7061
rect 28706 7058 28854 7068
rect 28913 7088 28950 7098
rect 28913 7068 28921 7088
rect 28941 7068 28950 7088
rect 28762 7057 28798 7058
rect 28610 6998 28647 6999
rect 28913 6998 28950 7068
rect 28985 7097 29016 7148
rect 29876 7135 30276 7153
rect 30294 7135 30315 7153
rect 29876 7129 30315 7135
rect 29882 7125 30315 7129
rect 30697 7158 30840 7179
rect 30884 7231 30918 7247
rect 31102 7237 31495 7257
rect 31515 7237 31518 7257
rect 31833 7250 31864 7271
rect 32051 7250 32087 7360
rect 32106 7359 32143 7360
rect 32202 7359 32239 7360
rect 32162 7300 32252 7306
rect 32162 7280 32171 7300
rect 32191 7298 32252 7300
rect 32191 7280 32216 7298
rect 32162 7278 32216 7280
rect 32236 7278 32252 7298
rect 32162 7272 32252 7278
rect 31676 7249 31713 7250
rect 31102 7232 31518 7237
rect 31675 7240 31713 7249
rect 31102 7231 31443 7232
rect 30884 7161 30921 7231
rect 31036 7171 31067 7172
rect 30697 7156 30834 7158
rect 30261 7123 30313 7125
rect 30697 7114 30740 7156
rect 30884 7141 30893 7161
rect 30913 7141 30921 7161
rect 30884 7131 30921 7141
rect 30980 7161 31067 7171
rect 30980 7141 30989 7161
rect 31009 7141 31067 7161
rect 30980 7132 31067 7141
rect 30980 7131 31017 7132
rect 30695 7104 30740 7114
rect 29035 7097 29072 7098
rect 28985 7088 29072 7097
rect 28985 7068 29043 7088
rect 29063 7068 29072 7088
rect 28985 7058 29072 7068
rect 29131 7088 29168 7098
rect 29131 7068 29139 7088
rect 29159 7068 29168 7088
rect 30695 7086 30704 7104
rect 30722 7086 30740 7104
rect 30695 7080 30740 7086
rect 31036 7081 31067 7132
rect 31102 7161 31139 7231
rect 31405 7230 31442 7231
rect 31675 7220 31684 7240
rect 31704 7220 31713 7240
rect 31675 7212 31713 7220
rect 31779 7244 31864 7250
rect 31894 7249 31931 7250
rect 31779 7224 31787 7244
rect 31807 7224 31864 7244
rect 31779 7216 31864 7224
rect 31893 7240 31931 7249
rect 31893 7220 31902 7240
rect 31922 7220 31931 7240
rect 31779 7215 31815 7216
rect 31893 7212 31931 7220
rect 31997 7244 32141 7250
rect 31997 7224 32005 7244
rect 32025 7241 32113 7244
rect 32025 7224 32060 7241
rect 31997 7223 32060 7224
rect 32079 7224 32113 7241
rect 32133 7224 32141 7244
rect 32079 7223 32141 7224
rect 31997 7216 32141 7223
rect 31997 7215 32033 7216
rect 32105 7215 32141 7216
rect 32207 7249 32244 7250
rect 32207 7248 32245 7249
rect 32267 7248 32294 7252
rect 32207 7246 32294 7248
rect 32207 7240 32271 7246
rect 32207 7220 32216 7240
rect 32236 7226 32271 7240
rect 32291 7226 32294 7246
rect 32236 7221 32294 7226
rect 32236 7220 32271 7221
rect 31676 7183 31713 7212
rect 31677 7181 31713 7183
rect 31254 7171 31290 7172
rect 31102 7141 31111 7161
rect 31131 7141 31139 7161
rect 31102 7131 31139 7141
rect 31198 7161 31346 7171
rect 31446 7168 31542 7170
rect 31198 7141 31207 7161
rect 31227 7141 31317 7161
rect 31337 7141 31346 7161
rect 31198 7132 31346 7141
rect 31404 7161 31542 7168
rect 31404 7141 31413 7161
rect 31433 7141 31542 7161
rect 31677 7159 31868 7181
rect 31894 7180 31931 7212
rect 32207 7208 32271 7220
rect 32311 7182 32338 7360
rect 32170 7180 32338 7182
rect 31894 7154 32338 7180
rect 31404 7132 31542 7141
rect 31198 7131 31235 7132
rect 30695 7077 30732 7080
rect 30928 7078 30969 7079
rect 28985 7057 29016 7058
rect 28609 6997 28950 6998
rect 29131 6997 29168 7068
rect 30820 7071 30969 7078
rect 30264 7058 30301 7063
rect 28534 6992 28950 6997
rect 28534 6972 28537 6992
rect 28557 6972 28950 6992
rect 28981 6973 29168 6997
rect 30255 7054 30302 7058
rect 30255 7036 30274 7054
rect 30292 7036 30302 7054
rect 30820 7051 30879 7071
rect 30899 7051 30938 7071
rect 30958 7051 30969 7071
rect 30820 7043 30969 7051
rect 31036 7074 31193 7081
rect 31036 7054 31156 7074
rect 31176 7054 31193 7074
rect 31036 7044 31193 7054
rect 31036 7043 31071 7044
rect 30255 6988 30302 7036
rect 31036 7022 31067 7043
rect 31254 7022 31290 7132
rect 31309 7131 31346 7132
rect 31405 7131 31442 7132
rect 31365 7072 31455 7078
rect 31365 7052 31374 7072
rect 31394 7070 31455 7072
rect 31394 7052 31419 7070
rect 31365 7050 31419 7052
rect 31439 7050 31455 7070
rect 31365 7044 31455 7050
rect 30879 7021 30916 7022
rect 29879 6985 30302 6988
rect 28754 6971 28819 6972
rect 29857 6955 30302 6985
rect 30691 7013 30729 7015
rect 30691 7005 30734 7013
rect 30691 6987 30702 7005
rect 30720 6987 30734 7005
rect 30691 6960 30734 6987
rect 30878 7012 30916 7021
rect 30878 6992 30887 7012
rect 30907 6992 30916 7012
rect 30878 6984 30916 6992
rect 30982 7016 31067 7022
rect 31097 7021 31134 7022
rect 30982 6996 30990 7016
rect 31010 6996 31067 7016
rect 30982 6988 31067 6996
rect 31096 7012 31134 7021
rect 31096 6992 31105 7012
rect 31125 6992 31134 7012
rect 30982 6987 31018 6988
rect 31096 6984 31134 6992
rect 31200 7020 31344 7022
rect 31200 7016 31252 7020
rect 31200 6996 31208 7016
rect 31228 7000 31252 7016
rect 31272 7016 31344 7020
rect 31272 7000 31316 7016
rect 31228 6996 31316 7000
rect 31336 6996 31344 7016
rect 31200 6988 31344 6996
rect 31200 6987 31236 6988
rect 31308 6987 31344 6988
rect 31410 7021 31447 7022
rect 31410 7020 31448 7021
rect 31410 7012 31474 7020
rect 31410 6992 31419 7012
rect 31439 6998 31474 7012
rect 31494 6998 31497 7018
rect 31439 6993 31497 6998
rect 31439 6992 31474 6993
rect 28950 6939 28990 6947
rect 28950 6917 28958 6939
rect 28982 6917 28990 6939
rect 28555 6688 28592 6694
rect 28555 6669 28563 6688
rect 28584 6669 28592 6688
rect 28555 6661 28592 6669
rect 28559 6328 28592 6661
rect 28656 6693 28824 6694
rect 28950 6693 28990 6917
rect 29453 6921 29621 6922
rect 29857 6921 29898 6955
rect 30255 6934 30302 6955
rect 29453 6911 29898 6921
rect 29970 6919 30113 6920
rect 29453 6895 29897 6911
rect 29453 6893 29621 6895
rect 29817 6894 29897 6895
rect 29970 6894 30115 6919
rect 30257 6894 30302 6934
rect 29453 6715 29480 6893
rect 29520 6855 29584 6867
rect 29860 6863 29897 6894
rect 30078 6863 30115 6894
rect 30260 6887 30302 6894
rect 30692 6953 30734 6960
rect 30879 6953 30916 6984
rect 31097 6953 31134 6984
rect 31410 6980 31474 6992
rect 31514 6954 31541 7132
rect 30692 6913 30737 6953
rect 30879 6928 31024 6953
rect 31097 6952 31177 6953
rect 31373 6952 31541 6954
rect 31097 6936 31541 6952
rect 30881 6927 31024 6928
rect 31096 6926 31541 6936
rect 30692 6892 30739 6913
rect 31096 6892 31137 6926
rect 31373 6925 31541 6926
rect 32004 6930 32044 7154
rect 32170 7153 32338 7154
rect 32402 7186 32435 7519
rect 33040 7518 33067 7696
rect 33107 7658 33171 7670
rect 33447 7666 33484 7698
rect 33510 7697 33701 7719
rect 33836 7717 33945 7737
rect 33965 7717 33974 7737
rect 33836 7710 33974 7717
rect 34032 7737 34180 7746
rect 34032 7717 34041 7737
rect 34061 7717 34151 7737
rect 34171 7717 34180 7737
rect 33836 7708 33932 7710
rect 34032 7707 34180 7717
rect 34239 7737 34276 7747
rect 34239 7717 34247 7737
rect 34267 7717 34276 7737
rect 34088 7706 34124 7707
rect 33665 7695 33701 7697
rect 33665 7666 33702 7695
rect 33107 7657 33142 7658
rect 33084 7652 33142 7657
rect 33084 7632 33087 7652
rect 33107 7638 33142 7652
rect 33162 7638 33171 7658
rect 33107 7630 33171 7638
rect 33133 7629 33171 7630
rect 33134 7628 33171 7629
rect 33237 7662 33273 7663
rect 33345 7662 33381 7663
rect 33237 7654 33381 7662
rect 33237 7634 33245 7654
rect 33265 7653 33353 7654
rect 33265 7634 33300 7653
rect 33321 7634 33353 7653
rect 33373 7634 33381 7654
rect 33237 7628 33381 7634
rect 33447 7658 33485 7666
rect 33563 7662 33599 7663
rect 33447 7638 33456 7658
rect 33476 7638 33485 7658
rect 33447 7629 33485 7638
rect 33514 7654 33599 7662
rect 33514 7634 33571 7654
rect 33591 7634 33599 7654
rect 33447 7628 33484 7629
rect 33514 7628 33599 7634
rect 33665 7658 33703 7666
rect 33665 7638 33674 7658
rect 33694 7638 33703 7658
rect 33936 7647 33973 7648
rect 34239 7647 34276 7717
rect 34311 7746 34342 7797
rect 34638 7792 34683 7798
rect 34638 7774 34656 7792
rect 34674 7774 34683 7792
rect 34638 7764 34683 7774
rect 34361 7746 34398 7747
rect 34311 7737 34398 7746
rect 34311 7717 34369 7737
rect 34389 7717 34398 7737
rect 34311 7707 34398 7717
rect 34457 7737 34494 7747
rect 34457 7717 34465 7737
rect 34485 7717 34494 7737
rect 34638 7722 34681 7764
rect 34544 7720 34681 7722
rect 34311 7706 34342 7707
rect 34457 7647 34494 7717
rect 33935 7646 34276 7647
rect 33665 7629 33703 7638
rect 33860 7641 34276 7646
rect 33665 7628 33702 7629
rect 33126 7600 33216 7606
rect 33126 7580 33142 7600
rect 33162 7598 33216 7600
rect 33162 7580 33187 7598
rect 33126 7578 33187 7580
rect 33207 7578 33216 7598
rect 33126 7572 33216 7578
rect 33139 7518 33176 7519
rect 33235 7518 33272 7519
rect 33291 7518 33327 7628
rect 33514 7607 33545 7628
rect 33860 7621 33863 7641
rect 33883 7621 34276 7641
rect 34460 7631 34494 7647
rect 34538 7699 34681 7720
rect 34236 7612 34276 7621
rect 34538 7612 34565 7699
rect 34638 7673 34681 7699
rect 34638 7655 34651 7673
rect 34669 7655 34681 7673
rect 34638 7644 34681 7655
rect 33510 7606 33545 7607
rect 33388 7596 33545 7606
rect 33388 7576 33405 7596
rect 33425 7576 33545 7596
rect 33388 7569 33545 7576
rect 33612 7599 33761 7607
rect 33612 7579 33623 7599
rect 33643 7579 33682 7599
rect 33702 7579 33761 7599
rect 34236 7595 34565 7612
rect 34236 7594 34276 7595
rect 33612 7572 33761 7579
rect 34633 7583 34673 7586
rect 34633 7577 34676 7583
rect 34258 7574 34676 7577
rect 33612 7571 33653 7572
rect 33346 7518 33383 7519
rect 33039 7509 33177 7518
rect 32902 7499 32938 7505
rect 32902 7481 32907 7499
rect 32929 7481 32938 7499
rect 32902 7477 32938 7481
rect 33039 7489 33148 7509
rect 33168 7489 33177 7509
rect 33039 7482 33177 7489
rect 33235 7509 33383 7518
rect 33235 7489 33244 7509
rect 33264 7489 33354 7509
rect 33374 7489 33383 7509
rect 33039 7480 33135 7482
rect 33235 7479 33383 7489
rect 33442 7509 33479 7519
rect 33442 7489 33450 7509
rect 33470 7489 33479 7509
rect 33291 7478 33327 7479
rect 32905 7318 32938 7477
rect 33139 7419 33176 7420
rect 33442 7419 33479 7489
rect 33514 7518 33545 7569
rect 34258 7556 34649 7574
rect 34667 7556 34676 7574
rect 34258 7554 34676 7556
rect 34258 7546 34285 7554
rect 34526 7551 34676 7554
rect 33838 7540 34006 7541
rect 34257 7540 34285 7546
rect 33838 7524 34285 7540
rect 34633 7546 34676 7551
rect 33564 7518 33601 7519
rect 33514 7509 33601 7518
rect 33514 7489 33572 7509
rect 33592 7489 33601 7509
rect 33514 7479 33601 7489
rect 33660 7509 33697 7519
rect 33660 7489 33668 7509
rect 33688 7489 33697 7509
rect 33514 7478 33545 7479
rect 33138 7418 33479 7419
rect 33660 7418 33697 7489
rect 33063 7413 33479 7418
rect 33063 7393 33066 7413
rect 33086 7393 33479 7413
rect 33510 7394 33697 7418
rect 33838 7514 34282 7524
rect 33838 7512 34006 7514
rect 33838 7334 33865 7512
rect 33905 7474 33969 7486
rect 34245 7482 34282 7514
rect 34308 7513 34499 7535
rect 34463 7511 34499 7513
rect 34463 7482 34500 7511
rect 34633 7490 34673 7546
rect 33905 7473 33940 7474
rect 33882 7468 33940 7473
rect 33882 7448 33885 7468
rect 33905 7454 33940 7468
rect 33960 7454 33969 7474
rect 33905 7446 33969 7454
rect 33931 7445 33969 7446
rect 33932 7444 33969 7445
rect 34035 7478 34071 7479
rect 34143 7478 34179 7479
rect 34035 7470 34179 7478
rect 34035 7450 34043 7470
rect 34063 7450 34098 7470
rect 34118 7450 34151 7470
rect 34171 7450 34179 7470
rect 34035 7444 34179 7450
rect 34245 7474 34283 7482
rect 34361 7478 34397 7479
rect 34245 7454 34254 7474
rect 34274 7454 34283 7474
rect 34245 7445 34283 7454
rect 34312 7470 34397 7478
rect 34312 7450 34369 7470
rect 34389 7450 34397 7470
rect 34245 7444 34282 7445
rect 34312 7444 34397 7450
rect 34463 7474 34501 7482
rect 34463 7454 34472 7474
rect 34492 7454 34501 7474
rect 34633 7472 34645 7490
rect 34663 7472 34673 7490
rect 34633 7462 34673 7472
rect 34463 7445 34501 7454
rect 34463 7444 34500 7445
rect 33924 7416 34014 7422
rect 33924 7396 33940 7416
rect 33960 7414 34014 7416
rect 33960 7396 33985 7414
rect 33924 7394 33985 7396
rect 34005 7394 34014 7414
rect 33924 7388 34014 7394
rect 33937 7334 33974 7335
rect 34033 7334 34070 7335
rect 34089 7334 34125 7444
rect 34312 7423 34343 7444
rect 34308 7422 34343 7423
rect 34186 7412 34343 7422
rect 34186 7392 34203 7412
rect 34223 7392 34343 7412
rect 34186 7385 34343 7392
rect 34410 7415 34559 7423
rect 34410 7395 34421 7415
rect 34441 7395 34480 7415
rect 34500 7395 34559 7415
rect 34410 7388 34559 7395
rect 34625 7391 34677 7409
rect 34410 7387 34451 7388
rect 34144 7334 34181 7335
rect 33837 7325 33975 7334
rect 32904 7317 32941 7318
rect 32875 7316 33043 7317
rect 33169 7316 33209 7318
rect 32700 7307 32739 7313
rect 32700 7285 32708 7307
rect 32732 7285 32739 7307
rect 32402 7178 32439 7186
rect 32402 7159 32410 7178
rect 32431 7159 32439 7178
rect 32402 7153 32439 7159
rect 32004 6908 32012 6930
rect 32036 6908 32044 6930
rect 32004 6900 32044 6908
rect 29520 6854 29555 6855
rect 29497 6849 29555 6854
rect 29497 6829 29500 6849
rect 29520 6835 29555 6849
rect 29575 6835 29584 6855
rect 29520 6827 29584 6835
rect 29546 6826 29584 6827
rect 29547 6825 29584 6826
rect 29650 6859 29686 6860
rect 29758 6859 29794 6860
rect 29650 6851 29794 6859
rect 29650 6831 29658 6851
rect 29678 6847 29766 6851
rect 29678 6831 29722 6847
rect 29650 6827 29722 6831
rect 29742 6831 29766 6847
rect 29786 6831 29794 6851
rect 29742 6827 29794 6831
rect 29650 6825 29794 6827
rect 29860 6855 29898 6863
rect 29976 6859 30012 6860
rect 29860 6835 29869 6855
rect 29889 6835 29898 6855
rect 29860 6826 29898 6835
rect 29927 6851 30012 6859
rect 29927 6831 29984 6851
rect 30004 6831 30012 6851
rect 29860 6825 29897 6826
rect 29927 6825 30012 6831
rect 30078 6855 30116 6863
rect 30078 6835 30087 6855
rect 30107 6835 30116 6855
rect 30078 6826 30116 6835
rect 30260 6860 30303 6887
rect 30260 6842 30274 6860
rect 30292 6842 30303 6860
rect 30260 6834 30303 6842
rect 30265 6832 30303 6834
rect 30692 6862 31137 6892
rect 32175 6875 32240 6876
rect 30692 6859 31115 6862
rect 30078 6825 30115 6826
rect 29539 6797 29629 6803
rect 29539 6777 29555 6797
rect 29575 6795 29629 6797
rect 29575 6777 29600 6795
rect 29539 6775 29600 6777
rect 29620 6775 29629 6795
rect 29539 6769 29629 6775
rect 29552 6715 29589 6716
rect 29648 6715 29685 6716
rect 29704 6715 29740 6825
rect 29927 6804 29958 6825
rect 30692 6811 30739 6859
rect 29923 6803 29958 6804
rect 29801 6793 29958 6803
rect 29801 6773 29818 6793
rect 29838 6773 29958 6793
rect 29801 6766 29958 6773
rect 30025 6796 30174 6804
rect 30025 6776 30036 6796
rect 30056 6776 30095 6796
rect 30115 6776 30174 6796
rect 30692 6793 30702 6811
rect 30720 6793 30739 6811
rect 30692 6789 30739 6793
rect 31826 6850 32013 6874
rect 32044 6855 32437 6875
rect 32457 6855 32460 6875
rect 32044 6850 32460 6855
rect 30693 6784 30730 6789
rect 30025 6769 30174 6776
rect 31826 6779 31863 6850
rect 32044 6849 32385 6850
rect 31978 6789 32009 6790
rect 30025 6768 30066 6769
rect 30262 6767 30299 6770
rect 29759 6715 29796 6716
rect 29452 6706 29590 6715
rect 28656 6667 29100 6693
rect 28656 6665 28824 6667
rect 28656 6487 28683 6665
rect 28723 6627 28787 6639
rect 29063 6635 29100 6667
rect 29126 6666 29317 6688
rect 29452 6686 29561 6706
rect 29581 6686 29590 6706
rect 29452 6679 29590 6686
rect 29648 6706 29796 6715
rect 29648 6686 29657 6706
rect 29677 6686 29767 6706
rect 29787 6686 29796 6706
rect 29452 6677 29548 6679
rect 29648 6676 29796 6686
rect 29855 6706 29892 6716
rect 29855 6686 29863 6706
rect 29883 6686 29892 6706
rect 29704 6675 29740 6676
rect 29281 6664 29317 6666
rect 29281 6635 29318 6664
rect 28723 6626 28758 6627
rect 28700 6621 28758 6626
rect 28700 6601 28703 6621
rect 28723 6607 28758 6621
rect 28778 6607 28787 6627
rect 28723 6601 28787 6607
rect 28700 6599 28787 6601
rect 28700 6595 28727 6599
rect 28749 6598 28787 6599
rect 28750 6597 28787 6598
rect 28853 6631 28889 6632
rect 28961 6631 28997 6632
rect 28853 6624 28997 6631
rect 28853 6623 28915 6624
rect 28853 6603 28861 6623
rect 28881 6606 28915 6623
rect 28934 6623 28997 6624
rect 28934 6606 28969 6623
rect 28881 6603 28969 6606
rect 28989 6603 28997 6623
rect 28853 6597 28997 6603
rect 29063 6627 29101 6635
rect 29179 6631 29215 6632
rect 29063 6607 29072 6627
rect 29092 6607 29101 6627
rect 29063 6598 29101 6607
rect 29130 6623 29215 6631
rect 29130 6603 29187 6623
rect 29207 6603 29215 6623
rect 29063 6597 29100 6598
rect 29130 6597 29215 6603
rect 29281 6627 29319 6635
rect 29281 6607 29290 6627
rect 29310 6607 29319 6627
rect 29552 6616 29589 6617
rect 29855 6616 29892 6686
rect 29927 6715 29958 6766
rect 30254 6761 30299 6767
rect 30254 6743 30272 6761
rect 30290 6743 30299 6761
rect 31826 6759 31835 6779
rect 31855 6759 31863 6779
rect 31826 6749 31863 6759
rect 31922 6779 32009 6789
rect 31922 6759 31931 6779
rect 31951 6759 32009 6779
rect 31922 6750 32009 6759
rect 31922 6749 31959 6750
rect 30254 6733 30299 6743
rect 29977 6715 30014 6716
rect 29927 6706 30014 6715
rect 29927 6686 29985 6706
rect 30005 6686 30014 6706
rect 29927 6676 30014 6686
rect 30073 6706 30110 6716
rect 30073 6686 30081 6706
rect 30101 6686 30110 6706
rect 30254 6691 30297 6733
rect 30681 6722 30733 6724
rect 30160 6689 30297 6691
rect 29927 6675 29958 6676
rect 30073 6616 30110 6686
rect 29551 6615 29892 6616
rect 29281 6598 29319 6607
rect 29476 6610 29892 6615
rect 29281 6597 29318 6598
rect 28742 6569 28832 6575
rect 28742 6549 28758 6569
rect 28778 6567 28832 6569
rect 28778 6549 28803 6567
rect 28742 6547 28803 6549
rect 28823 6547 28832 6567
rect 28742 6541 28832 6547
rect 28755 6487 28792 6488
rect 28851 6487 28888 6488
rect 28907 6487 28943 6597
rect 29130 6576 29161 6597
rect 29476 6590 29479 6610
rect 29499 6590 29892 6610
rect 30076 6600 30110 6616
rect 30154 6668 30297 6689
rect 30679 6718 31112 6722
rect 30679 6712 31118 6718
rect 30679 6694 30700 6712
rect 30718 6694 31118 6712
rect 31978 6699 32009 6750
rect 32044 6779 32081 6849
rect 32347 6848 32384 6849
rect 32196 6789 32232 6790
rect 32044 6759 32053 6779
rect 32073 6759 32081 6779
rect 32044 6749 32081 6759
rect 32140 6779 32288 6789
rect 32388 6786 32484 6788
rect 32140 6759 32149 6779
rect 32169 6759 32259 6779
rect 32279 6759 32288 6779
rect 32140 6750 32288 6759
rect 32346 6779 32484 6786
rect 32346 6759 32355 6779
rect 32375 6759 32484 6779
rect 32346 6750 32484 6759
rect 32140 6749 32177 6750
rect 31870 6696 31911 6697
rect 30679 6676 31118 6694
rect 29852 6581 29892 6590
rect 30154 6581 30181 6668
rect 30254 6642 30297 6668
rect 30254 6624 30267 6642
rect 30285 6624 30297 6642
rect 30254 6613 30297 6624
rect 29126 6575 29161 6576
rect 29004 6565 29161 6575
rect 29004 6545 29021 6565
rect 29041 6545 29161 6565
rect 29004 6538 29161 6545
rect 29228 6568 29374 6576
rect 29228 6548 29239 6568
rect 29259 6548 29298 6568
rect 29318 6548 29374 6568
rect 29852 6564 30181 6581
rect 29852 6563 29892 6564
rect 29228 6541 29374 6548
rect 30249 6552 30289 6555
rect 30249 6546 30292 6552
rect 29874 6543 30292 6546
rect 29228 6540 29269 6541
rect 28962 6487 28999 6488
rect 28655 6478 28793 6487
rect 28655 6458 28764 6478
rect 28784 6458 28793 6478
rect 28655 6451 28793 6458
rect 28851 6478 28999 6487
rect 28851 6458 28860 6478
rect 28880 6458 28970 6478
rect 28990 6458 28999 6478
rect 28655 6449 28751 6451
rect 28851 6448 28999 6458
rect 29058 6478 29095 6488
rect 29058 6458 29066 6478
rect 29086 6458 29095 6478
rect 28907 6447 28943 6448
rect 28755 6388 28792 6389
rect 29058 6388 29095 6458
rect 29130 6487 29161 6538
rect 29874 6525 30265 6543
rect 30283 6525 30292 6543
rect 29874 6523 30292 6525
rect 29874 6515 29901 6523
rect 30142 6520 30292 6523
rect 29454 6509 29622 6510
rect 29873 6509 29901 6515
rect 29454 6493 29901 6509
rect 30249 6515 30292 6520
rect 29180 6487 29217 6488
rect 29130 6478 29217 6487
rect 29130 6458 29188 6478
rect 29208 6458 29217 6478
rect 29130 6448 29217 6458
rect 29276 6478 29313 6488
rect 29276 6458 29284 6478
rect 29304 6458 29313 6478
rect 29130 6447 29161 6448
rect 28754 6387 29095 6388
rect 29276 6387 29313 6458
rect 28679 6382 29095 6387
rect 28679 6362 28682 6382
rect 28702 6362 29095 6382
rect 29126 6363 29313 6387
rect 29454 6483 29898 6493
rect 29454 6481 29622 6483
rect 28554 6283 28596 6328
rect 29454 6303 29481 6481
rect 29521 6443 29585 6455
rect 29861 6451 29898 6483
rect 29924 6482 30115 6504
rect 30079 6480 30115 6482
rect 30079 6451 30116 6480
rect 30249 6459 30289 6515
rect 29521 6442 29556 6443
rect 29498 6437 29556 6442
rect 29498 6417 29501 6437
rect 29521 6423 29556 6437
rect 29576 6423 29585 6443
rect 29521 6415 29585 6423
rect 29547 6414 29585 6415
rect 29548 6413 29585 6414
rect 29651 6447 29687 6448
rect 29759 6447 29795 6448
rect 29651 6439 29795 6447
rect 29651 6419 29659 6439
rect 29679 6419 29714 6439
rect 29734 6419 29767 6439
rect 29787 6419 29795 6439
rect 29651 6413 29795 6419
rect 29861 6443 29899 6451
rect 29977 6447 30013 6448
rect 29861 6423 29870 6443
rect 29890 6423 29899 6443
rect 29861 6414 29899 6423
rect 29928 6439 30013 6447
rect 29928 6419 29985 6439
rect 30005 6419 30013 6439
rect 29861 6413 29898 6414
rect 29928 6413 30013 6419
rect 30079 6443 30117 6451
rect 30079 6423 30088 6443
rect 30108 6423 30117 6443
rect 30249 6441 30261 6459
rect 30279 6441 30289 6459
rect 30681 6487 30733 6676
rect 31079 6651 31118 6676
rect 31762 6689 31911 6696
rect 31762 6669 31821 6689
rect 31841 6669 31880 6689
rect 31900 6669 31911 6689
rect 31762 6661 31911 6669
rect 31978 6692 32135 6699
rect 31978 6672 32098 6692
rect 32118 6672 32135 6692
rect 31978 6662 32135 6672
rect 31978 6661 32013 6662
rect 30863 6626 31050 6650
rect 31079 6631 31474 6651
rect 31494 6631 31497 6651
rect 31978 6640 32009 6661
rect 32196 6640 32232 6750
rect 32251 6749 32288 6750
rect 32347 6749 32384 6750
rect 32307 6690 32397 6696
rect 32307 6670 32316 6690
rect 32336 6688 32397 6690
rect 32336 6670 32361 6688
rect 32307 6668 32361 6670
rect 32381 6668 32397 6688
rect 32307 6662 32397 6668
rect 31821 6639 31858 6640
rect 31079 6626 31497 6631
rect 31820 6630 31858 6639
rect 30863 6555 30900 6626
rect 31079 6625 31422 6626
rect 31079 6622 31118 6625
rect 31384 6624 31421 6625
rect 31015 6565 31046 6566
rect 30863 6535 30872 6555
rect 30892 6535 30900 6555
rect 30863 6525 30900 6535
rect 30959 6555 31046 6565
rect 30959 6535 30968 6555
rect 30988 6535 31046 6555
rect 30959 6526 31046 6535
rect 30959 6525 30996 6526
rect 30681 6469 30697 6487
rect 30715 6469 30733 6487
rect 31015 6475 31046 6526
rect 31081 6555 31118 6622
rect 31820 6610 31829 6630
rect 31849 6610 31858 6630
rect 31820 6602 31858 6610
rect 31924 6634 32009 6640
rect 32039 6639 32076 6640
rect 31924 6614 31932 6634
rect 31952 6614 32009 6634
rect 31924 6606 32009 6614
rect 32038 6630 32076 6639
rect 32038 6610 32047 6630
rect 32067 6610 32076 6630
rect 31924 6605 31960 6606
rect 32038 6602 32076 6610
rect 32142 6634 32286 6640
rect 32142 6614 32150 6634
rect 32170 6633 32258 6634
rect 32170 6615 32205 6633
rect 32223 6615 32258 6633
rect 32170 6614 32258 6615
rect 32278 6614 32286 6634
rect 32142 6606 32286 6614
rect 32142 6605 32178 6606
rect 32250 6605 32286 6606
rect 32352 6639 32389 6640
rect 32352 6638 32390 6639
rect 32352 6630 32416 6638
rect 32352 6610 32361 6630
rect 32381 6616 32416 6630
rect 32436 6616 32439 6636
rect 32381 6611 32439 6616
rect 32381 6610 32416 6611
rect 31821 6573 31858 6602
rect 31822 6571 31858 6573
rect 31233 6565 31269 6566
rect 31081 6535 31090 6555
rect 31110 6535 31118 6555
rect 31081 6525 31118 6535
rect 31177 6555 31325 6565
rect 31425 6562 31521 6564
rect 31177 6535 31186 6555
rect 31206 6535 31296 6555
rect 31316 6535 31325 6555
rect 31177 6526 31325 6535
rect 31383 6555 31521 6562
rect 31383 6535 31392 6555
rect 31412 6535 31521 6555
rect 31822 6549 32013 6571
rect 32039 6570 32076 6602
rect 32352 6598 32416 6610
rect 32456 6574 32483 6750
rect 32402 6572 32483 6574
rect 32315 6570 32483 6572
rect 32039 6544 32483 6570
rect 32149 6542 32189 6544
rect 32315 6543 32483 6544
rect 31383 6526 31521 6535
rect 32424 6541 32483 6543
rect 31177 6525 31214 6526
rect 30907 6472 30948 6473
rect 30681 6451 30733 6469
rect 30799 6465 30948 6472
rect 30249 6431 30289 6441
rect 30799 6445 30858 6465
rect 30878 6445 30917 6465
rect 30937 6445 30948 6465
rect 30799 6437 30948 6445
rect 31015 6468 31172 6475
rect 31015 6448 31135 6468
rect 31155 6448 31172 6468
rect 31015 6438 31172 6448
rect 31015 6437 31050 6438
rect 30079 6414 30117 6423
rect 31015 6416 31046 6437
rect 31233 6416 31269 6526
rect 31288 6525 31325 6526
rect 31384 6525 31421 6526
rect 31344 6466 31434 6472
rect 31344 6446 31353 6466
rect 31373 6464 31434 6466
rect 31373 6446 31398 6464
rect 31344 6444 31398 6446
rect 31418 6444 31434 6464
rect 31344 6438 31434 6444
rect 30858 6415 30895 6416
rect 30079 6413 30116 6414
rect 29540 6385 29630 6391
rect 29540 6365 29556 6385
rect 29576 6383 29630 6385
rect 29576 6365 29601 6383
rect 29540 6363 29601 6365
rect 29621 6363 29630 6383
rect 29540 6357 29630 6363
rect 29553 6303 29590 6304
rect 29649 6303 29686 6304
rect 29705 6303 29741 6413
rect 29928 6392 29959 6413
rect 30857 6406 30895 6415
rect 29924 6391 29959 6392
rect 29802 6381 29959 6391
rect 29802 6361 29819 6381
rect 29839 6361 29959 6381
rect 29802 6354 29959 6361
rect 30026 6384 30175 6392
rect 30026 6364 30037 6384
rect 30057 6364 30096 6384
rect 30116 6364 30175 6384
rect 30685 6388 30725 6398
rect 30026 6357 30175 6364
rect 30241 6360 30293 6378
rect 30026 6356 30067 6357
rect 29760 6303 29797 6304
rect 29453 6294 29591 6303
rect 28925 6283 28958 6285
rect 28554 6271 29001 6283
rect 28557 6257 29001 6271
rect 28557 6255 28725 6257
rect 28557 6077 28584 6255
rect 28624 6217 28688 6229
rect 28964 6225 29001 6257
rect 29027 6256 29218 6278
rect 29453 6274 29562 6294
rect 29582 6274 29591 6294
rect 29453 6267 29591 6274
rect 29649 6294 29797 6303
rect 29649 6274 29658 6294
rect 29678 6274 29768 6294
rect 29788 6274 29797 6294
rect 29453 6265 29549 6267
rect 29649 6264 29797 6274
rect 29856 6294 29893 6304
rect 29856 6274 29864 6294
rect 29884 6274 29893 6294
rect 29705 6263 29741 6264
rect 29182 6254 29218 6256
rect 29182 6225 29219 6254
rect 28624 6216 28659 6217
rect 28601 6211 28659 6216
rect 28601 6191 28604 6211
rect 28624 6197 28659 6211
rect 28679 6197 28688 6217
rect 28624 6189 28688 6197
rect 28650 6188 28688 6189
rect 28651 6187 28688 6188
rect 28754 6221 28790 6222
rect 28862 6221 28898 6222
rect 28754 6213 28898 6221
rect 28754 6193 28762 6213
rect 28782 6211 28870 6213
rect 28782 6193 28815 6211
rect 28754 6192 28815 6193
rect 28836 6193 28870 6211
rect 28890 6193 28898 6213
rect 28836 6192 28898 6193
rect 28754 6187 28898 6192
rect 28964 6217 29002 6225
rect 29080 6221 29116 6222
rect 28964 6197 28973 6217
rect 28993 6197 29002 6217
rect 28964 6188 29002 6197
rect 29031 6213 29116 6221
rect 29031 6193 29088 6213
rect 29108 6193 29116 6213
rect 28964 6187 29001 6188
rect 29031 6187 29116 6193
rect 29182 6217 29220 6225
rect 29182 6197 29191 6217
rect 29211 6197 29220 6217
rect 29856 6207 29893 6274
rect 29928 6303 29959 6354
rect 30241 6342 30259 6360
rect 30277 6342 30293 6360
rect 29978 6303 30015 6304
rect 29928 6294 30015 6303
rect 29928 6274 29986 6294
rect 30006 6274 30015 6294
rect 29928 6264 30015 6274
rect 30074 6294 30111 6304
rect 30074 6274 30082 6294
rect 30102 6274 30111 6294
rect 29928 6263 29959 6264
rect 29553 6204 29590 6205
rect 29856 6204 29895 6207
rect 29552 6203 29895 6204
rect 30074 6203 30111 6274
rect 29182 6188 29220 6197
rect 29477 6198 29895 6203
rect 29182 6187 29219 6188
rect 28643 6159 28733 6165
rect 28643 6139 28659 6159
rect 28679 6157 28733 6159
rect 28679 6139 28704 6157
rect 28643 6137 28704 6139
rect 28724 6137 28733 6157
rect 28643 6131 28733 6137
rect 28656 6077 28693 6078
rect 28752 6077 28789 6078
rect 28808 6077 28844 6187
rect 29031 6166 29062 6187
rect 29477 6178 29480 6198
rect 29500 6178 29895 6198
rect 29924 6179 30111 6203
rect 29027 6165 29062 6166
rect 28905 6155 29062 6165
rect 28905 6135 28922 6155
rect 28942 6135 29062 6155
rect 28905 6128 29062 6135
rect 29129 6158 29278 6166
rect 29129 6138 29140 6158
rect 29160 6138 29199 6158
rect 29219 6138 29278 6158
rect 29129 6131 29278 6138
rect 29856 6153 29895 6178
rect 30241 6153 30293 6342
rect 30685 6370 30695 6388
rect 30713 6370 30725 6388
rect 30857 6386 30866 6406
rect 30886 6386 30895 6406
rect 30857 6378 30895 6386
rect 30961 6410 31046 6416
rect 31076 6415 31113 6416
rect 30961 6390 30969 6410
rect 30989 6390 31046 6410
rect 30961 6382 31046 6390
rect 31075 6406 31113 6415
rect 31075 6386 31084 6406
rect 31104 6386 31113 6406
rect 30961 6381 30997 6382
rect 31075 6378 31113 6386
rect 31179 6410 31323 6416
rect 31179 6390 31187 6410
rect 31207 6390 31240 6410
rect 31260 6390 31295 6410
rect 31315 6390 31323 6410
rect 31179 6382 31323 6390
rect 31179 6381 31215 6382
rect 31287 6381 31323 6382
rect 31389 6415 31426 6416
rect 31389 6414 31427 6415
rect 31389 6406 31453 6414
rect 31389 6386 31398 6406
rect 31418 6392 31453 6406
rect 31473 6392 31476 6412
rect 31418 6387 31476 6392
rect 31418 6386 31453 6387
rect 30685 6314 30725 6370
rect 30858 6349 30895 6378
rect 30859 6347 30895 6349
rect 30859 6325 31050 6347
rect 31076 6346 31113 6378
rect 31389 6374 31453 6386
rect 31493 6348 31520 6526
rect 32424 6523 32453 6541
rect 31352 6346 31520 6348
rect 31076 6336 31520 6346
rect 31661 6442 31848 6466
rect 31879 6447 32272 6467
rect 32292 6447 32295 6467
rect 31879 6442 32295 6447
rect 31661 6371 31698 6442
rect 31879 6441 32220 6442
rect 31813 6381 31844 6382
rect 31661 6351 31670 6371
rect 31690 6351 31698 6371
rect 31661 6341 31698 6351
rect 31757 6371 31844 6381
rect 31757 6351 31766 6371
rect 31786 6351 31844 6371
rect 31757 6342 31844 6351
rect 31757 6341 31794 6342
rect 30682 6309 30725 6314
rect 31073 6320 31520 6336
rect 31073 6314 31101 6320
rect 31352 6319 31520 6320
rect 30682 6306 30832 6309
rect 31073 6306 31100 6314
rect 30682 6304 31100 6306
rect 30682 6286 30691 6304
rect 30709 6286 31100 6304
rect 31813 6291 31844 6342
rect 31879 6371 31916 6441
rect 32182 6440 32219 6441
rect 32031 6381 32067 6382
rect 31879 6351 31888 6371
rect 31908 6351 31916 6371
rect 31879 6341 31916 6351
rect 31975 6371 32123 6381
rect 32223 6378 32319 6380
rect 31975 6351 31984 6371
rect 32004 6351 32094 6371
rect 32114 6351 32123 6371
rect 31975 6342 32123 6351
rect 32181 6371 32319 6378
rect 32181 6351 32190 6371
rect 32210 6351 32319 6371
rect 32181 6342 32319 6351
rect 31975 6341 32012 6342
rect 31705 6288 31746 6289
rect 30682 6283 31100 6286
rect 30682 6277 30725 6283
rect 30685 6274 30725 6277
rect 31597 6281 31746 6288
rect 31082 6265 31122 6266
rect 30793 6248 31122 6265
rect 31597 6261 31656 6281
rect 31676 6261 31715 6281
rect 31735 6261 31746 6281
rect 31597 6253 31746 6261
rect 31813 6284 31970 6291
rect 31813 6264 31933 6284
rect 31953 6264 31970 6284
rect 31813 6254 31970 6264
rect 31813 6253 31848 6254
rect 30677 6205 30720 6216
rect 30677 6187 30689 6205
rect 30707 6187 30720 6205
rect 30677 6161 30720 6187
rect 30793 6161 30820 6248
rect 31082 6239 31122 6248
rect 29856 6135 30295 6153
rect 29129 6130 29170 6131
rect 28863 6077 28900 6078
rect 28556 6068 28694 6077
rect 28556 6048 28665 6068
rect 28685 6048 28694 6068
rect 28556 6041 28694 6048
rect 28752 6068 28900 6077
rect 28752 6048 28761 6068
rect 28781 6048 28871 6068
rect 28891 6048 28900 6068
rect 28556 6039 28652 6041
rect 28752 6038 28900 6048
rect 28959 6068 28996 6078
rect 28959 6048 28967 6068
rect 28987 6048 28996 6068
rect 28808 6037 28844 6038
rect 28656 5978 28693 5979
rect 28959 5978 28996 6048
rect 29031 6077 29062 6128
rect 29856 6117 30256 6135
rect 30274 6117 30295 6135
rect 29856 6111 30295 6117
rect 29862 6107 30295 6111
rect 30677 6140 30820 6161
rect 30864 6213 30898 6229
rect 31082 6219 31475 6239
rect 31495 6219 31498 6239
rect 31813 6232 31844 6253
rect 32031 6232 32067 6342
rect 32086 6341 32123 6342
rect 32182 6341 32219 6342
rect 32142 6282 32232 6288
rect 32142 6262 32151 6282
rect 32171 6280 32232 6282
rect 32171 6262 32196 6280
rect 32142 6260 32196 6262
rect 32216 6260 32232 6280
rect 32142 6254 32232 6260
rect 31656 6231 31693 6232
rect 31082 6214 31498 6219
rect 31655 6222 31693 6231
rect 31082 6213 31423 6214
rect 30864 6143 30901 6213
rect 31016 6153 31047 6154
rect 30677 6138 30814 6140
rect 30241 6105 30293 6107
rect 30677 6096 30720 6138
rect 30864 6123 30873 6143
rect 30893 6123 30901 6143
rect 30864 6113 30901 6123
rect 30960 6143 31047 6153
rect 30960 6123 30969 6143
rect 30989 6123 31047 6143
rect 30960 6114 31047 6123
rect 30960 6113 30997 6114
rect 30675 6086 30720 6096
rect 29081 6077 29118 6078
rect 29031 6068 29118 6077
rect 29031 6048 29089 6068
rect 29109 6048 29118 6068
rect 29031 6038 29118 6048
rect 29177 6068 29214 6078
rect 29177 6048 29185 6068
rect 29205 6048 29214 6068
rect 30675 6068 30684 6086
rect 30702 6068 30720 6086
rect 30675 6062 30720 6068
rect 31016 6063 31047 6114
rect 31082 6143 31119 6213
rect 31385 6212 31422 6213
rect 31655 6202 31664 6222
rect 31684 6202 31693 6222
rect 31655 6194 31693 6202
rect 31759 6226 31844 6232
rect 31874 6231 31911 6232
rect 31759 6206 31767 6226
rect 31787 6206 31844 6226
rect 31759 6198 31844 6206
rect 31873 6222 31911 6231
rect 31873 6202 31882 6222
rect 31902 6202 31911 6222
rect 31759 6197 31795 6198
rect 31873 6194 31911 6202
rect 31977 6226 32121 6232
rect 31977 6206 31985 6226
rect 32005 6207 32037 6226
rect 32058 6207 32093 6226
rect 32005 6206 32093 6207
rect 32113 6206 32121 6226
rect 31977 6198 32121 6206
rect 31977 6197 32013 6198
rect 32085 6197 32121 6198
rect 32187 6231 32224 6232
rect 32187 6230 32225 6231
rect 32187 6222 32251 6230
rect 32187 6202 32196 6222
rect 32216 6208 32251 6222
rect 32271 6208 32274 6228
rect 32216 6203 32274 6208
rect 32216 6202 32251 6203
rect 31656 6165 31693 6194
rect 31657 6163 31693 6165
rect 31234 6153 31270 6154
rect 31082 6123 31091 6143
rect 31111 6123 31119 6143
rect 31082 6113 31119 6123
rect 31178 6143 31326 6153
rect 31426 6150 31522 6152
rect 31178 6123 31187 6143
rect 31207 6123 31297 6143
rect 31317 6123 31326 6143
rect 31178 6114 31326 6123
rect 31384 6143 31522 6150
rect 31384 6123 31393 6143
rect 31413 6123 31522 6143
rect 31657 6141 31848 6163
rect 31874 6162 31911 6194
rect 32187 6190 32251 6202
rect 32291 6164 32318 6342
rect 32150 6162 32318 6164
rect 31874 6136 32318 6162
rect 31384 6114 31522 6123
rect 31178 6113 31215 6114
rect 30675 6059 30712 6062
rect 30908 6060 30949 6061
rect 29031 6037 29062 6038
rect 28655 5977 28996 5978
rect 29177 5977 29214 6048
rect 30800 6053 30949 6060
rect 30244 6040 30281 6045
rect 30235 6036 30282 6040
rect 30235 6018 30254 6036
rect 30272 6018 30282 6036
rect 30800 6033 30859 6053
rect 30879 6033 30918 6053
rect 30938 6033 30949 6053
rect 30800 6025 30949 6033
rect 31016 6056 31173 6063
rect 31016 6036 31136 6056
rect 31156 6036 31173 6056
rect 31016 6026 31173 6036
rect 31016 6025 31051 6026
rect 28580 5972 28996 5977
rect 28580 5952 28583 5972
rect 28603 5952 28996 5972
rect 29027 5953 29214 5977
rect 29839 5975 29879 5980
rect 30235 5975 30282 6018
rect 31016 6004 31047 6025
rect 31234 6004 31270 6114
rect 31289 6113 31326 6114
rect 31385 6113 31422 6114
rect 31345 6054 31435 6060
rect 31345 6034 31354 6054
rect 31374 6052 31435 6054
rect 31374 6034 31399 6052
rect 31345 6032 31399 6034
rect 31419 6032 31435 6052
rect 31345 6026 31435 6032
rect 30859 6003 30896 6004
rect 29839 5936 30282 5975
rect 30672 5995 30709 5997
rect 30672 5987 30714 5995
rect 30672 5969 30682 5987
rect 30700 5969 30714 5987
rect 30672 5960 30714 5969
rect 30858 5994 30896 6003
rect 30858 5974 30867 5994
rect 30887 5974 30896 5994
rect 30858 5966 30896 5974
rect 30962 5998 31047 6004
rect 31077 6003 31114 6004
rect 30962 5978 30970 5998
rect 30990 5978 31047 5998
rect 30962 5970 31047 5978
rect 31076 5994 31114 6003
rect 31076 5974 31085 5994
rect 31105 5974 31114 5994
rect 30962 5969 30998 5970
rect 31076 5966 31114 5974
rect 31180 6002 31324 6004
rect 31180 5998 31232 6002
rect 31180 5978 31188 5998
rect 31208 5982 31232 5998
rect 31252 5998 31324 6002
rect 31252 5982 31296 5998
rect 31208 5978 31296 5982
rect 31316 5978 31324 5998
rect 31180 5970 31324 5978
rect 31180 5969 31216 5970
rect 31288 5969 31324 5970
rect 31390 6003 31427 6004
rect 31390 6002 31428 6003
rect 31390 5994 31454 6002
rect 31390 5974 31399 5994
rect 31419 5980 31454 5994
rect 31474 5980 31477 6000
rect 31419 5975 31477 5980
rect 31419 5974 31454 5975
rect 28933 5921 28973 5929
rect 28933 5899 28941 5921
rect 28965 5899 28973 5921
rect 28639 5675 28807 5676
rect 28933 5675 28973 5899
rect 29436 5903 29604 5904
rect 29839 5903 29879 5936
rect 30235 5903 30282 5936
rect 30673 5935 30714 5960
rect 30859 5935 30896 5966
rect 31077 5935 31114 5966
rect 31390 5962 31454 5974
rect 31494 5936 31521 6114
rect 30673 5908 30722 5935
rect 30858 5909 30907 5935
rect 31076 5934 31157 5935
rect 31353 5934 31521 5936
rect 31076 5909 31521 5934
rect 31077 5908 31521 5909
rect 29436 5902 29880 5903
rect 29436 5877 29881 5902
rect 29436 5875 29604 5877
rect 29800 5876 29881 5877
rect 30050 5876 30099 5902
rect 30235 5876 30284 5903
rect 29436 5697 29463 5875
rect 29503 5837 29567 5849
rect 29843 5845 29880 5876
rect 30061 5845 30098 5876
rect 30243 5851 30284 5876
rect 30675 5875 30722 5908
rect 31078 5875 31118 5908
rect 31353 5907 31521 5908
rect 31984 5912 32024 6136
rect 32150 6135 32318 6136
rect 31984 5890 31992 5912
rect 32016 5890 32024 5912
rect 31984 5882 32024 5890
rect 29503 5836 29538 5837
rect 29480 5831 29538 5836
rect 29480 5811 29483 5831
rect 29503 5817 29538 5831
rect 29558 5817 29567 5837
rect 29503 5809 29567 5817
rect 29529 5808 29567 5809
rect 29530 5807 29567 5808
rect 29633 5841 29669 5842
rect 29741 5841 29777 5842
rect 29633 5833 29777 5841
rect 29633 5813 29641 5833
rect 29661 5829 29749 5833
rect 29661 5813 29705 5829
rect 29633 5809 29705 5813
rect 29725 5813 29749 5829
rect 29769 5813 29777 5833
rect 29725 5809 29777 5813
rect 29633 5807 29777 5809
rect 29843 5837 29881 5845
rect 29959 5841 29995 5842
rect 29843 5817 29852 5837
rect 29872 5817 29881 5837
rect 29843 5808 29881 5817
rect 29910 5833 29995 5841
rect 29910 5813 29967 5833
rect 29987 5813 29995 5833
rect 29843 5807 29880 5808
rect 29910 5807 29995 5813
rect 30061 5837 30099 5845
rect 30061 5817 30070 5837
rect 30090 5817 30099 5837
rect 30061 5808 30099 5817
rect 30243 5842 30285 5851
rect 30243 5824 30257 5842
rect 30275 5824 30285 5842
rect 30243 5816 30285 5824
rect 30248 5814 30285 5816
rect 30675 5836 31118 5875
rect 30061 5807 30098 5808
rect 29522 5779 29612 5785
rect 29522 5759 29538 5779
rect 29558 5777 29612 5779
rect 29558 5759 29583 5777
rect 29522 5757 29583 5759
rect 29603 5757 29612 5777
rect 29522 5751 29612 5757
rect 29535 5697 29572 5698
rect 29631 5697 29668 5698
rect 29687 5697 29723 5807
rect 29910 5786 29941 5807
rect 30675 5793 30722 5836
rect 31078 5831 31118 5836
rect 31743 5834 31930 5858
rect 31961 5839 32354 5859
rect 32374 5839 32377 5859
rect 31961 5834 32377 5839
rect 29906 5785 29941 5786
rect 29784 5775 29941 5785
rect 29784 5755 29801 5775
rect 29821 5755 29941 5775
rect 29784 5748 29941 5755
rect 30008 5778 30157 5786
rect 30008 5758 30019 5778
rect 30039 5758 30078 5778
rect 30098 5758 30157 5778
rect 30675 5775 30685 5793
rect 30703 5775 30722 5793
rect 30675 5771 30722 5775
rect 30676 5766 30713 5771
rect 30008 5751 30157 5758
rect 31743 5763 31780 5834
rect 31961 5833 32302 5834
rect 31895 5773 31926 5774
rect 30008 5750 30049 5751
rect 30245 5749 30282 5752
rect 29742 5697 29779 5698
rect 29435 5688 29573 5697
rect 28639 5649 29083 5675
rect 28639 5647 28807 5649
rect 28639 5469 28666 5647
rect 28706 5609 28770 5621
rect 29046 5617 29083 5649
rect 29109 5648 29300 5670
rect 29435 5668 29544 5688
rect 29564 5668 29573 5688
rect 29435 5661 29573 5668
rect 29631 5688 29779 5697
rect 29631 5668 29640 5688
rect 29660 5668 29750 5688
rect 29770 5668 29779 5688
rect 29435 5659 29531 5661
rect 29631 5658 29779 5668
rect 29838 5688 29875 5698
rect 29838 5668 29846 5688
rect 29866 5668 29875 5688
rect 29687 5657 29723 5658
rect 29264 5646 29300 5648
rect 29264 5617 29301 5646
rect 28706 5608 28741 5609
rect 28683 5603 28741 5608
rect 28683 5583 28686 5603
rect 28706 5589 28741 5603
rect 28761 5589 28770 5609
rect 28706 5581 28770 5589
rect 28732 5580 28770 5581
rect 28733 5579 28770 5580
rect 28836 5613 28872 5614
rect 28944 5613 28980 5614
rect 28836 5605 28980 5613
rect 28836 5585 28844 5605
rect 28864 5604 28952 5605
rect 28864 5585 28899 5604
rect 28920 5585 28952 5604
rect 28972 5585 28980 5605
rect 28836 5579 28980 5585
rect 29046 5609 29084 5617
rect 29162 5613 29198 5614
rect 29046 5589 29055 5609
rect 29075 5589 29084 5609
rect 29046 5580 29084 5589
rect 29113 5605 29198 5613
rect 29113 5585 29170 5605
rect 29190 5585 29198 5605
rect 29046 5579 29083 5580
rect 29113 5579 29198 5585
rect 29264 5609 29302 5617
rect 29264 5589 29273 5609
rect 29293 5589 29302 5609
rect 29535 5598 29572 5599
rect 29838 5598 29875 5668
rect 29910 5697 29941 5748
rect 30237 5743 30282 5749
rect 30237 5725 30255 5743
rect 30273 5725 30282 5743
rect 31743 5743 31752 5763
rect 31772 5743 31780 5763
rect 31743 5733 31780 5743
rect 31839 5763 31926 5773
rect 31839 5743 31848 5763
rect 31868 5743 31926 5763
rect 31839 5734 31926 5743
rect 31839 5733 31876 5734
rect 30237 5715 30282 5725
rect 29960 5697 29997 5698
rect 29910 5688 29997 5697
rect 29910 5668 29968 5688
rect 29988 5668 29997 5688
rect 29910 5658 29997 5668
rect 30056 5688 30093 5698
rect 30056 5668 30064 5688
rect 30084 5668 30093 5688
rect 30237 5673 30280 5715
rect 30664 5704 30716 5706
rect 30143 5671 30280 5673
rect 29910 5657 29941 5658
rect 30056 5598 30093 5668
rect 29534 5597 29875 5598
rect 29264 5580 29302 5589
rect 29459 5592 29875 5597
rect 29264 5579 29301 5580
rect 28725 5551 28815 5557
rect 28725 5531 28741 5551
rect 28761 5549 28815 5551
rect 28761 5531 28786 5549
rect 28725 5529 28786 5531
rect 28806 5529 28815 5549
rect 28725 5523 28815 5529
rect 28738 5469 28775 5470
rect 28834 5469 28871 5470
rect 28890 5469 28926 5579
rect 29113 5558 29144 5579
rect 29459 5572 29462 5592
rect 29482 5572 29875 5592
rect 30059 5582 30093 5598
rect 30137 5650 30280 5671
rect 30662 5700 31095 5704
rect 30662 5694 31101 5700
rect 30662 5676 30683 5694
rect 30701 5676 31101 5694
rect 31895 5683 31926 5734
rect 31961 5763 31998 5833
rect 32264 5832 32301 5833
rect 32113 5773 32149 5774
rect 31961 5743 31970 5763
rect 31990 5743 31998 5763
rect 31961 5733 31998 5743
rect 32057 5763 32205 5773
rect 32305 5770 32401 5772
rect 32057 5743 32066 5763
rect 32086 5743 32176 5763
rect 32196 5743 32205 5763
rect 32057 5734 32205 5743
rect 32263 5763 32401 5770
rect 32263 5743 32272 5763
rect 32292 5743 32401 5763
rect 32263 5734 32401 5743
rect 32057 5733 32094 5734
rect 31787 5680 31828 5681
rect 30662 5658 31101 5676
rect 29835 5563 29875 5572
rect 30137 5563 30164 5650
rect 30237 5624 30280 5650
rect 30237 5606 30250 5624
rect 30268 5606 30280 5624
rect 30237 5595 30280 5606
rect 29109 5557 29144 5558
rect 28987 5547 29144 5557
rect 28987 5527 29004 5547
rect 29024 5527 29144 5547
rect 28987 5520 29144 5527
rect 29211 5550 29360 5558
rect 29211 5530 29222 5550
rect 29242 5530 29281 5550
rect 29301 5530 29360 5550
rect 29835 5546 30164 5563
rect 29835 5545 29875 5546
rect 29211 5523 29360 5530
rect 30232 5534 30272 5537
rect 30232 5528 30275 5534
rect 29857 5525 30275 5528
rect 29211 5522 29252 5523
rect 28945 5469 28982 5470
rect 28638 5460 28776 5469
rect 28336 5285 28376 5457
rect 28638 5440 28747 5460
rect 28767 5440 28776 5460
rect 28638 5433 28776 5440
rect 28834 5460 28982 5469
rect 28834 5440 28843 5460
rect 28863 5440 28953 5460
rect 28973 5440 28982 5460
rect 28638 5431 28734 5433
rect 28834 5430 28982 5440
rect 29041 5460 29078 5470
rect 29041 5440 29049 5460
rect 29069 5440 29078 5460
rect 28890 5429 28926 5430
rect 28738 5370 28775 5371
rect 29041 5370 29078 5440
rect 29113 5469 29144 5520
rect 29857 5507 30248 5525
rect 30266 5507 30275 5525
rect 29857 5505 30275 5507
rect 29857 5497 29884 5505
rect 30125 5502 30275 5505
rect 29437 5491 29605 5492
rect 29856 5491 29884 5497
rect 29437 5475 29884 5491
rect 30232 5497 30275 5502
rect 29163 5469 29200 5470
rect 29113 5460 29200 5469
rect 29113 5440 29171 5460
rect 29191 5440 29200 5460
rect 29113 5430 29200 5440
rect 29259 5460 29296 5470
rect 29259 5440 29267 5460
rect 29287 5440 29296 5460
rect 29113 5429 29144 5430
rect 28737 5369 29078 5370
rect 29259 5369 29296 5440
rect 28662 5364 29078 5369
rect 28662 5344 28665 5364
rect 28685 5344 29078 5364
rect 29109 5345 29296 5369
rect 29437 5465 29881 5475
rect 29437 5463 29605 5465
rect 29437 5285 29464 5463
rect 29504 5425 29568 5437
rect 29844 5433 29881 5465
rect 29907 5464 30098 5486
rect 30062 5462 30098 5464
rect 30062 5433 30099 5462
rect 30232 5441 30272 5497
rect 29504 5424 29539 5425
rect 29481 5419 29539 5424
rect 29481 5399 29484 5419
rect 29504 5405 29539 5419
rect 29559 5405 29568 5425
rect 29504 5397 29568 5405
rect 29530 5396 29568 5397
rect 29531 5395 29568 5396
rect 29634 5429 29670 5430
rect 29742 5429 29778 5430
rect 29634 5421 29778 5429
rect 29634 5401 29642 5421
rect 29662 5401 29697 5421
rect 29717 5401 29750 5421
rect 29770 5401 29778 5421
rect 29634 5395 29778 5401
rect 29844 5425 29882 5433
rect 29960 5429 29996 5430
rect 29844 5405 29853 5425
rect 29873 5405 29882 5425
rect 29844 5396 29882 5405
rect 29911 5421 29996 5429
rect 29911 5401 29968 5421
rect 29988 5401 29996 5421
rect 29844 5395 29881 5396
rect 29911 5395 29996 5401
rect 30062 5425 30100 5433
rect 30062 5405 30071 5425
rect 30091 5405 30100 5425
rect 30232 5423 30244 5441
rect 30262 5423 30272 5441
rect 30664 5469 30716 5658
rect 31062 5633 31101 5658
rect 31679 5673 31828 5680
rect 31679 5653 31738 5673
rect 31758 5653 31797 5673
rect 31817 5653 31828 5673
rect 31679 5645 31828 5653
rect 31895 5676 32052 5683
rect 31895 5656 32015 5676
rect 32035 5656 32052 5676
rect 31895 5646 32052 5656
rect 31895 5645 31930 5646
rect 30846 5608 31033 5632
rect 31062 5613 31457 5633
rect 31477 5613 31480 5633
rect 31895 5624 31926 5645
rect 32113 5624 32149 5734
rect 32168 5733 32205 5734
rect 32264 5733 32301 5734
rect 32224 5674 32314 5680
rect 32224 5654 32233 5674
rect 32253 5672 32314 5674
rect 32253 5654 32278 5672
rect 32224 5652 32278 5654
rect 32298 5652 32314 5672
rect 32224 5646 32314 5652
rect 31738 5623 31775 5624
rect 31062 5608 31480 5613
rect 31737 5614 31775 5623
rect 30846 5537 30883 5608
rect 31062 5607 31405 5608
rect 31062 5604 31101 5607
rect 31367 5606 31404 5607
rect 30998 5547 31029 5548
rect 30846 5517 30855 5537
rect 30875 5517 30883 5537
rect 30846 5507 30883 5517
rect 30942 5537 31029 5547
rect 30942 5517 30951 5537
rect 30971 5517 31029 5537
rect 30942 5508 31029 5517
rect 30942 5507 30979 5508
rect 30664 5451 30680 5469
rect 30698 5451 30716 5469
rect 30998 5457 31029 5508
rect 31064 5537 31101 5604
rect 31737 5594 31746 5614
rect 31766 5594 31775 5614
rect 31737 5586 31775 5594
rect 31841 5618 31926 5624
rect 31956 5623 31993 5624
rect 31841 5598 31849 5618
rect 31869 5598 31926 5618
rect 31841 5590 31926 5598
rect 31955 5614 31993 5623
rect 31955 5594 31964 5614
rect 31984 5594 31993 5614
rect 31841 5589 31877 5590
rect 31955 5586 31993 5594
rect 32059 5618 32203 5624
rect 32059 5598 32067 5618
rect 32087 5613 32175 5618
rect 32087 5598 32123 5613
rect 32059 5596 32123 5598
rect 32142 5598 32175 5613
rect 32195 5598 32203 5618
rect 32142 5596 32203 5598
rect 32059 5590 32203 5596
rect 32059 5589 32095 5590
rect 32167 5589 32203 5590
rect 32269 5623 32306 5624
rect 32269 5622 32307 5623
rect 32269 5614 32333 5622
rect 32269 5594 32278 5614
rect 32298 5600 32333 5614
rect 32353 5600 32356 5620
rect 32298 5595 32356 5600
rect 32298 5594 32333 5595
rect 31738 5557 31775 5586
rect 31739 5555 31775 5557
rect 31216 5547 31252 5548
rect 31064 5517 31073 5537
rect 31093 5517 31101 5537
rect 31064 5507 31101 5517
rect 31160 5537 31308 5547
rect 31408 5544 31504 5546
rect 31160 5517 31169 5537
rect 31189 5517 31279 5537
rect 31299 5517 31308 5537
rect 31160 5508 31308 5517
rect 31366 5537 31504 5544
rect 31366 5517 31375 5537
rect 31395 5517 31504 5537
rect 31739 5533 31930 5555
rect 31956 5554 31993 5586
rect 32269 5582 32333 5594
rect 32373 5556 32400 5734
rect 32232 5554 32400 5556
rect 31956 5540 32400 5554
rect 32424 5577 32452 6523
rect 32424 5547 32469 5577
rect 31956 5528 32403 5540
rect 31999 5526 32032 5528
rect 31366 5508 31504 5517
rect 31160 5507 31197 5508
rect 30890 5454 30931 5455
rect 30664 5433 30716 5451
rect 30782 5447 30931 5454
rect 30232 5413 30272 5423
rect 30782 5427 30841 5447
rect 30861 5427 30900 5447
rect 30920 5427 30931 5447
rect 30782 5419 30931 5427
rect 30998 5450 31155 5457
rect 30998 5430 31118 5450
rect 31138 5430 31155 5450
rect 30998 5420 31155 5430
rect 30998 5419 31033 5420
rect 30062 5396 30100 5405
rect 30998 5398 31029 5419
rect 31216 5398 31252 5508
rect 31271 5507 31308 5508
rect 31367 5507 31404 5508
rect 31327 5448 31417 5454
rect 31327 5428 31336 5448
rect 31356 5446 31417 5448
rect 31356 5428 31381 5446
rect 31327 5426 31381 5428
rect 31401 5426 31417 5446
rect 31327 5420 31417 5426
rect 30841 5397 30878 5398
rect 30062 5395 30099 5396
rect 29523 5367 29613 5373
rect 29523 5347 29539 5367
rect 29559 5365 29613 5367
rect 29559 5347 29584 5365
rect 29523 5345 29584 5347
rect 29604 5345 29613 5365
rect 29523 5339 29613 5345
rect 29536 5285 29573 5286
rect 29632 5285 29669 5286
rect 29688 5285 29724 5395
rect 29911 5374 29942 5395
rect 30840 5388 30878 5397
rect 29907 5373 29942 5374
rect 29785 5363 29942 5373
rect 29785 5343 29802 5363
rect 29822 5343 29942 5363
rect 29785 5336 29942 5343
rect 30009 5366 30158 5374
rect 30009 5346 30020 5366
rect 30040 5346 30079 5366
rect 30099 5346 30158 5366
rect 30668 5370 30708 5380
rect 30009 5339 30158 5346
rect 30224 5342 30276 5360
rect 30009 5338 30050 5339
rect 29743 5285 29780 5286
rect 28337 5270 28376 5285
rect 29436 5276 29574 5285
rect 28337 5269 28503 5270
rect 28629 5269 28669 5271
rect 28337 5243 28779 5269
rect 28337 5241 28503 5243
rect 28001 5129 28038 5137
rect 28001 5110 28009 5129
rect 28030 5110 28038 5129
rect 28001 5104 28038 5110
rect 28337 5063 28362 5241
rect 28402 5203 28466 5215
rect 28742 5211 28779 5243
rect 28805 5242 28996 5264
rect 29436 5256 29545 5276
rect 29565 5256 29574 5276
rect 29436 5249 29574 5256
rect 29632 5276 29780 5285
rect 29632 5256 29641 5276
rect 29661 5256 29751 5276
rect 29771 5256 29780 5276
rect 29436 5247 29532 5249
rect 29632 5246 29780 5256
rect 29839 5276 29876 5286
rect 29839 5256 29847 5276
rect 29867 5256 29876 5276
rect 29688 5245 29724 5246
rect 28960 5240 28996 5242
rect 28960 5211 28997 5240
rect 28402 5202 28437 5203
rect 28379 5197 28437 5202
rect 28379 5177 28382 5197
rect 28402 5183 28437 5197
rect 28457 5183 28466 5203
rect 28402 5175 28466 5183
rect 28428 5174 28466 5175
rect 28429 5173 28466 5174
rect 28532 5207 28568 5208
rect 28640 5207 28676 5208
rect 28532 5202 28676 5207
rect 28532 5199 28594 5202
rect 28532 5179 28540 5199
rect 28560 5179 28594 5199
rect 28532 5176 28594 5179
rect 28620 5199 28676 5202
rect 28620 5179 28648 5199
rect 28668 5179 28676 5199
rect 28620 5176 28676 5179
rect 28532 5173 28676 5176
rect 28742 5203 28780 5211
rect 28858 5207 28894 5208
rect 28742 5183 28751 5203
rect 28771 5183 28780 5203
rect 28742 5174 28780 5183
rect 28809 5199 28894 5207
rect 28809 5179 28866 5199
rect 28886 5179 28894 5199
rect 28742 5173 28779 5174
rect 28809 5173 28894 5179
rect 28960 5203 28998 5211
rect 28960 5183 28969 5203
rect 28989 5183 28998 5203
rect 29839 5189 29876 5256
rect 29911 5285 29942 5336
rect 30224 5324 30242 5342
rect 30260 5324 30276 5342
rect 29961 5285 29998 5286
rect 29911 5276 29998 5285
rect 29911 5256 29969 5276
rect 29989 5256 29998 5276
rect 29911 5246 29998 5256
rect 30057 5276 30094 5286
rect 30057 5256 30065 5276
rect 30085 5256 30094 5276
rect 29911 5245 29942 5246
rect 29536 5186 29573 5187
rect 29839 5186 29878 5189
rect 29535 5185 29878 5186
rect 30057 5185 30094 5256
rect 28960 5174 28998 5183
rect 29460 5180 29878 5185
rect 28960 5173 28997 5174
rect 28421 5145 28511 5151
rect 28421 5125 28437 5145
rect 28457 5143 28511 5145
rect 28457 5125 28482 5143
rect 28421 5123 28482 5125
rect 28502 5123 28511 5143
rect 28421 5117 28511 5123
rect 28434 5063 28471 5064
rect 28530 5063 28567 5064
rect 28586 5063 28622 5173
rect 28809 5152 28840 5173
rect 29460 5160 29463 5180
rect 29483 5160 29878 5180
rect 29907 5161 30094 5185
rect 28805 5151 28840 5152
rect 28683 5141 28840 5151
rect 28683 5121 28700 5141
rect 28720 5121 28840 5141
rect 28683 5114 28840 5121
rect 28907 5144 29056 5152
rect 28907 5124 28918 5144
rect 28938 5124 28977 5144
rect 28997 5124 29056 5144
rect 28907 5117 29056 5124
rect 29839 5135 29878 5160
rect 30224 5135 30276 5324
rect 30668 5352 30678 5370
rect 30696 5352 30708 5370
rect 30840 5368 30849 5388
rect 30869 5368 30878 5388
rect 30840 5360 30878 5368
rect 30944 5392 31029 5398
rect 31059 5397 31096 5398
rect 30944 5372 30952 5392
rect 30972 5372 31029 5392
rect 30944 5364 31029 5372
rect 31058 5388 31096 5397
rect 31058 5368 31067 5388
rect 31087 5368 31096 5388
rect 30944 5363 30980 5364
rect 31058 5360 31096 5368
rect 31162 5392 31306 5398
rect 31162 5372 31170 5392
rect 31190 5372 31223 5392
rect 31243 5372 31278 5392
rect 31298 5372 31306 5392
rect 31162 5364 31306 5372
rect 31162 5363 31198 5364
rect 31270 5363 31306 5364
rect 31372 5397 31409 5398
rect 31372 5396 31410 5397
rect 31372 5388 31436 5396
rect 31372 5368 31381 5388
rect 31401 5374 31436 5388
rect 31456 5374 31459 5394
rect 31401 5369 31459 5374
rect 31401 5368 31436 5369
rect 30668 5296 30708 5352
rect 30841 5331 30878 5360
rect 30842 5329 30878 5331
rect 30842 5307 31033 5329
rect 31059 5328 31096 5360
rect 31372 5356 31436 5368
rect 31476 5330 31503 5508
rect 32361 5483 32403 5528
rect 32424 5529 32435 5547
rect 32457 5529 32469 5547
rect 32424 5523 32469 5529
rect 32425 5522 32469 5523
rect 31335 5328 31503 5330
rect 31059 5318 31503 5328
rect 31644 5424 31831 5448
rect 31862 5429 32255 5449
rect 32275 5429 32278 5449
rect 31862 5424 32278 5429
rect 31644 5353 31681 5424
rect 31862 5423 32203 5424
rect 31796 5363 31827 5364
rect 31644 5333 31653 5353
rect 31673 5333 31681 5353
rect 31644 5323 31681 5333
rect 31740 5353 31827 5363
rect 31740 5333 31749 5353
rect 31769 5333 31827 5353
rect 31740 5324 31827 5333
rect 31740 5323 31777 5324
rect 30665 5291 30708 5296
rect 31056 5302 31503 5318
rect 31056 5296 31084 5302
rect 31335 5301 31503 5302
rect 30665 5288 30815 5291
rect 31056 5288 31083 5296
rect 30665 5286 31083 5288
rect 30665 5268 30674 5286
rect 30692 5268 31083 5286
rect 31796 5273 31827 5324
rect 31862 5353 31899 5423
rect 32165 5422 32202 5423
rect 32014 5363 32050 5364
rect 31862 5333 31871 5353
rect 31891 5333 31899 5353
rect 31862 5323 31899 5333
rect 31958 5353 32106 5363
rect 32206 5360 32302 5362
rect 31958 5333 31967 5353
rect 31987 5333 32077 5353
rect 32097 5333 32106 5353
rect 31958 5324 32106 5333
rect 32164 5353 32302 5360
rect 32164 5333 32173 5353
rect 32193 5333 32302 5353
rect 32164 5324 32302 5333
rect 31958 5323 31995 5324
rect 31688 5270 31729 5271
rect 30665 5265 31083 5268
rect 30665 5259 30708 5265
rect 30668 5256 30708 5259
rect 31583 5263 31729 5270
rect 31065 5247 31105 5248
rect 30776 5230 31105 5247
rect 31583 5243 31639 5263
rect 31659 5243 31698 5263
rect 31718 5243 31729 5263
rect 31583 5235 31729 5243
rect 31796 5266 31953 5273
rect 31796 5246 31916 5266
rect 31936 5246 31953 5266
rect 31796 5236 31953 5246
rect 31796 5235 31831 5236
rect 30660 5187 30703 5198
rect 30660 5169 30672 5187
rect 30690 5169 30703 5187
rect 30660 5143 30703 5169
rect 30776 5143 30803 5230
rect 31065 5221 31105 5230
rect 29839 5117 30278 5135
rect 28907 5116 28948 5117
rect 28641 5063 28678 5064
rect 28337 5054 28472 5063
rect 28337 5034 28443 5054
rect 28463 5034 28472 5054
rect 28337 5027 28472 5034
rect 28530 5054 28678 5063
rect 28530 5034 28539 5054
rect 28559 5034 28649 5054
rect 28669 5034 28678 5054
rect 28337 5025 28430 5027
rect 28530 5024 28678 5034
rect 28737 5054 28774 5064
rect 28737 5034 28745 5054
rect 28765 5034 28774 5054
rect 28586 5023 28622 5024
rect 28434 4964 28471 4965
rect 28737 4964 28774 5034
rect 28809 5063 28840 5114
rect 29839 5099 30239 5117
rect 30257 5099 30278 5117
rect 29839 5093 30278 5099
rect 29845 5089 30278 5093
rect 30660 5122 30803 5143
rect 30847 5195 30881 5211
rect 31065 5201 31458 5221
rect 31478 5201 31481 5221
rect 31796 5214 31827 5235
rect 32014 5214 32050 5324
rect 32069 5323 32106 5324
rect 32165 5323 32202 5324
rect 32125 5264 32215 5270
rect 32125 5244 32134 5264
rect 32154 5262 32215 5264
rect 32154 5244 32179 5262
rect 32125 5242 32179 5244
rect 32199 5242 32215 5262
rect 32125 5236 32215 5242
rect 31639 5213 31676 5214
rect 31065 5196 31481 5201
rect 31638 5204 31676 5213
rect 31065 5195 31406 5196
rect 30847 5125 30884 5195
rect 30999 5135 31030 5136
rect 30660 5120 30797 5122
rect 30224 5087 30276 5089
rect 30660 5078 30703 5120
rect 30847 5105 30856 5125
rect 30876 5105 30884 5125
rect 30847 5095 30884 5105
rect 30943 5125 31030 5135
rect 30943 5105 30952 5125
rect 30972 5105 31030 5125
rect 30943 5096 31030 5105
rect 30943 5095 30980 5096
rect 30658 5068 30703 5078
rect 28859 5063 28896 5064
rect 28809 5054 28896 5063
rect 28809 5034 28867 5054
rect 28887 5034 28896 5054
rect 28809 5024 28896 5034
rect 28955 5054 28992 5064
rect 28955 5034 28963 5054
rect 28983 5034 28992 5054
rect 30658 5050 30667 5068
rect 30685 5050 30703 5068
rect 30658 5044 30703 5050
rect 30999 5045 31030 5096
rect 31065 5125 31102 5195
rect 31368 5194 31405 5195
rect 31638 5184 31647 5204
rect 31667 5184 31676 5204
rect 31638 5176 31676 5184
rect 31742 5208 31827 5214
rect 31857 5213 31894 5214
rect 31742 5188 31750 5208
rect 31770 5188 31827 5208
rect 31742 5180 31827 5188
rect 31856 5204 31894 5213
rect 31856 5184 31865 5204
rect 31885 5184 31894 5204
rect 31742 5179 31778 5180
rect 31856 5176 31894 5184
rect 31960 5208 32104 5214
rect 31960 5188 31968 5208
rect 31988 5205 32076 5208
rect 31988 5188 32023 5205
rect 31960 5187 32023 5188
rect 32042 5188 32076 5205
rect 32096 5188 32104 5208
rect 32042 5187 32104 5188
rect 31960 5180 32104 5187
rect 31960 5179 31996 5180
rect 32068 5179 32104 5180
rect 32170 5213 32207 5214
rect 32170 5212 32208 5213
rect 32230 5212 32257 5216
rect 32170 5210 32257 5212
rect 32170 5204 32234 5210
rect 32170 5184 32179 5204
rect 32199 5190 32234 5204
rect 32254 5190 32257 5210
rect 32199 5185 32257 5190
rect 32199 5184 32234 5185
rect 31639 5147 31676 5176
rect 31640 5145 31676 5147
rect 31217 5135 31253 5136
rect 31065 5105 31074 5125
rect 31094 5105 31102 5125
rect 31065 5095 31102 5105
rect 31161 5125 31309 5135
rect 31409 5132 31505 5134
rect 31161 5105 31170 5125
rect 31190 5105 31280 5125
rect 31300 5105 31309 5125
rect 31161 5096 31309 5105
rect 31367 5125 31505 5132
rect 31367 5105 31376 5125
rect 31396 5105 31505 5125
rect 31640 5123 31831 5145
rect 31857 5144 31894 5176
rect 32170 5172 32234 5184
rect 32274 5146 32301 5324
rect 32133 5144 32301 5146
rect 31857 5118 32301 5144
rect 31367 5096 31505 5105
rect 31161 5095 31198 5096
rect 30658 5041 30695 5044
rect 30891 5042 30932 5043
rect 28809 5023 28840 5024
rect 28433 4963 28774 4964
rect 28955 4963 28992 5034
rect 30783 5035 30932 5042
rect 30227 5022 30264 5027
rect 28358 4958 28774 4963
rect 28358 4938 28361 4958
rect 28381 4938 28774 4958
rect 28805 4939 28992 4963
rect 30218 5018 30265 5022
rect 30218 5000 30237 5018
rect 30255 5000 30265 5018
rect 30783 5015 30842 5035
rect 30862 5015 30901 5035
rect 30921 5015 30932 5035
rect 30783 5007 30932 5015
rect 30999 5038 31156 5045
rect 30999 5018 31119 5038
rect 31139 5018 31156 5038
rect 30999 5008 31156 5018
rect 30999 5007 31034 5008
rect 29826 4941 29864 4942
rect 30218 4941 30265 5000
rect 30999 4986 31030 5007
rect 31217 4986 31253 5096
rect 31272 5095 31309 5096
rect 31368 5095 31405 5096
rect 31328 5036 31418 5042
rect 31328 5016 31337 5036
rect 31357 5034 31418 5036
rect 31357 5016 31382 5034
rect 31328 5014 31382 5016
rect 31402 5014 31418 5034
rect 31328 5008 31418 5014
rect 30842 4985 30879 4986
rect 30655 4977 30692 4979
rect 30655 4969 30697 4977
rect 30655 4951 30665 4969
rect 30683 4951 30697 4969
rect 30655 4942 30697 4951
rect 30841 4976 30879 4985
rect 30841 4956 30850 4976
rect 30870 4956 30879 4976
rect 30841 4948 30879 4956
rect 30945 4980 31030 4986
rect 31060 4985 31097 4986
rect 30945 4960 30953 4980
rect 30973 4960 31030 4980
rect 30945 4952 31030 4960
rect 31059 4976 31097 4985
rect 31059 4956 31068 4976
rect 31088 4956 31097 4976
rect 30945 4951 30981 4952
rect 31059 4948 31097 4956
rect 31163 4984 31307 4986
rect 31163 4980 31215 4984
rect 31163 4960 31171 4980
rect 31191 4964 31215 4980
rect 31235 4980 31307 4984
rect 31235 4964 31279 4980
rect 31191 4960 31279 4964
rect 31299 4960 31307 4980
rect 31163 4952 31307 4960
rect 31163 4951 31199 4952
rect 31271 4951 31307 4952
rect 31373 4985 31410 4986
rect 31373 4984 31411 4985
rect 31373 4976 31437 4984
rect 31373 4956 31382 4976
rect 31402 4962 31437 4976
rect 31457 4962 31460 4982
rect 31402 4957 31460 4962
rect 31402 4956 31437 4957
rect 28578 4937 28643 4938
rect 26693 4859 26731 4860
rect 26292 4821 26731 4859
rect 27603 4859 27611 4881
rect 27635 4859 27643 4881
rect 27603 4851 27643 4859
rect 28914 4903 28954 4911
rect 28914 4881 28922 4903
rect 28946 4881 28954 4903
rect 29826 4903 30265 4941
rect 29826 4902 29864 4903
rect 27914 4824 27979 4825
rect 25107 4806 25142 4807
rect 25084 4801 25142 4806
rect 25084 4781 25087 4801
rect 25107 4787 25142 4801
rect 25162 4787 25171 4807
rect 25107 4779 25171 4787
rect 25133 4778 25171 4779
rect 25134 4777 25171 4778
rect 25237 4811 25273 4812
rect 25345 4811 25381 4812
rect 25237 4803 25381 4811
rect 25237 4783 25245 4803
rect 25265 4799 25353 4803
rect 25265 4783 25309 4799
rect 25237 4779 25309 4783
rect 25329 4783 25353 4799
rect 25373 4783 25381 4803
rect 25329 4779 25381 4783
rect 25237 4777 25381 4779
rect 25447 4807 25485 4815
rect 25563 4811 25599 4812
rect 25447 4787 25456 4807
rect 25476 4787 25485 4807
rect 25447 4778 25485 4787
rect 25514 4803 25599 4811
rect 25514 4783 25571 4803
rect 25591 4783 25599 4803
rect 25447 4777 25484 4778
rect 25514 4777 25599 4783
rect 25665 4807 25703 4815
rect 25665 4787 25674 4807
rect 25694 4787 25703 4807
rect 25665 4778 25703 4787
rect 25847 4812 25889 4821
rect 25847 4794 25861 4812
rect 25879 4794 25889 4812
rect 25847 4786 25889 4794
rect 25852 4784 25889 4786
rect 25665 4777 25702 4778
rect 25126 4749 25216 4755
rect 25126 4729 25142 4749
rect 25162 4747 25216 4749
rect 25162 4729 25187 4747
rect 25126 4727 25187 4729
rect 25207 4727 25216 4747
rect 25126 4721 25216 4727
rect 25139 4667 25176 4668
rect 25235 4667 25272 4668
rect 25291 4667 25327 4777
rect 25514 4756 25545 4777
rect 26292 4762 26339 4821
rect 26693 4820 26731 4821
rect 25510 4755 25545 4756
rect 25388 4745 25545 4755
rect 25388 4725 25405 4745
rect 25425 4725 25545 4745
rect 25388 4718 25545 4725
rect 25612 4748 25761 4756
rect 25612 4728 25623 4748
rect 25643 4728 25682 4748
rect 25702 4728 25761 4748
rect 26292 4744 26302 4762
rect 26320 4744 26339 4762
rect 26292 4740 26339 4744
rect 27565 4799 27752 4823
rect 27783 4804 28176 4824
rect 28196 4804 28199 4824
rect 27783 4799 28199 4804
rect 26293 4735 26330 4740
rect 25612 4721 25761 4728
rect 27565 4728 27602 4799
rect 27783 4798 28124 4799
rect 27717 4738 27748 4739
rect 25612 4720 25653 4721
rect 25849 4719 25886 4722
rect 25346 4667 25383 4668
rect 25039 4658 25177 4667
rect 24243 4619 24687 4645
rect 24243 4617 24411 4619
rect 24243 4439 24270 4617
rect 24310 4579 24374 4591
rect 24650 4587 24687 4619
rect 24713 4618 24904 4640
rect 25039 4638 25148 4658
rect 25168 4638 25177 4658
rect 25039 4631 25177 4638
rect 25235 4658 25383 4667
rect 25235 4638 25244 4658
rect 25264 4638 25354 4658
rect 25374 4638 25383 4658
rect 25039 4629 25135 4631
rect 25235 4628 25383 4638
rect 25442 4658 25479 4668
rect 25442 4638 25450 4658
rect 25470 4638 25479 4658
rect 25291 4627 25327 4628
rect 24868 4616 24904 4618
rect 24868 4587 24905 4616
rect 24310 4578 24345 4579
rect 24287 4573 24345 4578
rect 24287 4553 24290 4573
rect 24310 4559 24345 4573
rect 24365 4559 24374 4579
rect 24310 4553 24374 4559
rect 24287 4551 24374 4553
rect 24287 4547 24314 4551
rect 24336 4550 24374 4551
rect 24337 4549 24374 4550
rect 24440 4583 24476 4584
rect 24548 4583 24584 4584
rect 24440 4576 24584 4583
rect 24440 4575 24502 4576
rect 24440 4555 24448 4575
rect 24468 4558 24502 4575
rect 24521 4575 24584 4576
rect 24521 4558 24556 4575
rect 24468 4555 24556 4558
rect 24576 4555 24584 4575
rect 24440 4549 24584 4555
rect 24650 4579 24688 4587
rect 24766 4583 24802 4584
rect 24650 4559 24659 4579
rect 24679 4559 24688 4579
rect 24650 4550 24688 4559
rect 24717 4575 24802 4583
rect 24717 4555 24774 4575
rect 24794 4555 24802 4575
rect 24650 4549 24687 4550
rect 24717 4549 24802 4555
rect 24868 4579 24906 4587
rect 24868 4559 24877 4579
rect 24897 4559 24906 4579
rect 25139 4568 25176 4569
rect 25442 4568 25479 4638
rect 25514 4667 25545 4718
rect 25841 4713 25886 4719
rect 25841 4695 25859 4713
rect 25877 4695 25886 4713
rect 27565 4708 27574 4728
rect 27594 4708 27602 4728
rect 27565 4698 27602 4708
rect 27661 4728 27748 4738
rect 27661 4708 27670 4728
rect 27690 4708 27748 4728
rect 27661 4699 27748 4708
rect 27661 4698 27698 4699
rect 25841 4685 25886 4695
rect 25564 4667 25601 4668
rect 25514 4658 25601 4667
rect 25514 4638 25572 4658
rect 25592 4638 25601 4658
rect 25514 4628 25601 4638
rect 25660 4658 25697 4668
rect 25660 4638 25668 4658
rect 25688 4638 25697 4658
rect 25841 4643 25884 4685
rect 26281 4673 26333 4675
rect 25747 4641 25884 4643
rect 25514 4627 25545 4628
rect 25660 4568 25697 4638
rect 25138 4567 25479 4568
rect 24868 4550 24906 4559
rect 25063 4562 25479 4567
rect 24868 4549 24905 4550
rect 24329 4521 24419 4527
rect 24329 4501 24345 4521
rect 24365 4519 24419 4521
rect 24365 4501 24390 4519
rect 24329 4499 24390 4501
rect 24410 4499 24419 4519
rect 24329 4493 24419 4499
rect 24342 4439 24379 4440
rect 24438 4439 24475 4440
rect 24494 4439 24530 4549
rect 24717 4528 24748 4549
rect 25063 4542 25066 4562
rect 25086 4542 25479 4562
rect 25663 4552 25697 4568
rect 25741 4620 25884 4641
rect 26279 4669 26712 4673
rect 26279 4663 26718 4669
rect 26279 4645 26300 4663
rect 26318 4645 26718 4663
rect 27717 4648 27748 4699
rect 27783 4728 27820 4798
rect 28086 4797 28123 4798
rect 27935 4738 27971 4739
rect 27783 4708 27792 4728
rect 27812 4708 27820 4728
rect 27783 4698 27820 4708
rect 27879 4728 28027 4738
rect 28127 4735 28223 4737
rect 27879 4708 27888 4728
rect 27908 4708 27998 4728
rect 28018 4708 28027 4728
rect 27879 4699 28027 4708
rect 28085 4728 28223 4735
rect 28085 4708 28094 4728
rect 28114 4708 28223 4728
rect 28085 4699 28223 4708
rect 27879 4698 27916 4699
rect 27609 4645 27650 4646
rect 26279 4627 26718 4645
rect 25439 4533 25479 4542
rect 25741 4533 25768 4620
rect 25841 4594 25884 4620
rect 25841 4576 25854 4594
rect 25872 4576 25884 4594
rect 25841 4565 25884 4576
rect 24713 4527 24748 4528
rect 24591 4517 24748 4527
rect 24591 4497 24608 4517
rect 24628 4497 24748 4517
rect 24591 4490 24748 4497
rect 24815 4520 24961 4528
rect 24815 4500 24826 4520
rect 24846 4500 24885 4520
rect 24905 4500 24961 4520
rect 25439 4516 25768 4533
rect 25439 4515 25479 4516
rect 24815 4493 24961 4500
rect 25836 4504 25876 4507
rect 25836 4498 25879 4504
rect 25461 4495 25879 4498
rect 24815 4492 24856 4493
rect 24549 4439 24586 4440
rect 24242 4430 24380 4439
rect 24242 4410 24351 4430
rect 24371 4410 24380 4430
rect 24242 4403 24380 4410
rect 24438 4430 24586 4439
rect 24438 4410 24447 4430
rect 24467 4410 24557 4430
rect 24577 4410 24586 4430
rect 24242 4401 24338 4403
rect 24438 4400 24586 4410
rect 24645 4430 24682 4440
rect 24645 4410 24653 4430
rect 24673 4410 24682 4430
rect 24494 4399 24530 4400
rect 24342 4340 24379 4341
rect 24645 4340 24682 4410
rect 24717 4439 24748 4490
rect 25461 4477 25852 4495
rect 25870 4477 25879 4495
rect 25461 4475 25879 4477
rect 25461 4467 25488 4475
rect 25729 4472 25879 4475
rect 25041 4461 25209 4462
rect 25460 4461 25488 4467
rect 25041 4445 25488 4461
rect 25836 4467 25879 4472
rect 24767 4439 24804 4440
rect 24717 4430 24804 4439
rect 24717 4410 24775 4430
rect 24795 4410 24804 4430
rect 24717 4400 24804 4410
rect 24863 4430 24900 4440
rect 24863 4410 24871 4430
rect 24891 4410 24900 4430
rect 24717 4399 24748 4400
rect 24341 4339 24682 4340
rect 24863 4339 24900 4410
rect 24266 4334 24682 4339
rect 24266 4314 24269 4334
rect 24289 4314 24682 4334
rect 24713 4315 24900 4339
rect 25041 4435 25485 4445
rect 25041 4433 25209 4435
rect 24075 4240 24119 4241
rect 24075 4234 24120 4240
rect 24075 4216 24087 4234
rect 24109 4216 24120 4234
rect 24141 4235 24183 4280
rect 25041 4255 25068 4433
rect 25108 4395 25172 4407
rect 25448 4403 25485 4435
rect 25511 4434 25702 4456
rect 25666 4432 25702 4434
rect 25666 4403 25703 4432
rect 25836 4411 25876 4467
rect 25108 4394 25143 4395
rect 25085 4389 25143 4394
rect 25085 4369 25088 4389
rect 25108 4375 25143 4389
rect 25163 4375 25172 4395
rect 25108 4367 25172 4375
rect 25134 4366 25172 4367
rect 25135 4365 25172 4366
rect 25238 4399 25274 4400
rect 25346 4399 25382 4400
rect 25238 4391 25382 4399
rect 25238 4371 25246 4391
rect 25266 4371 25301 4391
rect 25321 4371 25354 4391
rect 25374 4371 25382 4391
rect 25238 4365 25382 4371
rect 25448 4395 25486 4403
rect 25564 4399 25600 4400
rect 25448 4375 25457 4395
rect 25477 4375 25486 4395
rect 25448 4366 25486 4375
rect 25515 4391 25600 4399
rect 25515 4371 25572 4391
rect 25592 4371 25600 4391
rect 25448 4365 25485 4366
rect 25515 4365 25600 4371
rect 25666 4395 25704 4403
rect 25666 4375 25675 4395
rect 25695 4375 25704 4395
rect 25836 4393 25848 4411
rect 25866 4393 25876 4411
rect 26281 4438 26333 4627
rect 26679 4602 26718 4627
rect 27501 4638 27650 4645
rect 27501 4618 27560 4638
rect 27580 4618 27619 4638
rect 27639 4618 27650 4638
rect 27501 4610 27650 4618
rect 27717 4641 27874 4648
rect 27717 4621 27837 4641
rect 27857 4621 27874 4641
rect 27717 4611 27874 4621
rect 27717 4610 27752 4611
rect 26463 4577 26650 4601
rect 26679 4582 27074 4602
rect 27094 4582 27097 4602
rect 27717 4589 27748 4610
rect 27935 4589 27971 4699
rect 27990 4698 28027 4699
rect 28086 4698 28123 4699
rect 28046 4639 28136 4645
rect 28046 4619 28055 4639
rect 28075 4637 28136 4639
rect 28075 4619 28100 4637
rect 28046 4617 28100 4619
rect 28120 4617 28136 4637
rect 28046 4611 28136 4617
rect 27560 4588 27597 4589
rect 26679 4577 27097 4582
rect 27559 4579 27597 4588
rect 26463 4506 26500 4577
rect 26679 4576 27022 4577
rect 26679 4573 26718 4576
rect 26984 4575 27021 4576
rect 26615 4516 26646 4517
rect 26463 4486 26472 4506
rect 26492 4486 26500 4506
rect 26463 4476 26500 4486
rect 26559 4506 26646 4516
rect 26559 4486 26568 4506
rect 26588 4486 26646 4506
rect 26559 4477 26646 4486
rect 26559 4476 26596 4477
rect 26281 4420 26297 4438
rect 26315 4420 26333 4438
rect 26615 4426 26646 4477
rect 26681 4506 26718 4573
rect 27559 4559 27568 4579
rect 27588 4559 27597 4579
rect 27559 4551 27597 4559
rect 27663 4583 27748 4589
rect 27778 4588 27815 4589
rect 27663 4563 27671 4583
rect 27691 4563 27748 4583
rect 27663 4555 27748 4563
rect 27777 4579 27815 4588
rect 27777 4559 27786 4579
rect 27806 4559 27815 4579
rect 27663 4554 27699 4555
rect 27777 4551 27815 4559
rect 27881 4583 28025 4589
rect 27881 4563 27889 4583
rect 27909 4577 27997 4583
rect 27909 4563 27938 4577
rect 27881 4555 27938 4563
rect 27881 4554 27917 4555
rect 27961 4563 27997 4577
rect 28017 4563 28025 4583
rect 27961 4555 28025 4563
rect 27989 4554 28025 4555
rect 28091 4588 28128 4589
rect 28091 4587 28129 4588
rect 28091 4579 28155 4587
rect 28091 4559 28100 4579
rect 28120 4565 28155 4579
rect 28175 4565 28178 4585
rect 28120 4560 28178 4565
rect 28120 4559 28155 4560
rect 27560 4522 27597 4551
rect 27561 4520 27597 4522
rect 26833 4516 26869 4517
rect 26681 4486 26690 4506
rect 26710 4486 26718 4506
rect 26681 4476 26718 4486
rect 26777 4506 26925 4516
rect 27025 4513 27121 4515
rect 26777 4486 26786 4506
rect 26806 4486 26896 4506
rect 26916 4486 26925 4506
rect 26777 4477 26925 4486
rect 26983 4506 27121 4513
rect 26983 4486 26992 4506
rect 27012 4486 27121 4506
rect 27561 4498 27752 4520
rect 27778 4519 27815 4551
rect 28091 4547 28155 4559
rect 28195 4521 28222 4699
rect 28519 4652 28556 4658
rect 28519 4633 28527 4652
rect 28548 4633 28556 4652
rect 28519 4625 28556 4633
rect 28054 4519 28222 4521
rect 27778 4493 28222 4519
rect 27888 4491 27928 4493
rect 28054 4492 28222 4493
rect 26983 4477 27121 4486
rect 28181 4487 28222 4492
rect 26777 4476 26814 4477
rect 26507 4423 26548 4424
rect 26281 4402 26333 4420
rect 26399 4416 26548 4423
rect 25836 4383 25876 4393
rect 26399 4396 26458 4416
rect 26478 4396 26517 4416
rect 26537 4396 26548 4416
rect 26399 4388 26548 4396
rect 26615 4419 26772 4426
rect 26615 4399 26735 4419
rect 26755 4399 26772 4419
rect 26615 4389 26772 4399
rect 26615 4388 26650 4389
rect 25666 4366 25704 4375
rect 26615 4367 26646 4388
rect 26833 4367 26869 4477
rect 26888 4476 26925 4477
rect 26984 4476 27021 4477
rect 26944 4417 27034 4423
rect 26944 4397 26953 4417
rect 26973 4415 27034 4417
rect 26973 4397 26998 4415
rect 26944 4395 26998 4397
rect 27018 4395 27034 4415
rect 26944 4389 27034 4395
rect 26458 4366 26495 4367
rect 25666 4365 25703 4366
rect 25127 4337 25217 4343
rect 25127 4317 25143 4337
rect 25163 4335 25217 4337
rect 25163 4317 25188 4335
rect 25127 4315 25188 4317
rect 25208 4315 25217 4335
rect 25127 4309 25217 4315
rect 25140 4255 25177 4256
rect 25236 4255 25273 4256
rect 25292 4255 25328 4365
rect 25515 4344 25546 4365
rect 26457 4357 26495 4366
rect 25511 4343 25546 4344
rect 25389 4333 25546 4343
rect 25389 4313 25406 4333
rect 25426 4313 25546 4333
rect 25389 4306 25546 4313
rect 25613 4336 25762 4344
rect 25613 4316 25624 4336
rect 25644 4316 25683 4336
rect 25703 4316 25762 4336
rect 26285 4339 26325 4349
rect 25613 4309 25762 4316
rect 25828 4312 25880 4330
rect 25613 4308 25654 4309
rect 25347 4255 25384 4256
rect 25040 4246 25178 4255
rect 24512 4235 24545 4237
rect 24141 4223 24588 4235
rect 24075 4186 24120 4216
rect 24092 3240 24120 4186
rect 24144 4209 24588 4223
rect 24144 4207 24312 4209
rect 24144 4029 24171 4207
rect 24211 4169 24275 4181
rect 24551 4177 24588 4209
rect 24614 4208 24805 4230
rect 25040 4226 25149 4246
rect 25169 4226 25178 4246
rect 25040 4219 25178 4226
rect 25236 4246 25384 4255
rect 25236 4226 25245 4246
rect 25265 4226 25355 4246
rect 25375 4226 25384 4246
rect 25040 4217 25136 4219
rect 25236 4216 25384 4226
rect 25443 4246 25480 4256
rect 25443 4226 25451 4246
rect 25471 4226 25480 4246
rect 25292 4215 25328 4216
rect 24769 4206 24805 4208
rect 24769 4177 24806 4206
rect 24211 4168 24246 4169
rect 24188 4163 24246 4168
rect 24188 4143 24191 4163
rect 24211 4149 24246 4163
rect 24266 4149 24275 4169
rect 24211 4141 24275 4149
rect 24237 4140 24275 4141
rect 24238 4139 24275 4140
rect 24341 4173 24377 4174
rect 24449 4173 24485 4174
rect 24341 4167 24485 4173
rect 24341 4165 24402 4167
rect 24341 4145 24349 4165
rect 24369 4150 24402 4165
rect 24421 4165 24485 4167
rect 24421 4150 24457 4165
rect 24369 4145 24457 4150
rect 24477 4145 24485 4165
rect 24341 4139 24485 4145
rect 24551 4169 24589 4177
rect 24667 4173 24703 4174
rect 24551 4149 24560 4169
rect 24580 4149 24589 4169
rect 24551 4140 24589 4149
rect 24618 4165 24703 4173
rect 24618 4145 24675 4165
rect 24695 4145 24703 4165
rect 24551 4139 24588 4140
rect 24618 4139 24703 4145
rect 24769 4169 24807 4177
rect 24769 4149 24778 4169
rect 24798 4149 24807 4169
rect 25443 4159 25480 4226
rect 25515 4255 25546 4306
rect 25828 4294 25846 4312
rect 25864 4294 25880 4312
rect 25565 4255 25602 4256
rect 25515 4246 25602 4255
rect 25515 4226 25573 4246
rect 25593 4226 25602 4246
rect 25515 4216 25602 4226
rect 25661 4246 25698 4256
rect 25661 4226 25669 4246
rect 25689 4226 25698 4246
rect 25515 4215 25546 4216
rect 25140 4156 25177 4157
rect 25443 4156 25482 4159
rect 25139 4155 25482 4156
rect 25661 4155 25698 4226
rect 24769 4140 24807 4149
rect 25064 4150 25482 4155
rect 24769 4139 24806 4140
rect 24230 4111 24320 4117
rect 24230 4091 24246 4111
rect 24266 4109 24320 4111
rect 24266 4091 24291 4109
rect 24230 4089 24291 4091
rect 24311 4089 24320 4109
rect 24230 4083 24320 4089
rect 24243 4029 24280 4030
rect 24339 4029 24376 4030
rect 24395 4029 24431 4139
rect 24618 4118 24649 4139
rect 25064 4130 25067 4150
rect 25087 4130 25482 4150
rect 25511 4131 25698 4155
rect 24614 4117 24649 4118
rect 24492 4107 24649 4117
rect 24492 4087 24509 4107
rect 24529 4087 24649 4107
rect 24492 4080 24649 4087
rect 24716 4110 24865 4118
rect 24716 4090 24727 4110
rect 24747 4090 24786 4110
rect 24806 4090 24865 4110
rect 24716 4083 24865 4090
rect 25443 4105 25482 4130
rect 25828 4105 25880 4294
rect 26285 4321 26295 4339
rect 26313 4321 26325 4339
rect 26457 4337 26466 4357
rect 26486 4337 26495 4357
rect 26457 4329 26495 4337
rect 26561 4361 26646 4367
rect 26676 4366 26713 4367
rect 26561 4341 26569 4361
rect 26589 4341 26646 4361
rect 26561 4333 26646 4341
rect 26675 4357 26713 4366
rect 26675 4337 26684 4357
rect 26704 4337 26713 4357
rect 26561 4332 26597 4333
rect 26675 4329 26713 4337
rect 26779 4361 26923 4367
rect 26779 4341 26787 4361
rect 26807 4341 26840 4361
rect 26860 4341 26895 4361
rect 26915 4341 26923 4361
rect 26779 4333 26923 4341
rect 26779 4332 26815 4333
rect 26887 4332 26923 4333
rect 26989 4366 27026 4367
rect 26989 4365 27027 4366
rect 26989 4357 27053 4365
rect 26989 4337 26998 4357
rect 27018 4343 27053 4357
rect 27073 4343 27076 4363
rect 27018 4338 27076 4343
rect 27018 4337 27053 4338
rect 26285 4265 26325 4321
rect 26458 4300 26495 4329
rect 26459 4298 26495 4300
rect 26459 4276 26650 4298
rect 26676 4297 26713 4329
rect 26989 4325 27053 4337
rect 27093 4299 27120 4477
rect 26952 4297 27120 4299
rect 26676 4287 27120 4297
rect 27261 4393 27448 4417
rect 27479 4398 27872 4418
rect 27892 4398 27895 4418
rect 27479 4393 27895 4398
rect 27261 4322 27298 4393
rect 27479 4392 27820 4393
rect 27413 4332 27444 4333
rect 27261 4302 27270 4322
rect 27290 4302 27298 4322
rect 27261 4292 27298 4302
rect 27357 4322 27444 4332
rect 27357 4302 27366 4322
rect 27386 4302 27444 4322
rect 27357 4293 27444 4302
rect 27357 4292 27394 4293
rect 26282 4260 26325 4265
rect 26673 4271 27120 4287
rect 26673 4265 26701 4271
rect 26952 4270 27120 4271
rect 26282 4257 26432 4260
rect 26673 4257 26700 4265
rect 26282 4255 26700 4257
rect 26282 4237 26291 4255
rect 26309 4237 26700 4255
rect 27413 4242 27444 4293
rect 27479 4322 27516 4392
rect 27782 4391 27819 4392
rect 27631 4332 27667 4333
rect 27479 4302 27488 4322
rect 27508 4302 27516 4322
rect 27479 4292 27516 4302
rect 27575 4322 27723 4332
rect 27823 4329 27919 4331
rect 27575 4302 27584 4322
rect 27604 4302 27694 4322
rect 27714 4302 27723 4322
rect 27575 4293 27723 4302
rect 27781 4322 27919 4329
rect 27781 4302 27790 4322
rect 27810 4302 27919 4322
rect 28181 4305 28221 4487
rect 27781 4293 27919 4302
rect 27575 4292 27612 4293
rect 27305 4239 27346 4240
rect 26282 4234 26700 4237
rect 26282 4228 26325 4234
rect 26285 4225 26325 4228
rect 27197 4232 27346 4239
rect 26682 4216 26722 4217
rect 26393 4199 26722 4216
rect 27197 4212 27256 4232
rect 27276 4212 27315 4232
rect 27335 4212 27346 4232
rect 27197 4204 27346 4212
rect 27413 4235 27570 4242
rect 27413 4215 27533 4235
rect 27553 4215 27570 4235
rect 27413 4205 27570 4215
rect 27413 4204 27448 4205
rect 26277 4156 26320 4167
rect 26277 4138 26289 4156
rect 26307 4138 26320 4156
rect 26277 4112 26320 4138
rect 26393 4112 26420 4199
rect 26682 4190 26722 4199
rect 25443 4087 25882 4105
rect 24716 4082 24757 4083
rect 24450 4029 24487 4030
rect 24143 4020 24281 4029
rect 24143 4000 24252 4020
rect 24272 4000 24281 4020
rect 24143 3993 24281 4000
rect 24339 4020 24487 4029
rect 24339 4000 24348 4020
rect 24368 4000 24458 4020
rect 24478 4000 24487 4020
rect 24143 3991 24239 3993
rect 24339 3990 24487 4000
rect 24546 4020 24583 4030
rect 24546 4000 24554 4020
rect 24574 4000 24583 4020
rect 24395 3989 24431 3990
rect 24243 3930 24280 3931
rect 24546 3930 24583 4000
rect 24618 4029 24649 4080
rect 25443 4069 25843 4087
rect 25861 4069 25882 4087
rect 25443 4063 25882 4069
rect 25449 4059 25882 4063
rect 26277 4091 26420 4112
rect 26464 4164 26498 4180
rect 26682 4170 27075 4190
rect 27095 4170 27098 4190
rect 27413 4183 27444 4204
rect 27631 4183 27667 4293
rect 27686 4292 27723 4293
rect 27782 4292 27819 4293
rect 27742 4233 27832 4239
rect 27742 4213 27751 4233
rect 27771 4231 27832 4233
rect 27771 4213 27796 4231
rect 27742 4211 27796 4213
rect 27816 4211 27832 4231
rect 27742 4205 27832 4211
rect 27256 4182 27293 4183
rect 26682 4165 27098 4170
rect 27255 4173 27293 4182
rect 26682 4164 27023 4165
rect 26464 4094 26501 4164
rect 26616 4104 26647 4105
rect 26277 4089 26414 4091
rect 25828 4057 25880 4059
rect 26277 4047 26320 4089
rect 26464 4074 26473 4094
rect 26493 4074 26501 4094
rect 26464 4064 26501 4074
rect 26560 4094 26647 4104
rect 26560 4074 26569 4094
rect 26589 4074 26647 4094
rect 26560 4065 26647 4074
rect 26560 4064 26597 4065
rect 26275 4037 26320 4047
rect 24668 4029 24705 4030
rect 24618 4020 24705 4029
rect 24618 4000 24676 4020
rect 24696 4000 24705 4020
rect 24618 3990 24705 4000
rect 24764 4020 24801 4030
rect 24764 4000 24772 4020
rect 24792 4000 24801 4020
rect 26275 4019 26284 4037
rect 26302 4019 26320 4037
rect 26275 4013 26320 4019
rect 26616 4014 26647 4065
rect 26682 4094 26719 4164
rect 26985 4163 27022 4164
rect 27255 4153 27264 4173
rect 27284 4153 27293 4173
rect 27255 4145 27293 4153
rect 27359 4177 27444 4183
rect 27474 4182 27511 4183
rect 27359 4157 27367 4177
rect 27387 4157 27444 4177
rect 27359 4149 27444 4157
rect 27473 4173 27511 4182
rect 27473 4153 27482 4173
rect 27502 4153 27511 4173
rect 27359 4148 27395 4149
rect 27473 4145 27511 4153
rect 27577 4177 27721 4183
rect 27577 4157 27585 4177
rect 27605 4158 27637 4177
rect 27658 4158 27693 4177
rect 27605 4157 27693 4158
rect 27713 4157 27721 4177
rect 27577 4149 27721 4157
rect 27577 4148 27613 4149
rect 27685 4148 27721 4149
rect 27787 4182 27824 4183
rect 27787 4181 27825 4182
rect 27787 4173 27851 4181
rect 27787 4153 27796 4173
rect 27816 4159 27851 4173
rect 27871 4159 27874 4179
rect 27816 4154 27874 4159
rect 27816 4153 27851 4154
rect 27256 4116 27293 4145
rect 27257 4114 27293 4116
rect 26834 4104 26870 4105
rect 26682 4074 26691 4094
rect 26711 4074 26719 4094
rect 26682 4064 26719 4074
rect 26778 4094 26926 4104
rect 27026 4101 27122 4103
rect 26778 4074 26787 4094
rect 26807 4074 26897 4094
rect 26917 4074 26926 4094
rect 26778 4065 26926 4074
rect 26984 4094 27122 4101
rect 26984 4074 26993 4094
rect 27013 4074 27122 4094
rect 27257 4092 27448 4114
rect 27474 4113 27511 4145
rect 27787 4141 27851 4153
rect 27891 4115 27918 4293
rect 27750 4113 27918 4115
rect 27474 4087 27918 4113
rect 26984 4065 27122 4074
rect 26778 4064 26815 4065
rect 26275 4010 26312 4013
rect 26508 4011 26549 4012
rect 24618 3989 24649 3990
rect 24242 3929 24583 3930
rect 24764 3929 24801 4000
rect 26400 4004 26549 4011
rect 25831 3992 25868 3997
rect 25822 3988 25869 3992
rect 25822 3970 25841 3988
rect 25859 3970 25869 3988
rect 26400 3984 26459 4004
rect 26479 3984 26518 4004
rect 26538 3984 26549 4004
rect 26400 3976 26549 3984
rect 26616 4007 26773 4014
rect 26616 3987 26736 4007
rect 26756 3987 26773 4007
rect 26616 3977 26773 3987
rect 26616 3976 26651 3977
rect 24167 3924 24583 3929
rect 24167 3904 24170 3924
rect 24190 3904 24583 3924
rect 24614 3905 24801 3929
rect 25426 3927 25466 3932
rect 25822 3927 25869 3970
rect 26616 3955 26647 3976
rect 26834 3955 26870 4065
rect 26889 4064 26926 4065
rect 26985 4064 27022 4065
rect 26945 4005 27035 4011
rect 26945 3985 26954 4005
rect 26974 4003 27035 4005
rect 26974 3985 26999 4003
rect 26945 3983 26999 3985
rect 27019 3983 27035 4003
rect 26945 3977 27035 3983
rect 26459 3954 26496 3955
rect 25426 3888 25869 3927
rect 26272 3946 26309 3948
rect 26272 3938 26314 3946
rect 26272 3920 26282 3938
rect 26300 3920 26314 3938
rect 26272 3911 26314 3920
rect 26458 3945 26496 3954
rect 26458 3925 26467 3945
rect 26487 3925 26496 3945
rect 26458 3917 26496 3925
rect 26562 3949 26647 3955
rect 26677 3954 26714 3955
rect 26562 3929 26570 3949
rect 26590 3929 26647 3949
rect 26562 3921 26647 3929
rect 26676 3945 26714 3954
rect 26676 3925 26685 3945
rect 26705 3925 26714 3945
rect 26562 3920 26598 3921
rect 26676 3917 26714 3925
rect 26780 3953 26924 3955
rect 26780 3949 26832 3953
rect 26780 3929 26788 3949
rect 26808 3933 26832 3949
rect 26852 3949 26924 3953
rect 26852 3933 26896 3949
rect 26808 3929 26896 3933
rect 26916 3929 26924 3949
rect 26780 3921 26924 3929
rect 26780 3920 26816 3921
rect 26888 3920 26924 3921
rect 26990 3954 27027 3955
rect 26990 3953 27028 3954
rect 26990 3945 27054 3953
rect 26990 3925 26999 3945
rect 27019 3931 27054 3945
rect 27074 3931 27077 3951
rect 27019 3926 27077 3931
rect 27019 3925 27054 3926
rect 24520 3873 24560 3881
rect 24520 3851 24528 3873
rect 24552 3851 24560 3873
rect 24226 3627 24394 3628
rect 24520 3627 24560 3851
rect 25023 3855 25191 3856
rect 25426 3855 25466 3888
rect 25822 3855 25869 3888
rect 26273 3886 26314 3911
rect 26459 3886 26496 3917
rect 26677 3886 26714 3917
rect 26990 3913 27054 3925
rect 27094 3887 27121 4065
rect 26273 3859 26322 3886
rect 26458 3860 26507 3886
rect 26676 3885 26757 3886
rect 26953 3885 27121 3887
rect 26676 3860 27121 3885
rect 26677 3859 27121 3860
rect 25023 3854 25467 3855
rect 25023 3829 25468 3854
rect 25023 3827 25191 3829
rect 25387 3828 25468 3829
rect 25637 3828 25686 3854
rect 25822 3828 25871 3855
rect 25023 3649 25050 3827
rect 25090 3789 25154 3801
rect 25430 3797 25467 3828
rect 25648 3797 25685 3828
rect 25830 3803 25871 3828
rect 26275 3826 26322 3859
rect 26678 3826 26718 3859
rect 26953 3858 27121 3859
rect 27584 3863 27624 4087
rect 27750 4086 27918 4087
rect 27584 3841 27592 3863
rect 27616 3841 27624 3863
rect 27584 3833 27624 3841
rect 25090 3788 25125 3789
rect 25067 3783 25125 3788
rect 25067 3763 25070 3783
rect 25090 3769 25125 3783
rect 25145 3769 25154 3789
rect 25090 3761 25154 3769
rect 25116 3760 25154 3761
rect 25117 3759 25154 3760
rect 25220 3793 25256 3794
rect 25328 3793 25364 3794
rect 25220 3785 25364 3793
rect 25220 3765 25228 3785
rect 25248 3781 25336 3785
rect 25248 3765 25292 3781
rect 25220 3761 25292 3765
rect 25312 3765 25336 3781
rect 25356 3765 25364 3785
rect 25312 3761 25364 3765
rect 25220 3759 25364 3761
rect 25430 3789 25468 3797
rect 25546 3793 25582 3794
rect 25430 3769 25439 3789
rect 25459 3769 25468 3789
rect 25430 3760 25468 3769
rect 25497 3785 25582 3793
rect 25497 3765 25554 3785
rect 25574 3765 25582 3785
rect 25430 3759 25467 3760
rect 25497 3759 25582 3765
rect 25648 3789 25686 3797
rect 25648 3769 25657 3789
rect 25677 3769 25686 3789
rect 25648 3760 25686 3769
rect 25830 3794 25872 3803
rect 25830 3776 25844 3794
rect 25862 3776 25872 3794
rect 25830 3768 25872 3776
rect 25835 3766 25872 3768
rect 26275 3787 26718 3826
rect 25648 3759 25685 3760
rect 25109 3731 25199 3737
rect 25109 3711 25125 3731
rect 25145 3729 25199 3731
rect 25145 3711 25170 3729
rect 25109 3709 25170 3711
rect 25190 3709 25199 3729
rect 25109 3703 25199 3709
rect 25122 3649 25159 3650
rect 25218 3649 25255 3650
rect 25274 3649 25310 3759
rect 25497 3738 25528 3759
rect 26275 3744 26322 3787
rect 26678 3782 26718 3787
rect 27343 3785 27530 3809
rect 27561 3790 27954 3810
rect 27974 3790 27977 3810
rect 27561 3785 27977 3790
rect 25493 3737 25528 3738
rect 25371 3727 25528 3737
rect 25371 3707 25388 3727
rect 25408 3707 25528 3727
rect 25371 3700 25528 3707
rect 25595 3730 25744 3738
rect 25595 3710 25606 3730
rect 25626 3710 25665 3730
rect 25685 3710 25744 3730
rect 26275 3726 26285 3744
rect 26303 3726 26322 3744
rect 26275 3722 26322 3726
rect 26276 3717 26313 3722
rect 25595 3703 25744 3710
rect 27343 3714 27380 3785
rect 27561 3784 27902 3785
rect 27495 3724 27526 3725
rect 25595 3702 25636 3703
rect 25832 3701 25869 3704
rect 25329 3649 25366 3650
rect 25022 3640 25160 3649
rect 24226 3601 24670 3627
rect 24226 3599 24394 3601
rect 24226 3421 24253 3599
rect 24293 3561 24357 3573
rect 24633 3569 24670 3601
rect 24696 3600 24887 3622
rect 25022 3620 25131 3640
rect 25151 3620 25160 3640
rect 25022 3613 25160 3620
rect 25218 3640 25366 3649
rect 25218 3620 25227 3640
rect 25247 3620 25337 3640
rect 25357 3620 25366 3640
rect 25022 3611 25118 3613
rect 25218 3610 25366 3620
rect 25425 3640 25462 3650
rect 25425 3620 25433 3640
rect 25453 3620 25462 3640
rect 25274 3609 25310 3610
rect 24851 3598 24887 3600
rect 24851 3569 24888 3598
rect 24293 3560 24328 3561
rect 24270 3555 24328 3560
rect 24270 3535 24273 3555
rect 24293 3541 24328 3555
rect 24348 3541 24357 3561
rect 24293 3533 24357 3541
rect 24319 3532 24357 3533
rect 24320 3531 24357 3532
rect 24423 3565 24459 3566
rect 24531 3565 24567 3566
rect 24423 3557 24567 3565
rect 24423 3537 24431 3557
rect 24451 3556 24539 3557
rect 24451 3537 24486 3556
rect 24507 3537 24539 3556
rect 24559 3537 24567 3557
rect 24423 3531 24567 3537
rect 24633 3561 24671 3569
rect 24749 3565 24785 3566
rect 24633 3541 24642 3561
rect 24662 3541 24671 3561
rect 24633 3532 24671 3541
rect 24700 3557 24785 3565
rect 24700 3537 24757 3557
rect 24777 3537 24785 3557
rect 24633 3531 24670 3532
rect 24700 3531 24785 3537
rect 24851 3561 24889 3569
rect 24851 3541 24860 3561
rect 24880 3541 24889 3561
rect 25122 3550 25159 3551
rect 25425 3550 25462 3620
rect 25497 3649 25528 3700
rect 25824 3695 25869 3701
rect 25824 3677 25842 3695
rect 25860 3677 25869 3695
rect 27343 3694 27352 3714
rect 27372 3694 27380 3714
rect 27343 3684 27380 3694
rect 27439 3714 27526 3724
rect 27439 3694 27448 3714
rect 27468 3694 27526 3714
rect 27439 3685 27526 3694
rect 27439 3684 27476 3685
rect 25824 3667 25869 3677
rect 25547 3649 25584 3650
rect 25497 3640 25584 3649
rect 25497 3620 25555 3640
rect 25575 3620 25584 3640
rect 25497 3610 25584 3620
rect 25643 3640 25680 3650
rect 25643 3620 25651 3640
rect 25671 3620 25680 3640
rect 25824 3625 25867 3667
rect 26264 3655 26316 3657
rect 25730 3623 25867 3625
rect 25497 3609 25528 3610
rect 25643 3550 25680 3620
rect 25121 3549 25462 3550
rect 24851 3532 24889 3541
rect 25046 3544 25462 3549
rect 24851 3531 24888 3532
rect 24312 3503 24402 3509
rect 24312 3483 24328 3503
rect 24348 3501 24402 3503
rect 24348 3483 24373 3501
rect 24312 3481 24373 3483
rect 24393 3481 24402 3501
rect 24312 3475 24402 3481
rect 24325 3421 24362 3422
rect 24421 3421 24458 3422
rect 24477 3421 24513 3531
rect 24700 3510 24731 3531
rect 25046 3524 25049 3544
rect 25069 3524 25462 3544
rect 25646 3534 25680 3550
rect 25724 3602 25867 3623
rect 26262 3651 26695 3655
rect 26262 3645 26701 3651
rect 26262 3627 26283 3645
rect 26301 3627 26701 3645
rect 27495 3634 27526 3685
rect 27561 3714 27598 3784
rect 27864 3783 27901 3784
rect 27713 3724 27749 3725
rect 27561 3694 27570 3714
rect 27590 3694 27598 3714
rect 27561 3684 27598 3694
rect 27657 3714 27805 3724
rect 27905 3721 28001 3723
rect 27657 3694 27666 3714
rect 27686 3694 27776 3714
rect 27796 3694 27805 3714
rect 27657 3685 27805 3694
rect 27863 3714 28001 3721
rect 27863 3694 27872 3714
rect 27892 3694 28001 3714
rect 27863 3685 28001 3694
rect 27657 3684 27694 3685
rect 27387 3631 27428 3632
rect 26262 3609 26701 3627
rect 25422 3515 25462 3524
rect 25724 3515 25751 3602
rect 25824 3576 25867 3602
rect 25824 3558 25837 3576
rect 25855 3558 25867 3576
rect 25824 3547 25867 3558
rect 24696 3509 24731 3510
rect 24574 3499 24731 3509
rect 24574 3479 24591 3499
rect 24611 3479 24731 3499
rect 24574 3472 24731 3479
rect 24798 3502 24947 3510
rect 24798 3482 24809 3502
rect 24829 3482 24868 3502
rect 24888 3482 24947 3502
rect 25422 3498 25751 3515
rect 25422 3497 25462 3498
rect 24798 3475 24947 3482
rect 25819 3486 25859 3489
rect 25819 3480 25862 3486
rect 25444 3477 25862 3480
rect 24798 3474 24839 3475
rect 24532 3421 24569 3422
rect 24225 3412 24363 3421
rect 24225 3392 24334 3412
rect 24354 3392 24363 3412
rect 24225 3385 24363 3392
rect 24421 3412 24569 3421
rect 24421 3392 24430 3412
rect 24450 3392 24540 3412
rect 24560 3392 24569 3412
rect 24225 3383 24321 3385
rect 24421 3382 24569 3392
rect 24628 3412 24665 3422
rect 24628 3392 24636 3412
rect 24656 3392 24665 3412
rect 24477 3381 24513 3382
rect 24325 3322 24362 3323
rect 24628 3322 24665 3392
rect 24700 3421 24731 3472
rect 25444 3459 25835 3477
rect 25853 3459 25862 3477
rect 25444 3457 25862 3459
rect 25444 3449 25471 3457
rect 25712 3454 25862 3457
rect 25024 3443 25192 3444
rect 25443 3443 25471 3449
rect 25024 3427 25471 3443
rect 25819 3449 25862 3454
rect 24750 3421 24787 3422
rect 24700 3412 24787 3421
rect 24700 3392 24758 3412
rect 24778 3392 24787 3412
rect 24700 3382 24787 3392
rect 24846 3412 24883 3422
rect 24846 3392 24854 3412
rect 24874 3392 24883 3412
rect 24700 3381 24731 3382
rect 24324 3321 24665 3322
rect 24846 3321 24883 3392
rect 24249 3316 24665 3321
rect 24249 3296 24252 3316
rect 24272 3296 24665 3316
rect 24696 3297 24883 3321
rect 25024 3417 25468 3427
rect 25024 3415 25192 3417
rect 24091 3222 24120 3240
rect 25024 3237 25051 3415
rect 25091 3377 25155 3389
rect 25431 3385 25468 3417
rect 25494 3416 25685 3438
rect 25649 3414 25685 3416
rect 25649 3385 25686 3414
rect 25819 3393 25859 3449
rect 25091 3376 25126 3377
rect 25068 3371 25126 3376
rect 25068 3351 25071 3371
rect 25091 3357 25126 3371
rect 25146 3357 25155 3377
rect 25091 3349 25155 3357
rect 25117 3348 25155 3349
rect 25118 3347 25155 3348
rect 25221 3381 25257 3382
rect 25329 3381 25365 3382
rect 25221 3373 25365 3381
rect 25221 3353 25229 3373
rect 25249 3353 25284 3373
rect 25304 3353 25337 3373
rect 25357 3353 25365 3373
rect 25221 3347 25365 3353
rect 25431 3377 25469 3385
rect 25547 3381 25583 3382
rect 25431 3357 25440 3377
rect 25460 3357 25469 3377
rect 25431 3348 25469 3357
rect 25498 3373 25583 3381
rect 25498 3353 25555 3373
rect 25575 3353 25583 3373
rect 25431 3347 25468 3348
rect 25498 3347 25583 3353
rect 25649 3377 25687 3385
rect 25649 3357 25658 3377
rect 25678 3357 25687 3377
rect 25819 3375 25831 3393
rect 25849 3375 25859 3393
rect 26264 3420 26316 3609
rect 26662 3584 26701 3609
rect 27279 3624 27428 3631
rect 27279 3604 27338 3624
rect 27358 3604 27397 3624
rect 27417 3604 27428 3624
rect 27279 3596 27428 3604
rect 27495 3627 27652 3634
rect 27495 3607 27615 3627
rect 27635 3607 27652 3627
rect 27495 3597 27652 3607
rect 27495 3596 27530 3597
rect 26446 3559 26633 3583
rect 26662 3564 27057 3584
rect 27077 3564 27080 3584
rect 27495 3575 27526 3596
rect 27713 3575 27749 3685
rect 27768 3684 27805 3685
rect 27864 3684 27901 3685
rect 27824 3625 27914 3631
rect 27824 3605 27833 3625
rect 27853 3623 27914 3625
rect 27853 3605 27878 3623
rect 27824 3603 27878 3605
rect 27898 3603 27914 3623
rect 27824 3597 27914 3603
rect 27338 3574 27375 3575
rect 26662 3559 27080 3564
rect 27337 3565 27375 3574
rect 26446 3488 26483 3559
rect 26662 3558 27005 3559
rect 26662 3555 26701 3558
rect 26967 3557 27004 3558
rect 26598 3498 26629 3499
rect 26446 3468 26455 3488
rect 26475 3468 26483 3488
rect 26446 3458 26483 3468
rect 26542 3488 26629 3498
rect 26542 3468 26551 3488
rect 26571 3468 26629 3488
rect 26542 3459 26629 3468
rect 26542 3458 26579 3459
rect 26264 3402 26280 3420
rect 26298 3402 26316 3420
rect 26598 3408 26629 3459
rect 26664 3488 26701 3555
rect 27337 3545 27346 3565
rect 27366 3545 27375 3565
rect 27337 3537 27375 3545
rect 27441 3569 27526 3575
rect 27556 3574 27593 3575
rect 27441 3549 27449 3569
rect 27469 3549 27526 3569
rect 27441 3541 27526 3549
rect 27555 3565 27593 3574
rect 27555 3545 27564 3565
rect 27584 3545 27593 3565
rect 27441 3540 27477 3541
rect 27555 3537 27593 3545
rect 27659 3570 27803 3575
rect 27659 3569 27721 3570
rect 27659 3549 27667 3569
rect 27687 3551 27721 3569
rect 27742 3569 27803 3570
rect 27742 3551 27775 3569
rect 27687 3549 27775 3551
rect 27795 3549 27803 3569
rect 27659 3541 27803 3549
rect 27659 3540 27695 3541
rect 27767 3540 27803 3541
rect 27869 3574 27906 3575
rect 27869 3573 27907 3574
rect 27869 3565 27933 3573
rect 27869 3545 27878 3565
rect 27898 3551 27933 3565
rect 27953 3551 27956 3571
rect 27898 3546 27956 3551
rect 27898 3545 27933 3546
rect 27338 3508 27375 3537
rect 27339 3506 27375 3508
rect 26816 3498 26852 3499
rect 26664 3468 26673 3488
rect 26693 3468 26701 3488
rect 26664 3458 26701 3468
rect 26760 3488 26908 3498
rect 27008 3495 27104 3497
rect 26760 3468 26769 3488
rect 26789 3468 26879 3488
rect 26899 3468 26908 3488
rect 26760 3459 26908 3468
rect 26966 3488 27104 3495
rect 26966 3468 26975 3488
rect 26995 3468 27104 3488
rect 27339 3484 27530 3506
rect 27556 3505 27593 3537
rect 27869 3533 27933 3545
rect 27973 3507 28000 3685
rect 27832 3505 28000 3507
rect 27556 3491 28000 3505
rect 27556 3479 28003 3491
rect 27599 3477 27632 3479
rect 26966 3459 27104 3468
rect 26760 3458 26797 3459
rect 26490 3405 26531 3406
rect 26264 3384 26316 3402
rect 26382 3398 26531 3405
rect 25819 3365 25859 3375
rect 26382 3378 26441 3398
rect 26461 3378 26500 3398
rect 26520 3378 26531 3398
rect 26382 3370 26531 3378
rect 26598 3401 26755 3408
rect 26598 3381 26718 3401
rect 26738 3381 26755 3401
rect 26598 3371 26755 3381
rect 26598 3370 26633 3371
rect 25649 3348 25687 3357
rect 26598 3349 26629 3370
rect 26816 3349 26852 3459
rect 26871 3458 26908 3459
rect 26967 3458 27004 3459
rect 26927 3399 27017 3405
rect 26927 3379 26936 3399
rect 26956 3397 27017 3399
rect 26956 3379 26981 3397
rect 26927 3377 26981 3379
rect 27001 3377 27017 3397
rect 26927 3371 27017 3377
rect 26441 3348 26478 3349
rect 25649 3347 25686 3348
rect 25110 3319 25200 3325
rect 25110 3299 25126 3319
rect 25146 3317 25200 3319
rect 25146 3299 25171 3317
rect 25110 3297 25171 3299
rect 25191 3297 25200 3317
rect 25110 3291 25200 3297
rect 25123 3237 25160 3238
rect 25219 3237 25256 3238
rect 25275 3237 25311 3347
rect 25498 3326 25529 3347
rect 26440 3339 26478 3348
rect 25494 3325 25529 3326
rect 25372 3315 25529 3325
rect 25372 3295 25389 3315
rect 25409 3295 25529 3315
rect 25372 3288 25529 3295
rect 25596 3318 25745 3326
rect 25596 3298 25607 3318
rect 25627 3298 25666 3318
rect 25686 3298 25745 3318
rect 26268 3321 26308 3331
rect 25596 3291 25745 3298
rect 25811 3294 25863 3312
rect 25596 3290 25637 3291
rect 25330 3237 25367 3238
rect 24061 3220 24120 3222
rect 25023 3228 25161 3237
rect 24061 3219 24229 3220
rect 24355 3219 24395 3221
rect 24061 3193 24505 3219
rect 24061 3191 24229 3193
rect 24061 3189 24142 3191
rect 24061 3013 24088 3189
rect 24128 3153 24192 3165
rect 24468 3161 24505 3193
rect 24531 3192 24722 3214
rect 25023 3208 25132 3228
rect 25152 3208 25161 3228
rect 25023 3201 25161 3208
rect 25219 3228 25367 3237
rect 25219 3208 25228 3228
rect 25248 3208 25338 3228
rect 25358 3208 25367 3228
rect 25023 3199 25119 3201
rect 25219 3198 25367 3208
rect 25426 3228 25463 3238
rect 25426 3208 25434 3228
rect 25454 3208 25463 3228
rect 25275 3197 25311 3198
rect 24686 3190 24722 3192
rect 24686 3161 24723 3190
rect 24128 3152 24163 3153
rect 24105 3147 24163 3152
rect 24105 3127 24108 3147
rect 24128 3133 24163 3147
rect 24183 3133 24192 3153
rect 24128 3125 24192 3133
rect 24154 3124 24192 3125
rect 24155 3123 24192 3124
rect 24258 3157 24294 3158
rect 24366 3157 24402 3158
rect 24258 3149 24402 3157
rect 24258 3129 24266 3149
rect 24286 3148 24374 3149
rect 24286 3130 24321 3148
rect 24339 3130 24374 3148
rect 24286 3129 24374 3130
rect 24394 3129 24402 3149
rect 24258 3123 24402 3129
rect 24468 3153 24506 3161
rect 24584 3157 24620 3158
rect 24468 3133 24477 3153
rect 24497 3133 24506 3153
rect 24468 3124 24506 3133
rect 24535 3149 24620 3157
rect 24535 3129 24592 3149
rect 24612 3129 24620 3149
rect 24468 3123 24505 3124
rect 24535 3123 24620 3129
rect 24686 3153 24724 3161
rect 24686 3133 24695 3153
rect 24715 3133 24724 3153
rect 25426 3141 25463 3208
rect 25498 3237 25529 3288
rect 25811 3276 25829 3294
rect 25847 3276 25863 3294
rect 25548 3237 25585 3238
rect 25498 3228 25585 3237
rect 25498 3208 25556 3228
rect 25576 3208 25585 3228
rect 25498 3198 25585 3208
rect 25644 3228 25681 3238
rect 25644 3208 25652 3228
rect 25672 3208 25681 3228
rect 25498 3197 25529 3198
rect 25123 3138 25160 3139
rect 25426 3138 25465 3141
rect 25122 3137 25465 3138
rect 25644 3137 25681 3208
rect 24686 3124 24724 3133
rect 25047 3132 25465 3137
rect 24686 3123 24723 3124
rect 24147 3095 24237 3101
rect 24147 3075 24163 3095
rect 24183 3093 24237 3095
rect 24183 3075 24208 3093
rect 24147 3073 24208 3075
rect 24228 3073 24237 3093
rect 24147 3067 24237 3073
rect 24160 3013 24197 3014
rect 24256 3013 24293 3014
rect 24312 3013 24348 3123
rect 24535 3102 24566 3123
rect 25047 3112 25050 3132
rect 25070 3112 25465 3132
rect 25494 3113 25681 3137
rect 24531 3101 24566 3102
rect 24409 3091 24566 3101
rect 24409 3071 24426 3091
rect 24446 3071 24566 3091
rect 24409 3064 24566 3071
rect 24633 3094 24782 3102
rect 24633 3074 24644 3094
rect 24664 3074 24703 3094
rect 24723 3074 24782 3094
rect 24633 3067 24782 3074
rect 25426 3087 25465 3112
rect 25811 3087 25863 3276
rect 26268 3303 26278 3321
rect 26296 3303 26308 3321
rect 26440 3319 26449 3339
rect 26469 3319 26478 3339
rect 26440 3311 26478 3319
rect 26544 3343 26629 3349
rect 26659 3348 26696 3349
rect 26544 3323 26552 3343
rect 26572 3323 26629 3343
rect 26544 3315 26629 3323
rect 26658 3339 26696 3348
rect 26658 3319 26667 3339
rect 26687 3319 26696 3339
rect 26544 3314 26580 3315
rect 26658 3311 26696 3319
rect 26762 3343 26906 3349
rect 26762 3323 26770 3343
rect 26790 3323 26823 3343
rect 26843 3323 26878 3343
rect 26898 3323 26906 3343
rect 26762 3315 26906 3323
rect 26762 3314 26798 3315
rect 26870 3314 26906 3315
rect 26972 3348 27009 3349
rect 26972 3347 27010 3348
rect 26972 3339 27036 3347
rect 26972 3319 26981 3339
rect 27001 3325 27036 3339
rect 27056 3325 27059 3345
rect 27001 3320 27059 3325
rect 27001 3319 27036 3320
rect 26268 3247 26308 3303
rect 26441 3282 26478 3311
rect 26442 3280 26478 3282
rect 26442 3258 26633 3280
rect 26659 3279 26696 3311
rect 26972 3307 27036 3319
rect 27076 3281 27103 3459
rect 27961 3434 28003 3479
rect 26935 3279 27103 3281
rect 26659 3269 27103 3279
rect 27244 3375 27431 3399
rect 27462 3380 27855 3400
rect 27875 3380 27878 3400
rect 27462 3375 27878 3380
rect 27244 3304 27281 3375
rect 27462 3374 27803 3375
rect 27396 3314 27427 3315
rect 27244 3284 27253 3304
rect 27273 3284 27281 3304
rect 27244 3274 27281 3284
rect 27340 3304 27427 3314
rect 27340 3284 27349 3304
rect 27369 3284 27427 3304
rect 27340 3275 27427 3284
rect 27340 3274 27377 3275
rect 26265 3242 26308 3247
rect 26656 3253 27103 3269
rect 26656 3247 26684 3253
rect 26935 3252 27103 3253
rect 26265 3239 26415 3242
rect 26656 3239 26683 3247
rect 26265 3237 26683 3239
rect 26265 3219 26274 3237
rect 26292 3219 26683 3237
rect 27396 3224 27427 3275
rect 27462 3304 27499 3374
rect 27765 3373 27802 3374
rect 27614 3314 27650 3315
rect 27462 3284 27471 3304
rect 27491 3284 27499 3304
rect 27462 3274 27499 3284
rect 27558 3304 27706 3314
rect 27806 3311 27902 3313
rect 27558 3284 27567 3304
rect 27587 3284 27677 3304
rect 27697 3284 27706 3304
rect 27558 3275 27706 3284
rect 27764 3304 27902 3311
rect 27764 3284 27773 3304
rect 27793 3284 27902 3304
rect 27764 3275 27902 3284
rect 27558 3274 27595 3275
rect 27288 3221 27329 3222
rect 26265 3216 26683 3219
rect 26265 3210 26308 3216
rect 26268 3207 26308 3210
rect 27183 3214 27329 3221
rect 26665 3198 26705 3199
rect 26376 3181 26705 3198
rect 27183 3194 27239 3214
rect 27259 3194 27298 3214
rect 27318 3194 27329 3214
rect 27183 3186 27329 3194
rect 27396 3217 27553 3224
rect 27396 3197 27516 3217
rect 27536 3197 27553 3217
rect 27396 3187 27553 3197
rect 27396 3186 27431 3187
rect 26260 3138 26303 3149
rect 26260 3120 26272 3138
rect 26290 3120 26303 3138
rect 26260 3094 26303 3120
rect 26376 3094 26403 3181
rect 26665 3172 26705 3181
rect 25426 3069 25865 3087
rect 24633 3066 24674 3067
rect 24367 3013 24404 3014
rect 24060 3004 24198 3013
rect 24060 2984 24169 3004
rect 24189 2984 24198 3004
rect 24060 2977 24198 2984
rect 24256 3004 24404 3013
rect 24256 2984 24265 3004
rect 24285 2984 24375 3004
rect 24395 2984 24404 3004
rect 24060 2975 24156 2977
rect 24256 2974 24404 2984
rect 24463 3004 24500 3014
rect 24463 2984 24471 3004
rect 24491 2984 24500 3004
rect 24312 2973 24348 2974
rect 24160 2914 24197 2915
rect 24463 2914 24500 2984
rect 24535 3013 24566 3064
rect 25426 3051 25826 3069
rect 25844 3051 25865 3069
rect 25426 3045 25865 3051
rect 25432 3041 25865 3045
rect 26260 3073 26403 3094
rect 26447 3146 26481 3162
rect 26665 3152 27058 3172
rect 27078 3152 27081 3172
rect 27396 3165 27427 3186
rect 27614 3165 27650 3275
rect 27669 3274 27706 3275
rect 27765 3274 27802 3275
rect 27725 3215 27815 3221
rect 27725 3195 27734 3215
rect 27754 3213 27815 3215
rect 27754 3195 27779 3213
rect 27725 3193 27779 3195
rect 27799 3193 27815 3213
rect 27725 3187 27815 3193
rect 27239 3164 27276 3165
rect 26665 3147 27081 3152
rect 27238 3155 27276 3164
rect 26665 3146 27006 3147
rect 26447 3076 26484 3146
rect 26599 3086 26630 3087
rect 26260 3071 26397 3073
rect 25811 3039 25863 3041
rect 26260 3029 26303 3071
rect 26447 3056 26456 3076
rect 26476 3056 26484 3076
rect 26447 3046 26484 3056
rect 26543 3076 26630 3086
rect 26543 3056 26552 3076
rect 26572 3056 26630 3076
rect 26543 3047 26630 3056
rect 26543 3046 26580 3047
rect 26258 3019 26303 3029
rect 24585 3013 24622 3014
rect 24535 3004 24622 3013
rect 24535 2984 24593 3004
rect 24613 2984 24622 3004
rect 24535 2974 24622 2984
rect 24681 3004 24718 3014
rect 24681 2984 24689 3004
rect 24709 2984 24718 3004
rect 26258 3001 26267 3019
rect 26285 3001 26303 3019
rect 26258 2995 26303 3001
rect 26599 2996 26630 3047
rect 26665 3076 26702 3146
rect 26968 3145 27005 3146
rect 27238 3135 27247 3155
rect 27267 3135 27276 3155
rect 27238 3127 27276 3135
rect 27342 3159 27427 3165
rect 27457 3164 27494 3165
rect 27342 3139 27350 3159
rect 27370 3139 27427 3159
rect 27342 3131 27427 3139
rect 27456 3155 27494 3164
rect 27456 3135 27465 3155
rect 27485 3135 27494 3155
rect 27342 3130 27378 3131
rect 27456 3127 27494 3135
rect 27560 3159 27704 3165
rect 27560 3139 27568 3159
rect 27588 3156 27676 3159
rect 27588 3139 27623 3156
rect 27560 3138 27623 3139
rect 27642 3139 27676 3156
rect 27696 3139 27704 3159
rect 27642 3138 27704 3139
rect 27560 3131 27704 3138
rect 27560 3130 27596 3131
rect 27668 3130 27704 3131
rect 27770 3164 27807 3165
rect 27770 3163 27808 3164
rect 27830 3163 27857 3167
rect 27770 3161 27857 3163
rect 27770 3155 27834 3161
rect 27770 3135 27779 3155
rect 27799 3141 27834 3155
rect 27854 3141 27857 3161
rect 27799 3136 27857 3141
rect 27799 3135 27834 3136
rect 27239 3098 27276 3127
rect 27240 3096 27276 3098
rect 26817 3086 26853 3087
rect 26665 3056 26674 3076
rect 26694 3056 26702 3076
rect 26665 3046 26702 3056
rect 26761 3076 26909 3086
rect 27009 3083 27105 3085
rect 26761 3056 26770 3076
rect 26790 3056 26880 3076
rect 26900 3056 26909 3076
rect 26761 3047 26909 3056
rect 26967 3076 27105 3083
rect 26967 3056 26976 3076
rect 26996 3056 27105 3076
rect 27240 3074 27431 3096
rect 27457 3095 27494 3127
rect 27770 3123 27834 3135
rect 27874 3097 27901 3275
rect 27733 3095 27901 3097
rect 27457 3069 27901 3095
rect 26967 3047 27105 3056
rect 26761 3046 26798 3047
rect 26258 2992 26295 2995
rect 26491 2993 26532 2994
rect 24535 2973 24566 2974
rect 24159 2913 24500 2914
rect 24681 2913 24718 2984
rect 26383 2986 26532 2993
rect 25814 2974 25851 2979
rect 24084 2908 24500 2913
rect 24084 2888 24087 2908
rect 24107 2888 24500 2908
rect 24531 2889 24718 2913
rect 25805 2970 25852 2974
rect 25805 2952 25824 2970
rect 25842 2952 25852 2970
rect 26383 2966 26442 2986
rect 26462 2966 26501 2986
rect 26521 2966 26532 2986
rect 26383 2958 26532 2966
rect 26599 2989 26756 2996
rect 26599 2969 26719 2989
rect 26739 2969 26756 2989
rect 26599 2959 26756 2969
rect 26599 2958 26634 2959
rect 25805 2904 25852 2952
rect 26599 2937 26630 2958
rect 26817 2937 26853 3047
rect 26872 3046 26909 3047
rect 26968 3046 27005 3047
rect 26928 2987 27018 2993
rect 26928 2967 26937 2987
rect 26957 2985 27018 2987
rect 26957 2967 26982 2985
rect 26928 2965 26982 2967
rect 27002 2965 27018 2985
rect 26928 2959 27018 2965
rect 26442 2936 26479 2937
rect 25429 2901 25852 2904
rect 24304 2887 24369 2888
rect 25407 2871 25852 2901
rect 26254 2928 26292 2930
rect 26254 2920 26297 2928
rect 26254 2902 26265 2920
rect 26283 2902 26297 2920
rect 26254 2875 26297 2902
rect 26441 2927 26479 2936
rect 26441 2907 26450 2927
rect 26470 2907 26479 2927
rect 26441 2899 26479 2907
rect 26545 2931 26630 2937
rect 26660 2936 26697 2937
rect 26545 2911 26553 2931
rect 26573 2911 26630 2931
rect 26545 2903 26630 2911
rect 26659 2927 26697 2936
rect 26659 2907 26668 2927
rect 26688 2907 26697 2927
rect 26545 2902 26581 2903
rect 26659 2899 26697 2907
rect 26763 2935 26907 2937
rect 26763 2931 26815 2935
rect 26763 2911 26771 2931
rect 26791 2915 26815 2931
rect 26835 2931 26907 2935
rect 26835 2915 26879 2931
rect 26791 2911 26879 2915
rect 26899 2911 26907 2931
rect 26763 2903 26907 2911
rect 26763 2902 26799 2903
rect 26871 2902 26907 2903
rect 26973 2936 27010 2937
rect 26973 2935 27011 2936
rect 26973 2927 27037 2935
rect 26973 2907 26982 2927
rect 27002 2913 27037 2927
rect 27057 2913 27060 2933
rect 27002 2908 27060 2913
rect 27002 2907 27037 2908
rect 24500 2855 24540 2863
rect 24500 2833 24508 2855
rect 24532 2833 24540 2855
rect 24105 2604 24142 2610
rect 24105 2585 24113 2604
rect 24134 2585 24142 2604
rect 24105 2577 24142 2585
rect 23805 2456 23812 2478
rect 23836 2456 23844 2478
rect 23805 2450 23844 2456
rect 23335 2445 23375 2447
rect 23501 2446 23669 2447
rect 23603 2445 23640 2446
rect 22569 2429 22707 2438
rect 22363 2428 22400 2429
rect 22093 2375 22134 2376
rect 21867 2354 21919 2372
rect 21985 2368 22134 2375
rect 21435 2334 21475 2344
rect 21985 2348 22044 2368
rect 22064 2348 22103 2368
rect 22123 2348 22134 2368
rect 21985 2340 22134 2348
rect 22201 2371 22358 2378
rect 22201 2351 22321 2371
rect 22341 2351 22358 2371
rect 22201 2341 22358 2351
rect 22201 2340 22236 2341
rect 21265 2317 21303 2326
rect 22201 2319 22232 2340
rect 22419 2319 22455 2429
rect 22474 2428 22511 2429
rect 22570 2428 22607 2429
rect 22530 2369 22620 2375
rect 22530 2349 22539 2369
rect 22559 2367 22620 2369
rect 22559 2349 22584 2367
rect 22530 2347 22584 2349
rect 22604 2347 22620 2367
rect 22530 2341 22620 2347
rect 22044 2318 22081 2319
rect 21265 2316 21302 2317
rect 20726 2288 20816 2294
rect 20726 2268 20742 2288
rect 20762 2286 20816 2288
rect 20762 2268 20787 2286
rect 20726 2266 20787 2268
rect 20807 2266 20816 2286
rect 20726 2260 20816 2266
rect 20739 2206 20776 2207
rect 20835 2206 20872 2207
rect 20891 2206 20927 2316
rect 21114 2295 21145 2316
rect 22043 2309 22081 2318
rect 21110 2294 21145 2295
rect 20988 2284 21145 2294
rect 20988 2264 21005 2284
rect 21025 2264 21145 2284
rect 20988 2257 21145 2264
rect 21212 2287 21361 2295
rect 21212 2267 21223 2287
rect 21243 2267 21282 2287
rect 21302 2267 21361 2287
rect 21871 2291 21911 2301
rect 21212 2260 21361 2267
rect 21427 2263 21479 2281
rect 21212 2259 21253 2260
rect 20946 2206 20983 2207
rect 20639 2197 20777 2206
rect 20111 2186 20144 2188
rect 19740 2174 20187 2186
rect 18972 2052 19140 2054
rect 18696 2026 19140 2052
rect 18206 2004 18344 2013
rect 18000 2003 18037 2004
rect 17497 1949 17534 1952
rect 17730 1950 17771 1951
rect 15500 1901 15916 1906
rect 15500 1881 15503 1901
rect 15523 1881 15916 1901
rect 15947 1882 16134 1906
rect 16759 1904 16799 1909
rect 17155 1904 17202 1947
rect 17622 1943 17771 1950
rect 17622 1923 17681 1943
rect 17701 1923 17740 1943
rect 17760 1923 17771 1943
rect 17622 1915 17771 1923
rect 17838 1946 17995 1953
rect 17838 1926 17958 1946
rect 17978 1926 17995 1946
rect 17838 1916 17995 1926
rect 17838 1915 17873 1916
rect 16759 1865 17202 1904
rect 17838 1894 17869 1915
rect 18056 1894 18092 2004
rect 18111 2003 18148 2004
rect 18207 2003 18244 2004
rect 18167 1944 18257 1950
rect 18167 1924 18176 1944
rect 18196 1942 18257 1944
rect 18196 1924 18221 1942
rect 18167 1922 18221 1924
rect 18241 1922 18257 1942
rect 18167 1916 18257 1922
rect 17681 1893 17718 1894
rect 14540 1806 14548 1828
rect 14572 1806 14580 1828
rect 14540 1798 14580 1806
rect 15853 1850 15893 1858
rect 15853 1828 15861 1850
rect 15885 1828 15893 1850
rect 12059 1752 12094 1753
rect 12036 1747 12094 1752
rect 12036 1727 12039 1747
rect 12059 1733 12094 1747
rect 12114 1733 12123 1753
rect 12059 1725 12123 1733
rect 12085 1724 12123 1725
rect 12086 1723 12123 1724
rect 12189 1757 12225 1758
rect 12297 1757 12333 1758
rect 12189 1749 12333 1757
rect 12189 1729 12197 1749
rect 12217 1745 12305 1749
rect 12217 1729 12261 1745
rect 12189 1725 12261 1729
rect 12281 1729 12305 1745
rect 12325 1729 12333 1749
rect 12281 1725 12333 1729
rect 12189 1723 12333 1725
rect 12399 1753 12437 1761
rect 12515 1757 12551 1758
rect 12399 1733 12408 1753
rect 12428 1733 12437 1753
rect 12399 1724 12437 1733
rect 12466 1749 12551 1757
rect 12466 1729 12523 1749
rect 12543 1729 12551 1749
rect 12399 1723 12436 1724
rect 12466 1723 12551 1729
rect 12617 1753 12655 1761
rect 12617 1733 12626 1753
rect 12646 1733 12655 1753
rect 12617 1724 12655 1733
rect 12799 1758 12841 1767
rect 12799 1740 12813 1758
rect 12831 1740 12841 1758
rect 12799 1732 12841 1740
rect 12804 1730 12841 1732
rect 13231 1752 13674 1791
rect 12617 1723 12654 1724
rect 12078 1695 12168 1701
rect 12078 1675 12094 1695
rect 12114 1693 12168 1695
rect 12114 1675 12139 1693
rect 12078 1673 12139 1675
rect 12159 1673 12168 1693
rect 12078 1667 12168 1673
rect 12091 1613 12128 1614
rect 12187 1613 12224 1614
rect 12243 1613 12279 1723
rect 12466 1702 12497 1723
rect 13231 1709 13278 1752
rect 13634 1747 13674 1752
rect 14299 1750 14486 1774
rect 14517 1755 14910 1775
rect 14930 1755 14933 1775
rect 14517 1750 14933 1755
rect 12462 1701 12497 1702
rect 12340 1691 12497 1701
rect 12340 1671 12357 1691
rect 12377 1671 12497 1691
rect 12340 1664 12497 1671
rect 12564 1694 12713 1702
rect 12564 1674 12575 1694
rect 12595 1674 12634 1694
rect 12654 1674 12713 1694
rect 13231 1691 13241 1709
rect 13259 1691 13278 1709
rect 13231 1687 13278 1691
rect 13232 1682 13269 1687
rect 12564 1667 12713 1674
rect 14299 1679 14336 1750
rect 14517 1749 14858 1750
rect 14451 1689 14482 1690
rect 12564 1666 12605 1667
rect 12801 1665 12838 1668
rect 12298 1613 12335 1614
rect 11991 1604 12129 1613
rect 11195 1565 11639 1591
rect 11195 1563 11363 1565
rect 10148 1431 10595 1443
rect 10191 1429 10224 1431
rect 9558 1411 9696 1420
rect 9352 1410 9389 1411
rect 9082 1357 9123 1358
rect 8856 1336 8908 1354
rect 8974 1350 9123 1357
rect 8411 1317 8451 1327
rect 8974 1330 9033 1350
rect 9053 1330 9092 1350
rect 9112 1330 9123 1350
rect 8974 1322 9123 1330
rect 9190 1353 9347 1360
rect 9190 1333 9310 1353
rect 9330 1333 9347 1353
rect 9190 1323 9347 1333
rect 9190 1322 9225 1323
rect 8241 1300 8279 1309
rect 9190 1301 9221 1322
rect 9408 1301 9444 1411
rect 9463 1410 9500 1411
rect 9559 1410 9596 1411
rect 9519 1351 9609 1357
rect 9519 1331 9528 1351
rect 9548 1349 9609 1351
rect 9548 1331 9573 1349
rect 9519 1329 9573 1331
rect 9593 1329 9609 1349
rect 9519 1323 9609 1329
rect 9033 1300 9070 1301
rect 8241 1299 8278 1300
rect 7702 1271 7792 1277
rect 7702 1251 7718 1271
rect 7738 1269 7792 1271
rect 7738 1251 7763 1269
rect 7702 1249 7763 1251
rect 7783 1249 7792 1269
rect 7702 1243 7792 1249
rect 7715 1189 7752 1190
rect 7811 1189 7848 1190
rect 7867 1189 7903 1299
rect 8090 1278 8121 1299
rect 9032 1291 9070 1300
rect 8086 1277 8121 1278
rect 7964 1267 8121 1277
rect 7964 1247 7981 1267
rect 8001 1247 8121 1267
rect 7964 1240 8121 1247
rect 8188 1270 8337 1278
rect 8188 1250 8199 1270
rect 8219 1250 8258 1270
rect 8278 1250 8337 1270
rect 8860 1273 8900 1283
rect 8188 1243 8337 1250
rect 8403 1246 8455 1264
rect 8188 1242 8229 1243
rect 7922 1189 7959 1190
rect 7615 1180 7753 1189
rect 7615 1160 7724 1180
rect 7744 1160 7753 1180
rect 7615 1153 7753 1160
rect 7811 1180 7959 1189
rect 7811 1160 7820 1180
rect 7840 1160 7930 1180
rect 7950 1160 7959 1180
rect 7615 1151 7711 1153
rect 7811 1150 7959 1160
rect 8018 1180 8055 1190
rect 8018 1160 8026 1180
rect 8046 1160 8055 1180
rect 7867 1149 7903 1150
rect 8018 1093 8055 1160
rect 8090 1189 8121 1240
rect 8403 1228 8421 1246
rect 8439 1228 8455 1246
rect 8140 1189 8177 1190
rect 8090 1180 8177 1189
rect 8090 1160 8148 1180
rect 8168 1160 8177 1180
rect 8090 1150 8177 1160
rect 8236 1180 8273 1190
rect 8236 1160 8244 1180
rect 8264 1160 8273 1180
rect 8090 1149 8121 1150
rect 7715 1090 7752 1091
rect 8018 1090 8057 1093
rect 7714 1089 8057 1090
rect 8236 1089 8273 1160
rect 7639 1084 8057 1089
rect 7639 1064 7642 1084
rect 7662 1064 8057 1084
rect 8086 1065 8273 1089
rect 6180 1033 6217 1041
rect 6180 1014 6188 1033
rect 6209 1014 6217 1033
rect 6180 1008 6217 1014
rect 8018 1039 8057 1064
rect 8403 1039 8455 1228
rect 8860 1255 8870 1273
rect 8888 1255 8900 1273
rect 9032 1271 9041 1291
rect 9061 1271 9070 1291
rect 9032 1263 9070 1271
rect 9136 1295 9221 1301
rect 9251 1300 9288 1301
rect 9136 1275 9144 1295
rect 9164 1275 9221 1295
rect 9136 1267 9221 1275
rect 9250 1291 9288 1300
rect 9250 1271 9259 1291
rect 9279 1271 9288 1291
rect 9136 1266 9172 1267
rect 9250 1263 9288 1271
rect 9354 1295 9498 1301
rect 9354 1275 9362 1295
rect 9382 1275 9415 1295
rect 9435 1275 9470 1295
rect 9490 1275 9498 1295
rect 9354 1267 9498 1275
rect 9354 1266 9390 1267
rect 9462 1266 9498 1267
rect 9564 1300 9601 1301
rect 9564 1299 9602 1300
rect 9564 1291 9628 1299
rect 9564 1271 9573 1291
rect 9593 1277 9628 1291
rect 9648 1277 9651 1297
rect 9593 1272 9651 1277
rect 9593 1271 9628 1272
rect 8860 1199 8900 1255
rect 9033 1234 9070 1263
rect 9034 1232 9070 1234
rect 9034 1210 9225 1232
rect 9251 1231 9288 1263
rect 9564 1259 9628 1271
rect 9668 1233 9695 1411
rect 10553 1386 10595 1431
rect 9527 1231 9695 1233
rect 9251 1221 9695 1231
rect 9836 1327 10023 1351
rect 10054 1332 10447 1352
rect 10467 1332 10470 1352
rect 10054 1327 10470 1332
rect 9836 1256 9873 1327
rect 10054 1326 10395 1327
rect 9988 1266 10019 1267
rect 9836 1236 9845 1256
rect 9865 1236 9873 1256
rect 9836 1226 9873 1236
rect 9932 1256 10019 1266
rect 9932 1236 9941 1256
rect 9961 1236 10019 1256
rect 9932 1227 10019 1236
rect 9932 1226 9969 1227
rect 8857 1194 8900 1199
rect 9248 1205 9695 1221
rect 9248 1199 9276 1205
rect 9527 1204 9695 1205
rect 8857 1191 9007 1194
rect 9248 1191 9275 1199
rect 8857 1189 9275 1191
rect 8857 1171 8866 1189
rect 8884 1171 9275 1189
rect 9988 1176 10019 1227
rect 10054 1256 10091 1326
rect 10357 1325 10394 1326
rect 10206 1266 10242 1267
rect 10054 1236 10063 1256
rect 10083 1236 10091 1256
rect 10054 1226 10091 1236
rect 10150 1256 10298 1266
rect 10398 1263 10494 1265
rect 10150 1236 10159 1256
rect 10179 1236 10269 1256
rect 10289 1236 10298 1256
rect 10150 1227 10298 1236
rect 10356 1256 10494 1263
rect 10356 1236 10365 1256
rect 10385 1236 10494 1256
rect 10356 1227 10494 1236
rect 10150 1226 10187 1227
rect 9880 1173 9921 1174
rect 8857 1168 9275 1171
rect 8857 1162 8900 1168
rect 8860 1159 8900 1162
rect 9775 1166 9921 1173
rect 9257 1150 9297 1151
rect 8968 1133 9297 1150
rect 9775 1146 9831 1166
rect 9851 1146 9890 1166
rect 9910 1146 9921 1166
rect 9775 1138 9921 1146
rect 9988 1169 10145 1176
rect 9988 1149 10108 1169
rect 10128 1149 10145 1169
rect 9988 1139 10145 1149
rect 9988 1138 10023 1139
rect 8852 1090 8895 1101
rect 8852 1072 8864 1090
rect 8882 1072 8895 1090
rect 8852 1046 8895 1072
rect 8968 1046 8995 1133
rect 9257 1124 9297 1133
rect 8018 1021 8457 1039
rect 8018 1003 8418 1021
rect 8436 1003 8457 1021
rect 8018 997 8457 1003
rect 8024 993 8457 997
rect 8852 1025 8995 1046
rect 9039 1098 9073 1114
rect 9257 1104 9650 1124
rect 9670 1104 9673 1124
rect 9988 1117 10019 1138
rect 10206 1117 10242 1227
rect 10261 1226 10298 1227
rect 10357 1226 10394 1227
rect 10317 1167 10407 1173
rect 10317 1147 10326 1167
rect 10346 1165 10407 1167
rect 10346 1147 10371 1165
rect 10317 1145 10371 1147
rect 10391 1145 10407 1165
rect 10317 1139 10407 1145
rect 9831 1116 9868 1117
rect 9257 1099 9673 1104
rect 9830 1107 9868 1116
rect 9257 1098 9598 1099
rect 9039 1028 9076 1098
rect 9191 1038 9222 1039
rect 8852 1023 8989 1025
rect 8403 991 8455 993
rect 8852 981 8895 1023
rect 9039 1008 9048 1028
rect 9068 1008 9076 1028
rect 9039 998 9076 1008
rect 9135 1028 9222 1038
rect 9135 1008 9144 1028
rect 9164 1008 9222 1028
rect 9135 999 9222 1008
rect 9135 998 9172 999
rect 8850 971 8895 981
rect 8850 953 8859 971
rect 8877 953 8895 971
rect 8850 947 8895 953
rect 9191 948 9222 999
rect 9257 1028 9294 1098
rect 9560 1097 9597 1098
rect 9830 1087 9839 1107
rect 9859 1087 9868 1107
rect 9830 1079 9868 1087
rect 9934 1111 10019 1117
rect 10049 1116 10086 1117
rect 9934 1091 9942 1111
rect 9962 1091 10019 1111
rect 9934 1083 10019 1091
rect 10048 1107 10086 1116
rect 10048 1087 10057 1107
rect 10077 1087 10086 1107
rect 9934 1082 9970 1083
rect 10048 1079 10086 1087
rect 10152 1111 10296 1117
rect 10152 1091 10160 1111
rect 10180 1108 10268 1111
rect 10180 1091 10215 1108
rect 10152 1090 10215 1091
rect 10234 1091 10268 1108
rect 10288 1091 10296 1111
rect 10234 1090 10296 1091
rect 10152 1083 10296 1090
rect 10152 1082 10188 1083
rect 10260 1082 10296 1083
rect 10362 1116 10399 1117
rect 10362 1115 10400 1116
rect 10422 1115 10449 1119
rect 10362 1113 10449 1115
rect 10362 1107 10426 1113
rect 10362 1087 10371 1107
rect 10391 1093 10426 1107
rect 10446 1093 10449 1113
rect 10391 1088 10449 1093
rect 10391 1087 10426 1088
rect 9831 1050 9868 1079
rect 9832 1048 9868 1050
rect 9409 1038 9445 1039
rect 9257 1008 9266 1028
rect 9286 1008 9294 1028
rect 9257 998 9294 1008
rect 9353 1028 9501 1038
rect 9601 1035 9697 1037
rect 9353 1008 9362 1028
rect 9382 1008 9472 1028
rect 9492 1008 9501 1028
rect 9353 999 9501 1008
rect 9559 1028 9697 1035
rect 9559 1008 9568 1028
rect 9588 1008 9697 1028
rect 9832 1026 10023 1048
rect 10049 1047 10086 1079
rect 10362 1075 10426 1087
rect 10466 1049 10493 1227
rect 10325 1047 10493 1049
rect 10049 1021 10493 1047
rect 9559 999 9697 1008
rect 9353 998 9390 999
rect 8850 944 8887 947
rect 9083 945 9124 946
rect 8975 938 9124 945
rect 8406 926 8443 931
rect 8397 922 8444 926
rect 8397 904 8416 922
rect 8434 904 8444 922
rect 8975 918 9034 938
rect 9054 918 9093 938
rect 9113 918 9124 938
rect 8975 910 9124 918
rect 9191 941 9348 948
rect 9191 921 9311 941
rect 9331 921 9348 941
rect 9191 911 9348 921
rect 9191 910 9226 911
rect 8397 841 8444 904
rect 9191 889 9222 910
rect 9409 889 9445 999
rect 9464 998 9501 999
rect 9560 998 9597 999
rect 9520 939 9610 945
rect 9520 919 9529 939
rect 9549 937 9610 939
rect 9549 919 9574 937
rect 9520 917 9574 919
rect 9594 917 9610 937
rect 9520 911 9610 917
rect 9034 888 9071 889
rect 8847 880 8884 882
rect 8847 872 8889 880
rect 8847 854 8857 872
rect 8875 854 8889 872
rect 8847 845 8889 854
rect 9033 879 9071 888
rect 9033 859 9042 879
rect 9062 859 9071 879
rect 9033 851 9071 859
rect 9137 883 9222 889
rect 9252 888 9289 889
rect 9137 863 9145 883
rect 9165 863 9222 883
rect 9137 855 9222 863
rect 9251 879 9289 888
rect 9251 859 9260 879
rect 9280 859 9289 879
rect 9137 854 9173 855
rect 9251 851 9289 859
rect 9355 887 9499 889
rect 9355 883 9407 887
rect 9355 863 9363 883
rect 9383 867 9407 883
rect 9427 883 9499 887
rect 9427 867 9471 883
rect 9383 863 9471 867
rect 9491 863 9499 883
rect 9355 855 9499 863
rect 9355 854 9391 855
rect 9463 854 9499 855
rect 9565 888 9602 889
rect 9565 887 9603 888
rect 9565 879 9629 887
rect 9565 859 9574 879
rect 9594 865 9629 879
rect 9649 865 9652 885
rect 9594 860 9652 865
rect 9594 859 9629 860
rect 8397 826 8447 841
rect 8397 801 8411 826
rect 8443 801 8447 826
rect 8848 820 8889 845
rect 9034 820 9071 851
rect 9252 829 9289 851
rect 9565 847 9629 859
rect 9247 820 9289 829
rect 9669 821 9696 999
rect 8848 808 8893 820
rect 8397 788 8444 801
rect 5782 763 5790 785
rect 5814 763 5822 785
rect 5782 755 5822 763
rect 8844 750 8893 808
rect 9034 794 9096 820
rect 9247 819 9332 820
rect 9528 819 9696 821
rect 9247 793 9696 819
rect 9247 750 9286 793
rect 9528 792 9696 793
rect 10159 797 10199 1021
rect 10325 1020 10493 1021
rect 10557 1053 10590 1386
rect 11195 1385 11222 1563
rect 11262 1525 11326 1537
rect 11602 1533 11639 1565
rect 11665 1564 11856 1586
rect 11991 1584 12100 1604
rect 12120 1584 12129 1604
rect 11991 1577 12129 1584
rect 12187 1604 12335 1613
rect 12187 1584 12196 1604
rect 12216 1584 12306 1604
rect 12326 1584 12335 1604
rect 11991 1575 12087 1577
rect 12187 1574 12335 1584
rect 12394 1604 12431 1614
rect 12394 1584 12402 1604
rect 12422 1584 12431 1604
rect 12243 1573 12279 1574
rect 11820 1562 11856 1564
rect 11820 1533 11857 1562
rect 11262 1524 11297 1525
rect 11239 1519 11297 1524
rect 11239 1499 11242 1519
rect 11262 1505 11297 1519
rect 11317 1505 11326 1525
rect 11262 1497 11326 1505
rect 11288 1496 11326 1497
rect 11289 1495 11326 1496
rect 11392 1529 11428 1530
rect 11500 1529 11536 1530
rect 11392 1521 11536 1529
rect 11392 1501 11400 1521
rect 11420 1520 11508 1521
rect 11420 1501 11455 1520
rect 11476 1501 11508 1520
rect 11528 1501 11536 1521
rect 11392 1495 11536 1501
rect 11602 1525 11640 1533
rect 11718 1529 11754 1530
rect 11602 1505 11611 1525
rect 11631 1505 11640 1525
rect 11602 1496 11640 1505
rect 11669 1521 11754 1529
rect 11669 1501 11726 1521
rect 11746 1501 11754 1521
rect 11602 1495 11639 1496
rect 11669 1495 11754 1501
rect 11820 1525 11858 1533
rect 11820 1505 11829 1525
rect 11849 1505 11858 1525
rect 12091 1514 12128 1515
rect 12394 1514 12431 1584
rect 12466 1613 12497 1664
rect 12793 1659 12838 1665
rect 12793 1641 12811 1659
rect 12829 1641 12838 1659
rect 14299 1659 14308 1679
rect 14328 1659 14336 1679
rect 14299 1649 14336 1659
rect 14395 1679 14482 1689
rect 14395 1659 14404 1679
rect 14424 1659 14482 1679
rect 14395 1650 14482 1659
rect 14395 1649 14432 1650
rect 12793 1631 12838 1641
rect 12516 1613 12553 1614
rect 12466 1604 12553 1613
rect 12466 1584 12524 1604
rect 12544 1584 12553 1604
rect 12466 1574 12553 1584
rect 12612 1604 12649 1614
rect 12612 1584 12620 1604
rect 12640 1584 12649 1604
rect 12793 1589 12836 1631
rect 13220 1620 13272 1622
rect 12699 1587 12836 1589
rect 12466 1573 12497 1574
rect 12612 1514 12649 1584
rect 12090 1513 12431 1514
rect 11820 1496 11858 1505
rect 12015 1508 12431 1513
rect 11820 1495 11857 1496
rect 11281 1467 11371 1473
rect 11281 1447 11297 1467
rect 11317 1465 11371 1467
rect 11317 1447 11342 1465
rect 11281 1445 11342 1447
rect 11362 1445 11371 1465
rect 11281 1439 11371 1445
rect 11294 1385 11331 1386
rect 11390 1385 11427 1386
rect 11446 1385 11482 1495
rect 11669 1474 11700 1495
rect 12015 1488 12018 1508
rect 12038 1488 12431 1508
rect 12615 1498 12649 1514
rect 12693 1566 12836 1587
rect 13218 1616 13651 1620
rect 13218 1610 13657 1616
rect 13218 1592 13239 1610
rect 13257 1592 13657 1610
rect 14451 1599 14482 1650
rect 14517 1679 14554 1749
rect 14820 1748 14857 1749
rect 14669 1689 14705 1690
rect 14517 1659 14526 1679
rect 14546 1659 14554 1679
rect 14517 1649 14554 1659
rect 14613 1679 14761 1689
rect 14861 1686 14957 1688
rect 14613 1659 14622 1679
rect 14642 1659 14732 1679
rect 14752 1659 14761 1679
rect 14613 1650 14761 1659
rect 14819 1679 14957 1686
rect 14819 1659 14828 1679
rect 14848 1659 14957 1679
rect 14819 1650 14957 1659
rect 14613 1649 14650 1650
rect 14343 1596 14384 1597
rect 13218 1574 13657 1592
rect 12391 1479 12431 1488
rect 12693 1479 12720 1566
rect 12793 1540 12836 1566
rect 12793 1522 12806 1540
rect 12824 1522 12836 1540
rect 12793 1511 12836 1522
rect 11665 1473 11700 1474
rect 11543 1463 11700 1473
rect 11543 1443 11560 1463
rect 11580 1443 11700 1463
rect 11543 1436 11700 1443
rect 11767 1466 11916 1474
rect 11767 1446 11778 1466
rect 11798 1446 11837 1466
rect 11857 1446 11916 1466
rect 12391 1462 12720 1479
rect 12391 1461 12431 1462
rect 11767 1439 11916 1446
rect 12788 1450 12828 1453
rect 12788 1444 12831 1450
rect 12413 1441 12831 1444
rect 11767 1438 11808 1439
rect 11501 1385 11538 1386
rect 11194 1376 11332 1385
rect 11194 1356 11303 1376
rect 11323 1356 11332 1376
rect 11194 1349 11332 1356
rect 11390 1376 11538 1385
rect 11390 1356 11399 1376
rect 11419 1356 11509 1376
rect 11529 1356 11538 1376
rect 11194 1347 11290 1349
rect 11390 1346 11538 1356
rect 11597 1376 11634 1386
rect 11597 1356 11605 1376
rect 11625 1356 11634 1376
rect 11446 1345 11482 1346
rect 11294 1286 11331 1287
rect 11597 1286 11634 1356
rect 11669 1385 11700 1436
rect 12413 1423 12804 1441
rect 12822 1423 12831 1441
rect 12413 1421 12831 1423
rect 12413 1413 12440 1421
rect 12681 1418 12831 1421
rect 11993 1407 12161 1408
rect 12412 1407 12440 1413
rect 11993 1391 12440 1407
rect 12788 1413 12831 1418
rect 11719 1385 11756 1386
rect 11669 1376 11756 1385
rect 11669 1356 11727 1376
rect 11747 1356 11756 1376
rect 11669 1346 11756 1356
rect 11815 1376 11852 1386
rect 11815 1356 11823 1376
rect 11843 1356 11852 1376
rect 11669 1345 11700 1346
rect 11293 1285 11634 1286
rect 11815 1285 11852 1356
rect 11218 1280 11634 1285
rect 11218 1260 11221 1280
rect 11241 1260 11634 1280
rect 11665 1261 11852 1285
rect 11993 1381 12437 1391
rect 11993 1379 12161 1381
rect 11993 1201 12020 1379
rect 12060 1341 12124 1353
rect 12400 1349 12437 1381
rect 12463 1380 12654 1402
rect 12618 1378 12654 1380
rect 12618 1349 12655 1378
rect 12788 1357 12828 1413
rect 12060 1340 12095 1341
rect 12037 1335 12095 1340
rect 12037 1315 12040 1335
rect 12060 1321 12095 1335
rect 12115 1321 12124 1341
rect 12060 1313 12124 1321
rect 12086 1312 12124 1313
rect 12087 1311 12124 1312
rect 12190 1345 12226 1346
rect 12298 1345 12334 1346
rect 12190 1337 12334 1345
rect 12190 1317 12198 1337
rect 12218 1317 12253 1337
rect 12273 1317 12306 1337
rect 12326 1317 12334 1337
rect 12190 1311 12334 1317
rect 12400 1341 12438 1349
rect 12516 1345 12552 1346
rect 12400 1321 12409 1341
rect 12429 1321 12438 1341
rect 12400 1312 12438 1321
rect 12467 1337 12552 1345
rect 12467 1317 12524 1337
rect 12544 1317 12552 1337
rect 12400 1311 12437 1312
rect 12467 1311 12552 1317
rect 12618 1341 12656 1349
rect 12618 1321 12627 1341
rect 12647 1321 12656 1341
rect 12788 1339 12800 1357
rect 12818 1339 12828 1357
rect 13220 1385 13272 1574
rect 13618 1549 13657 1574
rect 14235 1589 14384 1596
rect 14235 1569 14294 1589
rect 14314 1569 14353 1589
rect 14373 1569 14384 1589
rect 14235 1561 14384 1569
rect 14451 1592 14608 1599
rect 14451 1572 14571 1592
rect 14591 1572 14608 1592
rect 14451 1562 14608 1572
rect 14451 1561 14486 1562
rect 13402 1524 13589 1548
rect 13618 1529 14013 1549
rect 14033 1529 14036 1549
rect 14451 1540 14482 1561
rect 14669 1540 14705 1650
rect 14724 1649 14761 1650
rect 14820 1649 14857 1650
rect 14780 1590 14870 1596
rect 14780 1570 14789 1590
rect 14809 1588 14870 1590
rect 14809 1570 14834 1588
rect 14780 1568 14834 1570
rect 14854 1568 14870 1588
rect 14780 1562 14870 1568
rect 14294 1539 14331 1540
rect 13618 1524 14036 1529
rect 14293 1530 14331 1539
rect 13402 1453 13439 1524
rect 13618 1523 13961 1524
rect 13618 1520 13657 1523
rect 13923 1522 13960 1523
rect 13554 1463 13585 1464
rect 13402 1433 13411 1453
rect 13431 1433 13439 1453
rect 13402 1423 13439 1433
rect 13498 1453 13585 1463
rect 13498 1433 13507 1453
rect 13527 1433 13585 1453
rect 13498 1424 13585 1433
rect 13498 1423 13535 1424
rect 13220 1367 13236 1385
rect 13254 1367 13272 1385
rect 13554 1373 13585 1424
rect 13620 1453 13657 1520
rect 14293 1510 14302 1530
rect 14322 1510 14331 1530
rect 14293 1502 14331 1510
rect 14397 1534 14482 1540
rect 14512 1539 14549 1540
rect 14397 1514 14405 1534
rect 14425 1514 14482 1534
rect 14397 1506 14482 1514
rect 14511 1530 14549 1539
rect 14511 1510 14520 1530
rect 14540 1510 14549 1530
rect 14397 1505 14433 1506
rect 14511 1502 14549 1510
rect 14615 1534 14759 1540
rect 14615 1514 14623 1534
rect 14643 1529 14731 1534
rect 14643 1514 14679 1529
rect 14615 1512 14679 1514
rect 14698 1514 14731 1529
rect 14751 1514 14759 1534
rect 14698 1512 14759 1514
rect 14615 1506 14759 1512
rect 14615 1505 14651 1506
rect 14723 1505 14759 1506
rect 14825 1539 14862 1540
rect 14825 1538 14863 1539
rect 14825 1530 14889 1538
rect 14825 1510 14834 1530
rect 14854 1516 14889 1530
rect 14909 1516 14912 1536
rect 14854 1511 14912 1516
rect 14854 1510 14889 1511
rect 14294 1473 14331 1502
rect 14295 1471 14331 1473
rect 13772 1463 13808 1464
rect 13620 1433 13629 1453
rect 13649 1433 13657 1453
rect 13620 1423 13657 1433
rect 13716 1453 13864 1463
rect 13964 1460 14060 1462
rect 13716 1433 13725 1453
rect 13745 1433 13835 1453
rect 13855 1433 13864 1453
rect 13716 1424 13864 1433
rect 13922 1453 14060 1460
rect 13922 1433 13931 1453
rect 13951 1433 14060 1453
rect 14295 1449 14486 1471
rect 14512 1470 14549 1502
rect 14825 1498 14889 1510
rect 14929 1472 14956 1650
rect 14788 1470 14956 1472
rect 14512 1456 14956 1470
rect 15559 1604 15727 1605
rect 15853 1604 15893 1828
rect 16356 1832 16524 1833
rect 16759 1832 16799 1865
rect 17155 1832 17202 1865
rect 17494 1885 17531 1887
rect 17494 1877 17536 1885
rect 17494 1859 17504 1877
rect 17522 1859 17536 1877
rect 17494 1850 17536 1859
rect 17680 1884 17718 1893
rect 17680 1864 17689 1884
rect 17709 1864 17718 1884
rect 17680 1856 17718 1864
rect 17784 1888 17869 1894
rect 17899 1893 17936 1894
rect 17784 1868 17792 1888
rect 17812 1868 17869 1888
rect 17784 1860 17869 1868
rect 17898 1884 17936 1893
rect 17898 1864 17907 1884
rect 17927 1864 17936 1884
rect 17784 1859 17820 1860
rect 17898 1856 17936 1864
rect 18002 1892 18146 1894
rect 18002 1888 18054 1892
rect 18002 1868 18010 1888
rect 18030 1872 18054 1888
rect 18074 1888 18146 1892
rect 18074 1872 18118 1888
rect 18030 1868 18118 1872
rect 18138 1868 18146 1888
rect 18002 1860 18146 1868
rect 18002 1859 18038 1860
rect 18110 1859 18146 1860
rect 18212 1893 18249 1894
rect 18212 1892 18250 1893
rect 18212 1884 18276 1892
rect 18212 1864 18221 1884
rect 18241 1870 18276 1884
rect 18296 1870 18299 1890
rect 18241 1865 18299 1870
rect 18241 1864 18276 1865
rect 16356 1831 16800 1832
rect 16356 1806 16801 1831
rect 16356 1804 16524 1806
rect 16720 1805 16801 1806
rect 16970 1805 17019 1831
rect 17155 1805 17204 1832
rect 16356 1626 16383 1804
rect 16423 1766 16487 1778
rect 16763 1774 16800 1805
rect 16981 1774 17018 1805
rect 17163 1780 17204 1805
rect 17495 1825 17536 1850
rect 17681 1825 17718 1856
rect 17899 1825 17936 1856
rect 18212 1852 18276 1864
rect 18316 1826 18343 2004
rect 17495 1798 17544 1825
rect 17680 1799 17729 1825
rect 17898 1824 17979 1825
rect 18175 1824 18343 1826
rect 17898 1799 18343 1824
rect 17899 1798 18343 1799
rect 16423 1765 16458 1766
rect 16400 1760 16458 1765
rect 16400 1740 16403 1760
rect 16423 1746 16458 1760
rect 16478 1746 16487 1766
rect 16423 1738 16487 1746
rect 16449 1737 16487 1738
rect 16450 1736 16487 1737
rect 16553 1770 16589 1771
rect 16661 1770 16697 1771
rect 16553 1762 16697 1770
rect 16553 1742 16561 1762
rect 16581 1758 16669 1762
rect 16581 1742 16625 1758
rect 16553 1738 16625 1742
rect 16645 1742 16669 1758
rect 16689 1742 16697 1762
rect 16645 1738 16697 1742
rect 16553 1736 16697 1738
rect 16763 1766 16801 1774
rect 16879 1770 16915 1771
rect 16763 1746 16772 1766
rect 16792 1746 16801 1766
rect 16763 1737 16801 1746
rect 16830 1762 16915 1770
rect 16830 1742 16887 1762
rect 16907 1742 16915 1762
rect 16763 1736 16800 1737
rect 16830 1736 16915 1742
rect 16981 1766 17019 1774
rect 16981 1746 16990 1766
rect 17010 1746 17019 1766
rect 16981 1737 17019 1746
rect 17163 1771 17205 1780
rect 17163 1753 17177 1771
rect 17195 1753 17205 1771
rect 17163 1745 17205 1753
rect 17168 1743 17205 1745
rect 17497 1765 17544 1798
rect 17900 1765 17940 1798
rect 18175 1797 18343 1798
rect 18806 1802 18846 2026
rect 18972 2025 19140 2026
rect 19743 2160 20187 2174
rect 19743 2158 19911 2160
rect 19743 1980 19770 2158
rect 19810 2120 19874 2132
rect 20150 2128 20187 2160
rect 20213 2159 20404 2181
rect 20639 2177 20748 2197
rect 20768 2177 20777 2197
rect 20639 2170 20777 2177
rect 20835 2197 20983 2206
rect 20835 2177 20844 2197
rect 20864 2177 20954 2197
rect 20974 2177 20983 2197
rect 20639 2168 20735 2170
rect 20835 2167 20983 2177
rect 21042 2197 21079 2207
rect 21042 2177 21050 2197
rect 21070 2177 21079 2197
rect 20891 2166 20927 2167
rect 20368 2157 20404 2159
rect 20368 2128 20405 2157
rect 19810 2119 19845 2120
rect 19787 2114 19845 2119
rect 19787 2094 19790 2114
rect 19810 2100 19845 2114
rect 19865 2100 19874 2120
rect 19810 2092 19874 2100
rect 19836 2091 19874 2092
rect 19837 2090 19874 2091
rect 19940 2124 19976 2125
rect 20048 2124 20084 2125
rect 19940 2116 20084 2124
rect 19940 2096 19948 2116
rect 19968 2114 20056 2116
rect 19968 2096 20001 2114
rect 19940 2095 20001 2096
rect 20022 2096 20056 2114
rect 20076 2096 20084 2116
rect 20022 2095 20084 2096
rect 19940 2090 20084 2095
rect 20150 2120 20188 2128
rect 20266 2124 20302 2125
rect 20150 2100 20159 2120
rect 20179 2100 20188 2120
rect 20150 2091 20188 2100
rect 20217 2116 20302 2124
rect 20217 2096 20274 2116
rect 20294 2096 20302 2116
rect 20150 2090 20187 2091
rect 20217 2090 20302 2096
rect 20368 2120 20406 2128
rect 20368 2100 20377 2120
rect 20397 2100 20406 2120
rect 21042 2110 21079 2177
rect 21114 2206 21145 2257
rect 21427 2245 21445 2263
rect 21463 2245 21479 2263
rect 21164 2206 21201 2207
rect 21114 2197 21201 2206
rect 21114 2177 21172 2197
rect 21192 2177 21201 2197
rect 21114 2167 21201 2177
rect 21260 2197 21297 2207
rect 21260 2177 21268 2197
rect 21288 2177 21297 2197
rect 21114 2166 21145 2167
rect 20739 2107 20776 2108
rect 21042 2107 21081 2110
rect 20738 2106 21081 2107
rect 21260 2106 21297 2177
rect 20368 2091 20406 2100
rect 20663 2101 21081 2106
rect 20368 2090 20405 2091
rect 19829 2062 19919 2068
rect 19829 2042 19845 2062
rect 19865 2060 19919 2062
rect 19865 2042 19890 2060
rect 19829 2040 19890 2042
rect 19910 2040 19919 2060
rect 19829 2034 19919 2040
rect 19842 1980 19879 1981
rect 19938 1980 19975 1981
rect 19994 1980 20030 2090
rect 20217 2069 20248 2090
rect 20663 2081 20666 2101
rect 20686 2081 21081 2101
rect 21110 2082 21297 2106
rect 20213 2068 20248 2069
rect 20091 2058 20248 2068
rect 20091 2038 20108 2058
rect 20128 2038 20248 2058
rect 20091 2031 20248 2038
rect 20315 2061 20464 2069
rect 20315 2041 20326 2061
rect 20346 2041 20385 2061
rect 20405 2041 20464 2061
rect 20315 2034 20464 2041
rect 21042 2056 21081 2081
rect 21427 2056 21479 2245
rect 21871 2273 21881 2291
rect 21899 2273 21911 2291
rect 22043 2289 22052 2309
rect 22072 2289 22081 2309
rect 22043 2281 22081 2289
rect 22147 2313 22232 2319
rect 22262 2318 22299 2319
rect 22147 2293 22155 2313
rect 22175 2293 22232 2313
rect 22147 2285 22232 2293
rect 22261 2309 22299 2318
rect 22261 2289 22270 2309
rect 22290 2289 22299 2309
rect 22147 2284 22183 2285
rect 22261 2281 22299 2289
rect 22365 2313 22509 2319
rect 22365 2293 22373 2313
rect 22393 2293 22426 2313
rect 22446 2293 22481 2313
rect 22501 2293 22509 2313
rect 22365 2285 22509 2293
rect 22365 2284 22401 2285
rect 22473 2284 22509 2285
rect 22575 2318 22612 2319
rect 22575 2317 22613 2318
rect 22575 2309 22639 2317
rect 22575 2289 22584 2309
rect 22604 2295 22639 2309
rect 22659 2295 22662 2315
rect 22604 2290 22662 2295
rect 22604 2289 22639 2290
rect 21871 2217 21911 2273
rect 22044 2252 22081 2281
rect 22045 2250 22081 2252
rect 22045 2228 22236 2250
rect 22262 2249 22299 2281
rect 22575 2277 22639 2289
rect 22679 2251 22706 2429
rect 22538 2249 22706 2251
rect 22262 2239 22706 2249
rect 22847 2345 23034 2369
rect 23065 2350 23458 2370
rect 23478 2350 23481 2370
rect 23065 2345 23481 2350
rect 22847 2274 22884 2345
rect 23065 2344 23406 2345
rect 22999 2284 23030 2285
rect 22847 2254 22856 2274
rect 22876 2254 22884 2274
rect 22847 2244 22884 2254
rect 22943 2274 23030 2284
rect 22943 2254 22952 2274
rect 22972 2254 23030 2274
rect 22943 2245 23030 2254
rect 22943 2244 22980 2245
rect 21868 2212 21911 2217
rect 22259 2223 22706 2239
rect 22259 2217 22287 2223
rect 22538 2222 22706 2223
rect 21868 2209 22018 2212
rect 22259 2209 22286 2217
rect 21868 2207 22286 2209
rect 21868 2189 21877 2207
rect 21895 2189 22286 2207
rect 22999 2194 23030 2245
rect 23065 2274 23102 2344
rect 23368 2343 23405 2344
rect 23606 2286 23639 2445
rect 23217 2284 23253 2285
rect 23065 2254 23074 2274
rect 23094 2254 23102 2274
rect 23065 2244 23102 2254
rect 23161 2274 23309 2284
rect 23409 2281 23505 2283
rect 23161 2254 23170 2274
rect 23190 2254 23280 2274
rect 23300 2254 23309 2274
rect 23161 2245 23309 2254
rect 23367 2274 23505 2281
rect 23367 2254 23376 2274
rect 23396 2254 23505 2274
rect 23606 2282 23642 2286
rect 23606 2264 23615 2282
rect 23637 2264 23642 2282
rect 23606 2258 23642 2264
rect 23367 2245 23505 2254
rect 23161 2244 23198 2245
rect 22891 2191 22932 2192
rect 21868 2186 22286 2189
rect 21868 2180 21911 2186
rect 21871 2177 21911 2180
rect 22783 2184 22932 2191
rect 22268 2168 22308 2169
rect 21979 2151 22308 2168
rect 22783 2164 22842 2184
rect 22862 2164 22901 2184
rect 22921 2164 22932 2184
rect 22783 2156 22932 2164
rect 22999 2187 23156 2194
rect 22999 2167 23119 2187
rect 23139 2167 23156 2187
rect 22999 2157 23156 2167
rect 22999 2156 23034 2157
rect 21863 2108 21906 2119
rect 21863 2090 21875 2108
rect 21893 2090 21906 2108
rect 21863 2064 21906 2090
rect 21979 2064 22006 2151
rect 22268 2142 22308 2151
rect 21042 2038 21481 2056
rect 20315 2033 20356 2034
rect 20049 1980 20086 1981
rect 19742 1971 19880 1980
rect 19742 1951 19851 1971
rect 19871 1951 19880 1971
rect 19742 1944 19880 1951
rect 19938 1971 20086 1980
rect 19938 1951 19947 1971
rect 19967 1951 20057 1971
rect 20077 1951 20086 1971
rect 19742 1942 19838 1944
rect 19938 1941 20086 1951
rect 20145 1971 20182 1981
rect 20145 1951 20153 1971
rect 20173 1951 20182 1971
rect 19994 1940 20030 1941
rect 19842 1881 19879 1882
rect 20145 1881 20182 1951
rect 20217 1980 20248 2031
rect 21042 2020 21442 2038
rect 21460 2020 21481 2038
rect 21042 2014 21481 2020
rect 21048 2010 21481 2014
rect 21863 2043 22006 2064
rect 22050 2116 22084 2132
rect 22268 2122 22661 2142
rect 22681 2122 22684 2142
rect 22999 2135 23030 2156
rect 23217 2135 23253 2245
rect 23272 2244 23309 2245
rect 23368 2244 23405 2245
rect 23328 2185 23418 2191
rect 23328 2165 23337 2185
rect 23357 2183 23418 2185
rect 23357 2165 23382 2183
rect 23328 2163 23382 2165
rect 23402 2163 23418 2183
rect 23328 2157 23418 2163
rect 22842 2134 22879 2135
rect 22268 2117 22684 2122
rect 22841 2125 22879 2134
rect 22268 2116 22609 2117
rect 22050 2046 22087 2116
rect 22202 2056 22233 2057
rect 21863 2041 22000 2043
rect 21427 2008 21479 2010
rect 21863 1999 21906 2041
rect 22050 2026 22059 2046
rect 22079 2026 22087 2046
rect 22050 2016 22087 2026
rect 22146 2046 22233 2056
rect 22146 2026 22155 2046
rect 22175 2026 22233 2046
rect 22146 2017 22233 2026
rect 22146 2016 22183 2017
rect 21861 1989 21906 1999
rect 20267 1980 20304 1981
rect 20217 1971 20304 1980
rect 20217 1951 20275 1971
rect 20295 1951 20304 1971
rect 20217 1941 20304 1951
rect 20363 1971 20400 1981
rect 20363 1951 20371 1971
rect 20391 1951 20400 1971
rect 21861 1971 21870 1989
rect 21888 1971 21906 1989
rect 21861 1965 21906 1971
rect 22202 1966 22233 2017
rect 22268 2046 22305 2116
rect 22571 2115 22608 2116
rect 22841 2105 22850 2125
rect 22870 2105 22879 2125
rect 22841 2097 22879 2105
rect 22945 2129 23030 2135
rect 23060 2134 23097 2135
rect 22945 2109 22953 2129
rect 22973 2109 23030 2129
rect 22945 2101 23030 2109
rect 23059 2125 23097 2134
rect 23059 2105 23068 2125
rect 23088 2105 23097 2125
rect 22945 2100 22981 2101
rect 23059 2097 23097 2105
rect 23163 2129 23307 2135
rect 23163 2109 23171 2129
rect 23191 2110 23223 2129
rect 23244 2110 23279 2129
rect 23191 2109 23279 2110
rect 23299 2109 23307 2129
rect 23163 2101 23307 2109
rect 23163 2100 23199 2101
rect 23271 2100 23307 2101
rect 23373 2134 23410 2135
rect 23373 2133 23411 2134
rect 23373 2125 23437 2133
rect 23373 2105 23382 2125
rect 23402 2111 23437 2125
rect 23457 2111 23460 2131
rect 23402 2106 23460 2111
rect 23402 2105 23437 2106
rect 22842 2068 22879 2097
rect 22843 2066 22879 2068
rect 22420 2056 22456 2057
rect 22268 2026 22277 2046
rect 22297 2026 22305 2046
rect 22268 2016 22305 2026
rect 22364 2046 22512 2056
rect 22612 2053 22708 2055
rect 22364 2026 22373 2046
rect 22393 2026 22483 2046
rect 22503 2026 22512 2046
rect 22364 2017 22512 2026
rect 22570 2046 22708 2053
rect 22570 2026 22579 2046
rect 22599 2026 22708 2046
rect 22843 2044 23034 2066
rect 23060 2065 23097 2097
rect 23373 2093 23437 2105
rect 23477 2067 23504 2245
rect 24109 2244 24142 2577
rect 24206 2609 24374 2610
rect 24500 2609 24540 2833
rect 25003 2837 25171 2838
rect 25407 2837 25448 2871
rect 25805 2850 25852 2871
rect 25003 2827 25448 2837
rect 25520 2835 25663 2836
rect 25003 2811 25447 2827
rect 25003 2809 25171 2811
rect 25367 2810 25447 2811
rect 25520 2810 25665 2835
rect 25807 2810 25852 2850
rect 25003 2631 25030 2809
rect 25070 2771 25134 2783
rect 25410 2779 25447 2810
rect 25628 2779 25665 2810
rect 25810 2803 25852 2810
rect 26255 2868 26297 2875
rect 26442 2868 26479 2899
rect 26660 2868 26697 2899
rect 26973 2895 27037 2907
rect 27077 2869 27104 3047
rect 26255 2828 26300 2868
rect 26442 2843 26587 2868
rect 26660 2867 26740 2868
rect 26936 2867 27104 2869
rect 26660 2851 27104 2867
rect 26444 2842 26587 2843
rect 26659 2841 27104 2851
rect 26255 2807 26302 2828
rect 26659 2807 26700 2841
rect 26936 2840 27104 2841
rect 27567 2845 27607 3069
rect 27733 3068 27901 3069
rect 27965 3101 27998 3434
rect 27965 3093 28002 3101
rect 27965 3074 27973 3093
rect 27994 3074 28002 3093
rect 27965 3068 28002 3074
rect 27567 2823 27575 2845
rect 27599 2823 27607 2845
rect 27567 2815 27607 2823
rect 25070 2770 25105 2771
rect 25047 2765 25105 2770
rect 25047 2745 25050 2765
rect 25070 2751 25105 2765
rect 25125 2751 25134 2771
rect 25070 2743 25134 2751
rect 25096 2742 25134 2743
rect 25097 2741 25134 2742
rect 25200 2775 25236 2776
rect 25308 2775 25344 2776
rect 25200 2767 25344 2775
rect 25200 2747 25208 2767
rect 25228 2763 25316 2767
rect 25228 2747 25272 2763
rect 25200 2743 25272 2747
rect 25292 2747 25316 2763
rect 25336 2747 25344 2767
rect 25292 2743 25344 2747
rect 25200 2741 25344 2743
rect 25410 2771 25448 2779
rect 25526 2775 25562 2776
rect 25410 2751 25419 2771
rect 25439 2751 25448 2771
rect 25410 2742 25448 2751
rect 25477 2767 25562 2775
rect 25477 2747 25534 2767
rect 25554 2747 25562 2767
rect 25410 2741 25447 2742
rect 25477 2741 25562 2747
rect 25628 2771 25666 2779
rect 25628 2751 25637 2771
rect 25657 2751 25666 2771
rect 25628 2742 25666 2751
rect 25810 2776 25853 2803
rect 25810 2758 25824 2776
rect 25842 2758 25853 2776
rect 25810 2750 25853 2758
rect 25815 2748 25853 2750
rect 26255 2777 26700 2807
rect 27738 2790 27803 2791
rect 26255 2774 26678 2777
rect 25628 2741 25665 2742
rect 25089 2713 25179 2719
rect 25089 2693 25105 2713
rect 25125 2711 25179 2713
rect 25125 2693 25150 2711
rect 25089 2691 25150 2693
rect 25170 2691 25179 2711
rect 25089 2685 25179 2691
rect 25102 2631 25139 2632
rect 25198 2631 25235 2632
rect 25254 2631 25290 2741
rect 25477 2720 25508 2741
rect 26255 2726 26302 2774
rect 25473 2719 25508 2720
rect 25351 2709 25508 2719
rect 25351 2689 25368 2709
rect 25388 2689 25508 2709
rect 25351 2682 25508 2689
rect 25575 2712 25724 2720
rect 25575 2692 25586 2712
rect 25606 2692 25645 2712
rect 25665 2692 25724 2712
rect 26255 2708 26265 2726
rect 26283 2708 26302 2726
rect 26255 2704 26302 2708
rect 27389 2765 27576 2789
rect 27607 2770 28000 2790
rect 28020 2770 28023 2790
rect 27607 2765 28023 2770
rect 26256 2699 26293 2704
rect 25575 2685 25724 2692
rect 27389 2694 27426 2765
rect 27607 2764 27948 2765
rect 27541 2704 27572 2705
rect 25575 2684 25616 2685
rect 25812 2683 25849 2686
rect 25309 2631 25346 2632
rect 25002 2622 25140 2631
rect 24206 2583 24650 2609
rect 24206 2581 24374 2583
rect 24206 2403 24233 2581
rect 24273 2543 24337 2555
rect 24613 2551 24650 2583
rect 24676 2582 24867 2604
rect 25002 2602 25111 2622
rect 25131 2602 25140 2622
rect 25002 2595 25140 2602
rect 25198 2622 25346 2631
rect 25198 2602 25207 2622
rect 25227 2602 25317 2622
rect 25337 2602 25346 2622
rect 25002 2593 25098 2595
rect 25198 2592 25346 2602
rect 25405 2622 25442 2632
rect 25405 2602 25413 2622
rect 25433 2602 25442 2622
rect 25254 2591 25290 2592
rect 24831 2580 24867 2582
rect 24831 2551 24868 2580
rect 24273 2542 24308 2543
rect 24250 2537 24308 2542
rect 24250 2517 24253 2537
rect 24273 2523 24308 2537
rect 24328 2523 24337 2543
rect 24273 2517 24337 2523
rect 24250 2515 24337 2517
rect 24250 2511 24277 2515
rect 24299 2514 24337 2515
rect 24300 2513 24337 2514
rect 24403 2547 24439 2548
rect 24511 2547 24547 2548
rect 24403 2540 24547 2547
rect 24403 2539 24465 2540
rect 24403 2519 24411 2539
rect 24431 2522 24465 2539
rect 24484 2539 24547 2540
rect 24484 2522 24519 2539
rect 24431 2519 24519 2522
rect 24539 2519 24547 2539
rect 24403 2513 24547 2519
rect 24613 2543 24651 2551
rect 24729 2547 24765 2548
rect 24613 2523 24622 2543
rect 24642 2523 24651 2543
rect 24613 2514 24651 2523
rect 24680 2539 24765 2547
rect 24680 2519 24737 2539
rect 24757 2519 24765 2539
rect 24613 2513 24650 2514
rect 24680 2513 24765 2519
rect 24831 2543 24869 2551
rect 24831 2523 24840 2543
rect 24860 2523 24869 2543
rect 25102 2532 25139 2533
rect 25405 2532 25442 2602
rect 25477 2631 25508 2682
rect 25804 2677 25849 2683
rect 25804 2659 25822 2677
rect 25840 2659 25849 2677
rect 27389 2674 27398 2694
rect 27418 2674 27426 2694
rect 27389 2664 27426 2674
rect 27485 2694 27572 2704
rect 27485 2674 27494 2694
rect 27514 2674 27572 2694
rect 27485 2665 27572 2674
rect 27485 2664 27522 2665
rect 25804 2649 25849 2659
rect 25527 2631 25564 2632
rect 25477 2622 25564 2631
rect 25477 2602 25535 2622
rect 25555 2602 25564 2622
rect 25477 2592 25564 2602
rect 25623 2622 25660 2632
rect 25623 2602 25631 2622
rect 25651 2602 25660 2622
rect 25804 2607 25847 2649
rect 26244 2637 26296 2639
rect 25710 2605 25847 2607
rect 25477 2591 25508 2592
rect 25623 2532 25660 2602
rect 25101 2531 25442 2532
rect 24831 2514 24869 2523
rect 25026 2526 25442 2531
rect 24831 2513 24868 2514
rect 24292 2485 24382 2491
rect 24292 2465 24308 2485
rect 24328 2483 24382 2485
rect 24328 2465 24353 2483
rect 24292 2463 24353 2465
rect 24373 2463 24382 2483
rect 24292 2457 24382 2463
rect 24305 2403 24342 2404
rect 24401 2403 24438 2404
rect 24457 2403 24493 2513
rect 24680 2492 24711 2513
rect 25026 2506 25029 2526
rect 25049 2506 25442 2526
rect 25626 2516 25660 2532
rect 25704 2584 25847 2605
rect 26242 2633 26675 2637
rect 26242 2627 26681 2633
rect 26242 2609 26263 2627
rect 26281 2609 26681 2627
rect 27541 2614 27572 2665
rect 27607 2694 27644 2764
rect 27910 2763 27947 2764
rect 27759 2704 27795 2705
rect 27607 2674 27616 2694
rect 27636 2674 27644 2694
rect 27607 2664 27644 2674
rect 27703 2694 27851 2704
rect 27951 2701 28047 2703
rect 27703 2674 27712 2694
rect 27732 2674 27822 2694
rect 27842 2674 27851 2694
rect 27703 2665 27851 2674
rect 27909 2694 28047 2701
rect 27909 2674 27918 2694
rect 27938 2674 28047 2694
rect 27909 2665 28047 2674
rect 27703 2664 27740 2665
rect 27433 2611 27474 2612
rect 26242 2591 26681 2609
rect 25402 2497 25442 2506
rect 25704 2497 25731 2584
rect 25804 2558 25847 2584
rect 25804 2540 25817 2558
rect 25835 2540 25847 2558
rect 25804 2529 25847 2540
rect 24676 2491 24711 2492
rect 24554 2481 24711 2491
rect 24554 2461 24571 2481
rect 24591 2461 24711 2481
rect 24554 2454 24711 2461
rect 24778 2484 24924 2492
rect 24778 2464 24789 2484
rect 24809 2464 24848 2484
rect 24868 2464 24924 2484
rect 25402 2480 25731 2497
rect 25402 2479 25442 2480
rect 24778 2457 24924 2464
rect 25799 2468 25839 2471
rect 25799 2462 25842 2468
rect 25424 2459 25842 2462
rect 24778 2456 24819 2457
rect 24512 2403 24549 2404
rect 24205 2394 24343 2403
rect 24205 2374 24314 2394
rect 24334 2374 24343 2394
rect 24205 2367 24343 2374
rect 24401 2394 24549 2403
rect 24401 2374 24410 2394
rect 24430 2374 24520 2394
rect 24540 2374 24549 2394
rect 24205 2365 24301 2367
rect 24401 2364 24549 2374
rect 24608 2394 24645 2404
rect 24608 2374 24616 2394
rect 24636 2374 24645 2394
rect 24457 2363 24493 2364
rect 24305 2304 24342 2305
rect 24608 2304 24645 2374
rect 24680 2403 24711 2454
rect 25424 2441 25815 2459
rect 25833 2441 25842 2459
rect 25424 2439 25842 2441
rect 25424 2431 25451 2439
rect 25692 2436 25842 2439
rect 25004 2425 25172 2426
rect 25423 2425 25451 2431
rect 25004 2409 25451 2425
rect 25799 2431 25842 2436
rect 24730 2403 24767 2404
rect 24680 2394 24767 2403
rect 24680 2374 24738 2394
rect 24758 2374 24767 2394
rect 24680 2364 24767 2374
rect 24826 2394 24863 2404
rect 24826 2374 24834 2394
rect 24854 2374 24863 2394
rect 24680 2363 24711 2364
rect 24304 2303 24645 2304
rect 24826 2303 24863 2374
rect 24229 2298 24645 2303
rect 24229 2278 24232 2298
rect 24252 2278 24645 2298
rect 24676 2279 24863 2303
rect 25004 2399 25448 2409
rect 25004 2397 25172 2399
rect 24104 2199 24146 2244
rect 25004 2219 25031 2397
rect 25071 2359 25135 2371
rect 25411 2367 25448 2399
rect 25474 2398 25665 2420
rect 25629 2396 25665 2398
rect 25629 2367 25666 2396
rect 25799 2375 25839 2431
rect 25071 2358 25106 2359
rect 25048 2353 25106 2358
rect 25048 2333 25051 2353
rect 25071 2339 25106 2353
rect 25126 2339 25135 2359
rect 25071 2331 25135 2339
rect 25097 2330 25135 2331
rect 25098 2329 25135 2330
rect 25201 2363 25237 2364
rect 25309 2363 25345 2364
rect 25201 2355 25345 2363
rect 25201 2335 25209 2355
rect 25229 2335 25264 2355
rect 25284 2335 25317 2355
rect 25337 2335 25345 2355
rect 25201 2329 25345 2335
rect 25411 2359 25449 2367
rect 25527 2363 25563 2364
rect 25411 2339 25420 2359
rect 25440 2339 25449 2359
rect 25411 2330 25449 2339
rect 25478 2355 25563 2363
rect 25478 2335 25535 2355
rect 25555 2335 25563 2355
rect 25411 2329 25448 2330
rect 25478 2329 25563 2335
rect 25629 2359 25667 2367
rect 25629 2339 25638 2359
rect 25658 2339 25667 2359
rect 25799 2357 25811 2375
rect 25829 2357 25839 2375
rect 26244 2402 26296 2591
rect 26642 2566 26681 2591
rect 27325 2604 27474 2611
rect 27325 2584 27384 2604
rect 27404 2584 27443 2604
rect 27463 2584 27474 2604
rect 27325 2576 27474 2584
rect 27541 2607 27698 2614
rect 27541 2587 27661 2607
rect 27681 2587 27698 2607
rect 27541 2577 27698 2587
rect 27541 2576 27576 2577
rect 26426 2541 26613 2565
rect 26642 2546 27037 2566
rect 27057 2546 27060 2566
rect 27541 2555 27572 2576
rect 27759 2555 27795 2665
rect 27814 2664 27851 2665
rect 27910 2664 27947 2665
rect 27870 2605 27960 2611
rect 27870 2585 27879 2605
rect 27899 2603 27960 2605
rect 27899 2585 27924 2603
rect 27870 2583 27924 2585
rect 27944 2583 27960 2603
rect 27870 2577 27960 2583
rect 27384 2554 27421 2555
rect 26642 2541 27060 2546
rect 27383 2545 27421 2554
rect 26426 2470 26463 2541
rect 26642 2540 26985 2541
rect 26642 2537 26681 2540
rect 26947 2539 26984 2540
rect 26578 2480 26609 2481
rect 26426 2450 26435 2470
rect 26455 2450 26463 2470
rect 26426 2440 26463 2450
rect 26522 2470 26609 2480
rect 26522 2450 26531 2470
rect 26551 2450 26609 2470
rect 26522 2441 26609 2450
rect 26522 2440 26559 2441
rect 26244 2384 26260 2402
rect 26278 2384 26296 2402
rect 26578 2390 26609 2441
rect 26644 2470 26681 2537
rect 27383 2525 27392 2545
rect 27412 2525 27421 2545
rect 27383 2517 27421 2525
rect 27487 2549 27572 2555
rect 27602 2554 27639 2555
rect 27487 2529 27495 2549
rect 27515 2529 27572 2549
rect 27487 2521 27572 2529
rect 27601 2545 27639 2554
rect 27601 2525 27610 2545
rect 27630 2525 27639 2545
rect 27487 2520 27523 2521
rect 27601 2517 27639 2525
rect 27705 2553 27849 2555
rect 27705 2549 27765 2553
rect 27705 2529 27713 2549
rect 27733 2531 27765 2549
rect 27788 2549 27849 2553
rect 27788 2531 27821 2549
rect 27733 2529 27821 2531
rect 27841 2529 27849 2549
rect 27705 2521 27849 2529
rect 27705 2520 27741 2521
rect 27813 2520 27849 2521
rect 27915 2554 27952 2555
rect 27915 2553 27953 2554
rect 27915 2545 27979 2553
rect 27915 2525 27924 2545
rect 27944 2531 27979 2545
rect 27999 2531 28002 2551
rect 27944 2526 28002 2531
rect 27944 2525 27979 2526
rect 27384 2488 27421 2517
rect 27385 2486 27421 2488
rect 26796 2480 26832 2481
rect 26644 2450 26653 2470
rect 26673 2450 26681 2470
rect 26644 2440 26681 2450
rect 26740 2470 26888 2480
rect 26988 2477 27084 2479
rect 26740 2450 26749 2470
rect 26769 2450 26859 2470
rect 26879 2450 26888 2470
rect 26740 2441 26888 2450
rect 26946 2470 27084 2477
rect 26946 2450 26955 2470
rect 26975 2450 27084 2470
rect 27385 2464 27576 2486
rect 27602 2485 27639 2517
rect 27915 2513 27979 2525
rect 27602 2484 27877 2485
rect 28019 2484 28046 2665
rect 27602 2459 28046 2484
rect 28182 2490 28221 4305
rect 28523 4292 28556 4625
rect 28620 4657 28788 4658
rect 28914 4657 28954 4881
rect 29417 4885 29585 4886
rect 29826 4885 29861 4902
rect 30218 4892 30265 4903
rect 29417 4859 29861 4885
rect 29417 4857 29585 4859
rect 29781 4858 29861 4859
rect 30016 4858 30083 4884
rect 30222 4858 30265 4892
rect 29417 4679 29444 4857
rect 29484 4819 29548 4831
rect 29824 4827 29861 4858
rect 30042 4827 30079 4858
rect 30224 4833 30265 4858
rect 30656 4917 30697 4942
rect 30842 4917 30879 4948
rect 31060 4917 31097 4948
rect 31373 4944 31437 4956
rect 31477 4918 31504 5096
rect 30656 4883 30699 4917
rect 30838 4891 30905 4917
rect 31060 4916 31140 4917
rect 31336 4916 31504 4918
rect 31060 4890 31504 4916
rect 30656 4872 30703 4883
rect 31060 4873 31095 4890
rect 31336 4889 31504 4890
rect 31967 4894 32007 5118
rect 32133 5117 32301 5118
rect 32365 5150 32398 5483
rect 32700 5470 32739 7285
rect 32875 7291 33319 7316
rect 32875 7110 32902 7291
rect 33044 7290 33319 7291
rect 32942 7250 33006 7262
rect 33282 7258 33319 7290
rect 33345 7289 33536 7311
rect 33837 7305 33946 7325
rect 33966 7305 33975 7325
rect 33837 7298 33975 7305
rect 34033 7325 34181 7334
rect 34033 7305 34042 7325
rect 34062 7305 34152 7325
rect 34172 7305 34181 7325
rect 33837 7296 33933 7298
rect 34033 7295 34181 7305
rect 34240 7325 34277 7335
rect 34240 7305 34248 7325
rect 34268 7305 34277 7325
rect 34089 7294 34125 7295
rect 33500 7287 33536 7289
rect 33500 7258 33537 7287
rect 32942 7249 32977 7250
rect 32919 7244 32977 7249
rect 32919 7224 32922 7244
rect 32942 7230 32977 7244
rect 32997 7230 33006 7250
rect 32942 7222 33006 7230
rect 32968 7221 33006 7222
rect 32969 7220 33006 7221
rect 33072 7254 33108 7255
rect 33180 7254 33216 7255
rect 33072 7246 33216 7254
rect 33072 7226 33080 7246
rect 33100 7244 33188 7246
rect 33100 7226 33133 7244
rect 33072 7222 33133 7226
rect 33156 7226 33188 7244
rect 33208 7226 33216 7246
rect 33156 7222 33216 7226
rect 33072 7220 33216 7222
rect 33282 7250 33320 7258
rect 33398 7254 33434 7255
rect 33282 7230 33291 7250
rect 33311 7230 33320 7250
rect 33282 7221 33320 7230
rect 33349 7246 33434 7254
rect 33349 7226 33406 7246
rect 33426 7226 33434 7246
rect 33282 7220 33319 7221
rect 33349 7220 33434 7226
rect 33500 7250 33538 7258
rect 33500 7230 33509 7250
rect 33529 7230 33538 7250
rect 34240 7238 34277 7305
rect 34312 7334 34343 7385
rect 34625 7373 34643 7391
rect 34661 7373 34677 7391
rect 34362 7334 34399 7335
rect 34312 7325 34399 7334
rect 34312 7305 34370 7325
rect 34390 7305 34399 7325
rect 34312 7295 34399 7305
rect 34458 7325 34495 7335
rect 34458 7305 34466 7325
rect 34486 7305 34495 7325
rect 34312 7294 34343 7295
rect 33937 7235 33974 7236
rect 34240 7235 34279 7238
rect 33936 7234 34279 7235
rect 34458 7234 34495 7305
rect 33500 7221 33538 7230
rect 33861 7229 34279 7234
rect 33500 7220 33537 7221
rect 32961 7192 33051 7198
rect 32961 7172 32977 7192
rect 32997 7190 33051 7192
rect 32997 7172 33022 7190
rect 32961 7170 33022 7172
rect 33042 7170 33051 7190
rect 32961 7164 33051 7170
rect 32974 7110 33011 7111
rect 33070 7110 33107 7111
rect 33126 7110 33162 7220
rect 33349 7199 33380 7220
rect 33861 7209 33864 7229
rect 33884 7209 34279 7229
rect 34308 7210 34495 7234
rect 33345 7198 33380 7199
rect 33223 7188 33380 7198
rect 33223 7168 33240 7188
rect 33260 7168 33380 7188
rect 33223 7161 33380 7168
rect 33447 7191 33596 7199
rect 33447 7171 33458 7191
rect 33478 7171 33517 7191
rect 33537 7171 33596 7191
rect 33447 7164 33596 7171
rect 34240 7184 34279 7209
rect 34625 7184 34677 7373
rect 34240 7166 34679 7184
rect 33447 7163 33488 7164
rect 33181 7110 33218 7111
rect 32874 7101 33012 7110
rect 32874 7081 32983 7101
rect 33003 7081 33012 7101
rect 32874 7074 33012 7081
rect 33070 7101 33218 7110
rect 33070 7081 33079 7101
rect 33099 7081 33189 7101
rect 33209 7081 33218 7101
rect 32874 7072 32970 7074
rect 33070 7071 33218 7081
rect 33277 7101 33314 7111
rect 33277 7081 33285 7101
rect 33305 7081 33314 7101
rect 33126 7070 33162 7071
rect 32974 7011 33011 7012
rect 33277 7011 33314 7081
rect 33349 7110 33380 7161
rect 34240 7148 34640 7166
rect 34658 7148 34679 7166
rect 34240 7142 34679 7148
rect 34246 7138 34679 7142
rect 34625 7136 34677 7138
rect 33399 7110 33436 7111
rect 33349 7101 33436 7110
rect 33349 7081 33407 7101
rect 33427 7081 33436 7101
rect 33349 7071 33436 7081
rect 33495 7101 33532 7111
rect 33495 7081 33503 7101
rect 33523 7081 33532 7101
rect 33349 7070 33380 7071
rect 32973 7010 33314 7011
rect 33495 7010 33532 7081
rect 34628 7071 34665 7076
rect 32898 7005 33314 7010
rect 32898 6985 32901 7005
rect 32921 6985 33314 7005
rect 33345 6986 33532 7010
rect 34619 7067 34666 7071
rect 34619 7049 34638 7067
rect 34656 7049 34666 7067
rect 34619 7001 34666 7049
rect 34243 6998 34666 7001
rect 33118 6984 33183 6985
rect 34221 6968 34666 6998
rect 33314 6952 33354 6960
rect 33314 6930 33322 6952
rect 33346 6930 33354 6952
rect 32919 6701 32956 6707
rect 32919 6682 32927 6701
rect 32948 6682 32956 6701
rect 32919 6674 32956 6682
rect 32923 6341 32956 6674
rect 33020 6706 33188 6707
rect 33314 6706 33354 6930
rect 33817 6934 33985 6935
rect 34221 6934 34262 6968
rect 34619 6947 34666 6968
rect 33817 6924 34262 6934
rect 34334 6932 34477 6933
rect 33817 6908 34261 6924
rect 33817 6906 33985 6908
rect 34181 6907 34261 6908
rect 34334 6907 34479 6932
rect 34621 6907 34666 6947
rect 33817 6728 33844 6906
rect 33884 6868 33948 6880
rect 34224 6876 34261 6907
rect 34442 6876 34479 6907
rect 34624 6900 34666 6907
rect 33884 6867 33919 6868
rect 33861 6862 33919 6867
rect 33861 6842 33864 6862
rect 33884 6848 33919 6862
rect 33939 6848 33948 6868
rect 33884 6840 33948 6848
rect 33910 6839 33948 6840
rect 33911 6838 33948 6839
rect 34014 6872 34050 6873
rect 34122 6872 34158 6873
rect 34014 6864 34158 6872
rect 34014 6844 34022 6864
rect 34042 6860 34130 6864
rect 34042 6844 34086 6860
rect 34014 6840 34086 6844
rect 34106 6844 34130 6860
rect 34150 6844 34158 6864
rect 34106 6840 34158 6844
rect 34014 6838 34158 6840
rect 34224 6868 34262 6876
rect 34340 6872 34376 6873
rect 34224 6848 34233 6868
rect 34253 6848 34262 6868
rect 34224 6839 34262 6848
rect 34291 6864 34376 6872
rect 34291 6844 34348 6864
rect 34368 6844 34376 6864
rect 34224 6838 34261 6839
rect 34291 6838 34376 6844
rect 34442 6868 34480 6876
rect 34442 6848 34451 6868
rect 34471 6848 34480 6868
rect 34442 6839 34480 6848
rect 34624 6873 34667 6900
rect 34624 6855 34638 6873
rect 34656 6855 34667 6873
rect 34624 6847 34667 6855
rect 34629 6845 34667 6847
rect 34442 6838 34479 6839
rect 33903 6810 33993 6816
rect 33903 6790 33919 6810
rect 33939 6808 33993 6810
rect 33939 6790 33964 6808
rect 33903 6788 33964 6790
rect 33984 6788 33993 6808
rect 33903 6782 33993 6788
rect 33916 6728 33953 6729
rect 34012 6728 34049 6729
rect 34068 6728 34104 6838
rect 34291 6817 34322 6838
rect 34287 6816 34322 6817
rect 34165 6806 34322 6816
rect 34165 6786 34182 6806
rect 34202 6786 34322 6806
rect 34165 6779 34322 6786
rect 34389 6809 34538 6817
rect 34389 6789 34400 6809
rect 34420 6789 34459 6809
rect 34479 6789 34538 6809
rect 34389 6782 34538 6789
rect 34389 6781 34430 6782
rect 34626 6780 34663 6783
rect 34123 6728 34160 6729
rect 33816 6719 33954 6728
rect 33020 6680 33464 6706
rect 33020 6678 33188 6680
rect 33020 6500 33047 6678
rect 33087 6640 33151 6652
rect 33427 6648 33464 6680
rect 33490 6679 33681 6701
rect 33816 6699 33925 6719
rect 33945 6699 33954 6719
rect 33816 6692 33954 6699
rect 34012 6719 34160 6728
rect 34012 6699 34021 6719
rect 34041 6699 34131 6719
rect 34151 6699 34160 6719
rect 33816 6690 33912 6692
rect 34012 6689 34160 6699
rect 34219 6719 34256 6729
rect 34219 6699 34227 6719
rect 34247 6699 34256 6719
rect 34068 6688 34104 6689
rect 33645 6677 33681 6679
rect 33645 6648 33682 6677
rect 33087 6639 33122 6640
rect 33064 6634 33122 6639
rect 33064 6614 33067 6634
rect 33087 6620 33122 6634
rect 33142 6620 33151 6640
rect 33087 6614 33151 6620
rect 33064 6612 33151 6614
rect 33064 6608 33091 6612
rect 33113 6611 33151 6612
rect 33114 6610 33151 6611
rect 33217 6644 33253 6645
rect 33325 6644 33361 6645
rect 33217 6637 33361 6644
rect 33217 6636 33279 6637
rect 33217 6616 33225 6636
rect 33245 6619 33279 6636
rect 33298 6636 33361 6637
rect 33298 6619 33333 6636
rect 33245 6616 33333 6619
rect 33353 6616 33361 6636
rect 33217 6610 33361 6616
rect 33427 6640 33465 6648
rect 33543 6644 33579 6645
rect 33427 6620 33436 6640
rect 33456 6620 33465 6640
rect 33427 6611 33465 6620
rect 33494 6636 33579 6644
rect 33494 6616 33551 6636
rect 33571 6616 33579 6636
rect 33427 6610 33464 6611
rect 33494 6610 33579 6616
rect 33645 6640 33683 6648
rect 33645 6620 33654 6640
rect 33674 6620 33683 6640
rect 33916 6629 33953 6630
rect 34219 6629 34256 6699
rect 34291 6728 34322 6779
rect 34618 6774 34663 6780
rect 34618 6756 34636 6774
rect 34654 6756 34663 6774
rect 34618 6746 34663 6756
rect 34341 6728 34378 6729
rect 34291 6719 34378 6728
rect 34291 6699 34349 6719
rect 34369 6699 34378 6719
rect 34291 6689 34378 6699
rect 34437 6719 34474 6729
rect 34437 6699 34445 6719
rect 34465 6699 34474 6719
rect 34618 6704 34661 6746
rect 34524 6702 34661 6704
rect 34291 6688 34322 6689
rect 34437 6629 34474 6699
rect 33915 6628 34256 6629
rect 33645 6611 33683 6620
rect 33840 6623 34256 6628
rect 33645 6610 33682 6611
rect 33106 6582 33196 6588
rect 33106 6562 33122 6582
rect 33142 6580 33196 6582
rect 33142 6562 33167 6580
rect 33106 6560 33167 6562
rect 33187 6560 33196 6580
rect 33106 6554 33196 6560
rect 33119 6500 33156 6501
rect 33215 6500 33252 6501
rect 33271 6500 33307 6610
rect 33494 6589 33525 6610
rect 33840 6603 33843 6623
rect 33863 6603 34256 6623
rect 34440 6613 34474 6629
rect 34518 6681 34661 6702
rect 34216 6594 34256 6603
rect 34518 6594 34545 6681
rect 34618 6655 34661 6681
rect 34618 6637 34631 6655
rect 34649 6637 34661 6655
rect 34618 6626 34661 6637
rect 33490 6588 33525 6589
rect 33368 6578 33525 6588
rect 33368 6558 33385 6578
rect 33405 6558 33525 6578
rect 33368 6551 33525 6558
rect 33592 6581 33738 6589
rect 33592 6561 33603 6581
rect 33623 6561 33662 6581
rect 33682 6561 33738 6581
rect 34216 6577 34545 6594
rect 34216 6576 34256 6577
rect 33592 6554 33738 6561
rect 34613 6565 34653 6568
rect 34613 6559 34656 6565
rect 34238 6556 34656 6559
rect 33592 6553 33633 6554
rect 33326 6500 33363 6501
rect 33019 6491 33157 6500
rect 33019 6471 33128 6491
rect 33148 6471 33157 6491
rect 33019 6464 33157 6471
rect 33215 6491 33363 6500
rect 33215 6471 33224 6491
rect 33244 6471 33334 6491
rect 33354 6471 33363 6491
rect 33019 6462 33115 6464
rect 33215 6461 33363 6471
rect 33422 6491 33459 6501
rect 33422 6471 33430 6491
rect 33450 6471 33459 6491
rect 33271 6460 33307 6461
rect 33119 6401 33156 6402
rect 33422 6401 33459 6471
rect 33494 6500 33525 6551
rect 34238 6538 34629 6556
rect 34647 6538 34656 6556
rect 34238 6536 34656 6538
rect 34238 6528 34265 6536
rect 34506 6533 34656 6536
rect 33818 6522 33986 6523
rect 34237 6522 34265 6528
rect 33818 6506 34265 6522
rect 34613 6528 34656 6533
rect 33544 6500 33581 6501
rect 33494 6491 33581 6500
rect 33494 6471 33552 6491
rect 33572 6471 33581 6491
rect 33494 6461 33581 6471
rect 33640 6491 33677 6501
rect 33640 6471 33648 6491
rect 33668 6471 33677 6491
rect 33494 6460 33525 6461
rect 33118 6400 33459 6401
rect 33640 6400 33677 6471
rect 33043 6395 33459 6400
rect 33043 6375 33046 6395
rect 33066 6375 33459 6395
rect 33490 6376 33677 6400
rect 33818 6496 34262 6506
rect 33818 6494 33986 6496
rect 32918 6296 32960 6341
rect 33818 6316 33845 6494
rect 33885 6456 33949 6468
rect 34225 6464 34262 6496
rect 34288 6495 34479 6517
rect 34443 6493 34479 6495
rect 34443 6464 34480 6493
rect 34613 6472 34653 6528
rect 33885 6455 33920 6456
rect 33862 6450 33920 6455
rect 33862 6430 33865 6450
rect 33885 6436 33920 6450
rect 33940 6436 33949 6456
rect 33885 6428 33949 6436
rect 33911 6427 33949 6428
rect 33912 6426 33949 6427
rect 34015 6460 34051 6461
rect 34123 6460 34159 6461
rect 34015 6452 34159 6460
rect 34015 6432 34023 6452
rect 34043 6432 34078 6452
rect 34098 6432 34131 6452
rect 34151 6432 34159 6452
rect 34015 6426 34159 6432
rect 34225 6456 34263 6464
rect 34341 6460 34377 6461
rect 34225 6436 34234 6456
rect 34254 6436 34263 6456
rect 34225 6427 34263 6436
rect 34292 6452 34377 6460
rect 34292 6432 34349 6452
rect 34369 6432 34377 6452
rect 34225 6426 34262 6427
rect 34292 6426 34377 6432
rect 34443 6456 34481 6464
rect 34443 6436 34452 6456
rect 34472 6436 34481 6456
rect 34613 6454 34625 6472
rect 34643 6454 34653 6472
rect 34613 6444 34653 6454
rect 34443 6427 34481 6436
rect 34443 6426 34480 6427
rect 33904 6398 33994 6404
rect 33904 6378 33920 6398
rect 33940 6396 33994 6398
rect 33940 6378 33965 6396
rect 33904 6376 33965 6378
rect 33985 6376 33994 6396
rect 33904 6370 33994 6376
rect 33917 6316 33954 6317
rect 34013 6316 34050 6317
rect 34069 6316 34105 6426
rect 34292 6405 34323 6426
rect 34288 6404 34323 6405
rect 34166 6394 34323 6404
rect 34166 6374 34183 6394
rect 34203 6374 34323 6394
rect 34166 6367 34323 6374
rect 34390 6397 34539 6405
rect 34390 6377 34401 6397
rect 34421 6377 34460 6397
rect 34480 6377 34539 6397
rect 34390 6370 34539 6377
rect 34605 6373 34657 6391
rect 34390 6369 34431 6370
rect 34124 6316 34161 6317
rect 33817 6307 33955 6316
rect 33289 6296 33322 6298
rect 32918 6284 33365 6296
rect 32921 6270 33365 6284
rect 32921 6268 33089 6270
rect 32921 6090 32948 6268
rect 32988 6230 33052 6242
rect 33328 6238 33365 6270
rect 33391 6269 33582 6291
rect 33817 6287 33926 6307
rect 33946 6287 33955 6307
rect 33817 6280 33955 6287
rect 34013 6307 34161 6316
rect 34013 6287 34022 6307
rect 34042 6287 34132 6307
rect 34152 6287 34161 6307
rect 33817 6278 33913 6280
rect 34013 6277 34161 6287
rect 34220 6307 34257 6317
rect 34220 6287 34228 6307
rect 34248 6287 34257 6307
rect 34069 6276 34105 6277
rect 33546 6267 33582 6269
rect 33546 6238 33583 6267
rect 32988 6229 33023 6230
rect 32965 6224 33023 6229
rect 32965 6204 32968 6224
rect 32988 6210 33023 6224
rect 33043 6210 33052 6230
rect 32988 6202 33052 6210
rect 33014 6201 33052 6202
rect 33015 6200 33052 6201
rect 33118 6234 33154 6235
rect 33226 6234 33262 6235
rect 33118 6226 33262 6234
rect 33118 6206 33126 6226
rect 33146 6224 33234 6226
rect 33146 6206 33179 6224
rect 33118 6205 33179 6206
rect 33200 6206 33234 6224
rect 33254 6206 33262 6226
rect 33200 6205 33262 6206
rect 33118 6200 33262 6205
rect 33328 6230 33366 6238
rect 33444 6234 33480 6235
rect 33328 6210 33337 6230
rect 33357 6210 33366 6230
rect 33328 6201 33366 6210
rect 33395 6226 33480 6234
rect 33395 6206 33452 6226
rect 33472 6206 33480 6226
rect 33328 6200 33365 6201
rect 33395 6200 33480 6206
rect 33546 6230 33584 6238
rect 33546 6210 33555 6230
rect 33575 6210 33584 6230
rect 34220 6220 34257 6287
rect 34292 6316 34323 6367
rect 34605 6355 34623 6373
rect 34641 6355 34657 6373
rect 34342 6316 34379 6317
rect 34292 6307 34379 6316
rect 34292 6287 34350 6307
rect 34370 6287 34379 6307
rect 34292 6277 34379 6287
rect 34438 6307 34475 6317
rect 34438 6287 34446 6307
rect 34466 6287 34475 6307
rect 34292 6276 34323 6277
rect 33917 6217 33954 6218
rect 34220 6217 34259 6220
rect 33916 6216 34259 6217
rect 34438 6216 34475 6287
rect 33546 6201 33584 6210
rect 33841 6211 34259 6216
rect 33546 6200 33583 6201
rect 33007 6172 33097 6178
rect 33007 6152 33023 6172
rect 33043 6170 33097 6172
rect 33043 6152 33068 6170
rect 33007 6150 33068 6152
rect 33088 6150 33097 6170
rect 33007 6144 33097 6150
rect 33020 6090 33057 6091
rect 33116 6090 33153 6091
rect 33172 6090 33208 6200
rect 33395 6179 33426 6200
rect 33841 6191 33844 6211
rect 33864 6191 34259 6211
rect 34288 6192 34475 6216
rect 33391 6178 33426 6179
rect 33269 6168 33426 6178
rect 33269 6148 33286 6168
rect 33306 6148 33426 6168
rect 33269 6141 33426 6148
rect 33493 6171 33642 6179
rect 33493 6151 33504 6171
rect 33524 6151 33563 6171
rect 33583 6151 33642 6171
rect 33493 6144 33642 6151
rect 34220 6166 34259 6191
rect 34605 6166 34657 6355
rect 34220 6148 34659 6166
rect 33493 6143 33534 6144
rect 33227 6090 33264 6091
rect 32920 6081 33058 6090
rect 32920 6061 33029 6081
rect 33049 6061 33058 6081
rect 32920 6054 33058 6061
rect 33116 6081 33264 6090
rect 33116 6061 33125 6081
rect 33145 6061 33235 6081
rect 33255 6061 33264 6081
rect 32920 6052 33016 6054
rect 33116 6051 33264 6061
rect 33323 6081 33360 6091
rect 33323 6061 33331 6081
rect 33351 6061 33360 6081
rect 33172 6050 33208 6051
rect 33020 5991 33057 5992
rect 33323 5991 33360 6061
rect 33395 6090 33426 6141
rect 34220 6130 34620 6148
rect 34638 6130 34659 6148
rect 34220 6124 34659 6130
rect 34226 6120 34659 6124
rect 34605 6118 34657 6120
rect 33445 6090 33482 6091
rect 33395 6081 33482 6090
rect 33395 6061 33453 6081
rect 33473 6061 33482 6081
rect 33395 6051 33482 6061
rect 33541 6081 33578 6091
rect 33541 6061 33549 6081
rect 33569 6061 33578 6081
rect 33395 6050 33426 6051
rect 33019 5990 33360 5991
rect 33541 5990 33578 6061
rect 34608 6053 34645 6058
rect 34599 6049 34646 6053
rect 34599 6031 34618 6049
rect 34636 6031 34646 6049
rect 32944 5985 33360 5990
rect 32944 5965 32947 5985
rect 32967 5965 33360 5985
rect 33391 5966 33578 5990
rect 34203 5988 34243 5993
rect 34599 5988 34646 6031
rect 34203 5949 34646 5988
rect 33297 5934 33337 5942
rect 33297 5912 33305 5934
rect 33329 5912 33337 5934
rect 33003 5688 33171 5689
rect 33297 5688 33337 5912
rect 33800 5916 33968 5917
rect 34203 5916 34243 5949
rect 34599 5916 34646 5949
rect 33800 5915 34244 5916
rect 33800 5890 34245 5915
rect 33800 5888 33968 5890
rect 34164 5889 34245 5890
rect 34414 5889 34463 5915
rect 34599 5889 34648 5916
rect 33800 5710 33827 5888
rect 33867 5850 33931 5862
rect 34207 5858 34244 5889
rect 34425 5858 34462 5889
rect 34607 5864 34648 5889
rect 33867 5849 33902 5850
rect 33844 5844 33902 5849
rect 33844 5824 33847 5844
rect 33867 5830 33902 5844
rect 33922 5830 33931 5850
rect 33867 5822 33931 5830
rect 33893 5821 33931 5822
rect 33894 5820 33931 5821
rect 33997 5854 34033 5855
rect 34105 5854 34141 5855
rect 33997 5846 34141 5854
rect 33997 5826 34005 5846
rect 34025 5842 34113 5846
rect 34025 5826 34069 5842
rect 33997 5822 34069 5826
rect 34089 5826 34113 5842
rect 34133 5826 34141 5846
rect 34089 5822 34141 5826
rect 33997 5820 34141 5822
rect 34207 5850 34245 5858
rect 34323 5854 34359 5855
rect 34207 5830 34216 5850
rect 34236 5830 34245 5850
rect 34207 5821 34245 5830
rect 34274 5846 34359 5854
rect 34274 5826 34331 5846
rect 34351 5826 34359 5846
rect 34207 5820 34244 5821
rect 34274 5820 34359 5826
rect 34425 5850 34463 5858
rect 34425 5830 34434 5850
rect 34454 5830 34463 5850
rect 34425 5821 34463 5830
rect 34607 5855 34649 5864
rect 34607 5837 34621 5855
rect 34639 5837 34649 5855
rect 34607 5829 34649 5837
rect 34612 5827 34649 5829
rect 34425 5820 34462 5821
rect 33886 5792 33976 5798
rect 33886 5772 33902 5792
rect 33922 5790 33976 5792
rect 33922 5772 33947 5790
rect 33886 5770 33947 5772
rect 33967 5770 33976 5790
rect 33886 5764 33976 5770
rect 33899 5710 33936 5711
rect 33995 5710 34032 5711
rect 34051 5710 34087 5820
rect 34274 5799 34305 5820
rect 34270 5798 34305 5799
rect 34148 5788 34305 5798
rect 34148 5768 34165 5788
rect 34185 5768 34305 5788
rect 34148 5761 34305 5768
rect 34372 5791 34521 5799
rect 34372 5771 34383 5791
rect 34403 5771 34442 5791
rect 34462 5771 34521 5791
rect 34372 5764 34521 5771
rect 34372 5763 34413 5764
rect 34609 5762 34646 5765
rect 34106 5710 34143 5711
rect 33799 5701 33937 5710
rect 33003 5662 33447 5688
rect 33003 5660 33171 5662
rect 33003 5482 33030 5660
rect 33070 5622 33134 5634
rect 33410 5630 33447 5662
rect 33473 5661 33664 5683
rect 33799 5681 33908 5701
rect 33928 5681 33937 5701
rect 33799 5674 33937 5681
rect 33995 5701 34143 5710
rect 33995 5681 34004 5701
rect 34024 5681 34114 5701
rect 34134 5681 34143 5701
rect 33799 5672 33895 5674
rect 33995 5671 34143 5681
rect 34202 5701 34239 5711
rect 34202 5681 34210 5701
rect 34230 5681 34239 5701
rect 34051 5670 34087 5671
rect 33628 5659 33664 5661
rect 33628 5630 33665 5659
rect 33070 5621 33105 5622
rect 33047 5616 33105 5621
rect 33047 5596 33050 5616
rect 33070 5602 33105 5616
rect 33125 5602 33134 5622
rect 33070 5594 33134 5602
rect 33096 5593 33134 5594
rect 33097 5592 33134 5593
rect 33200 5626 33236 5627
rect 33308 5626 33344 5627
rect 33200 5618 33344 5626
rect 33200 5598 33208 5618
rect 33228 5617 33316 5618
rect 33228 5598 33263 5617
rect 33284 5598 33316 5617
rect 33336 5598 33344 5618
rect 33200 5592 33344 5598
rect 33410 5622 33448 5630
rect 33526 5626 33562 5627
rect 33410 5602 33419 5622
rect 33439 5602 33448 5622
rect 33410 5593 33448 5602
rect 33477 5618 33562 5626
rect 33477 5598 33534 5618
rect 33554 5598 33562 5618
rect 33410 5592 33447 5593
rect 33477 5592 33562 5598
rect 33628 5622 33666 5630
rect 33628 5602 33637 5622
rect 33657 5602 33666 5622
rect 33899 5611 33936 5612
rect 34202 5611 34239 5681
rect 34274 5710 34305 5761
rect 34601 5756 34646 5762
rect 34601 5738 34619 5756
rect 34637 5738 34646 5756
rect 34601 5728 34646 5738
rect 34324 5710 34361 5711
rect 34274 5701 34361 5710
rect 34274 5681 34332 5701
rect 34352 5681 34361 5701
rect 34274 5671 34361 5681
rect 34420 5701 34457 5711
rect 34420 5681 34428 5701
rect 34448 5681 34457 5701
rect 34601 5686 34644 5728
rect 34507 5684 34644 5686
rect 34274 5670 34305 5671
rect 34420 5611 34457 5681
rect 33898 5610 34239 5611
rect 33628 5593 33666 5602
rect 33823 5605 34239 5610
rect 33628 5592 33665 5593
rect 33089 5564 33179 5570
rect 33089 5544 33105 5564
rect 33125 5562 33179 5564
rect 33125 5544 33150 5562
rect 33089 5542 33150 5544
rect 33170 5542 33179 5562
rect 33089 5536 33179 5542
rect 33102 5482 33139 5483
rect 33198 5482 33235 5483
rect 33254 5482 33290 5592
rect 33477 5571 33508 5592
rect 33823 5585 33826 5605
rect 33846 5585 34239 5605
rect 34423 5595 34457 5611
rect 34501 5663 34644 5684
rect 34199 5576 34239 5585
rect 34501 5576 34528 5663
rect 34601 5637 34644 5663
rect 34601 5619 34614 5637
rect 34632 5619 34644 5637
rect 34601 5608 34644 5619
rect 33473 5570 33508 5571
rect 33351 5560 33508 5570
rect 33351 5540 33368 5560
rect 33388 5540 33508 5560
rect 33351 5533 33508 5540
rect 33575 5563 33724 5571
rect 33575 5543 33586 5563
rect 33606 5543 33645 5563
rect 33665 5543 33724 5563
rect 34199 5559 34528 5576
rect 34199 5558 34239 5559
rect 33575 5536 33724 5543
rect 34596 5547 34636 5550
rect 34596 5541 34639 5547
rect 34221 5538 34639 5541
rect 33575 5535 33616 5536
rect 33309 5482 33346 5483
rect 33002 5473 33140 5482
rect 32700 5298 32740 5470
rect 33002 5453 33111 5473
rect 33131 5453 33140 5473
rect 33002 5446 33140 5453
rect 33198 5473 33346 5482
rect 33198 5453 33207 5473
rect 33227 5453 33317 5473
rect 33337 5453 33346 5473
rect 33002 5444 33098 5446
rect 33198 5443 33346 5453
rect 33405 5473 33442 5483
rect 33405 5453 33413 5473
rect 33433 5453 33442 5473
rect 33254 5442 33290 5443
rect 33102 5383 33139 5384
rect 33405 5383 33442 5453
rect 33477 5482 33508 5533
rect 34221 5520 34612 5538
rect 34630 5520 34639 5538
rect 34221 5518 34639 5520
rect 34221 5510 34248 5518
rect 34489 5515 34639 5518
rect 33801 5504 33969 5505
rect 34220 5504 34248 5510
rect 33801 5488 34248 5504
rect 34596 5510 34639 5515
rect 33527 5482 33564 5483
rect 33477 5473 33564 5482
rect 33477 5453 33535 5473
rect 33555 5453 33564 5473
rect 33477 5443 33564 5453
rect 33623 5473 33660 5483
rect 33623 5453 33631 5473
rect 33651 5453 33660 5473
rect 33477 5442 33508 5443
rect 33101 5382 33442 5383
rect 33623 5382 33660 5453
rect 33026 5377 33442 5382
rect 33026 5357 33029 5377
rect 33049 5357 33442 5377
rect 33473 5358 33660 5382
rect 33801 5478 34245 5488
rect 33801 5476 33969 5478
rect 33801 5298 33828 5476
rect 33868 5438 33932 5450
rect 34208 5446 34245 5478
rect 34271 5477 34462 5499
rect 34426 5475 34462 5477
rect 34426 5446 34463 5475
rect 34596 5454 34636 5510
rect 33868 5437 33903 5438
rect 33845 5432 33903 5437
rect 33845 5412 33848 5432
rect 33868 5418 33903 5432
rect 33923 5418 33932 5438
rect 33868 5410 33932 5418
rect 33894 5409 33932 5410
rect 33895 5408 33932 5409
rect 33998 5442 34034 5443
rect 34106 5442 34142 5443
rect 33998 5434 34142 5442
rect 33998 5414 34006 5434
rect 34026 5414 34061 5434
rect 34081 5414 34114 5434
rect 34134 5414 34142 5434
rect 33998 5408 34142 5414
rect 34208 5438 34246 5446
rect 34324 5442 34360 5443
rect 34208 5418 34217 5438
rect 34237 5418 34246 5438
rect 34208 5409 34246 5418
rect 34275 5434 34360 5442
rect 34275 5414 34332 5434
rect 34352 5414 34360 5434
rect 34208 5408 34245 5409
rect 34275 5408 34360 5414
rect 34426 5438 34464 5446
rect 34426 5418 34435 5438
rect 34455 5418 34464 5438
rect 34596 5436 34608 5454
rect 34626 5436 34636 5454
rect 34596 5426 34636 5436
rect 34426 5409 34464 5418
rect 34426 5408 34463 5409
rect 33887 5380 33977 5386
rect 33887 5360 33903 5380
rect 33923 5378 33977 5380
rect 33923 5360 33948 5378
rect 33887 5358 33948 5360
rect 33968 5358 33977 5378
rect 33887 5352 33977 5358
rect 33900 5298 33937 5299
rect 33996 5298 34033 5299
rect 34052 5298 34088 5408
rect 34275 5387 34306 5408
rect 34271 5386 34306 5387
rect 34149 5376 34306 5386
rect 34149 5356 34166 5376
rect 34186 5356 34306 5376
rect 34149 5349 34306 5356
rect 34373 5379 34522 5387
rect 34373 5359 34384 5379
rect 34404 5359 34443 5379
rect 34463 5359 34522 5379
rect 34373 5352 34522 5359
rect 34588 5355 34640 5373
rect 34373 5351 34414 5352
rect 34107 5298 34144 5299
rect 32701 5283 32740 5298
rect 33800 5289 33938 5298
rect 32701 5282 32867 5283
rect 32993 5282 33033 5284
rect 32701 5256 33143 5282
rect 32701 5254 32867 5256
rect 32365 5142 32402 5150
rect 32365 5123 32373 5142
rect 32394 5123 32402 5142
rect 32365 5117 32402 5123
rect 32701 5076 32726 5254
rect 32766 5216 32830 5228
rect 33106 5224 33143 5256
rect 33169 5255 33360 5277
rect 33800 5269 33909 5289
rect 33929 5269 33938 5289
rect 33800 5262 33938 5269
rect 33996 5289 34144 5298
rect 33996 5269 34005 5289
rect 34025 5269 34115 5289
rect 34135 5269 34144 5289
rect 33800 5260 33896 5262
rect 33996 5259 34144 5269
rect 34203 5289 34240 5299
rect 34203 5269 34211 5289
rect 34231 5269 34240 5289
rect 34052 5258 34088 5259
rect 33324 5253 33360 5255
rect 33324 5224 33361 5253
rect 32766 5215 32801 5216
rect 32743 5210 32801 5215
rect 32743 5190 32746 5210
rect 32766 5196 32801 5210
rect 32821 5196 32830 5216
rect 32766 5188 32830 5196
rect 32792 5187 32830 5188
rect 32793 5186 32830 5187
rect 32896 5220 32932 5221
rect 33004 5220 33040 5221
rect 32896 5215 33040 5220
rect 32896 5212 32958 5215
rect 32896 5192 32904 5212
rect 32924 5192 32958 5212
rect 32896 5189 32958 5192
rect 32984 5212 33040 5215
rect 32984 5192 33012 5212
rect 33032 5192 33040 5212
rect 32984 5189 33040 5192
rect 32896 5186 33040 5189
rect 33106 5216 33144 5224
rect 33222 5220 33258 5221
rect 33106 5196 33115 5216
rect 33135 5196 33144 5216
rect 33106 5187 33144 5196
rect 33173 5212 33258 5220
rect 33173 5192 33230 5212
rect 33250 5192 33258 5212
rect 33106 5186 33143 5187
rect 33173 5186 33258 5192
rect 33324 5216 33362 5224
rect 33324 5196 33333 5216
rect 33353 5196 33362 5216
rect 34203 5202 34240 5269
rect 34275 5298 34306 5349
rect 34588 5337 34606 5355
rect 34624 5337 34640 5355
rect 34325 5298 34362 5299
rect 34275 5289 34362 5298
rect 34275 5269 34333 5289
rect 34353 5269 34362 5289
rect 34275 5259 34362 5269
rect 34421 5289 34458 5299
rect 34421 5269 34429 5289
rect 34449 5269 34458 5289
rect 34275 5258 34306 5259
rect 33900 5199 33937 5200
rect 34203 5199 34242 5202
rect 33899 5198 34242 5199
rect 34421 5198 34458 5269
rect 33324 5187 33362 5196
rect 33824 5193 34242 5198
rect 33324 5186 33361 5187
rect 32785 5158 32875 5164
rect 32785 5138 32801 5158
rect 32821 5156 32875 5158
rect 32821 5138 32846 5156
rect 32785 5136 32846 5138
rect 32866 5136 32875 5156
rect 32785 5130 32875 5136
rect 32798 5076 32835 5077
rect 32894 5076 32931 5077
rect 32950 5076 32986 5186
rect 33173 5165 33204 5186
rect 33824 5173 33827 5193
rect 33847 5173 34242 5193
rect 34271 5174 34458 5198
rect 33169 5164 33204 5165
rect 33047 5154 33204 5164
rect 33047 5134 33064 5154
rect 33084 5134 33204 5154
rect 33047 5127 33204 5134
rect 33271 5157 33420 5165
rect 33271 5137 33282 5157
rect 33302 5137 33341 5157
rect 33361 5137 33420 5157
rect 33271 5130 33420 5137
rect 34203 5148 34242 5173
rect 34588 5148 34640 5337
rect 34203 5130 34642 5148
rect 33271 5129 33312 5130
rect 33005 5076 33042 5077
rect 32701 5067 32836 5076
rect 32701 5047 32807 5067
rect 32827 5047 32836 5067
rect 32701 5040 32836 5047
rect 32894 5067 33042 5076
rect 32894 5047 32903 5067
rect 32923 5047 33013 5067
rect 33033 5047 33042 5067
rect 32701 5038 32794 5040
rect 32894 5037 33042 5047
rect 33101 5067 33138 5077
rect 33101 5047 33109 5067
rect 33129 5047 33138 5067
rect 32950 5036 32986 5037
rect 32798 4977 32835 4978
rect 33101 4977 33138 5047
rect 33173 5076 33204 5127
rect 34203 5112 34603 5130
rect 34621 5112 34642 5130
rect 34203 5106 34642 5112
rect 34209 5102 34642 5106
rect 34588 5100 34640 5102
rect 33223 5076 33260 5077
rect 33173 5067 33260 5076
rect 33173 5047 33231 5067
rect 33251 5047 33260 5067
rect 33173 5037 33260 5047
rect 33319 5067 33356 5077
rect 33319 5047 33327 5067
rect 33347 5047 33356 5067
rect 33173 5036 33204 5037
rect 32797 4976 33138 4977
rect 33319 4976 33356 5047
rect 34591 5035 34628 5040
rect 32722 4971 33138 4976
rect 32722 4951 32725 4971
rect 32745 4951 33138 4971
rect 33169 4952 33356 4976
rect 34582 5031 34629 5035
rect 34582 5013 34601 5031
rect 34619 5013 34629 5031
rect 34190 4954 34228 4955
rect 34582 4954 34629 5013
rect 32942 4950 33007 4951
rect 31057 4872 31095 4873
rect 30656 4834 31095 4872
rect 31967 4872 31975 4894
rect 31999 4872 32007 4894
rect 31967 4864 32007 4872
rect 33278 4916 33318 4924
rect 33278 4894 33286 4916
rect 33310 4894 33318 4916
rect 34190 4916 34629 4954
rect 34190 4915 34228 4916
rect 32278 4837 32343 4838
rect 29484 4818 29519 4819
rect 29461 4813 29519 4818
rect 29461 4793 29464 4813
rect 29484 4799 29519 4813
rect 29539 4799 29548 4819
rect 29484 4791 29548 4799
rect 29510 4790 29548 4791
rect 29511 4789 29548 4790
rect 29614 4823 29650 4824
rect 29722 4823 29758 4824
rect 29614 4815 29758 4823
rect 29614 4795 29622 4815
rect 29642 4811 29730 4815
rect 29642 4795 29686 4811
rect 29614 4791 29686 4795
rect 29706 4795 29730 4811
rect 29750 4795 29758 4815
rect 29706 4791 29758 4795
rect 29614 4789 29758 4791
rect 29824 4819 29862 4827
rect 29940 4823 29976 4824
rect 29824 4799 29833 4819
rect 29853 4799 29862 4819
rect 29824 4790 29862 4799
rect 29891 4815 29976 4823
rect 29891 4795 29948 4815
rect 29968 4795 29976 4815
rect 29824 4789 29861 4790
rect 29891 4789 29976 4795
rect 30042 4819 30080 4827
rect 30042 4799 30051 4819
rect 30071 4799 30080 4819
rect 30042 4790 30080 4799
rect 30224 4824 30266 4833
rect 30224 4806 30238 4824
rect 30256 4806 30266 4824
rect 30224 4798 30266 4806
rect 30229 4796 30266 4798
rect 30042 4789 30079 4790
rect 29503 4761 29593 4767
rect 29503 4741 29519 4761
rect 29539 4759 29593 4761
rect 29539 4741 29564 4759
rect 29503 4739 29564 4741
rect 29584 4739 29593 4759
rect 29503 4733 29593 4739
rect 29516 4679 29553 4680
rect 29612 4679 29649 4680
rect 29668 4679 29704 4789
rect 29891 4768 29922 4789
rect 30656 4775 30703 4834
rect 31057 4833 31095 4834
rect 29887 4767 29922 4768
rect 29765 4757 29922 4767
rect 29765 4737 29782 4757
rect 29802 4737 29922 4757
rect 29765 4730 29922 4737
rect 29989 4760 30138 4768
rect 29989 4740 30000 4760
rect 30020 4740 30059 4760
rect 30079 4740 30138 4760
rect 30656 4757 30666 4775
rect 30684 4757 30703 4775
rect 30656 4753 30703 4757
rect 31929 4812 32116 4836
rect 32147 4817 32540 4837
rect 32560 4817 32563 4837
rect 32147 4812 32563 4817
rect 30657 4748 30694 4753
rect 29989 4733 30138 4740
rect 31929 4741 31966 4812
rect 32147 4811 32488 4812
rect 32081 4751 32112 4752
rect 29989 4732 30030 4733
rect 30226 4731 30263 4734
rect 29723 4679 29760 4680
rect 29416 4670 29554 4679
rect 28620 4631 29064 4657
rect 28620 4629 28788 4631
rect 28620 4451 28647 4629
rect 28687 4591 28751 4603
rect 29027 4599 29064 4631
rect 29090 4630 29281 4652
rect 29416 4650 29525 4670
rect 29545 4650 29554 4670
rect 29416 4643 29554 4650
rect 29612 4670 29760 4679
rect 29612 4650 29621 4670
rect 29641 4650 29731 4670
rect 29751 4650 29760 4670
rect 29416 4641 29512 4643
rect 29612 4640 29760 4650
rect 29819 4670 29856 4680
rect 29819 4650 29827 4670
rect 29847 4650 29856 4670
rect 29668 4639 29704 4640
rect 29245 4628 29281 4630
rect 29245 4599 29282 4628
rect 28687 4590 28722 4591
rect 28664 4585 28722 4590
rect 28664 4565 28667 4585
rect 28687 4571 28722 4585
rect 28742 4571 28751 4591
rect 28687 4565 28751 4571
rect 28664 4563 28751 4565
rect 28664 4559 28691 4563
rect 28713 4562 28751 4563
rect 28714 4561 28751 4562
rect 28817 4595 28853 4596
rect 28925 4595 28961 4596
rect 28817 4588 28961 4595
rect 28817 4587 28879 4588
rect 28817 4567 28825 4587
rect 28845 4570 28879 4587
rect 28898 4587 28961 4588
rect 28898 4570 28933 4587
rect 28845 4567 28933 4570
rect 28953 4567 28961 4587
rect 28817 4561 28961 4567
rect 29027 4591 29065 4599
rect 29143 4595 29179 4596
rect 29027 4571 29036 4591
rect 29056 4571 29065 4591
rect 29027 4562 29065 4571
rect 29094 4587 29179 4595
rect 29094 4567 29151 4587
rect 29171 4567 29179 4587
rect 29027 4561 29064 4562
rect 29094 4561 29179 4567
rect 29245 4591 29283 4599
rect 29245 4571 29254 4591
rect 29274 4571 29283 4591
rect 29516 4580 29553 4581
rect 29819 4580 29856 4650
rect 29891 4679 29922 4730
rect 30218 4725 30263 4731
rect 30218 4707 30236 4725
rect 30254 4707 30263 4725
rect 31929 4721 31938 4741
rect 31958 4721 31966 4741
rect 31929 4711 31966 4721
rect 32025 4741 32112 4751
rect 32025 4721 32034 4741
rect 32054 4721 32112 4741
rect 32025 4712 32112 4721
rect 32025 4711 32062 4712
rect 30218 4697 30263 4707
rect 29941 4679 29978 4680
rect 29891 4670 29978 4679
rect 29891 4650 29949 4670
rect 29969 4650 29978 4670
rect 29891 4640 29978 4650
rect 30037 4670 30074 4680
rect 30037 4650 30045 4670
rect 30065 4650 30074 4670
rect 30218 4655 30261 4697
rect 30645 4686 30697 4688
rect 30124 4653 30261 4655
rect 29891 4639 29922 4640
rect 30037 4580 30074 4650
rect 29515 4579 29856 4580
rect 29245 4562 29283 4571
rect 29440 4574 29856 4579
rect 29245 4561 29282 4562
rect 28706 4533 28796 4539
rect 28706 4513 28722 4533
rect 28742 4531 28796 4533
rect 28742 4513 28767 4531
rect 28706 4511 28767 4513
rect 28787 4511 28796 4531
rect 28706 4505 28796 4511
rect 28719 4451 28756 4452
rect 28815 4451 28852 4452
rect 28871 4451 28907 4561
rect 29094 4540 29125 4561
rect 29440 4554 29443 4574
rect 29463 4554 29856 4574
rect 30040 4564 30074 4580
rect 30118 4632 30261 4653
rect 30643 4682 31076 4686
rect 30643 4676 31082 4682
rect 30643 4658 30664 4676
rect 30682 4658 31082 4676
rect 32081 4661 32112 4712
rect 32147 4741 32184 4811
rect 32450 4810 32487 4811
rect 32299 4751 32335 4752
rect 32147 4721 32156 4741
rect 32176 4721 32184 4741
rect 32147 4711 32184 4721
rect 32243 4741 32391 4751
rect 32491 4748 32587 4750
rect 32243 4721 32252 4741
rect 32272 4721 32362 4741
rect 32382 4721 32391 4741
rect 32243 4712 32391 4721
rect 32449 4741 32587 4748
rect 32449 4721 32458 4741
rect 32478 4721 32587 4741
rect 32449 4712 32587 4721
rect 32243 4711 32280 4712
rect 31973 4658 32014 4659
rect 30643 4640 31082 4658
rect 29816 4545 29856 4554
rect 30118 4545 30145 4632
rect 30218 4606 30261 4632
rect 30218 4588 30231 4606
rect 30249 4588 30261 4606
rect 30218 4577 30261 4588
rect 29090 4539 29125 4540
rect 28968 4529 29125 4539
rect 28968 4509 28985 4529
rect 29005 4509 29125 4529
rect 28968 4502 29125 4509
rect 29192 4532 29338 4540
rect 29192 4512 29203 4532
rect 29223 4512 29262 4532
rect 29282 4512 29338 4532
rect 29816 4528 30145 4545
rect 29816 4527 29856 4528
rect 29192 4505 29338 4512
rect 30213 4516 30253 4519
rect 30213 4510 30256 4516
rect 29838 4507 30256 4510
rect 29192 4504 29233 4505
rect 28926 4451 28963 4452
rect 28619 4442 28757 4451
rect 28619 4422 28728 4442
rect 28748 4422 28757 4442
rect 28619 4415 28757 4422
rect 28815 4442 28963 4451
rect 28815 4422 28824 4442
rect 28844 4422 28934 4442
rect 28954 4422 28963 4442
rect 28619 4413 28715 4415
rect 28815 4412 28963 4422
rect 29022 4442 29059 4452
rect 29022 4422 29030 4442
rect 29050 4422 29059 4442
rect 28871 4411 28907 4412
rect 28719 4352 28756 4353
rect 29022 4352 29059 4422
rect 29094 4451 29125 4502
rect 29838 4489 30229 4507
rect 30247 4489 30256 4507
rect 29838 4487 30256 4489
rect 29838 4479 29865 4487
rect 30106 4484 30256 4487
rect 29418 4473 29586 4474
rect 29837 4473 29865 4479
rect 29418 4457 29865 4473
rect 30213 4479 30256 4484
rect 29144 4451 29181 4452
rect 29094 4442 29181 4451
rect 29094 4422 29152 4442
rect 29172 4422 29181 4442
rect 29094 4412 29181 4422
rect 29240 4442 29277 4452
rect 29240 4422 29248 4442
rect 29268 4422 29277 4442
rect 29094 4411 29125 4412
rect 28718 4351 29059 4352
rect 29240 4351 29277 4422
rect 28643 4346 29059 4351
rect 28643 4326 28646 4346
rect 28666 4326 29059 4346
rect 29090 4327 29277 4351
rect 29418 4447 29862 4457
rect 29418 4445 29586 4447
rect 28452 4252 28496 4253
rect 28452 4246 28497 4252
rect 28452 4228 28464 4246
rect 28486 4228 28497 4246
rect 28518 4247 28560 4292
rect 29418 4267 29445 4445
rect 29485 4407 29549 4419
rect 29825 4415 29862 4447
rect 29888 4446 30079 4468
rect 30043 4444 30079 4446
rect 30043 4415 30080 4444
rect 30213 4423 30253 4479
rect 29485 4406 29520 4407
rect 29462 4401 29520 4406
rect 29462 4381 29465 4401
rect 29485 4387 29520 4401
rect 29540 4387 29549 4407
rect 29485 4379 29549 4387
rect 29511 4378 29549 4379
rect 29512 4377 29549 4378
rect 29615 4411 29651 4412
rect 29723 4411 29759 4412
rect 29615 4403 29759 4411
rect 29615 4383 29623 4403
rect 29643 4383 29678 4403
rect 29698 4383 29731 4403
rect 29751 4383 29759 4403
rect 29615 4377 29759 4383
rect 29825 4407 29863 4415
rect 29941 4411 29977 4412
rect 29825 4387 29834 4407
rect 29854 4387 29863 4407
rect 29825 4378 29863 4387
rect 29892 4403 29977 4411
rect 29892 4383 29949 4403
rect 29969 4383 29977 4403
rect 29825 4377 29862 4378
rect 29892 4377 29977 4383
rect 30043 4407 30081 4415
rect 30043 4387 30052 4407
rect 30072 4387 30081 4407
rect 30213 4405 30225 4423
rect 30243 4405 30253 4423
rect 30645 4451 30697 4640
rect 31043 4615 31082 4640
rect 31865 4651 32014 4658
rect 31865 4631 31924 4651
rect 31944 4631 31983 4651
rect 32003 4631 32014 4651
rect 31865 4623 32014 4631
rect 32081 4654 32238 4661
rect 32081 4634 32201 4654
rect 32221 4634 32238 4654
rect 32081 4624 32238 4634
rect 32081 4623 32116 4624
rect 30827 4590 31014 4614
rect 31043 4595 31438 4615
rect 31458 4595 31461 4615
rect 32081 4602 32112 4623
rect 32299 4602 32335 4712
rect 32354 4711 32391 4712
rect 32450 4711 32487 4712
rect 32410 4652 32500 4658
rect 32410 4632 32419 4652
rect 32439 4650 32500 4652
rect 32439 4632 32464 4650
rect 32410 4630 32464 4632
rect 32484 4630 32500 4650
rect 32410 4624 32500 4630
rect 31924 4601 31961 4602
rect 31043 4590 31461 4595
rect 31923 4592 31961 4601
rect 30827 4519 30864 4590
rect 31043 4589 31386 4590
rect 31043 4586 31082 4589
rect 31348 4588 31385 4589
rect 30979 4529 31010 4530
rect 30827 4499 30836 4519
rect 30856 4499 30864 4519
rect 30827 4489 30864 4499
rect 30923 4519 31010 4529
rect 30923 4499 30932 4519
rect 30952 4499 31010 4519
rect 30923 4490 31010 4499
rect 30923 4489 30960 4490
rect 30645 4433 30661 4451
rect 30679 4433 30697 4451
rect 30979 4439 31010 4490
rect 31045 4519 31082 4586
rect 31923 4572 31932 4592
rect 31952 4572 31961 4592
rect 31923 4564 31961 4572
rect 32027 4596 32112 4602
rect 32142 4601 32179 4602
rect 32027 4576 32035 4596
rect 32055 4576 32112 4596
rect 32027 4568 32112 4576
rect 32141 4592 32179 4601
rect 32141 4572 32150 4592
rect 32170 4572 32179 4592
rect 32027 4567 32063 4568
rect 32141 4564 32179 4572
rect 32245 4596 32389 4602
rect 32245 4576 32253 4596
rect 32273 4590 32361 4596
rect 32273 4576 32302 4590
rect 32245 4568 32302 4576
rect 32245 4567 32281 4568
rect 32325 4576 32361 4590
rect 32381 4576 32389 4596
rect 32325 4568 32389 4576
rect 32353 4567 32389 4568
rect 32455 4601 32492 4602
rect 32455 4600 32493 4601
rect 32455 4592 32519 4600
rect 32455 4572 32464 4592
rect 32484 4578 32519 4592
rect 32539 4578 32542 4598
rect 32484 4573 32542 4578
rect 32484 4572 32519 4573
rect 31924 4535 31961 4564
rect 31925 4533 31961 4535
rect 31197 4529 31233 4530
rect 31045 4499 31054 4519
rect 31074 4499 31082 4519
rect 31045 4489 31082 4499
rect 31141 4519 31289 4529
rect 31389 4526 31485 4528
rect 31141 4499 31150 4519
rect 31170 4499 31260 4519
rect 31280 4499 31289 4519
rect 31141 4490 31289 4499
rect 31347 4519 31485 4526
rect 31347 4499 31356 4519
rect 31376 4499 31485 4519
rect 31925 4511 32116 4533
rect 32142 4532 32179 4564
rect 32455 4560 32519 4572
rect 32559 4534 32586 4712
rect 32883 4665 32920 4671
rect 32883 4646 32891 4665
rect 32912 4646 32920 4665
rect 32883 4638 32920 4646
rect 32418 4532 32586 4534
rect 32142 4506 32586 4532
rect 32252 4504 32292 4506
rect 32418 4505 32586 4506
rect 31347 4490 31485 4499
rect 32545 4500 32586 4505
rect 31141 4489 31178 4490
rect 30871 4436 30912 4437
rect 30645 4415 30697 4433
rect 30763 4429 30912 4436
rect 30213 4395 30253 4405
rect 30763 4409 30822 4429
rect 30842 4409 30881 4429
rect 30901 4409 30912 4429
rect 30763 4401 30912 4409
rect 30979 4432 31136 4439
rect 30979 4412 31099 4432
rect 31119 4412 31136 4432
rect 30979 4402 31136 4412
rect 30979 4401 31014 4402
rect 30043 4378 30081 4387
rect 30979 4380 31010 4401
rect 31197 4380 31233 4490
rect 31252 4489 31289 4490
rect 31348 4489 31385 4490
rect 31308 4430 31398 4436
rect 31308 4410 31317 4430
rect 31337 4428 31398 4430
rect 31337 4410 31362 4428
rect 31308 4408 31362 4410
rect 31382 4408 31398 4428
rect 31308 4402 31398 4408
rect 30822 4379 30859 4380
rect 30043 4377 30080 4378
rect 29504 4349 29594 4355
rect 29504 4329 29520 4349
rect 29540 4347 29594 4349
rect 29540 4329 29565 4347
rect 29504 4327 29565 4329
rect 29585 4327 29594 4347
rect 29504 4321 29594 4327
rect 29517 4267 29554 4268
rect 29613 4267 29650 4268
rect 29669 4267 29705 4377
rect 29892 4356 29923 4377
rect 30821 4370 30859 4379
rect 29888 4355 29923 4356
rect 29766 4345 29923 4355
rect 29766 4325 29783 4345
rect 29803 4325 29923 4345
rect 29766 4318 29923 4325
rect 29990 4348 30139 4356
rect 29990 4328 30001 4348
rect 30021 4328 30060 4348
rect 30080 4328 30139 4348
rect 30649 4352 30689 4362
rect 29990 4321 30139 4328
rect 30205 4324 30257 4342
rect 29990 4320 30031 4321
rect 29724 4267 29761 4268
rect 29417 4258 29555 4267
rect 28889 4247 28922 4249
rect 28518 4235 28965 4247
rect 28452 4198 28497 4228
rect 28469 3252 28497 4198
rect 28521 4221 28965 4235
rect 28521 4219 28689 4221
rect 28521 4041 28548 4219
rect 28588 4181 28652 4193
rect 28928 4189 28965 4221
rect 28991 4220 29182 4242
rect 29417 4238 29526 4258
rect 29546 4238 29555 4258
rect 29417 4231 29555 4238
rect 29613 4258 29761 4267
rect 29613 4238 29622 4258
rect 29642 4238 29732 4258
rect 29752 4238 29761 4258
rect 29417 4229 29513 4231
rect 29613 4228 29761 4238
rect 29820 4258 29857 4268
rect 29820 4238 29828 4258
rect 29848 4238 29857 4258
rect 29669 4227 29705 4228
rect 29146 4218 29182 4220
rect 29146 4189 29183 4218
rect 28588 4180 28623 4181
rect 28565 4175 28623 4180
rect 28565 4155 28568 4175
rect 28588 4161 28623 4175
rect 28643 4161 28652 4181
rect 28588 4153 28652 4161
rect 28614 4152 28652 4153
rect 28615 4151 28652 4152
rect 28718 4185 28754 4186
rect 28826 4185 28862 4186
rect 28718 4179 28862 4185
rect 28718 4177 28779 4179
rect 28718 4157 28726 4177
rect 28746 4162 28779 4177
rect 28798 4177 28862 4179
rect 28798 4162 28834 4177
rect 28746 4157 28834 4162
rect 28854 4157 28862 4177
rect 28718 4151 28862 4157
rect 28928 4181 28966 4189
rect 29044 4185 29080 4186
rect 28928 4161 28937 4181
rect 28957 4161 28966 4181
rect 28928 4152 28966 4161
rect 28995 4177 29080 4185
rect 28995 4157 29052 4177
rect 29072 4157 29080 4177
rect 28928 4151 28965 4152
rect 28995 4151 29080 4157
rect 29146 4181 29184 4189
rect 29146 4161 29155 4181
rect 29175 4161 29184 4181
rect 29820 4171 29857 4238
rect 29892 4267 29923 4318
rect 30205 4306 30223 4324
rect 30241 4306 30257 4324
rect 29942 4267 29979 4268
rect 29892 4258 29979 4267
rect 29892 4238 29950 4258
rect 29970 4238 29979 4258
rect 29892 4228 29979 4238
rect 30038 4258 30075 4268
rect 30038 4238 30046 4258
rect 30066 4238 30075 4258
rect 29892 4227 29923 4228
rect 29517 4168 29554 4169
rect 29820 4168 29859 4171
rect 29516 4167 29859 4168
rect 30038 4167 30075 4238
rect 29146 4152 29184 4161
rect 29441 4162 29859 4167
rect 29146 4151 29183 4152
rect 28607 4123 28697 4129
rect 28607 4103 28623 4123
rect 28643 4121 28697 4123
rect 28643 4103 28668 4121
rect 28607 4101 28668 4103
rect 28688 4101 28697 4121
rect 28607 4095 28697 4101
rect 28620 4041 28657 4042
rect 28716 4041 28753 4042
rect 28772 4041 28808 4151
rect 28995 4130 29026 4151
rect 29441 4142 29444 4162
rect 29464 4142 29859 4162
rect 29888 4143 30075 4167
rect 28991 4129 29026 4130
rect 28869 4119 29026 4129
rect 28869 4099 28886 4119
rect 28906 4099 29026 4119
rect 28869 4092 29026 4099
rect 29093 4122 29242 4130
rect 29093 4102 29104 4122
rect 29124 4102 29163 4122
rect 29183 4102 29242 4122
rect 29093 4095 29242 4102
rect 29820 4117 29859 4142
rect 30205 4117 30257 4306
rect 30649 4334 30659 4352
rect 30677 4334 30689 4352
rect 30821 4350 30830 4370
rect 30850 4350 30859 4370
rect 30821 4342 30859 4350
rect 30925 4374 31010 4380
rect 31040 4379 31077 4380
rect 30925 4354 30933 4374
rect 30953 4354 31010 4374
rect 30925 4346 31010 4354
rect 31039 4370 31077 4379
rect 31039 4350 31048 4370
rect 31068 4350 31077 4370
rect 30925 4345 30961 4346
rect 31039 4342 31077 4350
rect 31143 4374 31287 4380
rect 31143 4354 31151 4374
rect 31171 4354 31204 4374
rect 31224 4354 31259 4374
rect 31279 4354 31287 4374
rect 31143 4346 31287 4354
rect 31143 4345 31179 4346
rect 31251 4345 31287 4346
rect 31353 4379 31390 4380
rect 31353 4378 31391 4379
rect 31353 4370 31417 4378
rect 31353 4350 31362 4370
rect 31382 4356 31417 4370
rect 31437 4356 31440 4376
rect 31382 4351 31440 4356
rect 31382 4350 31417 4351
rect 30649 4278 30689 4334
rect 30822 4313 30859 4342
rect 30823 4311 30859 4313
rect 30823 4289 31014 4311
rect 31040 4310 31077 4342
rect 31353 4338 31417 4350
rect 31457 4312 31484 4490
rect 31316 4310 31484 4312
rect 31040 4300 31484 4310
rect 31625 4406 31812 4430
rect 31843 4411 32236 4431
rect 32256 4411 32259 4431
rect 31843 4406 32259 4411
rect 31625 4335 31662 4406
rect 31843 4405 32184 4406
rect 31777 4345 31808 4346
rect 31625 4315 31634 4335
rect 31654 4315 31662 4335
rect 31625 4305 31662 4315
rect 31721 4335 31808 4345
rect 31721 4315 31730 4335
rect 31750 4315 31808 4335
rect 31721 4306 31808 4315
rect 31721 4305 31758 4306
rect 30646 4273 30689 4278
rect 31037 4284 31484 4300
rect 31037 4278 31065 4284
rect 31316 4283 31484 4284
rect 30646 4270 30796 4273
rect 31037 4270 31064 4278
rect 30646 4268 31064 4270
rect 30646 4250 30655 4268
rect 30673 4250 31064 4268
rect 31777 4255 31808 4306
rect 31843 4335 31880 4405
rect 32146 4404 32183 4405
rect 31995 4345 32031 4346
rect 31843 4315 31852 4335
rect 31872 4315 31880 4335
rect 31843 4305 31880 4315
rect 31939 4335 32087 4345
rect 32187 4342 32283 4344
rect 31939 4315 31948 4335
rect 31968 4315 32058 4335
rect 32078 4315 32087 4335
rect 31939 4306 32087 4315
rect 32145 4335 32283 4342
rect 32145 4315 32154 4335
rect 32174 4315 32283 4335
rect 32545 4318 32585 4500
rect 32145 4306 32283 4315
rect 31939 4305 31976 4306
rect 31669 4252 31710 4253
rect 30646 4247 31064 4250
rect 30646 4241 30689 4247
rect 30649 4238 30689 4241
rect 31561 4245 31710 4252
rect 31046 4229 31086 4230
rect 30757 4212 31086 4229
rect 31561 4225 31620 4245
rect 31640 4225 31679 4245
rect 31699 4225 31710 4245
rect 31561 4217 31710 4225
rect 31777 4248 31934 4255
rect 31777 4228 31897 4248
rect 31917 4228 31934 4248
rect 31777 4218 31934 4228
rect 31777 4217 31812 4218
rect 30641 4169 30684 4180
rect 30641 4151 30653 4169
rect 30671 4151 30684 4169
rect 30641 4125 30684 4151
rect 30757 4125 30784 4212
rect 31046 4203 31086 4212
rect 29820 4099 30259 4117
rect 29093 4094 29134 4095
rect 28827 4041 28864 4042
rect 28520 4032 28658 4041
rect 28520 4012 28629 4032
rect 28649 4012 28658 4032
rect 28520 4005 28658 4012
rect 28716 4032 28864 4041
rect 28716 4012 28725 4032
rect 28745 4012 28835 4032
rect 28855 4012 28864 4032
rect 28520 4003 28616 4005
rect 28716 4002 28864 4012
rect 28923 4032 28960 4042
rect 28923 4012 28931 4032
rect 28951 4012 28960 4032
rect 28772 4001 28808 4002
rect 28620 3942 28657 3943
rect 28923 3942 28960 4012
rect 28995 4041 29026 4092
rect 29820 4081 30220 4099
rect 30238 4081 30259 4099
rect 29820 4075 30259 4081
rect 29826 4071 30259 4075
rect 30641 4104 30784 4125
rect 30828 4177 30862 4193
rect 31046 4183 31439 4203
rect 31459 4183 31462 4203
rect 31777 4196 31808 4217
rect 31995 4196 32031 4306
rect 32050 4305 32087 4306
rect 32146 4305 32183 4306
rect 32106 4246 32196 4252
rect 32106 4226 32115 4246
rect 32135 4244 32196 4246
rect 32135 4226 32160 4244
rect 32106 4224 32160 4226
rect 32180 4224 32196 4244
rect 32106 4218 32196 4224
rect 31620 4195 31657 4196
rect 31046 4178 31462 4183
rect 31619 4186 31657 4195
rect 31046 4177 31387 4178
rect 30828 4107 30865 4177
rect 30980 4117 31011 4118
rect 30641 4102 30778 4104
rect 30205 4069 30257 4071
rect 30641 4060 30684 4102
rect 30828 4087 30837 4107
rect 30857 4087 30865 4107
rect 30828 4077 30865 4087
rect 30924 4107 31011 4117
rect 30924 4087 30933 4107
rect 30953 4087 31011 4107
rect 30924 4078 31011 4087
rect 30924 4077 30961 4078
rect 30639 4050 30684 4060
rect 29045 4041 29082 4042
rect 28995 4032 29082 4041
rect 28995 4012 29053 4032
rect 29073 4012 29082 4032
rect 28995 4002 29082 4012
rect 29141 4032 29178 4042
rect 29141 4012 29149 4032
rect 29169 4012 29178 4032
rect 30639 4032 30648 4050
rect 30666 4032 30684 4050
rect 30639 4026 30684 4032
rect 30980 4027 31011 4078
rect 31046 4107 31083 4177
rect 31349 4176 31386 4177
rect 31619 4166 31628 4186
rect 31648 4166 31657 4186
rect 31619 4158 31657 4166
rect 31723 4190 31808 4196
rect 31838 4195 31875 4196
rect 31723 4170 31731 4190
rect 31751 4170 31808 4190
rect 31723 4162 31808 4170
rect 31837 4186 31875 4195
rect 31837 4166 31846 4186
rect 31866 4166 31875 4186
rect 31723 4161 31759 4162
rect 31837 4158 31875 4166
rect 31941 4190 32085 4196
rect 31941 4170 31949 4190
rect 31969 4171 32001 4190
rect 32022 4171 32057 4190
rect 31969 4170 32057 4171
rect 32077 4170 32085 4190
rect 31941 4162 32085 4170
rect 31941 4161 31977 4162
rect 32049 4161 32085 4162
rect 32151 4195 32188 4196
rect 32151 4194 32189 4195
rect 32151 4186 32215 4194
rect 32151 4166 32160 4186
rect 32180 4172 32215 4186
rect 32235 4172 32238 4192
rect 32180 4167 32238 4172
rect 32180 4166 32215 4167
rect 31620 4129 31657 4158
rect 31621 4127 31657 4129
rect 31198 4117 31234 4118
rect 31046 4087 31055 4107
rect 31075 4087 31083 4107
rect 31046 4077 31083 4087
rect 31142 4107 31290 4117
rect 31390 4114 31486 4116
rect 31142 4087 31151 4107
rect 31171 4087 31261 4107
rect 31281 4087 31290 4107
rect 31142 4078 31290 4087
rect 31348 4107 31486 4114
rect 31348 4087 31357 4107
rect 31377 4087 31486 4107
rect 31621 4105 31812 4127
rect 31838 4126 31875 4158
rect 32151 4154 32215 4166
rect 32255 4128 32282 4306
rect 32114 4126 32282 4128
rect 31838 4100 32282 4126
rect 31348 4078 31486 4087
rect 31142 4077 31179 4078
rect 30639 4023 30676 4026
rect 30872 4024 30913 4025
rect 28995 4001 29026 4002
rect 28619 3941 28960 3942
rect 29141 3941 29178 4012
rect 30764 4017 30913 4024
rect 30208 4004 30245 4009
rect 30199 4000 30246 4004
rect 30199 3982 30218 4000
rect 30236 3982 30246 4000
rect 30764 3997 30823 4017
rect 30843 3997 30882 4017
rect 30902 3997 30913 4017
rect 30764 3989 30913 3997
rect 30980 4020 31137 4027
rect 30980 4000 31100 4020
rect 31120 4000 31137 4020
rect 30980 3990 31137 4000
rect 30980 3989 31015 3990
rect 28544 3936 28960 3941
rect 28544 3916 28547 3936
rect 28567 3916 28960 3936
rect 28991 3917 29178 3941
rect 29803 3939 29843 3944
rect 30199 3939 30246 3982
rect 30980 3968 31011 3989
rect 31198 3968 31234 4078
rect 31253 4077 31290 4078
rect 31349 4077 31386 4078
rect 31309 4018 31399 4024
rect 31309 3998 31318 4018
rect 31338 4016 31399 4018
rect 31338 3998 31363 4016
rect 31309 3996 31363 3998
rect 31383 3996 31399 4016
rect 31309 3990 31399 3996
rect 30823 3967 30860 3968
rect 29803 3900 30246 3939
rect 30636 3959 30673 3961
rect 30636 3951 30678 3959
rect 30636 3933 30646 3951
rect 30664 3933 30678 3951
rect 30636 3924 30678 3933
rect 30822 3958 30860 3967
rect 30822 3938 30831 3958
rect 30851 3938 30860 3958
rect 30822 3930 30860 3938
rect 30926 3962 31011 3968
rect 31041 3967 31078 3968
rect 30926 3942 30934 3962
rect 30954 3942 31011 3962
rect 30926 3934 31011 3942
rect 31040 3958 31078 3967
rect 31040 3938 31049 3958
rect 31069 3938 31078 3958
rect 30926 3933 30962 3934
rect 31040 3930 31078 3938
rect 31144 3966 31288 3968
rect 31144 3962 31196 3966
rect 31144 3942 31152 3962
rect 31172 3946 31196 3962
rect 31216 3962 31288 3966
rect 31216 3946 31260 3962
rect 31172 3942 31260 3946
rect 31280 3942 31288 3962
rect 31144 3934 31288 3942
rect 31144 3933 31180 3934
rect 31252 3933 31288 3934
rect 31354 3967 31391 3968
rect 31354 3966 31392 3967
rect 31354 3958 31418 3966
rect 31354 3938 31363 3958
rect 31383 3944 31418 3958
rect 31438 3944 31441 3964
rect 31383 3939 31441 3944
rect 31383 3938 31418 3939
rect 28897 3885 28937 3893
rect 28897 3863 28905 3885
rect 28929 3863 28937 3885
rect 28603 3639 28771 3640
rect 28897 3639 28937 3863
rect 29400 3867 29568 3868
rect 29803 3867 29843 3900
rect 30199 3867 30246 3900
rect 30637 3899 30678 3924
rect 30823 3899 30860 3930
rect 31041 3899 31078 3930
rect 31354 3926 31418 3938
rect 31458 3900 31485 4078
rect 30637 3872 30686 3899
rect 30822 3873 30871 3899
rect 31040 3898 31121 3899
rect 31317 3898 31485 3900
rect 31040 3873 31485 3898
rect 31041 3872 31485 3873
rect 29400 3866 29844 3867
rect 29400 3841 29845 3866
rect 29400 3839 29568 3841
rect 29764 3840 29845 3841
rect 30014 3840 30063 3866
rect 30199 3840 30248 3867
rect 29400 3661 29427 3839
rect 29467 3801 29531 3813
rect 29807 3809 29844 3840
rect 30025 3809 30062 3840
rect 30207 3815 30248 3840
rect 30639 3839 30686 3872
rect 31042 3839 31082 3872
rect 31317 3871 31485 3872
rect 31948 3876 31988 4100
rect 32114 4099 32282 4100
rect 31948 3854 31956 3876
rect 31980 3854 31988 3876
rect 31948 3846 31988 3854
rect 29467 3800 29502 3801
rect 29444 3795 29502 3800
rect 29444 3775 29447 3795
rect 29467 3781 29502 3795
rect 29522 3781 29531 3801
rect 29467 3773 29531 3781
rect 29493 3772 29531 3773
rect 29494 3771 29531 3772
rect 29597 3805 29633 3806
rect 29705 3805 29741 3806
rect 29597 3797 29741 3805
rect 29597 3777 29605 3797
rect 29625 3793 29713 3797
rect 29625 3777 29669 3793
rect 29597 3773 29669 3777
rect 29689 3777 29713 3793
rect 29733 3777 29741 3797
rect 29689 3773 29741 3777
rect 29597 3771 29741 3773
rect 29807 3801 29845 3809
rect 29923 3805 29959 3806
rect 29807 3781 29816 3801
rect 29836 3781 29845 3801
rect 29807 3772 29845 3781
rect 29874 3797 29959 3805
rect 29874 3777 29931 3797
rect 29951 3777 29959 3797
rect 29807 3771 29844 3772
rect 29874 3771 29959 3777
rect 30025 3801 30063 3809
rect 30025 3781 30034 3801
rect 30054 3781 30063 3801
rect 30025 3772 30063 3781
rect 30207 3806 30249 3815
rect 30207 3788 30221 3806
rect 30239 3788 30249 3806
rect 30207 3780 30249 3788
rect 30212 3778 30249 3780
rect 30639 3800 31082 3839
rect 30025 3771 30062 3772
rect 29486 3743 29576 3749
rect 29486 3723 29502 3743
rect 29522 3741 29576 3743
rect 29522 3723 29547 3741
rect 29486 3721 29547 3723
rect 29567 3721 29576 3741
rect 29486 3715 29576 3721
rect 29499 3661 29536 3662
rect 29595 3661 29632 3662
rect 29651 3661 29687 3771
rect 29874 3750 29905 3771
rect 30639 3757 30686 3800
rect 31042 3795 31082 3800
rect 31707 3798 31894 3822
rect 31925 3803 32318 3823
rect 32338 3803 32341 3823
rect 31925 3798 32341 3803
rect 29870 3749 29905 3750
rect 29748 3739 29905 3749
rect 29748 3719 29765 3739
rect 29785 3719 29905 3739
rect 29748 3712 29905 3719
rect 29972 3742 30121 3750
rect 29972 3722 29983 3742
rect 30003 3722 30042 3742
rect 30062 3722 30121 3742
rect 30639 3739 30649 3757
rect 30667 3739 30686 3757
rect 30639 3735 30686 3739
rect 30640 3730 30677 3735
rect 29972 3715 30121 3722
rect 31707 3727 31744 3798
rect 31925 3797 32266 3798
rect 31859 3737 31890 3738
rect 29972 3714 30013 3715
rect 30209 3713 30246 3716
rect 29706 3661 29743 3662
rect 29399 3652 29537 3661
rect 28603 3613 29047 3639
rect 28603 3611 28771 3613
rect 28603 3433 28630 3611
rect 28670 3573 28734 3585
rect 29010 3581 29047 3613
rect 29073 3612 29264 3634
rect 29399 3632 29508 3652
rect 29528 3632 29537 3652
rect 29399 3625 29537 3632
rect 29595 3652 29743 3661
rect 29595 3632 29604 3652
rect 29624 3632 29714 3652
rect 29734 3632 29743 3652
rect 29399 3623 29495 3625
rect 29595 3622 29743 3632
rect 29802 3652 29839 3662
rect 29802 3632 29810 3652
rect 29830 3632 29839 3652
rect 29651 3621 29687 3622
rect 29228 3610 29264 3612
rect 29228 3581 29265 3610
rect 28670 3572 28705 3573
rect 28647 3567 28705 3572
rect 28647 3547 28650 3567
rect 28670 3553 28705 3567
rect 28725 3553 28734 3573
rect 28670 3545 28734 3553
rect 28696 3544 28734 3545
rect 28697 3543 28734 3544
rect 28800 3577 28836 3578
rect 28908 3577 28944 3578
rect 28800 3569 28944 3577
rect 28800 3549 28808 3569
rect 28828 3568 28916 3569
rect 28828 3549 28863 3568
rect 28884 3549 28916 3568
rect 28936 3549 28944 3569
rect 28800 3543 28944 3549
rect 29010 3573 29048 3581
rect 29126 3577 29162 3578
rect 29010 3553 29019 3573
rect 29039 3553 29048 3573
rect 29010 3544 29048 3553
rect 29077 3569 29162 3577
rect 29077 3549 29134 3569
rect 29154 3549 29162 3569
rect 29010 3543 29047 3544
rect 29077 3543 29162 3549
rect 29228 3573 29266 3581
rect 29228 3553 29237 3573
rect 29257 3553 29266 3573
rect 29499 3562 29536 3563
rect 29802 3562 29839 3632
rect 29874 3661 29905 3712
rect 30201 3707 30246 3713
rect 30201 3689 30219 3707
rect 30237 3689 30246 3707
rect 31707 3707 31716 3727
rect 31736 3707 31744 3727
rect 31707 3697 31744 3707
rect 31803 3727 31890 3737
rect 31803 3707 31812 3727
rect 31832 3707 31890 3727
rect 31803 3698 31890 3707
rect 31803 3697 31840 3698
rect 30201 3679 30246 3689
rect 29924 3661 29961 3662
rect 29874 3652 29961 3661
rect 29874 3632 29932 3652
rect 29952 3632 29961 3652
rect 29874 3622 29961 3632
rect 30020 3652 30057 3662
rect 30020 3632 30028 3652
rect 30048 3632 30057 3652
rect 30201 3637 30244 3679
rect 30628 3668 30680 3670
rect 30107 3635 30244 3637
rect 29874 3621 29905 3622
rect 30020 3562 30057 3632
rect 29498 3561 29839 3562
rect 29228 3544 29266 3553
rect 29423 3556 29839 3561
rect 29228 3543 29265 3544
rect 28689 3515 28779 3521
rect 28689 3495 28705 3515
rect 28725 3513 28779 3515
rect 28725 3495 28750 3513
rect 28689 3493 28750 3495
rect 28770 3493 28779 3513
rect 28689 3487 28779 3493
rect 28702 3433 28739 3434
rect 28798 3433 28835 3434
rect 28854 3433 28890 3543
rect 29077 3522 29108 3543
rect 29423 3536 29426 3556
rect 29446 3536 29839 3556
rect 30023 3546 30057 3562
rect 30101 3614 30244 3635
rect 30626 3664 31059 3668
rect 30626 3658 31065 3664
rect 30626 3640 30647 3658
rect 30665 3640 31065 3658
rect 31859 3647 31890 3698
rect 31925 3727 31962 3797
rect 32228 3796 32265 3797
rect 32077 3737 32113 3738
rect 31925 3707 31934 3727
rect 31954 3707 31962 3727
rect 31925 3697 31962 3707
rect 32021 3727 32169 3737
rect 32269 3734 32365 3736
rect 32021 3707 32030 3727
rect 32050 3707 32140 3727
rect 32160 3707 32169 3727
rect 32021 3698 32169 3707
rect 32227 3727 32365 3734
rect 32227 3707 32236 3727
rect 32256 3707 32365 3727
rect 32227 3698 32365 3707
rect 32021 3697 32058 3698
rect 31751 3644 31792 3645
rect 30626 3622 31065 3640
rect 29799 3527 29839 3536
rect 30101 3527 30128 3614
rect 30201 3588 30244 3614
rect 30201 3570 30214 3588
rect 30232 3570 30244 3588
rect 30201 3559 30244 3570
rect 29073 3521 29108 3522
rect 28951 3511 29108 3521
rect 28951 3491 28968 3511
rect 28988 3491 29108 3511
rect 28951 3484 29108 3491
rect 29175 3514 29324 3522
rect 29175 3494 29186 3514
rect 29206 3494 29245 3514
rect 29265 3494 29324 3514
rect 29799 3510 30128 3527
rect 29799 3509 29839 3510
rect 29175 3487 29324 3494
rect 30196 3498 30236 3501
rect 30196 3492 30239 3498
rect 29821 3489 30239 3492
rect 29175 3486 29216 3487
rect 28909 3433 28946 3434
rect 28602 3424 28740 3433
rect 28602 3404 28711 3424
rect 28731 3404 28740 3424
rect 28602 3397 28740 3404
rect 28798 3424 28946 3433
rect 28798 3404 28807 3424
rect 28827 3404 28917 3424
rect 28937 3404 28946 3424
rect 28602 3395 28698 3397
rect 28798 3394 28946 3404
rect 29005 3424 29042 3434
rect 29005 3404 29013 3424
rect 29033 3404 29042 3424
rect 28854 3393 28890 3394
rect 28702 3334 28739 3335
rect 29005 3334 29042 3404
rect 29077 3433 29108 3484
rect 29821 3471 30212 3489
rect 30230 3471 30239 3489
rect 29821 3469 30239 3471
rect 29821 3461 29848 3469
rect 30089 3466 30239 3469
rect 29401 3455 29569 3456
rect 29820 3455 29848 3461
rect 29401 3439 29848 3455
rect 30196 3461 30239 3466
rect 29127 3433 29164 3434
rect 29077 3424 29164 3433
rect 29077 3404 29135 3424
rect 29155 3404 29164 3424
rect 29077 3394 29164 3404
rect 29223 3424 29260 3434
rect 29223 3404 29231 3424
rect 29251 3404 29260 3424
rect 29077 3393 29108 3394
rect 28701 3333 29042 3334
rect 29223 3333 29260 3404
rect 28626 3328 29042 3333
rect 28626 3308 28629 3328
rect 28649 3308 29042 3328
rect 29073 3309 29260 3333
rect 29401 3429 29845 3439
rect 29401 3427 29569 3429
rect 28468 3234 28497 3252
rect 29401 3249 29428 3427
rect 29468 3389 29532 3401
rect 29808 3397 29845 3429
rect 29871 3428 30062 3450
rect 30026 3426 30062 3428
rect 30026 3397 30063 3426
rect 30196 3405 30236 3461
rect 29468 3388 29503 3389
rect 29445 3383 29503 3388
rect 29445 3363 29448 3383
rect 29468 3369 29503 3383
rect 29523 3369 29532 3389
rect 29468 3361 29532 3369
rect 29494 3360 29532 3361
rect 29495 3359 29532 3360
rect 29598 3393 29634 3394
rect 29706 3393 29742 3394
rect 29598 3385 29742 3393
rect 29598 3365 29606 3385
rect 29626 3365 29661 3385
rect 29681 3365 29714 3385
rect 29734 3365 29742 3385
rect 29598 3359 29742 3365
rect 29808 3389 29846 3397
rect 29924 3393 29960 3394
rect 29808 3369 29817 3389
rect 29837 3369 29846 3389
rect 29808 3360 29846 3369
rect 29875 3385 29960 3393
rect 29875 3365 29932 3385
rect 29952 3365 29960 3385
rect 29808 3359 29845 3360
rect 29875 3359 29960 3365
rect 30026 3389 30064 3397
rect 30026 3369 30035 3389
rect 30055 3369 30064 3389
rect 30196 3387 30208 3405
rect 30226 3387 30236 3405
rect 30628 3433 30680 3622
rect 31026 3597 31065 3622
rect 31643 3637 31792 3644
rect 31643 3617 31702 3637
rect 31722 3617 31761 3637
rect 31781 3617 31792 3637
rect 31643 3609 31792 3617
rect 31859 3640 32016 3647
rect 31859 3620 31979 3640
rect 31999 3620 32016 3640
rect 31859 3610 32016 3620
rect 31859 3609 31894 3610
rect 30810 3572 30997 3596
rect 31026 3577 31421 3597
rect 31441 3577 31444 3597
rect 31859 3588 31890 3609
rect 32077 3588 32113 3698
rect 32132 3697 32169 3698
rect 32228 3697 32265 3698
rect 32188 3638 32278 3644
rect 32188 3618 32197 3638
rect 32217 3636 32278 3638
rect 32217 3618 32242 3636
rect 32188 3616 32242 3618
rect 32262 3616 32278 3636
rect 32188 3610 32278 3616
rect 31702 3587 31739 3588
rect 31026 3572 31444 3577
rect 31701 3578 31739 3587
rect 30810 3501 30847 3572
rect 31026 3571 31369 3572
rect 31026 3568 31065 3571
rect 31331 3570 31368 3571
rect 30962 3511 30993 3512
rect 30810 3481 30819 3501
rect 30839 3481 30847 3501
rect 30810 3471 30847 3481
rect 30906 3501 30993 3511
rect 30906 3481 30915 3501
rect 30935 3481 30993 3501
rect 30906 3472 30993 3481
rect 30906 3471 30943 3472
rect 30628 3415 30644 3433
rect 30662 3415 30680 3433
rect 30962 3421 30993 3472
rect 31028 3501 31065 3568
rect 31701 3558 31710 3578
rect 31730 3558 31739 3578
rect 31701 3550 31739 3558
rect 31805 3582 31890 3588
rect 31920 3587 31957 3588
rect 31805 3562 31813 3582
rect 31833 3562 31890 3582
rect 31805 3554 31890 3562
rect 31919 3578 31957 3587
rect 31919 3558 31928 3578
rect 31948 3558 31957 3578
rect 31805 3553 31841 3554
rect 31919 3550 31957 3558
rect 32023 3583 32167 3588
rect 32023 3582 32085 3583
rect 32023 3562 32031 3582
rect 32051 3564 32085 3582
rect 32106 3582 32167 3583
rect 32106 3564 32139 3582
rect 32051 3562 32139 3564
rect 32159 3562 32167 3582
rect 32023 3554 32167 3562
rect 32023 3553 32059 3554
rect 32131 3553 32167 3554
rect 32233 3587 32270 3588
rect 32233 3586 32271 3587
rect 32233 3578 32297 3586
rect 32233 3558 32242 3578
rect 32262 3564 32297 3578
rect 32317 3564 32320 3584
rect 32262 3559 32320 3564
rect 32262 3558 32297 3559
rect 31702 3521 31739 3550
rect 31703 3519 31739 3521
rect 31180 3511 31216 3512
rect 31028 3481 31037 3501
rect 31057 3481 31065 3501
rect 31028 3471 31065 3481
rect 31124 3501 31272 3511
rect 31372 3508 31468 3510
rect 31124 3481 31133 3501
rect 31153 3481 31243 3501
rect 31263 3481 31272 3501
rect 31124 3472 31272 3481
rect 31330 3501 31468 3508
rect 31330 3481 31339 3501
rect 31359 3481 31468 3501
rect 31703 3497 31894 3519
rect 31920 3518 31957 3550
rect 32233 3546 32297 3558
rect 32337 3520 32364 3698
rect 32196 3518 32364 3520
rect 31920 3504 32364 3518
rect 31920 3492 32367 3504
rect 31963 3490 31996 3492
rect 31330 3472 31468 3481
rect 31124 3471 31161 3472
rect 30854 3418 30895 3419
rect 30628 3397 30680 3415
rect 30746 3411 30895 3418
rect 30196 3377 30236 3387
rect 30746 3391 30805 3411
rect 30825 3391 30864 3411
rect 30884 3391 30895 3411
rect 30746 3383 30895 3391
rect 30962 3414 31119 3421
rect 30962 3394 31082 3414
rect 31102 3394 31119 3414
rect 30962 3384 31119 3394
rect 30962 3383 30997 3384
rect 30026 3360 30064 3369
rect 30962 3362 30993 3383
rect 31180 3362 31216 3472
rect 31235 3471 31272 3472
rect 31331 3471 31368 3472
rect 31291 3412 31381 3418
rect 31291 3392 31300 3412
rect 31320 3410 31381 3412
rect 31320 3392 31345 3410
rect 31291 3390 31345 3392
rect 31365 3390 31381 3410
rect 31291 3384 31381 3390
rect 30805 3361 30842 3362
rect 30026 3359 30063 3360
rect 29487 3331 29577 3337
rect 29487 3311 29503 3331
rect 29523 3329 29577 3331
rect 29523 3311 29548 3329
rect 29487 3309 29548 3311
rect 29568 3309 29577 3329
rect 29487 3303 29577 3309
rect 29500 3249 29537 3250
rect 29596 3249 29633 3250
rect 29652 3249 29688 3359
rect 29875 3338 29906 3359
rect 30804 3352 30842 3361
rect 29871 3337 29906 3338
rect 29749 3327 29906 3337
rect 29749 3307 29766 3327
rect 29786 3307 29906 3327
rect 29749 3300 29906 3307
rect 29973 3330 30122 3338
rect 29973 3310 29984 3330
rect 30004 3310 30043 3330
rect 30063 3310 30122 3330
rect 30632 3334 30672 3344
rect 29973 3303 30122 3310
rect 30188 3306 30240 3324
rect 29973 3302 30014 3303
rect 29707 3249 29744 3250
rect 28438 3232 28497 3234
rect 29400 3240 29538 3249
rect 28438 3231 28606 3232
rect 28732 3231 28772 3233
rect 28438 3205 28882 3231
rect 28438 3203 28606 3205
rect 28438 3201 28519 3203
rect 28438 3025 28465 3201
rect 28505 3165 28569 3177
rect 28845 3173 28882 3205
rect 28908 3204 29099 3226
rect 29400 3220 29509 3240
rect 29529 3220 29538 3240
rect 29400 3213 29538 3220
rect 29596 3240 29744 3249
rect 29596 3220 29605 3240
rect 29625 3220 29715 3240
rect 29735 3220 29744 3240
rect 29400 3211 29496 3213
rect 29596 3210 29744 3220
rect 29803 3240 29840 3250
rect 29803 3220 29811 3240
rect 29831 3220 29840 3240
rect 29652 3209 29688 3210
rect 29063 3202 29099 3204
rect 29063 3173 29100 3202
rect 28505 3164 28540 3165
rect 28482 3159 28540 3164
rect 28482 3139 28485 3159
rect 28505 3145 28540 3159
rect 28560 3145 28569 3165
rect 28505 3137 28569 3145
rect 28531 3136 28569 3137
rect 28532 3135 28569 3136
rect 28635 3169 28671 3170
rect 28743 3169 28779 3170
rect 28635 3161 28779 3169
rect 28635 3141 28643 3161
rect 28663 3160 28751 3161
rect 28663 3142 28698 3160
rect 28716 3142 28751 3160
rect 28663 3141 28751 3142
rect 28771 3141 28779 3161
rect 28635 3135 28779 3141
rect 28845 3165 28883 3173
rect 28961 3169 28997 3170
rect 28845 3145 28854 3165
rect 28874 3145 28883 3165
rect 28845 3136 28883 3145
rect 28912 3161 28997 3169
rect 28912 3141 28969 3161
rect 28989 3141 28997 3161
rect 28845 3135 28882 3136
rect 28912 3135 28997 3141
rect 29063 3165 29101 3173
rect 29063 3145 29072 3165
rect 29092 3145 29101 3165
rect 29803 3153 29840 3220
rect 29875 3249 29906 3300
rect 30188 3288 30206 3306
rect 30224 3288 30240 3306
rect 29925 3249 29962 3250
rect 29875 3240 29962 3249
rect 29875 3220 29933 3240
rect 29953 3220 29962 3240
rect 29875 3210 29962 3220
rect 30021 3240 30058 3250
rect 30021 3220 30029 3240
rect 30049 3220 30058 3240
rect 29875 3209 29906 3210
rect 29500 3150 29537 3151
rect 29803 3150 29842 3153
rect 29499 3149 29842 3150
rect 30021 3149 30058 3220
rect 29063 3136 29101 3145
rect 29424 3144 29842 3149
rect 29063 3135 29100 3136
rect 28524 3107 28614 3113
rect 28524 3087 28540 3107
rect 28560 3105 28614 3107
rect 28560 3087 28585 3105
rect 28524 3085 28585 3087
rect 28605 3085 28614 3105
rect 28524 3079 28614 3085
rect 28537 3025 28574 3026
rect 28633 3025 28670 3026
rect 28689 3025 28725 3135
rect 28912 3114 28943 3135
rect 29424 3124 29427 3144
rect 29447 3124 29842 3144
rect 29871 3125 30058 3149
rect 28908 3113 28943 3114
rect 28786 3103 28943 3113
rect 28786 3083 28803 3103
rect 28823 3083 28943 3103
rect 28786 3076 28943 3083
rect 29010 3106 29159 3114
rect 29010 3086 29021 3106
rect 29041 3086 29080 3106
rect 29100 3086 29159 3106
rect 29010 3079 29159 3086
rect 29803 3099 29842 3124
rect 30188 3099 30240 3288
rect 30632 3316 30642 3334
rect 30660 3316 30672 3334
rect 30804 3332 30813 3352
rect 30833 3332 30842 3352
rect 30804 3324 30842 3332
rect 30908 3356 30993 3362
rect 31023 3361 31060 3362
rect 30908 3336 30916 3356
rect 30936 3336 30993 3356
rect 30908 3328 30993 3336
rect 31022 3352 31060 3361
rect 31022 3332 31031 3352
rect 31051 3332 31060 3352
rect 30908 3327 30944 3328
rect 31022 3324 31060 3332
rect 31126 3356 31270 3362
rect 31126 3336 31134 3356
rect 31154 3336 31187 3356
rect 31207 3336 31242 3356
rect 31262 3336 31270 3356
rect 31126 3328 31270 3336
rect 31126 3327 31162 3328
rect 31234 3327 31270 3328
rect 31336 3361 31373 3362
rect 31336 3360 31374 3361
rect 31336 3352 31400 3360
rect 31336 3332 31345 3352
rect 31365 3338 31400 3352
rect 31420 3338 31423 3358
rect 31365 3333 31423 3338
rect 31365 3332 31400 3333
rect 30632 3260 30672 3316
rect 30805 3295 30842 3324
rect 30806 3293 30842 3295
rect 30806 3271 30997 3293
rect 31023 3292 31060 3324
rect 31336 3320 31400 3332
rect 31440 3294 31467 3472
rect 32325 3447 32367 3492
rect 31299 3292 31467 3294
rect 31023 3282 31467 3292
rect 31608 3388 31795 3412
rect 31826 3393 32219 3413
rect 32239 3393 32242 3413
rect 31826 3388 32242 3393
rect 31608 3317 31645 3388
rect 31826 3387 32167 3388
rect 31760 3327 31791 3328
rect 31608 3297 31617 3317
rect 31637 3297 31645 3317
rect 31608 3287 31645 3297
rect 31704 3317 31791 3327
rect 31704 3297 31713 3317
rect 31733 3297 31791 3317
rect 31704 3288 31791 3297
rect 31704 3287 31741 3288
rect 30629 3255 30672 3260
rect 31020 3266 31467 3282
rect 31020 3260 31048 3266
rect 31299 3265 31467 3266
rect 30629 3252 30779 3255
rect 31020 3252 31047 3260
rect 30629 3250 31047 3252
rect 30629 3232 30638 3250
rect 30656 3232 31047 3250
rect 31760 3237 31791 3288
rect 31826 3317 31863 3387
rect 32129 3386 32166 3387
rect 31978 3327 32014 3328
rect 31826 3297 31835 3317
rect 31855 3297 31863 3317
rect 31826 3287 31863 3297
rect 31922 3317 32070 3327
rect 32170 3324 32266 3326
rect 31922 3297 31931 3317
rect 31951 3297 32041 3317
rect 32061 3297 32070 3317
rect 31922 3288 32070 3297
rect 32128 3317 32266 3324
rect 32128 3297 32137 3317
rect 32157 3297 32266 3317
rect 32128 3288 32266 3297
rect 31922 3287 31959 3288
rect 31652 3234 31693 3235
rect 30629 3229 31047 3232
rect 30629 3223 30672 3229
rect 30632 3220 30672 3223
rect 31547 3227 31693 3234
rect 31029 3211 31069 3212
rect 30740 3194 31069 3211
rect 31547 3207 31603 3227
rect 31623 3207 31662 3227
rect 31682 3207 31693 3227
rect 31547 3199 31693 3207
rect 31760 3230 31917 3237
rect 31760 3210 31880 3230
rect 31900 3210 31917 3230
rect 31760 3200 31917 3210
rect 31760 3199 31795 3200
rect 30624 3151 30667 3162
rect 30624 3133 30636 3151
rect 30654 3133 30667 3151
rect 30624 3107 30667 3133
rect 30740 3107 30767 3194
rect 31029 3185 31069 3194
rect 29803 3081 30242 3099
rect 29010 3078 29051 3079
rect 28744 3025 28781 3026
rect 28437 3016 28575 3025
rect 28437 2996 28546 3016
rect 28566 2996 28575 3016
rect 28437 2989 28575 2996
rect 28633 3016 28781 3025
rect 28633 2996 28642 3016
rect 28662 2996 28752 3016
rect 28772 2996 28781 3016
rect 28437 2987 28533 2989
rect 28633 2986 28781 2996
rect 28840 3016 28877 3026
rect 28840 2996 28848 3016
rect 28868 2996 28877 3016
rect 28689 2985 28725 2986
rect 28537 2926 28574 2927
rect 28840 2926 28877 2996
rect 28912 3025 28943 3076
rect 29803 3063 30203 3081
rect 30221 3063 30242 3081
rect 29803 3057 30242 3063
rect 29809 3053 30242 3057
rect 30624 3086 30767 3107
rect 30811 3159 30845 3175
rect 31029 3165 31422 3185
rect 31442 3165 31445 3185
rect 31760 3178 31791 3199
rect 31978 3178 32014 3288
rect 32033 3287 32070 3288
rect 32129 3287 32166 3288
rect 32089 3228 32179 3234
rect 32089 3208 32098 3228
rect 32118 3226 32179 3228
rect 32118 3208 32143 3226
rect 32089 3206 32143 3208
rect 32163 3206 32179 3226
rect 32089 3200 32179 3206
rect 31603 3177 31640 3178
rect 31029 3160 31445 3165
rect 31602 3168 31640 3177
rect 31029 3159 31370 3160
rect 30811 3089 30848 3159
rect 30963 3099 30994 3100
rect 30624 3084 30761 3086
rect 30188 3051 30240 3053
rect 30624 3042 30667 3084
rect 30811 3069 30820 3089
rect 30840 3069 30848 3089
rect 30811 3059 30848 3069
rect 30907 3089 30994 3099
rect 30907 3069 30916 3089
rect 30936 3069 30994 3089
rect 30907 3060 30994 3069
rect 30907 3059 30944 3060
rect 30622 3032 30667 3042
rect 28962 3025 28999 3026
rect 28912 3016 28999 3025
rect 28912 2996 28970 3016
rect 28990 2996 28999 3016
rect 28912 2986 28999 2996
rect 29058 3016 29095 3026
rect 29058 2996 29066 3016
rect 29086 2996 29095 3016
rect 30622 3014 30631 3032
rect 30649 3014 30667 3032
rect 30622 3008 30667 3014
rect 30963 3009 30994 3060
rect 31029 3089 31066 3159
rect 31332 3158 31369 3159
rect 31602 3148 31611 3168
rect 31631 3148 31640 3168
rect 31602 3140 31640 3148
rect 31706 3172 31791 3178
rect 31821 3177 31858 3178
rect 31706 3152 31714 3172
rect 31734 3152 31791 3172
rect 31706 3144 31791 3152
rect 31820 3168 31858 3177
rect 31820 3148 31829 3168
rect 31849 3148 31858 3168
rect 31706 3143 31742 3144
rect 31820 3140 31858 3148
rect 31924 3172 32068 3178
rect 31924 3152 31932 3172
rect 31952 3169 32040 3172
rect 31952 3152 31987 3169
rect 31924 3151 31987 3152
rect 32006 3152 32040 3169
rect 32060 3152 32068 3172
rect 32006 3151 32068 3152
rect 31924 3144 32068 3151
rect 31924 3143 31960 3144
rect 32032 3143 32068 3144
rect 32134 3177 32171 3178
rect 32134 3176 32172 3177
rect 32194 3176 32221 3180
rect 32134 3174 32221 3176
rect 32134 3168 32198 3174
rect 32134 3148 32143 3168
rect 32163 3154 32198 3168
rect 32218 3154 32221 3174
rect 32163 3149 32221 3154
rect 32163 3148 32198 3149
rect 31603 3111 31640 3140
rect 31604 3109 31640 3111
rect 31181 3099 31217 3100
rect 31029 3069 31038 3089
rect 31058 3069 31066 3089
rect 31029 3059 31066 3069
rect 31125 3089 31273 3099
rect 31373 3096 31469 3098
rect 31125 3069 31134 3089
rect 31154 3069 31244 3089
rect 31264 3069 31273 3089
rect 31125 3060 31273 3069
rect 31331 3089 31469 3096
rect 31331 3069 31340 3089
rect 31360 3069 31469 3089
rect 31604 3087 31795 3109
rect 31821 3108 31858 3140
rect 32134 3136 32198 3148
rect 32238 3110 32265 3288
rect 32097 3108 32265 3110
rect 31821 3082 32265 3108
rect 31331 3060 31469 3069
rect 31125 3059 31162 3060
rect 30622 3005 30659 3008
rect 30855 3006 30896 3007
rect 28912 2985 28943 2986
rect 28536 2925 28877 2926
rect 29058 2925 29095 2996
rect 30747 2999 30896 3006
rect 30191 2986 30228 2991
rect 28461 2920 28877 2925
rect 28461 2900 28464 2920
rect 28484 2900 28877 2920
rect 28908 2901 29095 2925
rect 30182 2982 30229 2986
rect 30182 2964 30201 2982
rect 30219 2964 30229 2982
rect 30747 2979 30806 2999
rect 30826 2979 30865 2999
rect 30885 2979 30896 2999
rect 30747 2971 30896 2979
rect 30963 3002 31120 3009
rect 30963 2982 31083 3002
rect 31103 2982 31120 3002
rect 30963 2972 31120 2982
rect 30963 2971 30998 2972
rect 30182 2916 30229 2964
rect 30963 2950 30994 2971
rect 31181 2950 31217 3060
rect 31236 3059 31273 3060
rect 31332 3059 31369 3060
rect 31292 3000 31382 3006
rect 31292 2980 31301 3000
rect 31321 2998 31382 3000
rect 31321 2980 31346 2998
rect 31292 2978 31346 2980
rect 31366 2978 31382 2998
rect 31292 2972 31382 2978
rect 30806 2949 30843 2950
rect 29806 2913 30229 2916
rect 28681 2899 28746 2900
rect 29784 2883 30229 2913
rect 30618 2941 30656 2943
rect 30618 2933 30661 2941
rect 30618 2915 30629 2933
rect 30647 2915 30661 2933
rect 30618 2888 30661 2915
rect 30805 2940 30843 2949
rect 30805 2920 30814 2940
rect 30834 2920 30843 2940
rect 30805 2912 30843 2920
rect 30909 2944 30994 2950
rect 31024 2949 31061 2950
rect 30909 2924 30917 2944
rect 30937 2924 30994 2944
rect 30909 2916 30994 2924
rect 31023 2940 31061 2949
rect 31023 2920 31032 2940
rect 31052 2920 31061 2940
rect 30909 2915 30945 2916
rect 31023 2912 31061 2920
rect 31127 2948 31271 2950
rect 31127 2944 31179 2948
rect 31127 2924 31135 2944
rect 31155 2928 31179 2944
rect 31199 2944 31271 2948
rect 31199 2928 31243 2944
rect 31155 2924 31243 2928
rect 31263 2924 31271 2944
rect 31127 2916 31271 2924
rect 31127 2915 31163 2916
rect 31235 2915 31271 2916
rect 31337 2949 31374 2950
rect 31337 2948 31375 2949
rect 31337 2940 31401 2948
rect 31337 2920 31346 2940
rect 31366 2926 31401 2940
rect 31421 2926 31424 2946
rect 31366 2921 31424 2926
rect 31366 2920 31401 2921
rect 28877 2867 28917 2875
rect 28877 2845 28885 2867
rect 28909 2845 28917 2867
rect 28482 2616 28519 2622
rect 28482 2597 28490 2616
rect 28511 2597 28519 2616
rect 28482 2589 28519 2597
rect 28182 2468 28189 2490
rect 28213 2468 28221 2490
rect 28182 2462 28221 2468
rect 27712 2457 27752 2459
rect 27878 2458 28046 2459
rect 27980 2457 28017 2458
rect 26946 2441 27084 2450
rect 26740 2440 26777 2441
rect 26470 2387 26511 2388
rect 26244 2366 26296 2384
rect 26362 2380 26511 2387
rect 25799 2347 25839 2357
rect 26362 2360 26421 2380
rect 26441 2360 26480 2380
rect 26500 2360 26511 2380
rect 26362 2352 26511 2360
rect 26578 2383 26735 2390
rect 26578 2363 26698 2383
rect 26718 2363 26735 2383
rect 26578 2353 26735 2363
rect 26578 2352 26613 2353
rect 25629 2330 25667 2339
rect 26578 2331 26609 2352
rect 26796 2331 26832 2441
rect 26851 2440 26888 2441
rect 26947 2440 26984 2441
rect 26907 2381 26997 2387
rect 26907 2361 26916 2381
rect 26936 2379 26997 2381
rect 26936 2361 26961 2379
rect 26907 2359 26961 2361
rect 26981 2359 26997 2379
rect 26907 2353 26997 2359
rect 26421 2330 26458 2331
rect 25629 2329 25666 2330
rect 25090 2301 25180 2307
rect 25090 2281 25106 2301
rect 25126 2299 25180 2301
rect 25126 2281 25151 2299
rect 25090 2279 25151 2281
rect 25171 2279 25180 2299
rect 25090 2273 25180 2279
rect 25103 2219 25140 2220
rect 25199 2219 25236 2220
rect 25255 2219 25291 2329
rect 25478 2308 25509 2329
rect 26420 2321 26458 2330
rect 25474 2307 25509 2308
rect 25352 2297 25509 2307
rect 25352 2277 25369 2297
rect 25389 2277 25509 2297
rect 25352 2270 25509 2277
rect 25576 2300 25725 2308
rect 25576 2280 25587 2300
rect 25607 2280 25646 2300
rect 25666 2280 25725 2300
rect 26248 2303 26288 2313
rect 25576 2273 25725 2280
rect 25791 2276 25843 2294
rect 25576 2272 25617 2273
rect 25310 2219 25347 2220
rect 25003 2210 25141 2219
rect 24475 2199 24508 2201
rect 24104 2187 24551 2199
rect 23336 2065 23504 2067
rect 23060 2039 23504 2065
rect 22570 2017 22708 2026
rect 22364 2016 22401 2017
rect 21861 1962 21898 1965
rect 22094 1963 22135 1964
rect 20217 1940 20248 1941
rect 19841 1880 20182 1881
rect 20363 1880 20400 1951
rect 21986 1956 22135 1963
rect 21430 1943 21467 1948
rect 21421 1939 21468 1943
rect 21421 1921 21440 1939
rect 21458 1921 21468 1939
rect 21986 1936 22045 1956
rect 22065 1936 22104 1956
rect 22124 1936 22135 1956
rect 21986 1928 22135 1936
rect 22202 1959 22359 1966
rect 22202 1939 22322 1959
rect 22342 1939 22359 1959
rect 22202 1929 22359 1939
rect 22202 1928 22237 1929
rect 19766 1875 20182 1880
rect 19766 1855 19769 1875
rect 19789 1855 20182 1875
rect 20213 1856 20400 1880
rect 21025 1878 21065 1883
rect 21421 1878 21468 1921
rect 22202 1907 22233 1928
rect 22420 1907 22456 2017
rect 22475 2016 22512 2017
rect 22571 2016 22608 2017
rect 22531 1957 22621 1963
rect 22531 1937 22540 1957
rect 22560 1955 22621 1957
rect 22560 1937 22585 1955
rect 22531 1935 22585 1937
rect 22605 1935 22621 1955
rect 22531 1929 22621 1935
rect 22045 1906 22082 1907
rect 21025 1839 21468 1878
rect 21858 1898 21895 1900
rect 21858 1890 21900 1898
rect 21858 1872 21868 1890
rect 21886 1872 21900 1890
rect 21858 1863 21900 1872
rect 22044 1897 22082 1906
rect 22044 1877 22053 1897
rect 22073 1877 22082 1897
rect 22044 1869 22082 1877
rect 22148 1901 22233 1907
rect 22263 1906 22300 1907
rect 22148 1881 22156 1901
rect 22176 1881 22233 1901
rect 22148 1873 22233 1881
rect 22262 1897 22300 1906
rect 22262 1877 22271 1897
rect 22291 1877 22300 1897
rect 22148 1872 22184 1873
rect 22262 1869 22300 1877
rect 22366 1905 22510 1907
rect 22366 1901 22418 1905
rect 22366 1881 22374 1901
rect 22394 1885 22418 1901
rect 22438 1901 22510 1905
rect 22438 1885 22482 1901
rect 22394 1881 22482 1885
rect 22502 1881 22510 1901
rect 22366 1873 22510 1881
rect 22366 1872 22402 1873
rect 22474 1872 22510 1873
rect 22576 1906 22613 1907
rect 22576 1905 22614 1906
rect 22576 1897 22640 1905
rect 22576 1877 22585 1897
rect 22605 1883 22640 1897
rect 22660 1883 22663 1903
rect 22605 1878 22663 1883
rect 22605 1877 22640 1878
rect 18806 1780 18814 1802
rect 18838 1780 18846 1802
rect 18806 1772 18846 1780
rect 20119 1824 20159 1832
rect 20119 1802 20127 1824
rect 20151 1802 20159 1824
rect 16981 1736 17018 1737
rect 16442 1708 16532 1714
rect 16442 1688 16458 1708
rect 16478 1706 16532 1708
rect 16478 1688 16503 1706
rect 16442 1686 16503 1688
rect 16523 1686 16532 1706
rect 16442 1680 16532 1686
rect 16455 1626 16492 1627
rect 16551 1626 16588 1627
rect 16607 1626 16643 1736
rect 16830 1715 16861 1736
rect 17497 1726 17940 1765
rect 16826 1714 16861 1715
rect 16704 1704 16861 1714
rect 16704 1684 16721 1704
rect 16741 1684 16861 1704
rect 16704 1677 16861 1684
rect 16928 1707 17077 1715
rect 16928 1687 16939 1707
rect 16959 1687 16998 1707
rect 17018 1687 17077 1707
rect 16928 1680 17077 1687
rect 17497 1683 17544 1726
rect 17900 1721 17940 1726
rect 18565 1724 18752 1748
rect 18783 1729 19176 1749
rect 19196 1729 19199 1749
rect 18783 1724 19199 1729
rect 16928 1679 16969 1680
rect 17165 1678 17202 1681
rect 16662 1626 16699 1627
rect 16355 1617 16493 1626
rect 15559 1578 16003 1604
rect 15559 1576 15727 1578
rect 14512 1444 14959 1456
rect 14555 1442 14588 1444
rect 13922 1424 14060 1433
rect 13716 1423 13753 1424
rect 13446 1370 13487 1371
rect 13220 1349 13272 1367
rect 13338 1363 13487 1370
rect 12788 1329 12828 1339
rect 13338 1343 13397 1363
rect 13417 1343 13456 1363
rect 13476 1343 13487 1363
rect 13338 1335 13487 1343
rect 13554 1366 13711 1373
rect 13554 1346 13674 1366
rect 13694 1346 13711 1366
rect 13554 1336 13711 1346
rect 13554 1335 13589 1336
rect 12618 1312 12656 1321
rect 13554 1314 13585 1335
rect 13772 1314 13808 1424
rect 13827 1423 13864 1424
rect 13923 1423 13960 1424
rect 13883 1364 13973 1370
rect 13883 1344 13892 1364
rect 13912 1362 13973 1364
rect 13912 1344 13937 1362
rect 13883 1342 13937 1344
rect 13957 1342 13973 1362
rect 13883 1336 13973 1342
rect 13397 1313 13434 1314
rect 12618 1311 12655 1312
rect 12079 1283 12169 1289
rect 12079 1263 12095 1283
rect 12115 1281 12169 1283
rect 12115 1263 12140 1281
rect 12079 1261 12140 1263
rect 12160 1261 12169 1281
rect 12079 1255 12169 1261
rect 12092 1201 12129 1202
rect 12188 1201 12225 1202
rect 12244 1201 12280 1311
rect 12467 1290 12498 1311
rect 13396 1304 13434 1313
rect 12463 1289 12498 1290
rect 12341 1279 12498 1289
rect 12341 1259 12358 1279
rect 12378 1259 12498 1279
rect 12341 1252 12498 1259
rect 12565 1282 12714 1290
rect 12565 1262 12576 1282
rect 12596 1262 12635 1282
rect 12655 1262 12714 1282
rect 13224 1286 13264 1296
rect 12565 1255 12714 1262
rect 12780 1258 12832 1276
rect 12565 1254 12606 1255
rect 12299 1201 12336 1202
rect 11992 1192 12130 1201
rect 11992 1172 12101 1192
rect 12121 1172 12130 1192
rect 11992 1165 12130 1172
rect 12188 1192 12336 1201
rect 12188 1172 12197 1192
rect 12217 1172 12307 1192
rect 12327 1172 12336 1192
rect 11992 1163 12088 1165
rect 12188 1162 12336 1172
rect 12395 1192 12432 1202
rect 12395 1172 12403 1192
rect 12423 1172 12432 1192
rect 12244 1161 12280 1162
rect 12395 1105 12432 1172
rect 12467 1201 12498 1252
rect 12780 1240 12798 1258
rect 12816 1240 12832 1258
rect 12517 1201 12554 1202
rect 12467 1192 12554 1201
rect 12467 1172 12525 1192
rect 12545 1172 12554 1192
rect 12467 1162 12554 1172
rect 12613 1192 12650 1202
rect 12613 1172 12621 1192
rect 12641 1172 12650 1192
rect 12467 1161 12498 1162
rect 12092 1102 12129 1103
rect 12395 1102 12434 1105
rect 12091 1101 12434 1102
rect 12613 1101 12650 1172
rect 12016 1096 12434 1101
rect 12016 1076 12019 1096
rect 12039 1076 12434 1096
rect 12463 1077 12650 1101
rect 10557 1045 10594 1053
rect 10557 1026 10565 1045
rect 10586 1026 10594 1045
rect 10557 1020 10594 1026
rect 12395 1051 12434 1076
rect 12780 1051 12832 1240
rect 13224 1268 13234 1286
rect 13252 1268 13264 1286
rect 13396 1284 13405 1304
rect 13425 1284 13434 1304
rect 13396 1276 13434 1284
rect 13500 1308 13585 1314
rect 13615 1313 13652 1314
rect 13500 1288 13508 1308
rect 13528 1288 13585 1308
rect 13500 1280 13585 1288
rect 13614 1304 13652 1313
rect 13614 1284 13623 1304
rect 13643 1284 13652 1304
rect 13500 1279 13536 1280
rect 13614 1276 13652 1284
rect 13718 1308 13862 1314
rect 13718 1288 13726 1308
rect 13746 1288 13779 1308
rect 13799 1288 13834 1308
rect 13854 1288 13862 1308
rect 13718 1280 13862 1288
rect 13718 1279 13754 1280
rect 13826 1279 13862 1280
rect 13928 1313 13965 1314
rect 13928 1312 13966 1313
rect 13928 1304 13992 1312
rect 13928 1284 13937 1304
rect 13957 1290 13992 1304
rect 14012 1290 14015 1310
rect 13957 1285 14015 1290
rect 13957 1284 13992 1285
rect 13224 1212 13264 1268
rect 13397 1247 13434 1276
rect 13398 1245 13434 1247
rect 13398 1223 13589 1245
rect 13615 1244 13652 1276
rect 13928 1272 13992 1284
rect 14032 1246 14059 1424
rect 14917 1399 14959 1444
rect 13891 1244 14059 1246
rect 13615 1234 14059 1244
rect 14200 1340 14387 1364
rect 14418 1345 14811 1365
rect 14831 1345 14834 1365
rect 14418 1340 14834 1345
rect 14200 1269 14237 1340
rect 14418 1339 14759 1340
rect 14352 1279 14383 1280
rect 14200 1249 14209 1269
rect 14229 1249 14237 1269
rect 14200 1239 14237 1249
rect 14296 1269 14383 1279
rect 14296 1249 14305 1269
rect 14325 1249 14383 1269
rect 14296 1240 14383 1249
rect 14296 1239 14333 1240
rect 13221 1207 13264 1212
rect 13612 1218 14059 1234
rect 13612 1212 13640 1218
rect 13891 1217 14059 1218
rect 13221 1204 13371 1207
rect 13612 1204 13639 1212
rect 13221 1202 13639 1204
rect 13221 1184 13230 1202
rect 13248 1184 13639 1202
rect 14352 1189 14383 1240
rect 14418 1269 14455 1339
rect 14721 1338 14758 1339
rect 14570 1279 14606 1280
rect 14418 1249 14427 1269
rect 14447 1249 14455 1269
rect 14418 1239 14455 1249
rect 14514 1269 14662 1279
rect 14762 1276 14858 1278
rect 14514 1249 14523 1269
rect 14543 1249 14633 1269
rect 14653 1249 14662 1269
rect 14514 1240 14662 1249
rect 14720 1269 14858 1276
rect 14720 1249 14729 1269
rect 14749 1249 14858 1269
rect 14720 1240 14858 1249
rect 14514 1239 14551 1240
rect 14244 1186 14285 1187
rect 13221 1181 13639 1184
rect 13221 1175 13264 1181
rect 13224 1172 13264 1175
rect 14139 1179 14285 1186
rect 13621 1163 13661 1164
rect 13332 1146 13661 1163
rect 14139 1159 14195 1179
rect 14215 1159 14254 1179
rect 14274 1159 14285 1179
rect 14139 1151 14285 1159
rect 14352 1182 14509 1189
rect 14352 1162 14472 1182
rect 14492 1162 14509 1182
rect 14352 1152 14509 1162
rect 14352 1151 14387 1152
rect 13216 1103 13259 1114
rect 13216 1085 13228 1103
rect 13246 1085 13259 1103
rect 13216 1059 13259 1085
rect 13332 1059 13359 1146
rect 13621 1137 13661 1146
rect 12395 1033 12834 1051
rect 12395 1015 12795 1033
rect 12813 1015 12834 1033
rect 12395 1009 12834 1015
rect 12401 1005 12834 1009
rect 13216 1038 13359 1059
rect 13403 1111 13437 1127
rect 13621 1117 14014 1137
rect 14034 1117 14037 1137
rect 14352 1130 14383 1151
rect 14570 1130 14606 1240
rect 14625 1239 14662 1240
rect 14721 1239 14758 1240
rect 14681 1180 14771 1186
rect 14681 1160 14690 1180
rect 14710 1178 14771 1180
rect 14710 1160 14735 1178
rect 14681 1158 14735 1160
rect 14755 1158 14771 1178
rect 14681 1152 14771 1158
rect 14195 1129 14232 1130
rect 13621 1112 14037 1117
rect 14194 1120 14232 1129
rect 13621 1111 13962 1112
rect 13403 1041 13440 1111
rect 13555 1051 13586 1052
rect 13216 1036 13353 1038
rect 12780 1003 12832 1005
rect 13216 994 13259 1036
rect 13403 1021 13412 1041
rect 13432 1021 13440 1041
rect 13403 1011 13440 1021
rect 13499 1041 13586 1051
rect 13499 1021 13508 1041
rect 13528 1021 13586 1041
rect 13499 1012 13586 1021
rect 13499 1011 13536 1012
rect 13214 984 13259 994
rect 13214 966 13223 984
rect 13241 966 13259 984
rect 13214 960 13259 966
rect 13555 961 13586 1012
rect 13621 1041 13658 1111
rect 13924 1110 13961 1111
rect 14194 1100 14203 1120
rect 14223 1100 14232 1120
rect 14194 1092 14232 1100
rect 14298 1124 14383 1130
rect 14413 1129 14450 1130
rect 14298 1104 14306 1124
rect 14326 1104 14383 1124
rect 14298 1096 14383 1104
rect 14412 1120 14450 1129
rect 14412 1100 14421 1120
rect 14441 1100 14450 1120
rect 14298 1095 14334 1096
rect 14412 1092 14450 1100
rect 14516 1124 14660 1130
rect 14516 1104 14524 1124
rect 14544 1121 14632 1124
rect 14544 1104 14579 1121
rect 14516 1103 14579 1104
rect 14598 1104 14632 1121
rect 14652 1104 14660 1124
rect 14598 1103 14660 1104
rect 14516 1096 14660 1103
rect 14516 1095 14552 1096
rect 14624 1095 14660 1096
rect 14726 1129 14763 1130
rect 14726 1128 14764 1129
rect 14786 1128 14813 1132
rect 14726 1126 14813 1128
rect 14726 1120 14790 1126
rect 14726 1100 14735 1120
rect 14755 1106 14790 1120
rect 14810 1106 14813 1126
rect 14755 1101 14813 1106
rect 14755 1100 14790 1101
rect 14195 1063 14232 1092
rect 14196 1061 14232 1063
rect 13773 1051 13809 1052
rect 13621 1021 13630 1041
rect 13650 1021 13658 1041
rect 13621 1011 13658 1021
rect 13717 1041 13865 1051
rect 13965 1048 14061 1050
rect 13717 1021 13726 1041
rect 13746 1021 13836 1041
rect 13856 1021 13865 1041
rect 13717 1012 13865 1021
rect 13923 1041 14061 1048
rect 13923 1021 13932 1041
rect 13952 1021 14061 1041
rect 14196 1039 14387 1061
rect 14413 1060 14450 1092
rect 14726 1088 14790 1100
rect 14830 1062 14857 1240
rect 14689 1060 14857 1062
rect 14413 1034 14857 1060
rect 13923 1012 14061 1021
rect 13717 1011 13754 1012
rect 13214 957 13251 960
rect 13447 958 13488 959
rect 13339 951 13488 958
rect 12783 938 12820 943
rect 12774 934 12821 938
rect 12774 916 12793 934
rect 12811 916 12821 934
rect 13339 931 13398 951
rect 13418 931 13457 951
rect 13477 931 13488 951
rect 13339 923 13488 931
rect 13555 954 13712 961
rect 13555 934 13675 954
rect 13695 934 13712 954
rect 13555 924 13712 934
rect 13555 923 13590 924
rect 12774 853 12821 916
rect 13555 902 13586 923
rect 13773 902 13809 1012
rect 13828 1011 13865 1012
rect 13924 1011 13961 1012
rect 13884 952 13974 958
rect 13884 932 13893 952
rect 13913 950 13974 952
rect 13913 932 13938 950
rect 13884 930 13938 932
rect 13958 930 13974 950
rect 13884 924 13974 930
rect 13398 901 13435 902
rect 13211 893 13248 895
rect 13211 885 13253 893
rect 13211 867 13221 885
rect 13239 867 13253 885
rect 13211 858 13253 867
rect 13397 892 13435 901
rect 13397 872 13406 892
rect 13426 872 13435 892
rect 13397 864 13435 872
rect 13501 896 13586 902
rect 13616 901 13653 902
rect 13501 876 13509 896
rect 13529 876 13586 896
rect 13501 868 13586 876
rect 13615 892 13653 901
rect 13615 872 13624 892
rect 13644 872 13653 892
rect 13501 867 13537 868
rect 13615 864 13653 872
rect 13719 900 13863 902
rect 13719 896 13771 900
rect 13719 876 13727 896
rect 13747 880 13771 896
rect 13791 896 13863 900
rect 13791 880 13835 896
rect 13747 876 13835 880
rect 13855 876 13863 896
rect 13719 868 13863 876
rect 13719 867 13755 868
rect 13827 867 13863 868
rect 13929 901 13966 902
rect 13929 900 13967 901
rect 13929 892 13993 900
rect 13929 872 13938 892
rect 13958 878 13993 892
rect 14013 878 14016 898
rect 13958 873 14016 878
rect 13958 872 13993 873
rect 12774 838 12824 853
rect 12774 813 12788 838
rect 12820 813 12824 838
rect 13212 833 13253 858
rect 13398 833 13435 864
rect 13616 842 13653 864
rect 13929 860 13993 872
rect 13611 833 13653 842
rect 14033 834 14060 1012
rect 13212 821 13257 833
rect 12774 800 12821 813
rect 10159 775 10167 797
rect 10191 775 10199 797
rect 10159 767 10199 775
rect 13208 763 13257 821
rect 13398 807 13460 833
rect 13611 832 13696 833
rect 13892 832 14060 834
rect 13611 806 14060 832
rect 13611 763 13650 806
rect 13892 805 14060 806
rect 14523 810 14563 1034
rect 14689 1033 14857 1034
rect 14921 1066 14954 1399
rect 15559 1398 15586 1576
rect 15626 1538 15690 1550
rect 15966 1546 16003 1578
rect 16029 1577 16220 1599
rect 16355 1597 16464 1617
rect 16484 1597 16493 1617
rect 16355 1590 16493 1597
rect 16551 1617 16699 1626
rect 16551 1597 16560 1617
rect 16580 1597 16670 1617
rect 16690 1597 16699 1617
rect 16355 1588 16451 1590
rect 16551 1587 16699 1597
rect 16758 1617 16795 1627
rect 16758 1597 16766 1617
rect 16786 1597 16795 1617
rect 16607 1586 16643 1587
rect 16184 1575 16220 1577
rect 16184 1546 16221 1575
rect 15626 1537 15661 1538
rect 15603 1532 15661 1537
rect 15603 1512 15606 1532
rect 15626 1518 15661 1532
rect 15681 1518 15690 1538
rect 15626 1510 15690 1518
rect 15652 1509 15690 1510
rect 15653 1508 15690 1509
rect 15756 1542 15792 1543
rect 15864 1542 15900 1543
rect 15756 1534 15900 1542
rect 15756 1514 15764 1534
rect 15784 1533 15872 1534
rect 15784 1514 15819 1533
rect 15840 1514 15872 1533
rect 15892 1514 15900 1534
rect 15756 1508 15900 1514
rect 15966 1538 16004 1546
rect 16082 1542 16118 1543
rect 15966 1518 15975 1538
rect 15995 1518 16004 1538
rect 15966 1509 16004 1518
rect 16033 1534 16118 1542
rect 16033 1514 16090 1534
rect 16110 1514 16118 1534
rect 15966 1508 16003 1509
rect 16033 1508 16118 1514
rect 16184 1538 16222 1546
rect 16184 1518 16193 1538
rect 16213 1518 16222 1538
rect 16455 1527 16492 1528
rect 16758 1527 16795 1597
rect 16830 1626 16861 1677
rect 17157 1672 17202 1678
rect 17157 1654 17175 1672
rect 17193 1654 17202 1672
rect 17497 1665 17507 1683
rect 17525 1665 17544 1683
rect 17497 1661 17544 1665
rect 17498 1656 17535 1661
rect 17157 1644 17202 1654
rect 18565 1653 18602 1724
rect 18783 1723 19124 1724
rect 18717 1663 18748 1664
rect 16880 1626 16917 1627
rect 16830 1617 16917 1626
rect 16830 1597 16888 1617
rect 16908 1597 16917 1617
rect 16830 1587 16917 1597
rect 16976 1617 17013 1627
rect 16976 1597 16984 1617
rect 17004 1597 17013 1617
rect 17157 1602 17200 1644
rect 18565 1633 18574 1653
rect 18594 1633 18602 1653
rect 18565 1623 18602 1633
rect 18661 1653 18748 1663
rect 18661 1633 18670 1653
rect 18690 1633 18748 1653
rect 18661 1624 18748 1633
rect 18661 1623 18698 1624
rect 17063 1600 17200 1602
rect 16830 1586 16861 1587
rect 16976 1527 17013 1597
rect 16454 1526 16795 1527
rect 16184 1509 16222 1518
rect 16379 1521 16795 1526
rect 16184 1508 16221 1509
rect 15645 1480 15735 1486
rect 15645 1460 15661 1480
rect 15681 1478 15735 1480
rect 15681 1460 15706 1478
rect 15645 1458 15706 1460
rect 15726 1458 15735 1478
rect 15645 1452 15735 1458
rect 15658 1398 15695 1399
rect 15754 1398 15791 1399
rect 15810 1398 15846 1508
rect 16033 1487 16064 1508
rect 16379 1501 16382 1521
rect 16402 1501 16795 1521
rect 16979 1511 17013 1527
rect 17057 1579 17200 1600
rect 17486 1594 17538 1596
rect 16755 1492 16795 1501
rect 17057 1492 17084 1579
rect 17157 1553 17200 1579
rect 17157 1535 17170 1553
rect 17188 1535 17200 1553
rect 17484 1590 17917 1594
rect 17484 1584 17923 1590
rect 17484 1566 17505 1584
rect 17523 1566 17923 1584
rect 18717 1573 18748 1624
rect 18783 1653 18820 1723
rect 19086 1722 19123 1723
rect 18935 1663 18971 1664
rect 18783 1633 18792 1653
rect 18812 1633 18820 1653
rect 18783 1623 18820 1633
rect 18879 1653 19027 1663
rect 19127 1660 19223 1662
rect 18879 1633 18888 1653
rect 18908 1633 18998 1653
rect 19018 1633 19027 1653
rect 18879 1624 19027 1633
rect 19085 1653 19223 1660
rect 19085 1633 19094 1653
rect 19114 1633 19223 1653
rect 19085 1624 19223 1633
rect 18879 1623 18916 1624
rect 18609 1570 18650 1571
rect 17484 1548 17923 1566
rect 17157 1524 17200 1535
rect 16029 1486 16064 1487
rect 15907 1476 16064 1486
rect 15907 1456 15924 1476
rect 15944 1456 16064 1476
rect 15907 1449 16064 1456
rect 16131 1479 16280 1487
rect 16131 1459 16142 1479
rect 16162 1459 16201 1479
rect 16221 1459 16280 1479
rect 16755 1475 17084 1492
rect 16755 1474 16795 1475
rect 16131 1452 16280 1459
rect 17152 1463 17192 1466
rect 17152 1457 17195 1463
rect 16777 1454 17195 1457
rect 16131 1451 16172 1452
rect 15865 1398 15902 1399
rect 15558 1389 15696 1398
rect 15558 1369 15667 1389
rect 15687 1369 15696 1389
rect 15558 1362 15696 1369
rect 15754 1389 15902 1398
rect 15754 1369 15763 1389
rect 15783 1369 15873 1389
rect 15893 1369 15902 1389
rect 15558 1360 15654 1362
rect 15754 1359 15902 1369
rect 15961 1389 15998 1399
rect 15961 1369 15969 1389
rect 15989 1369 15998 1389
rect 15810 1358 15846 1359
rect 15658 1299 15695 1300
rect 15961 1299 15998 1369
rect 16033 1398 16064 1449
rect 16777 1436 17168 1454
rect 17186 1436 17195 1454
rect 16777 1434 17195 1436
rect 16777 1426 16804 1434
rect 17045 1431 17195 1434
rect 16357 1420 16525 1421
rect 16776 1420 16804 1426
rect 16357 1404 16804 1420
rect 17152 1426 17195 1431
rect 16083 1398 16120 1399
rect 16033 1389 16120 1398
rect 16033 1369 16091 1389
rect 16111 1369 16120 1389
rect 16033 1359 16120 1369
rect 16179 1389 16216 1399
rect 16179 1369 16187 1389
rect 16207 1369 16216 1389
rect 16033 1358 16064 1359
rect 15657 1298 15998 1299
rect 16179 1298 16216 1369
rect 15582 1293 15998 1298
rect 15582 1273 15585 1293
rect 15605 1273 15998 1293
rect 16029 1274 16216 1298
rect 16357 1394 16801 1404
rect 16357 1392 16525 1394
rect 16357 1214 16384 1392
rect 16424 1354 16488 1366
rect 16764 1362 16801 1394
rect 16827 1393 17018 1415
rect 16982 1391 17018 1393
rect 16982 1362 17019 1391
rect 17152 1370 17192 1426
rect 16424 1353 16459 1354
rect 16401 1348 16459 1353
rect 16401 1328 16404 1348
rect 16424 1334 16459 1348
rect 16479 1334 16488 1354
rect 16424 1326 16488 1334
rect 16450 1325 16488 1326
rect 16451 1324 16488 1325
rect 16554 1358 16590 1359
rect 16662 1358 16698 1359
rect 16554 1350 16698 1358
rect 16554 1330 16562 1350
rect 16582 1330 16617 1350
rect 16637 1330 16670 1350
rect 16690 1330 16698 1350
rect 16554 1324 16698 1330
rect 16764 1354 16802 1362
rect 16880 1358 16916 1359
rect 16764 1334 16773 1354
rect 16793 1334 16802 1354
rect 16764 1325 16802 1334
rect 16831 1350 16916 1358
rect 16831 1330 16888 1350
rect 16908 1330 16916 1350
rect 16764 1324 16801 1325
rect 16831 1324 16916 1330
rect 16982 1354 17020 1362
rect 16982 1334 16991 1354
rect 17011 1334 17020 1354
rect 17152 1352 17164 1370
rect 17182 1352 17192 1370
rect 17152 1342 17192 1352
rect 17486 1359 17538 1548
rect 17884 1523 17923 1548
rect 18501 1563 18650 1570
rect 18501 1543 18560 1563
rect 18580 1543 18619 1563
rect 18639 1543 18650 1563
rect 18501 1535 18650 1543
rect 18717 1566 18874 1573
rect 18717 1546 18837 1566
rect 18857 1546 18874 1566
rect 18717 1536 18874 1546
rect 18717 1535 18752 1536
rect 17668 1498 17855 1522
rect 17884 1503 18279 1523
rect 18299 1503 18302 1523
rect 18717 1514 18748 1535
rect 18935 1514 18971 1624
rect 18990 1623 19027 1624
rect 19086 1623 19123 1624
rect 19046 1564 19136 1570
rect 19046 1544 19055 1564
rect 19075 1562 19136 1564
rect 19075 1544 19100 1562
rect 19046 1542 19100 1544
rect 19120 1542 19136 1562
rect 19046 1536 19136 1542
rect 18560 1513 18597 1514
rect 17884 1498 18302 1503
rect 18559 1504 18597 1513
rect 17668 1427 17705 1498
rect 17884 1497 18227 1498
rect 17884 1494 17923 1497
rect 18189 1496 18226 1497
rect 17820 1437 17851 1438
rect 17668 1407 17677 1427
rect 17697 1407 17705 1427
rect 17668 1397 17705 1407
rect 17764 1427 17851 1437
rect 17764 1407 17773 1427
rect 17793 1407 17851 1427
rect 17764 1398 17851 1407
rect 17764 1397 17801 1398
rect 16982 1325 17020 1334
rect 17486 1341 17502 1359
rect 17520 1341 17538 1359
rect 17820 1347 17851 1398
rect 17886 1427 17923 1494
rect 18559 1484 18568 1504
rect 18588 1484 18597 1504
rect 18559 1476 18597 1484
rect 18663 1508 18748 1514
rect 18778 1513 18815 1514
rect 18663 1488 18671 1508
rect 18691 1488 18748 1508
rect 18663 1480 18748 1488
rect 18777 1504 18815 1513
rect 18777 1484 18786 1504
rect 18806 1484 18815 1504
rect 18663 1479 18699 1480
rect 18777 1476 18815 1484
rect 18881 1508 19025 1514
rect 18881 1488 18889 1508
rect 18909 1503 18997 1508
rect 18909 1488 18945 1503
rect 18881 1486 18945 1488
rect 18964 1488 18997 1503
rect 19017 1488 19025 1508
rect 18964 1486 19025 1488
rect 18881 1480 19025 1486
rect 18881 1479 18917 1480
rect 18989 1479 19025 1480
rect 19091 1513 19128 1514
rect 19091 1512 19129 1513
rect 19091 1504 19155 1512
rect 19091 1484 19100 1504
rect 19120 1490 19155 1504
rect 19175 1490 19178 1510
rect 19120 1485 19178 1490
rect 19120 1484 19155 1485
rect 18560 1447 18597 1476
rect 18561 1445 18597 1447
rect 18038 1437 18074 1438
rect 17886 1407 17895 1427
rect 17915 1407 17923 1427
rect 17886 1397 17923 1407
rect 17982 1427 18130 1437
rect 18230 1434 18326 1436
rect 17982 1407 17991 1427
rect 18011 1407 18101 1427
rect 18121 1407 18130 1427
rect 17982 1398 18130 1407
rect 18188 1427 18326 1434
rect 18188 1407 18197 1427
rect 18217 1407 18326 1427
rect 18561 1423 18752 1445
rect 18778 1444 18815 1476
rect 19091 1472 19155 1484
rect 19195 1446 19222 1624
rect 19054 1444 19222 1446
rect 18778 1430 19222 1444
rect 19825 1578 19993 1579
rect 20119 1578 20159 1802
rect 20622 1806 20790 1807
rect 21025 1806 21065 1839
rect 21421 1806 21468 1839
rect 21859 1838 21900 1863
rect 22045 1838 22082 1869
rect 22263 1838 22300 1869
rect 22576 1865 22640 1877
rect 22680 1839 22707 2017
rect 21859 1811 21908 1838
rect 22044 1812 22093 1838
rect 22262 1837 22343 1838
rect 22539 1837 22707 1839
rect 22262 1812 22707 1837
rect 22263 1811 22707 1812
rect 20622 1805 21066 1806
rect 20622 1780 21067 1805
rect 20622 1778 20790 1780
rect 20986 1779 21067 1780
rect 21236 1779 21285 1805
rect 21421 1779 21470 1806
rect 20622 1600 20649 1778
rect 20689 1740 20753 1752
rect 21029 1748 21066 1779
rect 21247 1748 21284 1779
rect 21429 1754 21470 1779
rect 21861 1778 21908 1811
rect 22264 1778 22304 1811
rect 22539 1810 22707 1811
rect 23170 1815 23210 2039
rect 23336 2038 23504 2039
rect 24107 2173 24551 2187
rect 24107 2171 24275 2173
rect 24107 1993 24134 2171
rect 24174 2133 24238 2145
rect 24514 2141 24551 2173
rect 24577 2172 24768 2194
rect 25003 2190 25112 2210
rect 25132 2190 25141 2210
rect 25003 2183 25141 2190
rect 25199 2210 25347 2219
rect 25199 2190 25208 2210
rect 25228 2190 25318 2210
rect 25338 2190 25347 2210
rect 25003 2181 25099 2183
rect 25199 2180 25347 2190
rect 25406 2210 25443 2220
rect 25406 2190 25414 2210
rect 25434 2190 25443 2210
rect 25255 2179 25291 2180
rect 24732 2170 24768 2172
rect 24732 2141 24769 2170
rect 24174 2132 24209 2133
rect 24151 2127 24209 2132
rect 24151 2107 24154 2127
rect 24174 2113 24209 2127
rect 24229 2113 24238 2133
rect 24174 2105 24238 2113
rect 24200 2104 24238 2105
rect 24201 2103 24238 2104
rect 24304 2137 24340 2138
rect 24412 2137 24448 2138
rect 24304 2129 24448 2137
rect 24304 2109 24312 2129
rect 24332 2127 24420 2129
rect 24332 2109 24365 2127
rect 24304 2108 24365 2109
rect 24386 2109 24420 2127
rect 24440 2109 24448 2129
rect 24386 2108 24448 2109
rect 24304 2103 24448 2108
rect 24514 2133 24552 2141
rect 24630 2137 24666 2138
rect 24514 2113 24523 2133
rect 24543 2113 24552 2133
rect 24514 2104 24552 2113
rect 24581 2129 24666 2137
rect 24581 2109 24638 2129
rect 24658 2109 24666 2129
rect 24514 2103 24551 2104
rect 24581 2103 24666 2109
rect 24732 2133 24770 2141
rect 24732 2113 24741 2133
rect 24761 2113 24770 2133
rect 25406 2123 25443 2190
rect 25478 2219 25509 2270
rect 25791 2258 25809 2276
rect 25827 2258 25843 2276
rect 25528 2219 25565 2220
rect 25478 2210 25565 2219
rect 25478 2190 25536 2210
rect 25556 2190 25565 2210
rect 25478 2180 25565 2190
rect 25624 2210 25661 2220
rect 25624 2190 25632 2210
rect 25652 2190 25661 2210
rect 25478 2179 25509 2180
rect 25103 2120 25140 2121
rect 25406 2120 25445 2123
rect 25102 2119 25445 2120
rect 25624 2119 25661 2190
rect 24732 2104 24770 2113
rect 25027 2114 25445 2119
rect 24732 2103 24769 2104
rect 24193 2075 24283 2081
rect 24193 2055 24209 2075
rect 24229 2073 24283 2075
rect 24229 2055 24254 2073
rect 24193 2053 24254 2055
rect 24274 2053 24283 2073
rect 24193 2047 24283 2053
rect 24206 1993 24243 1994
rect 24302 1993 24339 1994
rect 24358 1993 24394 2103
rect 24581 2082 24612 2103
rect 25027 2094 25030 2114
rect 25050 2094 25445 2114
rect 25474 2095 25661 2119
rect 24577 2081 24612 2082
rect 24455 2071 24612 2081
rect 24455 2051 24472 2071
rect 24492 2051 24612 2071
rect 24455 2044 24612 2051
rect 24679 2074 24828 2082
rect 24679 2054 24690 2074
rect 24710 2054 24749 2074
rect 24769 2054 24828 2074
rect 24679 2047 24828 2054
rect 25406 2069 25445 2094
rect 25791 2069 25843 2258
rect 26248 2285 26258 2303
rect 26276 2285 26288 2303
rect 26420 2301 26429 2321
rect 26449 2301 26458 2321
rect 26420 2293 26458 2301
rect 26524 2325 26609 2331
rect 26639 2330 26676 2331
rect 26524 2305 26532 2325
rect 26552 2305 26609 2325
rect 26524 2297 26609 2305
rect 26638 2321 26676 2330
rect 26638 2301 26647 2321
rect 26667 2301 26676 2321
rect 26524 2296 26560 2297
rect 26638 2293 26676 2301
rect 26742 2325 26886 2331
rect 26742 2305 26750 2325
rect 26770 2305 26803 2325
rect 26823 2305 26858 2325
rect 26878 2305 26886 2325
rect 26742 2297 26886 2305
rect 26742 2296 26778 2297
rect 26850 2296 26886 2297
rect 26952 2330 26989 2331
rect 26952 2329 26990 2330
rect 26952 2321 27016 2329
rect 26952 2301 26961 2321
rect 26981 2307 27016 2321
rect 27036 2307 27039 2327
rect 26981 2302 27039 2307
rect 26981 2301 27016 2302
rect 26248 2229 26288 2285
rect 26421 2264 26458 2293
rect 26422 2262 26458 2264
rect 26422 2240 26613 2262
rect 26639 2261 26676 2293
rect 26952 2289 27016 2301
rect 27056 2263 27083 2441
rect 26915 2261 27083 2263
rect 26639 2251 27083 2261
rect 27224 2357 27411 2381
rect 27442 2362 27835 2382
rect 27855 2362 27858 2382
rect 27442 2357 27858 2362
rect 27224 2286 27261 2357
rect 27442 2356 27783 2357
rect 27376 2296 27407 2297
rect 27224 2266 27233 2286
rect 27253 2266 27261 2286
rect 27224 2256 27261 2266
rect 27320 2286 27407 2296
rect 27320 2266 27329 2286
rect 27349 2266 27407 2286
rect 27320 2257 27407 2266
rect 27320 2256 27357 2257
rect 26245 2224 26288 2229
rect 26636 2235 27083 2251
rect 26636 2229 26664 2235
rect 26915 2234 27083 2235
rect 26245 2221 26395 2224
rect 26636 2221 26663 2229
rect 26245 2219 26663 2221
rect 26245 2201 26254 2219
rect 26272 2201 26663 2219
rect 27376 2206 27407 2257
rect 27442 2286 27479 2356
rect 27745 2355 27782 2356
rect 27983 2298 28016 2457
rect 27594 2296 27630 2297
rect 27442 2266 27451 2286
rect 27471 2266 27479 2286
rect 27442 2256 27479 2266
rect 27538 2286 27686 2296
rect 27786 2293 27882 2295
rect 27538 2266 27547 2286
rect 27567 2266 27657 2286
rect 27677 2266 27686 2286
rect 27538 2257 27686 2266
rect 27744 2286 27882 2293
rect 27744 2266 27753 2286
rect 27773 2266 27882 2286
rect 27983 2294 28019 2298
rect 27983 2276 27992 2294
rect 28014 2276 28019 2294
rect 27983 2270 28019 2276
rect 27744 2257 27882 2266
rect 27538 2256 27575 2257
rect 27268 2203 27309 2204
rect 26245 2198 26663 2201
rect 26245 2192 26288 2198
rect 26248 2189 26288 2192
rect 27160 2196 27309 2203
rect 26645 2180 26685 2181
rect 26356 2163 26685 2180
rect 27160 2176 27219 2196
rect 27239 2176 27278 2196
rect 27298 2176 27309 2196
rect 27160 2168 27309 2176
rect 27376 2199 27533 2206
rect 27376 2179 27496 2199
rect 27516 2179 27533 2199
rect 27376 2169 27533 2179
rect 27376 2168 27411 2169
rect 26240 2120 26283 2131
rect 26240 2102 26252 2120
rect 26270 2102 26283 2120
rect 26240 2076 26283 2102
rect 26356 2076 26383 2163
rect 26645 2154 26685 2163
rect 25406 2051 25845 2069
rect 24679 2046 24720 2047
rect 24413 1993 24450 1994
rect 24106 1984 24244 1993
rect 24106 1964 24215 1984
rect 24235 1964 24244 1984
rect 24106 1957 24244 1964
rect 24302 1984 24450 1993
rect 24302 1964 24311 1984
rect 24331 1964 24421 1984
rect 24441 1964 24450 1984
rect 24106 1955 24202 1957
rect 24302 1954 24450 1964
rect 24509 1984 24546 1994
rect 24509 1964 24517 1984
rect 24537 1964 24546 1984
rect 24358 1953 24394 1954
rect 24206 1894 24243 1895
rect 24509 1894 24546 1964
rect 24581 1993 24612 2044
rect 25406 2033 25806 2051
rect 25824 2033 25845 2051
rect 25406 2027 25845 2033
rect 25412 2023 25845 2027
rect 26240 2055 26383 2076
rect 26427 2128 26461 2144
rect 26645 2134 27038 2154
rect 27058 2134 27061 2154
rect 27376 2147 27407 2168
rect 27594 2147 27630 2257
rect 27649 2256 27686 2257
rect 27745 2256 27782 2257
rect 27705 2197 27795 2203
rect 27705 2177 27714 2197
rect 27734 2195 27795 2197
rect 27734 2177 27759 2195
rect 27705 2175 27759 2177
rect 27779 2175 27795 2195
rect 27705 2169 27795 2175
rect 27219 2146 27256 2147
rect 26645 2129 27061 2134
rect 27218 2137 27256 2146
rect 26645 2128 26986 2129
rect 26427 2058 26464 2128
rect 26579 2068 26610 2069
rect 26240 2053 26377 2055
rect 25791 2021 25843 2023
rect 26240 2011 26283 2053
rect 26427 2038 26436 2058
rect 26456 2038 26464 2058
rect 26427 2028 26464 2038
rect 26523 2058 26610 2068
rect 26523 2038 26532 2058
rect 26552 2038 26610 2058
rect 26523 2029 26610 2038
rect 26523 2028 26560 2029
rect 26238 2001 26283 2011
rect 24631 1993 24668 1994
rect 24581 1984 24668 1993
rect 24581 1964 24639 1984
rect 24659 1964 24668 1984
rect 24581 1954 24668 1964
rect 24727 1984 24764 1994
rect 24727 1964 24735 1984
rect 24755 1964 24764 1984
rect 26238 1983 26247 2001
rect 26265 1983 26283 2001
rect 26238 1977 26283 1983
rect 26579 1978 26610 2029
rect 26645 2058 26682 2128
rect 26948 2127 26985 2128
rect 27218 2117 27227 2137
rect 27247 2117 27256 2137
rect 27218 2109 27256 2117
rect 27322 2141 27407 2147
rect 27437 2146 27474 2147
rect 27322 2121 27330 2141
rect 27350 2121 27407 2141
rect 27322 2113 27407 2121
rect 27436 2137 27474 2146
rect 27436 2117 27445 2137
rect 27465 2117 27474 2137
rect 27322 2112 27358 2113
rect 27436 2109 27474 2117
rect 27540 2141 27684 2147
rect 27540 2121 27548 2141
rect 27568 2122 27600 2141
rect 27621 2122 27656 2141
rect 27568 2121 27656 2122
rect 27676 2121 27684 2141
rect 27540 2113 27684 2121
rect 27540 2112 27576 2113
rect 27648 2112 27684 2113
rect 27750 2146 27787 2147
rect 27750 2145 27788 2146
rect 27750 2137 27814 2145
rect 27750 2117 27759 2137
rect 27779 2123 27814 2137
rect 27834 2123 27837 2143
rect 27779 2118 27837 2123
rect 27779 2117 27814 2118
rect 27219 2080 27256 2109
rect 27220 2078 27256 2080
rect 26797 2068 26833 2069
rect 26645 2038 26654 2058
rect 26674 2038 26682 2058
rect 26645 2028 26682 2038
rect 26741 2058 26889 2068
rect 26989 2065 27085 2067
rect 26741 2038 26750 2058
rect 26770 2038 26860 2058
rect 26880 2038 26889 2058
rect 26741 2029 26889 2038
rect 26947 2058 27085 2065
rect 26947 2038 26956 2058
rect 26976 2038 27085 2058
rect 27220 2056 27411 2078
rect 27437 2077 27474 2109
rect 27750 2105 27814 2117
rect 27854 2079 27881 2257
rect 28486 2256 28519 2589
rect 28583 2621 28751 2622
rect 28877 2621 28917 2845
rect 29380 2849 29548 2850
rect 29784 2849 29825 2883
rect 30182 2862 30229 2883
rect 29380 2839 29825 2849
rect 29897 2847 30040 2848
rect 29380 2823 29824 2839
rect 29380 2821 29548 2823
rect 29744 2822 29824 2823
rect 29897 2822 30042 2847
rect 30184 2822 30229 2862
rect 29380 2643 29407 2821
rect 29447 2783 29511 2795
rect 29787 2791 29824 2822
rect 30005 2791 30042 2822
rect 30187 2815 30229 2822
rect 30619 2881 30661 2888
rect 30806 2881 30843 2912
rect 31024 2881 31061 2912
rect 31337 2908 31401 2920
rect 31441 2882 31468 3060
rect 30619 2841 30664 2881
rect 30806 2856 30951 2881
rect 31024 2880 31104 2881
rect 31300 2880 31468 2882
rect 31024 2864 31468 2880
rect 30808 2855 30951 2856
rect 31023 2854 31468 2864
rect 30619 2820 30666 2841
rect 31023 2820 31064 2854
rect 31300 2853 31468 2854
rect 31931 2858 31971 3082
rect 32097 3081 32265 3082
rect 32329 3114 32362 3447
rect 32329 3106 32366 3114
rect 32329 3087 32337 3106
rect 32358 3087 32366 3106
rect 32329 3081 32366 3087
rect 31931 2836 31939 2858
rect 31963 2836 31971 2858
rect 31931 2828 31971 2836
rect 29447 2782 29482 2783
rect 29424 2777 29482 2782
rect 29424 2757 29427 2777
rect 29447 2763 29482 2777
rect 29502 2763 29511 2783
rect 29447 2755 29511 2763
rect 29473 2754 29511 2755
rect 29474 2753 29511 2754
rect 29577 2787 29613 2788
rect 29685 2787 29721 2788
rect 29577 2779 29721 2787
rect 29577 2759 29585 2779
rect 29605 2775 29693 2779
rect 29605 2759 29649 2775
rect 29577 2755 29649 2759
rect 29669 2759 29693 2775
rect 29713 2759 29721 2779
rect 29669 2755 29721 2759
rect 29577 2753 29721 2755
rect 29787 2783 29825 2791
rect 29903 2787 29939 2788
rect 29787 2763 29796 2783
rect 29816 2763 29825 2783
rect 29787 2754 29825 2763
rect 29854 2779 29939 2787
rect 29854 2759 29911 2779
rect 29931 2759 29939 2779
rect 29787 2753 29824 2754
rect 29854 2753 29939 2759
rect 30005 2783 30043 2791
rect 30005 2763 30014 2783
rect 30034 2763 30043 2783
rect 30005 2754 30043 2763
rect 30187 2788 30230 2815
rect 30187 2770 30201 2788
rect 30219 2770 30230 2788
rect 30187 2762 30230 2770
rect 30192 2760 30230 2762
rect 30619 2790 31064 2820
rect 32102 2803 32167 2804
rect 30619 2787 31042 2790
rect 30005 2753 30042 2754
rect 29466 2725 29556 2731
rect 29466 2705 29482 2725
rect 29502 2723 29556 2725
rect 29502 2705 29527 2723
rect 29466 2703 29527 2705
rect 29547 2703 29556 2723
rect 29466 2697 29556 2703
rect 29479 2643 29516 2644
rect 29575 2643 29612 2644
rect 29631 2643 29667 2753
rect 29854 2732 29885 2753
rect 30619 2739 30666 2787
rect 29850 2731 29885 2732
rect 29728 2721 29885 2731
rect 29728 2701 29745 2721
rect 29765 2701 29885 2721
rect 29728 2694 29885 2701
rect 29952 2724 30101 2732
rect 29952 2704 29963 2724
rect 29983 2704 30022 2724
rect 30042 2704 30101 2724
rect 30619 2721 30629 2739
rect 30647 2721 30666 2739
rect 30619 2717 30666 2721
rect 31753 2778 31940 2802
rect 31971 2783 32364 2803
rect 32384 2783 32387 2803
rect 31971 2778 32387 2783
rect 30620 2712 30657 2717
rect 29952 2697 30101 2704
rect 31753 2707 31790 2778
rect 31971 2777 32312 2778
rect 31905 2717 31936 2718
rect 29952 2696 29993 2697
rect 30189 2695 30226 2698
rect 29686 2643 29723 2644
rect 29379 2634 29517 2643
rect 28583 2595 29027 2621
rect 28583 2593 28751 2595
rect 28583 2415 28610 2593
rect 28650 2555 28714 2567
rect 28990 2563 29027 2595
rect 29053 2594 29244 2616
rect 29379 2614 29488 2634
rect 29508 2614 29517 2634
rect 29379 2607 29517 2614
rect 29575 2634 29723 2643
rect 29575 2614 29584 2634
rect 29604 2614 29694 2634
rect 29714 2614 29723 2634
rect 29379 2605 29475 2607
rect 29575 2604 29723 2614
rect 29782 2634 29819 2644
rect 29782 2614 29790 2634
rect 29810 2614 29819 2634
rect 29631 2603 29667 2604
rect 29208 2592 29244 2594
rect 29208 2563 29245 2592
rect 28650 2554 28685 2555
rect 28627 2549 28685 2554
rect 28627 2529 28630 2549
rect 28650 2535 28685 2549
rect 28705 2535 28714 2555
rect 28650 2529 28714 2535
rect 28627 2527 28714 2529
rect 28627 2523 28654 2527
rect 28676 2526 28714 2527
rect 28677 2525 28714 2526
rect 28780 2559 28816 2560
rect 28888 2559 28924 2560
rect 28780 2552 28924 2559
rect 28780 2551 28842 2552
rect 28780 2531 28788 2551
rect 28808 2534 28842 2551
rect 28861 2551 28924 2552
rect 28861 2534 28896 2551
rect 28808 2531 28896 2534
rect 28916 2531 28924 2551
rect 28780 2525 28924 2531
rect 28990 2555 29028 2563
rect 29106 2559 29142 2560
rect 28990 2535 28999 2555
rect 29019 2535 29028 2555
rect 28990 2526 29028 2535
rect 29057 2551 29142 2559
rect 29057 2531 29114 2551
rect 29134 2531 29142 2551
rect 28990 2525 29027 2526
rect 29057 2525 29142 2531
rect 29208 2555 29246 2563
rect 29208 2535 29217 2555
rect 29237 2535 29246 2555
rect 29479 2544 29516 2545
rect 29782 2544 29819 2614
rect 29854 2643 29885 2694
rect 30181 2689 30226 2695
rect 30181 2671 30199 2689
rect 30217 2671 30226 2689
rect 31753 2687 31762 2707
rect 31782 2687 31790 2707
rect 31753 2677 31790 2687
rect 31849 2707 31936 2717
rect 31849 2687 31858 2707
rect 31878 2687 31936 2707
rect 31849 2678 31936 2687
rect 31849 2677 31886 2678
rect 30181 2661 30226 2671
rect 29904 2643 29941 2644
rect 29854 2634 29941 2643
rect 29854 2614 29912 2634
rect 29932 2614 29941 2634
rect 29854 2604 29941 2614
rect 30000 2634 30037 2644
rect 30000 2614 30008 2634
rect 30028 2614 30037 2634
rect 30181 2619 30224 2661
rect 30608 2650 30660 2652
rect 30087 2617 30224 2619
rect 29854 2603 29885 2604
rect 30000 2544 30037 2614
rect 29478 2543 29819 2544
rect 29208 2526 29246 2535
rect 29403 2538 29819 2543
rect 29208 2525 29245 2526
rect 28669 2497 28759 2503
rect 28669 2477 28685 2497
rect 28705 2495 28759 2497
rect 28705 2477 28730 2495
rect 28669 2475 28730 2477
rect 28750 2475 28759 2495
rect 28669 2469 28759 2475
rect 28682 2415 28719 2416
rect 28778 2415 28815 2416
rect 28834 2415 28870 2525
rect 29057 2504 29088 2525
rect 29403 2518 29406 2538
rect 29426 2518 29819 2538
rect 30003 2528 30037 2544
rect 30081 2596 30224 2617
rect 30606 2646 31039 2650
rect 30606 2640 31045 2646
rect 30606 2622 30627 2640
rect 30645 2622 31045 2640
rect 31905 2627 31936 2678
rect 31971 2707 32008 2777
rect 32274 2776 32311 2777
rect 32123 2717 32159 2718
rect 31971 2687 31980 2707
rect 32000 2687 32008 2707
rect 31971 2677 32008 2687
rect 32067 2707 32215 2717
rect 32315 2714 32411 2716
rect 32067 2687 32076 2707
rect 32096 2687 32186 2707
rect 32206 2687 32215 2707
rect 32067 2678 32215 2687
rect 32273 2707 32411 2714
rect 32273 2687 32282 2707
rect 32302 2687 32411 2707
rect 32273 2678 32411 2687
rect 32067 2677 32104 2678
rect 31797 2624 31838 2625
rect 30606 2604 31045 2622
rect 29779 2509 29819 2518
rect 30081 2509 30108 2596
rect 30181 2570 30224 2596
rect 30181 2552 30194 2570
rect 30212 2552 30224 2570
rect 30181 2541 30224 2552
rect 29053 2503 29088 2504
rect 28931 2493 29088 2503
rect 28931 2473 28948 2493
rect 28968 2473 29088 2493
rect 28931 2466 29088 2473
rect 29155 2496 29301 2504
rect 29155 2476 29166 2496
rect 29186 2476 29225 2496
rect 29245 2476 29301 2496
rect 29779 2492 30108 2509
rect 29779 2491 29819 2492
rect 29155 2469 29301 2476
rect 30176 2480 30216 2483
rect 30176 2474 30219 2480
rect 29801 2471 30219 2474
rect 29155 2468 29196 2469
rect 28889 2415 28926 2416
rect 28582 2406 28720 2415
rect 28582 2386 28691 2406
rect 28711 2386 28720 2406
rect 28582 2379 28720 2386
rect 28778 2406 28926 2415
rect 28778 2386 28787 2406
rect 28807 2386 28897 2406
rect 28917 2386 28926 2406
rect 28582 2377 28678 2379
rect 28778 2376 28926 2386
rect 28985 2406 29022 2416
rect 28985 2386 28993 2406
rect 29013 2386 29022 2406
rect 28834 2375 28870 2376
rect 28682 2316 28719 2317
rect 28985 2316 29022 2386
rect 29057 2415 29088 2466
rect 29801 2453 30192 2471
rect 30210 2453 30219 2471
rect 29801 2451 30219 2453
rect 29801 2443 29828 2451
rect 30069 2448 30219 2451
rect 29381 2437 29549 2438
rect 29800 2437 29828 2443
rect 29381 2421 29828 2437
rect 30176 2443 30219 2448
rect 29107 2415 29144 2416
rect 29057 2406 29144 2415
rect 29057 2386 29115 2406
rect 29135 2386 29144 2406
rect 29057 2376 29144 2386
rect 29203 2406 29240 2416
rect 29203 2386 29211 2406
rect 29231 2386 29240 2406
rect 29057 2375 29088 2376
rect 28681 2315 29022 2316
rect 29203 2315 29240 2386
rect 28606 2310 29022 2315
rect 28606 2290 28609 2310
rect 28629 2290 29022 2310
rect 29053 2291 29240 2315
rect 29381 2411 29825 2421
rect 29381 2409 29549 2411
rect 28481 2211 28523 2256
rect 29381 2231 29408 2409
rect 29448 2371 29512 2383
rect 29788 2379 29825 2411
rect 29851 2410 30042 2432
rect 30006 2408 30042 2410
rect 30006 2379 30043 2408
rect 30176 2387 30216 2443
rect 29448 2370 29483 2371
rect 29425 2365 29483 2370
rect 29425 2345 29428 2365
rect 29448 2351 29483 2365
rect 29503 2351 29512 2371
rect 29448 2343 29512 2351
rect 29474 2342 29512 2343
rect 29475 2341 29512 2342
rect 29578 2375 29614 2376
rect 29686 2375 29722 2376
rect 29578 2367 29722 2375
rect 29578 2347 29586 2367
rect 29606 2347 29641 2367
rect 29661 2347 29694 2367
rect 29714 2347 29722 2367
rect 29578 2341 29722 2347
rect 29788 2371 29826 2379
rect 29904 2375 29940 2376
rect 29788 2351 29797 2371
rect 29817 2351 29826 2371
rect 29788 2342 29826 2351
rect 29855 2367 29940 2375
rect 29855 2347 29912 2367
rect 29932 2347 29940 2367
rect 29788 2341 29825 2342
rect 29855 2341 29940 2347
rect 30006 2371 30044 2379
rect 30006 2351 30015 2371
rect 30035 2351 30044 2371
rect 30176 2369 30188 2387
rect 30206 2369 30216 2387
rect 30608 2415 30660 2604
rect 31006 2579 31045 2604
rect 31689 2617 31838 2624
rect 31689 2597 31748 2617
rect 31768 2597 31807 2617
rect 31827 2597 31838 2617
rect 31689 2589 31838 2597
rect 31905 2620 32062 2627
rect 31905 2600 32025 2620
rect 32045 2600 32062 2620
rect 31905 2590 32062 2600
rect 31905 2589 31940 2590
rect 30790 2554 30977 2578
rect 31006 2559 31401 2579
rect 31421 2559 31424 2579
rect 31905 2568 31936 2589
rect 32123 2568 32159 2678
rect 32178 2677 32215 2678
rect 32274 2677 32311 2678
rect 32234 2618 32324 2624
rect 32234 2598 32243 2618
rect 32263 2616 32324 2618
rect 32263 2598 32288 2616
rect 32234 2596 32288 2598
rect 32308 2596 32324 2616
rect 32234 2590 32324 2596
rect 31748 2567 31785 2568
rect 31006 2554 31424 2559
rect 31747 2558 31785 2567
rect 30790 2483 30827 2554
rect 31006 2553 31349 2554
rect 31006 2550 31045 2553
rect 31311 2552 31348 2553
rect 30942 2493 30973 2494
rect 30790 2463 30799 2483
rect 30819 2463 30827 2483
rect 30790 2453 30827 2463
rect 30886 2483 30973 2493
rect 30886 2463 30895 2483
rect 30915 2463 30973 2483
rect 30886 2454 30973 2463
rect 30886 2453 30923 2454
rect 30608 2397 30624 2415
rect 30642 2397 30660 2415
rect 30942 2403 30973 2454
rect 31008 2483 31045 2550
rect 31747 2538 31756 2558
rect 31776 2538 31785 2558
rect 31747 2530 31785 2538
rect 31851 2562 31936 2568
rect 31966 2567 32003 2568
rect 31851 2542 31859 2562
rect 31879 2542 31936 2562
rect 31851 2534 31936 2542
rect 31965 2558 32003 2567
rect 31965 2538 31974 2558
rect 31994 2538 32003 2558
rect 31851 2533 31887 2534
rect 31965 2530 32003 2538
rect 32069 2566 32213 2568
rect 32069 2562 32129 2566
rect 32069 2542 32077 2562
rect 32097 2544 32129 2562
rect 32152 2562 32213 2566
rect 32152 2544 32185 2562
rect 32097 2542 32185 2544
rect 32205 2542 32213 2562
rect 32069 2534 32213 2542
rect 32069 2533 32105 2534
rect 32177 2533 32213 2534
rect 32279 2567 32316 2568
rect 32279 2566 32317 2567
rect 32279 2558 32343 2566
rect 32279 2538 32288 2558
rect 32308 2544 32343 2558
rect 32363 2544 32366 2564
rect 32308 2539 32366 2544
rect 32308 2538 32343 2539
rect 31748 2501 31785 2530
rect 31749 2499 31785 2501
rect 31160 2493 31196 2494
rect 31008 2463 31017 2483
rect 31037 2463 31045 2483
rect 31008 2453 31045 2463
rect 31104 2483 31252 2493
rect 31352 2490 31448 2492
rect 31104 2463 31113 2483
rect 31133 2463 31223 2483
rect 31243 2463 31252 2483
rect 31104 2454 31252 2463
rect 31310 2483 31448 2490
rect 31310 2463 31319 2483
rect 31339 2463 31448 2483
rect 31749 2477 31940 2499
rect 31966 2498 32003 2530
rect 32279 2526 32343 2538
rect 31966 2497 32241 2498
rect 32383 2497 32410 2678
rect 31966 2472 32410 2497
rect 32546 2503 32585 4318
rect 32887 4305 32920 4638
rect 32984 4670 33152 4671
rect 33278 4670 33318 4894
rect 33781 4898 33949 4899
rect 34190 4898 34225 4915
rect 34582 4905 34629 4916
rect 33781 4872 34225 4898
rect 33781 4870 33949 4872
rect 34145 4871 34225 4872
rect 34380 4871 34447 4897
rect 34586 4871 34629 4905
rect 33781 4692 33808 4870
rect 33848 4832 33912 4844
rect 34188 4840 34225 4871
rect 34406 4840 34443 4871
rect 34588 4846 34629 4871
rect 33848 4831 33883 4832
rect 33825 4826 33883 4831
rect 33825 4806 33828 4826
rect 33848 4812 33883 4826
rect 33903 4812 33912 4832
rect 33848 4804 33912 4812
rect 33874 4803 33912 4804
rect 33875 4802 33912 4803
rect 33978 4836 34014 4837
rect 34086 4836 34122 4837
rect 33978 4828 34122 4836
rect 33978 4808 33986 4828
rect 34006 4824 34094 4828
rect 34006 4808 34050 4824
rect 33978 4804 34050 4808
rect 34070 4808 34094 4824
rect 34114 4808 34122 4828
rect 34070 4804 34122 4808
rect 33978 4802 34122 4804
rect 34188 4832 34226 4840
rect 34304 4836 34340 4837
rect 34188 4812 34197 4832
rect 34217 4812 34226 4832
rect 34188 4803 34226 4812
rect 34255 4828 34340 4836
rect 34255 4808 34312 4828
rect 34332 4808 34340 4828
rect 34188 4802 34225 4803
rect 34255 4802 34340 4808
rect 34406 4832 34444 4840
rect 34406 4812 34415 4832
rect 34435 4812 34444 4832
rect 34406 4803 34444 4812
rect 34588 4837 34630 4846
rect 34588 4819 34602 4837
rect 34620 4819 34630 4837
rect 34588 4811 34630 4819
rect 34593 4809 34630 4811
rect 34406 4802 34443 4803
rect 33867 4774 33957 4780
rect 33867 4754 33883 4774
rect 33903 4772 33957 4774
rect 33903 4754 33928 4772
rect 33867 4752 33928 4754
rect 33948 4752 33957 4772
rect 33867 4746 33957 4752
rect 33880 4692 33917 4693
rect 33976 4692 34013 4693
rect 34032 4692 34068 4802
rect 34255 4781 34286 4802
rect 34251 4780 34286 4781
rect 34129 4770 34286 4780
rect 34129 4750 34146 4770
rect 34166 4750 34286 4770
rect 34129 4743 34286 4750
rect 34353 4773 34502 4781
rect 34353 4753 34364 4773
rect 34384 4753 34423 4773
rect 34443 4753 34502 4773
rect 34353 4746 34502 4753
rect 34353 4745 34394 4746
rect 34590 4744 34627 4747
rect 34087 4692 34124 4693
rect 33780 4683 33918 4692
rect 32984 4644 33428 4670
rect 32984 4642 33152 4644
rect 32984 4464 33011 4642
rect 33051 4604 33115 4616
rect 33391 4612 33428 4644
rect 33454 4643 33645 4665
rect 33780 4663 33889 4683
rect 33909 4663 33918 4683
rect 33780 4656 33918 4663
rect 33976 4683 34124 4692
rect 33976 4663 33985 4683
rect 34005 4663 34095 4683
rect 34115 4663 34124 4683
rect 33780 4654 33876 4656
rect 33976 4653 34124 4663
rect 34183 4683 34220 4693
rect 34183 4663 34191 4683
rect 34211 4663 34220 4683
rect 34032 4652 34068 4653
rect 33609 4641 33645 4643
rect 33609 4612 33646 4641
rect 33051 4603 33086 4604
rect 33028 4598 33086 4603
rect 33028 4578 33031 4598
rect 33051 4584 33086 4598
rect 33106 4584 33115 4604
rect 33051 4578 33115 4584
rect 33028 4576 33115 4578
rect 33028 4572 33055 4576
rect 33077 4575 33115 4576
rect 33078 4574 33115 4575
rect 33181 4608 33217 4609
rect 33289 4608 33325 4609
rect 33181 4601 33325 4608
rect 33181 4600 33243 4601
rect 33181 4580 33189 4600
rect 33209 4583 33243 4600
rect 33262 4600 33325 4601
rect 33262 4583 33297 4600
rect 33209 4580 33297 4583
rect 33317 4580 33325 4600
rect 33181 4574 33325 4580
rect 33391 4604 33429 4612
rect 33507 4608 33543 4609
rect 33391 4584 33400 4604
rect 33420 4584 33429 4604
rect 33391 4575 33429 4584
rect 33458 4600 33543 4608
rect 33458 4580 33515 4600
rect 33535 4580 33543 4600
rect 33391 4574 33428 4575
rect 33458 4574 33543 4580
rect 33609 4604 33647 4612
rect 33609 4584 33618 4604
rect 33638 4584 33647 4604
rect 33880 4593 33917 4594
rect 34183 4593 34220 4663
rect 34255 4692 34286 4743
rect 34582 4738 34627 4744
rect 34582 4720 34600 4738
rect 34618 4720 34627 4738
rect 34582 4710 34627 4720
rect 34305 4692 34342 4693
rect 34255 4683 34342 4692
rect 34255 4663 34313 4683
rect 34333 4663 34342 4683
rect 34255 4653 34342 4663
rect 34401 4683 34438 4693
rect 34401 4663 34409 4683
rect 34429 4663 34438 4683
rect 34582 4668 34625 4710
rect 34488 4666 34625 4668
rect 34255 4652 34286 4653
rect 34401 4593 34438 4663
rect 33879 4592 34220 4593
rect 33609 4575 33647 4584
rect 33804 4587 34220 4592
rect 33609 4574 33646 4575
rect 33070 4546 33160 4552
rect 33070 4526 33086 4546
rect 33106 4544 33160 4546
rect 33106 4526 33131 4544
rect 33070 4524 33131 4526
rect 33151 4524 33160 4544
rect 33070 4518 33160 4524
rect 33083 4464 33120 4465
rect 33179 4464 33216 4465
rect 33235 4464 33271 4574
rect 33458 4553 33489 4574
rect 33804 4567 33807 4587
rect 33827 4567 34220 4587
rect 34404 4577 34438 4593
rect 34482 4645 34625 4666
rect 34180 4558 34220 4567
rect 34482 4558 34509 4645
rect 34582 4619 34625 4645
rect 34582 4601 34595 4619
rect 34613 4601 34625 4619
rect 34582 4590 34625 4601
rect 33454 4552 33489 4553
rect 33332 4542 33489 4552
rect 33332 4522 33349 4542
rect 33369 4522 33489 4542
rect 33332 4515 33489 4522
rect 33556 4545 33702 4553
rect 33556 4525 33567 4545
rect 33587 4525 33626 4545
rect 33646 4525 33702 4545
rect 34180 4541 34509 4558
rect 34180 4540 34220 4541
rect 33556 4518 33702 4525
rect 34577 4529 34617 4532
rect 34577 4523 34620 4529
rect 34202 4520 34620 4523
rect 33556 4517 33597 4518
rect 33290 4464 33327 4465
rect 32983 4455 33121 4464
rect 32983 4435 33092 4455
rect 33112 4435 33121 4455
rect 32983 4428 33121 4435
rect 33179 4455 33327 4464
rect 33179 4435 33188 4455
rect 33208 4435 33298 4455
rect 33318 4435 33327 4455
rect 32983 4426 33079 4428
rect 33179 4425 33327 4435
rect 33386 4455 33423 4465
rect 33386 4435 33394 4455
rect 33414 4435 33423 4455
rect 33235 4424 33271 4425
rect 33083 4365 33120 4366
rect 33386 4365 33423 4435
rect 33458 4464 33489 4515
rect 34202 4502 34593 4520
rect 34611 4502 34620 4520
rect 34202 4500 34620 4502
rect 34202 4492 34229 4500
rect 34470 4497 34620 4500
rect 33782 4486 33950 4487
rect 34201 4486 34229 4492
rect 33782 4470 34229 4486
rect 34577 4492 34620 4497
rect 33508 4464 33545 4465
rect 33458 4455 33545 4464
rect 33458 4435 33516 4455
rect 33536 4435 33545 4455
rect 33458 4425 33545 4435
rect 33604 4455 33641 4465
rect 33604 4435 33612 4455
rect 33632 4435 33641 4455
rect 33458 4424 33489 4425
rect 33082 4364 33423 4365
rect 33604 4364 33641 4435
rect 33007 4359 33423 4364
rect 33007 4339 33010 4359
rect 33030 4339 33423 4359
rect 33454 4340 33641 4364
rect 33782 4460 34226 4470
rect 33782 4458 33950 4460
rect 32816 4265 32860 4266
rect 32816 4259 32861 4265
rect 32816 4241 32828 4259
rect 32850 4241 32861 4259
rect 32882 4260 32924 4305
rect 33782 4280 33809 4458
rect 33849 4420 33913 4432
rect 34189 4428 34226 4460
rect 34252 4459 34443 4481
rect 34407 4457 34443 4459
rect 34407 4428 34444 4457
rect 34577 4436 34617 4492
rect 33849 4419 33884 4420
rect 33826 4414 33884 4419
rect 33826 4394 33829 4414
rect 33849 4400 33884 4414
rect 33904 4400 33913 4420
rect 33849 4392 33913 4400
rect 33875 4391 33913 4392
rect 33876 4390 33913 4391
rect 33979 4424 34015 4425
rect 34087 4424 34123 4425
rect 33979 4416 34123 4424
rect 33979 4396 33987 4416
rect 34007 4396 34042 4416
rect 34062 4396 34095 4416
rect 34115 4396 34123 4416
rect 33979 4390 34123 4396
rect 34189 4420 34227 4428
rect 34305 4424 34341 4425
rect 34189 4400 34198 4420
rect 34218 4400 34227 4420
rect 34189 4391 34227 4400
rect 34256 4416 34341 4424
rect 34256 4396 34313 4416
rect 34333 4396 34341 4416
rect 34189 4390 34226 4391
rect 34256 4390 34341 4396
rect 34407 4420 34445 4428
rect 34407 4400 34416 4420
rect 34436 4400 34445 4420
rect 34577 4418 34589 4436
rect 34607 4418 34617 4436
rect 34577 4408 34617 4418
rect 34407 4391 34445 4400
rect 34407 4390 34444 4391
rect 33868 4362 33958 4368
rect 33868 4342 33884 4362
rect 33904 4360 33958 4362
rect 33904 4342 33929 4360
rect 33868 4340 33929 4342
rect 33949 4340 33958 4360
rect 33868 4334 33958 4340
rect 33881 4280 33918 4281
rect 33977 4280 34014 4281
rect 34033 4280 34069 4390
rect 34256 4369 34287 4390
rect 34252 4368 34287 4369
rect 34130 4358 34287 4368
rect 34130 4338 34147 4358
rect 34167 4338 34287 4358
rect 34130 4331 34287 4338
rect 34354 4361 34503 4369
rect 34354 4341 34365 4361
rect 34385 4341 34424 4361
rect 34444 4341 34503 4361
rect 34354 4334 34503 4341
rect 34569 4337 34621 4355
rect 34354 4333 34395 4334
rect 34088 4280 34125 4281
rect 33781 4271 33919 4280
rect 33253 4260 33286 4262
rect 32882 4248 33329 4260
rect 32816 4211 32861 4241
rect 32833 3265 32861 4211
rect 32885 4234 33329 4248
rect 32885 4232 33053 4234
rect 32885 4054 32912 4232
rect 32952 4194 33016 4206
rect 33292 4202 33329 4234
rect 33355 4233 33546 4255
rect 33781 4251 33890 4271
rect 33910 4251 33919 4271
rect 33781 4244 33919 4251
rect 33977 4271 34125 4280
rect 33977 4251 33986 4271
rect 34006 4251 34096 4271
rect 34116 4251 34125 4271
rect 33781 4242 33877 4244
rect 33977 4241 34125 4251
rect 34184 4271 34221 4281
rect 34184 4251 34192 4271
rect 34212 4251 34221 4271
rect 34033 4240 34069 4241
rect 33510 4231 33546 4233
rect 33510 4202 33547 4231
rect 32952 4193 32987 4194
rect 32929 4188 32987 4193
rect 32929 4168 32932 4188
rect 32952 4174 32987 4188
rect 33007 4174 33016 4194
rect 32952 4166 33016 4174
rect 32978 4165 33016 4166
rect 32979 4164 33016 4165
rect 33082 4198 33118 4199
rect 33190 4198 33226 4199
rect 33082 4192 33226 4198
rect 33082 4190 33143 4192
rect 33082 4170 33090 4190
rect 33110 4175 33143 4190
rect 33162 4190 33226 4192
rect 33162 4175 33198 4190
rect 33110 4170 33198 4175
rect 33218 4170 33226 4190
rect 33082 4164 33226 4170
rect 33292 4194 33330 4202
rect 33408 4198 33444 4199
rect 33292 4174 33301 4194
rect 33321 4174 33330 4194
rect 33292 4165 33330 4174
rect 33359 4190 33444 4198
rect 33359 4170 33416 4190
rect 33436 4170 33444 4190
rect 33292 4164 33329 4165
rect 33359 4164 33444 4170
rect 33510 4194 33548 4202
rect 33510 4174 33519 4194
rect 33539 4174 33548 4194
rect 34184 4184 34221 4251
rect 34256 4280 34287 4331
rect 34569 4319 34587 4337
rect 34605 4319 34621 4337
rect 34306 4280 34343 4281
rect 34256 4271 34343 4280
rect 34256 4251 34314 4271
rect 34334 4251 34343 4271
rect 34256 4241 34343 4251
rect 34402 4271 34439 4281
rect 34402 4251 34410 4271
rect 34430 4251 34439 4271
rect 34256 4240 34287 4241
rect 33881 4181 33918 4182
rect 34184 4181 34223 4184
rect 33880 4180 34223 4181
rect 34402 4180 34439 4251
rect 33510 4165 33548 4174
rect 33805 4175 34223 4180
rect 33510 4164 33547 4165
rect 32971 4136 33061 4142
rect 32971 4116 32987 4136
rect 33007 4134 33061 4136
rect 33007 4116 33032 4134
rect 32971 4114 33032 4116
rect 33052 4114 33061 4134
rect 32971 4108 33061 4114
rect 32984 4054 33021 4055
rect 33080 4054 33117 4055
rect 33136 4054 33172 4164
rect 33359 4143 33390 4164
rect 33805 4155 33808 4175
rect 33828 4155 34223 4175
rect 34252 4156 34439 4180
rect 33355 4142 33390 4143
rect 33233 4132 33390 4142
rect 33233 4112 33250 4132
rect 33270 4112 33390 4132
rect 33233 4105 33390 4112
rect 33457 4135 33606 4143
rect 33457 4115 33468 4135
rect 33488 4115 33527 4135
rect 33547 4115 33606 4135
rect 33457 4108 33606 4115
rect 34184 4130 34223 4155
rect 34569 4130 34621 4319
rect 34184 4112 34623 4130
rect 33457 4107 33498 4108
rect 33191 4054 33228 4055
rect 32884 4045 33022 4054
rect 32884 4025 32993 4045
rect 33013 4025 33022 4045
rect 32884 4018 33022 4025
rect 33080 4045 33228 4054
rect 33080 4025 33089 4045
rect 33109 4025 33199 4045
rect 33219 4025 33228 4045
rect 32884 4016 32980 4018
rect 33080 4015 33228 4025
rect 33287 4045 33324 4055
rect 33287 4025 33295 4045
rect 33315 4025 33324 4045
rect 33136 4014 33172 4015
rect 32984 3955 33021 3956
rect 33287 3955 33324 4025
rect 33359 4054 33390 4105
rect 34184 4094 34584 4112
rect 34602 4094 34623 4112
rect 34184 4088 34623 4094
rect 34190 4084 34623 4088
rect 34569 4082 34621 4084
rect 33409 4054 33446 4055
rect 33359 4045 33446 4054
rect 33359 4025 33417 4045
rect 33437 4025 33446 4045
rect 33359 4015 33446 4025
rect 33505 4045 33542 4055
rect 33505 4025 33513 4045
rect 33533 4025 33542 4045
rect 33359 4014 33390 4015
rect 32983 3954 33324 3955
rect 33505 3954 33542 4025
rect 34572 4017 34609 4022
rect 34563 4013 34610 4017
rect 34563 3995 34582 4013
rect 34600 3995 34610 4013
rect 32908 3949 33324 3954
rect 32908 3929 32911 3949
rect 32931 3929 33324 3949
rect 33355 3930 33542 3954
rect 34167 3952 34207 3957
rect 34563 3952 34610 3995
rect 34167 3913 34610 3952
rect 33261 3898 33301 3906
rect 33261 3876 33269 3898
rect 33293 3876 33301 3898
rect 32967 3652 33135 3653
rect 33261 3652 33301 3876
rect 33764 3880 33932 3881
rect 34167 3880 34207 3913
rect 34563 3880 34610 3913
rect 33764 3879 34208 3880
rect 33764 3854 34209 3879
rect 33764 3852 33932 3854
rect 34128 3853 34209 3854
rect 34378 3853 34427 3879
rect 34563 3853 34612 3880
rect 33764 3674 33791 3852
rect 33831 3814 33895 3826
rect 34171 3822 34208 3853
rect 34389 3822 34426 3853
rect 34571 3828 34612 3853
rect 33831 3813 33866 3814
rect 33808 3808 33866 3813
rect 33808 3788 33811 3808
rect 33831 3794 33866 3808
rect 33886 3794 33895 3814
rect 33831 3786 33895 3794
rect 33857 3785 33895 3786
rect 33858 3784 33895 3785
rect 33961 3818 33997 3819
rect 34069 3818 34105 3819
rect 33961 3810 34105 3818
rect 33961 3790 33969 3810
rect 33989 3806 34077 3810
rect 33989 3790 34033 3806
rect 33961 3786 34033 3790
rect 34053 3790 34077 3806
rect 34097 3790 34105 3810
rect 34053 3786 34105 3790
rect 33961 3784 34105 3786
rect 34171 3814 34209 3822
rect 34287 3818 34323 3819
rect 34171 3794 34180 3814
rect 34200 3794 34209 3814
rect 34171 3785 34209 3794
rect 34238 3810 34323 3818
rect 34238 3790 34295 3810
rect 34315 3790 34323 3810
rect 34171 3784 34208 3785
rect 34238 3784 34323 3790
rect 34389 3814 34427 3822
rect 34389 3794 34398 3814
rect 34418 3794 34427 3814
rect 34389 3785 34427 3794
rect 34571 3819 34613 3828
rect 34571 3801 34585 3819
rect 34603 3801 34613 3819
rect 34571 3793 34613 3801
rect 34576 3791 34613 3793
rect 34389 3784 34426 3785
rect 33850 3756 33940 3762
rect 33850 3736 33866 3756
rect 33886 3754 33940 3756
rect 33886 3736 33911 3754
rect 33850 3734 33911 3736
rect 33931 3734 33940 3754
rect 33850 3728 33940 3734
rect 33863 3674 33900 3675
rect 33959 3674 33996 3675
rect 34015 3674 34051 3784
rect 34238 3763 34269 3784
rect 34234 3762 34269 3763
rect 34112 3752 34269 3762
rect 34112 3732 34129 3752
rect 34149 3732 34269 3752
rect 34112 3725 34269 3732
rect 34336 3755 34485 3763
rect 34336 3735 34347 3755
rect 34367 3735 34406 3755
rect 34426 3735 34485 3755
rect 34336 3728 34485 3735
rect 34336 3727 34377 3728
rect 34573 3726 34610 3729
rect 34070 3674 34107 3675
rect 33763 3665 33901 3674
rect 32967 3626 33411 3652
rect 32967 3624 33135 3626
rect 32967 3446 32994 3624
rect 33034 3586 33098 3598
rect 33374 3594 33411 3626
rect 33437 3625 33628 3647
rect 33763 3645 33872 3665
rect 33892 3645 33901 3665
rect 33763 3638 33901 3645
rect 33959 3665 34107 3674
rect 33959 3645 33968 3665
rect 33988 3645 34078 3665
rect 34098 3645 34107 3665
rect 33763 3636 33859 3638
rect 33959 3635 34107 3645
rect 34166 3665 34203 3675
rect 34166 3645 34174 3665
rect 34194 3645 34203 3665
rect 34015 3634 34051 3635
rect 33592 3623 33628 3625
rect 33592 3594 33629 3623
rect 33034 3585 33069 3586
rect 33011 3580 33069 3585
rect 33011 3560 33014 3580
rect 33034 3566 33069 3580
rect 33089 3566 33098 3586
rect 33034 3558 33098 3566
rect 33060 3557 33098 3558
rect 33061 3556 33098 3557
rect 33164 3590 33200 3591
rect 33272 3590 33308 3591
rect 33164 3582 33308 3590
rect 33164 3562 33172 3582
rect 33192 3581 33280 3582
rect 33192 3562 33227 3581
rect 33248 3562 33280 3581
rect 33300 3562 33308 3582
rect 33164 3556 33308 3562
rect 33374 3586 33412 3594
rect 33490 3590 33526 3591
rect 33374 3566 33383 3586
rect 33403 3566 33412 3586
rect 33374 3557 33412 3566
rect 33441 3582 33526 3590
rect 33441 3562 33498 3582
rect 33518 3562 33526 3582
rect 33374 3556 33411 3557
rect 33441 3556 33526 3562
rect 33592 3586 33630 3594
rect 33592 3566 33601 3586
rect 33621 3566 33630 3586
rect 33863 3575 33900 3576
rect 34166 3575 34203 3645
rect 34238 3674 34269 3725
rect 34565 3720 34610 3726
rect 34565 3702 34583 3720
rect 34601 3702 34610 3720
rect 34565 3692 34610 3702
rect 34288 3674 34325 3675
rect 34238 3665 34325 3674
rect 34238 3645 34296 3665
rect 34316 3645 34325 3665
rect 34238 3635 34325 3645
rect 34384 3665 34421 3675
rect 34384 3645 34392 3665
rect 34412 3645 34421 3665
rect 34565 3650 34608 3692
rect 34471 3648 34608 3650
rect 34238 3634 34269 3635
rect 34384 3575 34421 3645
rect 33862 3574 34203 3575
rect 33592 3557 33630 3566
rect 33787 3569 34203 3574
rect 33592 3556 33629 3557
rect 33053 3528 33143 3534
rect 33053 3508 33069 3528
rect 33089 3526 33143 3528
rect 33089 3508 33114 3526
rect 33053 3506 33114 3508
rect 33134 3506 33143 3526
rect 33053 3500 33143 3506
rect 33066 3446 33103 3447
rect 33162 3446 33199 3447
rect 33218 3446 33254 3556
rect 33441 3535 33472 3556
rect 33787 3549 33790 3569
rect 33810 3549 34203 3569
rect 34387 3559 34421 3575
rect 34465 3627 34608 3648
rect 34163 3540 34203 3549
rect 34465 3540 34492 3627
rect 34565 3601 34608 3627
rect 34565 3583 34578 3601
rect 34596 3583 34608 3601
rect 34565 3572 34608 3583
rect 33437 3534 33472 3535
rect 33315 3524 33472 3534
rect 33315 3504 33332 3524
rect 33352 3504 33472 3524
rect 33315 3497 33472 3504
rect 33539 3527 33688 3535
rect 33539 3507 33550 3527
rect 33570 3507 33609 3527
rect 33629 3507 33688 3527
rect 34163 3523 34492 3540
rect 34163 3522 34203 3523
rect 33539 3500 33688 3507
rect 34560 3511 34600 3514
rect 34560 3505 34603 3511
rect 34185 3502 34603 3505
rect 33539 3499 33580 3500
rect 33273 3446 33310 3447
rect 32966 3437 33104 3446
rect 32966 3417 33075 3437
rect 33095 3417 33104 3437
rect 32966 3410 33104 3417
rect 33162 3437 33310 3446
rect 33162 3417 33171 3437
rect 33191 3417 33281 3437
rect 33301 3417 33310 3437
rect 32966 3408 33062 3410
rect 33162 3407 33310 3417
rect 33369 3437 33406 3447
rect 33369 3417 33377 3437
rect 33397 3417 33406 3437
rect 33218 3406 33254 3407
rect 33066 3347 33103 3348
rect 33369 3347 33406 3417
rect 33441 3446 33472 3497
rect 34185 3484 34576 3502
rect 34594 3484 34603 3502
rect 34185 3482 34603 3484
rect 34185 3474 34212 3482
rect 34453 3479 34603 3482
rect 33765 3468 33933 3469
rect 34184 3468 34212 3474
rect 33765 3452 34212 3468
rect 34560 3474 34603 3479
rect 33491 3446 33528 3447
rect 33441 3437 33528 3446
rect 33441 3417 33499 3437
rect 33519 3417 33528 3437
rect 33441 3407 33528 3417
rect 33587 3437 33624 3447
rect 33587 3417 33595 3437
rect 33615 3417 33624 3437
rect 33441 3406 33472 3407
rect 33065 3346 33406 3347
rect 33587 3346 33624 3417
rect 32990 3341 33406 3346
rect 32990 3321 32993 3341
rect 33013 3321 33406 3341
rect 33437 3322 33624 3346
rect 33765 3442 34209 3452
rect 33765 3440 33933 3442
rect 32832 3247 32861 3265
rect 33765 3262 33792 3440
rect 33832 3402 33896 3414
rect 34172 3410 34209 3442
rect 34235 3441 34426 3463
rect 34390 3439 34426 3441
rect 34390 3410 34427 3439
rect 34560 3418 34600 3474
rect 33832 3401 33867 3402
rect 33809 3396 33867 3401
rect 33809 3376 33812 3396
rect 33832 3382 33867 3396
rect 33887 3382 33896 3402
rect 33832 3374 33896 3382
rect 33858 3373 33896 3374
rect 33859 3372 33896 3373
rect 33962 3406 33998 3407
rect 34070 3406 34106 3407
rect 33962 3398 34106 3406
rect 33962 3378 33970 3398
rect 33990 3378 34025 3398
rect 34045 3378 34078 3398
rect 34098 3378 34106 3398
rect 33962 3372 34106 3378
rect 34172 3402 34210 3410
rect 34288 3406 34324 3407
rect 34172 3382 34181 3402
rect 34201 3382 34210 3402
rect 34172 3373 34210 3382
rect 34239 3398 34324 3406
rect 34239 3378 34296 3398
rect 34316 3378 34324 3398
rect 34172 3372 34209 3373
rect 34239 3372 34324 3378
rect 34390 3402 34428 3410
rect 34390 3382 34399 3402
rect 34419 3382 34428 3402
rect 34560 3400 34572 3418
rect 34590 3400 34600 3418
rect 34560 3390 34600 3400
rect 34390 3373 34428 3382
rect 34390 3372 34427 3373
rect 33851 3344 33941 3350
rect 33851 3324 33867 3344
rect 33887 3342 33941 3344
rect 33887 3324 33912 3342
rect 33851 3322 33912 3324
rect 33932 3322 33941 3342
rect 33851 3316 33941 3322
rect 33864 3262 33901 3263
rect 33960 3262 33997 3263
rect 34016 3262 34052 3372
rect 34239 3351 34270 3372
rect 34235 3350 34270 3351
rect 34113 3340 34270 3350
rect 34113 3320 34130 3340
rect 34150 3320 34270 3340
rect 34113 3313 34270 3320
rect 34337 3343 34486 3351
rect 34337 3323 34348 3343
rect 34368 3323 34407 3343
rect 34427 3323 34486 3343
rect 34337 3316 34486 3323
rect 34552 3319 34604 3337
rect 34337 3315 34378 3316
rect 34071 3262 34108 3263
rect 32802 3245 32861 3247
rect 33764 3253 33902 3262
rect 32802 3244 32970 3245
rect 33096 3244 33136 3246
rect 32802 3218 33246 3244
rect 32802 3216 32970 3218
rect 32802 3214 32883 3216
rect 32802 3038 32829 3214
rect 32869 3178 32933 3190
rect 33209 3186 33246 3218
rect 33272 3217 33463 3239
rect 33764 3233 33873 3253
rect 33893 3233 33902 3253
rect 33764 3226 33902 3233
rect 33960 3253 34108 3262
rect 33960 3233 33969 3253
rect 33989 3233 34079 3253
rect 34099 3233 34108 3253
rect 33764 3224 33860 3226
rect 33960 3223 34108 3233
rect 34167 3253 34204 3263
rect 34167 3233 34175 3253
rect 34195 3233 34204 3253
rect 34016 3222 34052 3223
rect 33427 3215 33463 3217
rect 33427 3186 33464 3215
rect 32869 3177 32904 3178
rect 32846 3172 32904 3177
rect 32846 3152 32849 3172
rect 32869 3158 32904 3172
rect 32924 3158 32933 3178
rect 32869 3150 32933 3158
rect 32895 3149 32933 3150
rect 32896 3148 32933 3149
rect 32999 3182 33035 3183
rect 33107 3182 33143 3183
rect 32999 3174 33143 3182
rect 32999 3154 33007 3174
rect 33027 3173 33115 3174
rect 33027 3155 33062 3173
rect 33080 3155 33115 3173
rect 33027 3154 33115 3155
rect 33135 3154 33143 3174
rect 32999 3148 33143 3154
rect 33209 3178 33247 3186
rect 33325 3182 33361 3183
rect 33209 3158 33218 3178
rect 33238 3158 33247 3178
rect 33209 3149 33247 3158
rect 33276 3174 33361 3182
rect 33276 3154 33333 3174
rect 33353 3154 33361 3174
rect 33209 3148 33246 3149
rect 33276 3148 33361 3154
rect 33427 3178 33465 3186
rect 33427 3158 33436 3178
rect 33456 3158 33465 3178
rect 34167 3166 34204 3233
rect 34239 3262 34270 3313
rect 34552 3301 34570 3319
rect 34588 3301 34604 3319
rect 34289 3262 34326 3263
rect 34239 3253 34326 3262
rect 34239 3233 34297 3253
rect 34317 3233 34326 3253
rect 34239 3223 34326 3233
rect 34385 3253 34422 3263
rect 34385 3233 34393 3253
rect 34413 3233 34422 3253
rect 34239 3222 34270 3223
rect 33864 3163 33901 3164
rect 34167 3163 34206 3166
rect 33863 3162 34206 3163
rect 34385 3162 34422 3233
rect 33427 3149 33465 3158
rect 33788 3157 34206 3162
rect 33427 3148 33464 3149
rect 32888 3120 32978 3126
rect 32888 3100 32904 3120
rect 32924 3118 32978 3120
rect 32924 3100 32949 3118
rect 32888 3098 32949 3100
rect 32969 3098 32978 3118
rect 32888 3092 32978 3098
rect 32901 3038 32938 3039
rect 32997 3038 33034 3039
rect 33053 3038 33089 3148
rect 33276 3127 33307 3148
rect 33788 3137 33791 3157
rect 33811 3137 34206 3157
rect 34235 3138 34422 3162
rect 33272 3126 33307 3127
rect 33150 3116 33307 3126
rect 33150 3096 33167 3116
rect 33187 3096 33307 3116
rect 33150 3089 33307 3096
rect 33374 3119 33523 3127
rect 33374 3099 33385 3119
rect 33405 3099 33444 3119
rect 33464 3099 33523 3119
rect 33374 3092 33523 3099
rect 34167 3112 34206 3137
rect 34552 3112 34604 3301
rect 34167 3094 34606 3112
rect 33374 3091 33415 3092
rect 33108 3038 33145 3039
rect 32801 3029 32939 3038
rect 32801 3009 32910 3029
rect 32930 3009 32939 3029
rect 32801 3002 32939 3009
rect 32997 3029 33145 3038
rect 32997 3009 33006 3029
rect 33026 3009 33116 3029
rect 33136 3009 33145 3029
rect 32801 3000 32897 3002
rect 32997 2999 33145 3009
rect 33204 3029 33241 3039
rect 33204 3009 33212 3029
rect 33232 3009 33241 3029
rect 33053 2998 33089 2999
rect 32901 2939 32938 2940
rect 33204 2939 33241 3009
rect 33276 3038 33307 3089
rect 34167 3076 34567 3094
rect 34585 3076 34606 3094
rect 34167 3070 34606 3076
rect 34173 3066 34606 3070
rect 34552 3064 34604 3066
rect 33326 3038 33363 3039
rect 33276 3029 33363 3038
rect 33276 3009 33334 3029
rect 33354 3009 33363 3029
rect 33276 2999 33363 3009
rect 33422 3029 33459 3039
rect 33422 3009 33430 3029
rect 33450 3009 33459 3029
rect 33276 2998 33307 2999
rect 32900 2938 33241 2939
rect 33422 2938 33459 3009
rect 34555 2999 34592 3004
rect 32825 2933 33241 2938
rect 32825 2913 32828 2933
rect 32848 2913 33241 2933
rect 33272 2914 33459 2938
rect 34546 2995 34593 2999
rect 34546 2977 34565 2995
rect 34583 2977 34593 2995
rect 34546 2929 34593 2977
rect 34170 2926 34593 2929
rect 33045 2912 33110 2913
rect 34148 2896 34593 2926
rect 33241 2880 33281 2888
rect 33241 2858 33249 2880
rect 33273 2858 33281 2880
rect 32846 2629 32883 2635
rect 32846 2610 32854 2629
rect 32875 2610 32883 2629
rect 32846 2602 32883 2610
rect 32546 2481 32553 2503
rect 32577 2481 32585 2503
rect 32546 2475 32585 2481
rect 32076 2470 32116 2472
rect 32242 2471 32410 2472
rect 32344 2470 32381 2471
rect 31310 2454 31448 2463
rect 31104 2453 31141 2454
rect 30834 2400 30875 2401
rect 30608 2379 30660 2397
rect 30726 2393 30875 2400
rect 30176 2359 30216 2369
rect 30726 2373 30785 2393
rect 30805 2373 30844 2393
rect 30864 2373 30875 2393
rect 30726 2365 30875 2373
rect 30942 2396 31099 2403
rect 30942 2376 31062 2396
rect 31082 2376 31099 2396
rect 30942 2366 31099 2376
rect 30942 2365 30977 2366
rect 30006 2342 30044 2351
rect 30942 2344 30973 2365
rect 31160 2344 31196 2454
rect 31215 2453 31252 2454
rect 31311 2453 31348 2454
rect 31271 2394 31361 2400
rect 31271 2374 31280 2394
rect 31300 2392 31361 2394
rect 31300 2374 31325 2392
rect 31271 2372 31325 2374
rect 31345 2372 31361 2392
rect 31271 2366 31361 2372
rect 30785 2343 30822 2344
rect 30006 2341 30043 2342
rect 29467 2313 29557 2319
rect 29467 2293 29483 2313
rect 29503 2311 29557 2313
rect 29503 2293 29528 2311
rect 29467 2291 29528 2293
rect 29548 2291 29557 2311
rect 29467 2285 29557 2291
rect 29480 2231 29517 2232
rect 29576 2231 29613 2232
rect 29632 2231 29668 2341
rect 29855 2320 29886 2341
rect 30784 2334 30822 2343
rect 29851 2319 29886 2320
rect 29729 2309 29886 2319
rect 29729 2289 29746 2309
rect 29766 2289 29886 2309
rect 29729 2282 29886 2289
rect 29953 2312 30102 2320
rect 29953 2292 29964 2312
rect 29984 2292 30023 2312
rect 30043 2292 30102 2312
rect 30612 2316 30652 2326
rect 29953 2285 30102 2292
rect 30168 2288 30220 2306
rect 29953 2284 29994 2285
rect 29687 2231 29724 2232
rect 29380 2222 29518 2231
rect 28852 2211 28885 2213
rect 28481 2199 28928 2211
rect 27713 2077 27881 2079
rect 27437 2051 27881 2077
rect 26947 2029 27085 2038
rect 26741 2028 26778 2029
rect 26238 1974 26275 1977
rect 26471 1975 26512 1976
rect 24581 1953 24612 1954
rect 24205 1893 24546 1894
rect 24727 1893 24764 1964
rect 26363 1968 26512 1975
rect 25794 1956 25831 1961
rect 25785 1952 25832 1956
rect 25785 1934 25804 1952
rect 25822 1934 25832 1952
rect 26363 1948 26422 1968
rect 26442 1948 26481 1968
rect 26501 1948 26512 1968
rect 26363 1940 26512 1948
rect 26579 1971 26736 1978
rect 26579 1951 26699 1971
rect 26719 1951 26736 1971
rect 26579 1941 26736 1951
rect 26579 1940 26614 1941
rect 24130 1888 24546 1893
rect 24130 1868 24133 1888
rect 24153 1868 24546 1888
rect 24577 1869 24764 1893
rect 25389 1891 25429 1896
rect 25785 1891 25832 1934
rect 26579 1919 26610 1940
rect 26797 1919 26833 2029
rect 26852 2028 26889 2029
rect 26948 2028 26985 2029
rect 26908 1969 26998 1975
rect 26908 1949 26917 1969
rect 26937 1967 26998 1969
rect 26937 1949 26962 1967
rect 26908 1947 26962 1949
rect 26982 1947 26998 1967
rect 26908 1941 26998 1947
rect 26422 1918 26459 1919
rect 25389 1852 25832 1891
rect 26235 1910 26272 1912
rect 26235 1902 26277 1910
rect 26235 1884 26245 1902
rect 26263 1884 26277 1902
rect 26235 1875 26277 1884
rect 26421 1909 26459 1918
rect 26421 1889 26430 1909
rect 26450 1889 26459 1909
rect 26421 1881 26459 1889
rect 26525 1913 26610 1919
rect 26640 1918 26677 1919
rect 26525 1893 26533 1913
rect 26553 1893 26610 1913
rect 26525 1885 26610 1893
rect 26639 1909 26677 1918
rect 26639 1889 26648 1909
rect 26668 1889 26677 1909
rect 26525 1884 26561 1885
rect 26639 1881 26677 1889
rect 26743 1917 26887 1919
rect 26743 1913 26795 1917
rect 26743 1893 26751 1913
rect 26771 1897 26795 1913
rect 26815 1913 26887 1917
rect 26815 1897 26859 1913
rect 26771 1893 26859 1897
rect 26879 1893 26887 1913
rect 26743 1885 26887 1893
rect 26743 1884 26779 1885
rect 26851 1884 26887 1885
rect 26953 1918 26990 1919
rect 26953 1917 26991 1918
rect 26953 1909 27017 1917
rect 26953 1889 26962 1909
rect 26982 1895 27017 1909
rect 27037 1895 27040 1915
rect 26982 1890 27040 1895
rect 26982 1889 27017 1890
rect 23170 1793 23178 1815
rect 23202 1793 23210 1815
rect 23170 1785 23210 1793
rect 24483 1837 24523 1845
rect 24483 1815 24491 1837
rect 24515 1815 24523 1837
rect 20689 1739 20724 1740
rect 20666 1734 20724 1739
rect 20666 1714 20669 1734
rect 20689 1720 20724 1734
rect 20744 1720 20753 1740
rect 20689 1712 20753 1720
rect 20715 1711 20753 1712
rect 20716 1710 20753 1711
rect 20819 1744 20855 1745
rect 20927 1744 20963 1745
rect 20819 1736 20963 1744
rect 20819 1716 20827 1736
rect 20847 1732 20935 1736
rect 20847 1716 20891 1732
rect 20819 1712 20891 1716
rect 20911 1716 20935 1732
rect 20955 1716 20963 1736
rect 20911 1712 20963 1716
rect 20819 1710 20963 1712
rect 21029 1740 21067 1748
rect 21145 1744 21181 1745
rect 21029 1720 21038 1740
rect 21058 1720 21067 1740
rect 21029 1711 21067 1720
rect 21096 1736 21181 1744
rect 21096 1716 21153 1736
rect 21173 1716 21181 1736
rect 21029 1710 21066 1711
rect 21096 1710 21181 1716
rect 21247 1740 21285 1748
rect 21247 1720 21256 1740
rect 21276 1720 21285 1740
rect 21247 1711 21285 1720
rect 21429 1745 21471 1754
rect 21429 1727 21443 1745
rect 21461 1727 21471 1745
rect 21429 1719 21471 1727
rect 21434 1717 21471 1719
rect 21861 1739 22304 1778
rect 21247 1710 21284 1711
rect 20708 1682 20798 1688
rect 20708 1662 20724 1682
rect 20744 1680 20798 1682
rect 20744 1662 20769 1680
rect 20708 1660 20769 1662
rect 20789 1660 20798 1680
rect 20708 1654 20798 1660
rect 20721 1600 20758 1601
rect 20817 1600 20854 1601
rect 20873 1600 20909 1710
rect 21096 1689 21127 1710
rect 21861 1696 21908 1739
rect 22264 1734 22304 1739
rect 22929 1737 23116 1761
rect 23147 1742 23540 1762
rect 23560 1742 23563 1762
rect 23147 1737 23563 1742
rect 21092 1688 21127 1689
rect 20970 1678 21127 1688
rect 20970 1658 20987 1678
rect 21007 1658 21127 1678
rect 20970 1651 21127 1658
rect 21194 1681 21343 1689
rect 21194 1661 21205 1681
rect 21225 1661 21264 1681
rect 21284 1661 21343 1681
rect 21861 1678 21871 1696
rect 21889 1678 21908 1696
rect 21861 1674 21908 1678
rect 21862 1669 21899 1674
rect 21194 1654 21343 1661
rect 22929 1666 22966 1737
rect 23147 1736 23488 1737
rect 23081 1676 23112 1677
rect 21194 1653 21235 1654
rect 21431 1652 21468 1655
rect 20928 1600 20965 1601
rect 20621 1591 20759 1600
rect 19825 1552 20269 1578
rect 19825 1550 19993 1552
rect 18778 1418 19225 1430
rect 18821 1416 18854 1418
rect 18188 1398 18326 1407
rect 17982 1397 18019 1398
rect 17712 1344 17753 1345
rect 16982 1324 17019 1325
rect 16443 1296 16533 1302
rect 16443 1276 16459 1296
rect 16479 1294 16533 1296
rect 16479 1276 16504 1294
rect 16443 1274 16504 1276
rect 16524 1274 16533 1294
rect 16443 1268 16533 1274
rect 16456 1214 16493 1215
rect 16552 1214 16589 1215
rect 16608 1214 16644 1324
rect 16831 1303 16862 1324
rect 17486 1323 17538 1341
rect 17604 1337 17753 1344
rect 17604 1317 17663 1337
rect 17683 1317 17722 1337
rect 17742 1317 17753 1337
rect 17604 1309 17753 1317
rect 17820 1340 17977 1347
rect 17820 1320 17940 1340
rect 17960 1320 17977 1340
rect 17820 1310 17977 1320
rect 17820 1309 17855 1310
rect 16827 1302 16862 1303
rect 16705 1292 16862 1302
rect 16705 1272 16722 1292
rect 16742 1272 16862 1292
rect 16705 1265 16862 1272
rect 16929 1295 17078 1303
rect 16929 1275 16940 1295
rect 16960 1275 16999 1295
rect 17019 1275 17078 1295
rect 16929 1268 17078 1275
rect 17144 1271 17196 1289
rect 17820 1288 17851 1309
rect 18038 1288 18074 1398
rect 18093 1397 18130 1398
rect 18189 1397 18226 1398
rect 18149 1338 18239 1344
rect 18149 1318 18158 1338
rect 18178 1336 18239 1338
rect 18178 1318 18203 1336
rect 18149 1316 18203 1318
rect 18223 1316 18239 1336
rect 18149 1310 18239 1316
rect 17663 1287 17700 1288
rect 16929 1267 16970 1268
rect 16663 1214 16700 1215
rect 16356 1205 16494 1214
rect 16356 1185 16465 1205
rect 16485 1185 16494 1205
rect 16356 1178 16494 1185
rect 16552 1205 16700 1214
rect 16552 1185 16561 1205
rect 16581 1185 16671 1205
rect 16691 1185 16700 1205
rect 16356 1176 16452 1178
rect 16552 1175 16700 1185
rect 16759 1205 16796 1215
rect 16759 1185 16767 1205
rect 16787 1185 16796 1205
rect 16608 1174 16644 1175
rect 16759 1118 16796 1185
rect 16831 1214 16862 1265
rect 17144 1253 17162 1271
rect 17180 1253 17196 1271
rect 17662 1278 17700 1287
rect 16881 1214 16918 1215
rect 16831 1205 16918 1214
rect 16831 1185 16889 1205
rect 16909 1185 16918 1205
rect 16831 1175 16918 1185
rect 16977 1205 17014 1215
rect 16977 1185 16985 1205
rect 17005 1185 17014 1205
rect 16831 1174 16862 1175
rect 16456 1115 16493 1116
rect 16759 1115 16798 1118
rect 16455 1114 16798 1115
rect 16977 1114 17014 1185
rect 16380 1109 16798 1114
rect 16380 1089 16383 1109
rect 16403 1089 16798 1109
rect 16827 1090 17014 1114
rect 14921 1058 14958 1066
rect 14921 1039 14929 1058
rect 14950 1039 14958 1058
rect 14921 1033 14958 1039
rect 16759 1064 16798 1089
rect 17144 1064 17196 1253
rect 17490 1260 17530 1270
rect 17490 1242 17500 1260
rect 17518 1242 17530 1260
rect 17662 1258 17671 1278
rect 17691 1258 17700 1278
rect 17662 1250 17700 1258
rect 17766 1282 17851 1288
rect 17881 1287 17918 1288
rect 17766 1262 17774 1282
rect 17794 1262 17851 1282
rect 17766 1254 17851 1262
rect 17880 1278 17918 1287
rect 17880 1258 17889 1278
rect 17909 1258 17918 1278
rect 17766 1253 17802 1254
rect 17880 1250 17918 1258
rect 17984 1282 18128 1288
rect 17984 1262 17992 1282
rect 18012 1262 18045 1282
rect 18065 1262 18100 1282
rect 18120 1262 18128 1282
rect 17984 1254 18128 1262
rect 17984 1253 18020 1254
rect 18092 1253 18128 1254
rect 18194 1287 18231 1288
rect 18194 1286 18232 1287
rect 18194 1278 18258 1286
rect 18194 1258 18203 1278
rect 18223 1264 18258 1278
rect 18278 1264 18281 1284
rect 18223 1259 18281 1264
rect 18223 1258 18258 1259
rect 17490 1186 17530 1242
rect 17663 1221 17700 1250
rect 17664 1219 17700 1221
rect 17664 1197 17855 1219
rect 17881 1218 17918 1250
rect 18194 1246 18258 1258
rect 18298 1220 18325 1398
rect 19183 1373 19225 1418
rect 18157 1218 18325 1220
rect 17881 1208 18325 1218
rect 18466 1314 18653 1338
rect 18684 1319 19077 1339
rect 19097 1319 19100 1339
rect 18684 1314 19100 1319
rect 18466 1243 18503 1314
rect 18684 1313 19025 1314
rect 18618 1253 18649 1254
rect 18466 1223 18475 1243
rect 18495 1223 18503 1243
rect 18466 1213 18503 1223
rect 18562 1243 18649 1253
rect 18562 1223 18571 1243
rect 18591 1223 18649 1243
rect 18562 1214 18649 1223
rect 18562 1213 18599 1214
rect 17487 1181 17530 1186
rect 17878 1192 18325 1208
rect 17878 1186 17906 1192
rect 18157 1191 18325 1192
rect 17487 1178 17637 1181
rect 17878 1178 17905 1186
rect 17487 1176 17905 1178
rect 17487 1158 17496 1176
rect 17514 1158 17905 1176
rect 18618 1163 18649 1214
rect 18684 1243 18721 1313
rect 18987 1312 19024 1313
rect 18836 1253 18872 1254
rect 18684 1223 18693 1243
rect 18713 1223 18721 1243
rect 18684 1213 18721 1223
rect 18780 1243 18928 1253
rect 19028 1250 19124 1252
rect 18780 1223 18789 1243
rect 18809 1223 18899 1243
rect 18919 1223 18928 1243
rect 18780 1214 18928 1223
rect 18986 1243 19124 1250
rect 18986 1223 18995 1243
rect 19015 1223 19124 1243
rect 18986 1214 19124 1223
rect 18780 1213 18817 1214
rect 18510 1160 18551 1161
rect 17487 1155 17905 1158
rect 17487 1149 17530 1155
rect 17490 1146 17530 1149
rect 18405 1153 18551 1160
rect 17887 1137 17927 1138
rect 17598 1120 17927 1137
rect 18405 1133 18461 1153
rect 18481 1133 18520 1153
rect 18540 1133 18551 1153
rect 18405 1125 18551 1133
rect 18618 1156 18775 1163
rect 18618 1136 18738 1156
rect 18758 1136 18775 1156
rect 18618 1126 18775 1136
rect 18618 1125 18653 1126
rect 17482 1077 17525 1088
rect 16759 1046 17198 1064
rect 16759 1028 17159 1046
rect 17177 1028 17198 1046
rect 16759 1022 17198 1028
rect 16765 1018 17198 1022
rect 17482 1059 17494 1077
rect 17512 1059 17525 1077
rect 17482 1033 17525 1059
rect 17598 1033 17625 1120
rect 17887 1111 17927 1120
rect 17144 1016 17196 1018
rect 17482 1012 17625 1033
rect 17669 1085 17703 1101
rect 17887 1091 18280 1111
rect 18300 1091 18303 1111
rect 18618 1104 18649 1125
rect 18836 1104 18872 1214
rect 18891 1213 18928 1214
rect 18987 1213 19024 1214
rect 18947 1154 19037 1160
rect 18947 1134 18956 1154
rect 18976 1152 19037 1154
rect 18976 1134 19001 1152
rect 18947 1132 19001 1134
rect 19021 1132 19037 1152
rect 18947 1126 19037 1132
rect 18461 1103 18498 1104
rect 17887 1086 18303 1091
rect 18460 1094 18498 1103
rect 17887 1085 18228 1086
rect 17669 1015 17706 1085
rect 17821 1025 17852 1026
rect 17482 1010 17619 1012
rect 17482 968 17525 1010
rect 17669 995 17678 1015
rect 17698 995 17706 1015
rect 17669 985 17706 995
rect 17765 1015 17852 1025
rect 17765 995 17774 1015
rect 17794 995 17852 1015
rect 17765 986 17852 995
rect 17765 985 17802 986
rect 17480 958 17525 968
rect 17147 951 17184 956
rect 17138 947 17185 951
rect 17138 929 17157 947
rect 17175 929 17185 947
rect 17480 940 17489 958
rect 17507 940 17525 958
rect 17480 934 17525 940
rect 17821 935 17852 986
rect 17887 1015 17924 1085
rect 18190 1084 18227 1085
rect 18460 1074 18469 1094
rect 18489 1074 18498 1094
rect 18460 1066 18498 1074
rect 18564 1098 18649 1104
rect 18679 1103 18716 1104
rect 18564 1078 18572 1098
rect 18592 1078 18649 1098
rect 18564 1070 18649 1078
rect 18678 1094 18716 1103
rect 18678 1074 18687 1094
rect 18707 1074 18716 1094
rect 18564 1069 18600 1070
rect 18678 1066 18716 1074
rect 18782 1098 18926 1104
rect 18782 1078 18790 1098
rect 18810 1095 18898 1098
rect 18810 1078 18845 1095
rect 18782 1077 18845 1078
rect 18864 1078 18898 1095
rect 18918 1078 18926 1098
rect 18864 1077 18926 1078
rect 18782 1070 18926 1077
rect 18782 1069 18818 1070
rect 18890 1069 18926 1070
rect 18992 1103 19029 1104
rect 18992 1102 19030 1103
rect 19052 1102 19079 1106
rect 18992 1100 19079 1102
rect 18992 1094 19056 1100
rect 18992 1074 19001 1094
rect 19021 1080 19056 1094
rect 19076 1080 19079 1100
rect 19021 1075 19079 1080
rect 19021 1074 19056 1075
rect 18461 1037 18498 1066
rect 18462 1035 18498 1037
rect 18039 1025 18075 1026
rect 17887 995 17896 1015
rect 17916 995 17924 1015
rect 17887 985 17924 995
rect 17983 1015 18131 1025
rect 18231 1022 18327 1024
rect 17983 995 17992 1015
rect 18012 995 18102 1015
rect 18122 995 18131 1015
rect 17983 986 18131 995
rect 18189 1015 18327 1022
rect 18189 995 18198 1015
rect 18218 995 18327 1015
rect 18462 1013 18653 1035
rect 18679 1034 18716 1066
rect 18992 1062 19056 1074
rect 19096 1036 19123 1214
rect 18955 1034 19123 1036
rect 18679 1008 19123 1034
rect 18189 986 18327 995
rect 17983 985 18020 986
rect 17480 931 17517 934
rect 17713 932 17754 933
rect 17138 866 17185 929
rect 17605 925 17754 932
rect 17605 905 17664 925
rect 17684 905 17723 925
rect 17743 905 17754 925
rect 17605 897 17754 905
rect 17821 928 17978 935
rect 17821 908 17941 928
rect 17961 908 17978 928
rect 17821 898 17978 908
rect 17821 897 17856 898
rect 17821 876 17852 897
rect 18039 876 18075 986
rect 18094 985 18131 986
rect 18190 985 18227 986
rect 18150 926 18240 932
rect 18150 906 18159 926
rect 18179 924 18240 926
rect 18179 906 18204 924
rect 18150 904 18204 906
rect 18224 904 18240 924
rect 18150 898 18240 904
rect 17664 875 17701 876
rect 17477 867 17514 869
rect 17138 851 17188 866
rect 17138 826 17152 851
rect 17184 826 17188 851
rect 17477 859 17519 867
rect 17477 841 17487 859
rect 17505 841 17519 859
rect 17477 832 17519 841
rect 17663 866 17701 875
rect 17663 846 17672 866
rect 17692 846 17701 866
rect 17663 838 17701 846
rect 17767 870 17852 876
rect 17882 875 17919 876
rect 17767 850 17775 870
rect 17795 850 17852 870
rect 17767 842 17852 850
rect 17881 866 17919 875
rect 17881 846 17890 866
rect 17910 846 17919 866
rect 17767 841 17803 842
rect 17881 838 17919 846
rect 17985 874 18129 876
rect 17985 870 18037 874
rect 17985 850 17993 870
rect 18013 854 18037 870
rect 18057 870 18129 874
rect 18057 854 18101 870
rect 18013 850 18101 854
rect 18121 850 18129 870
rect 17985 842 18129 850
rect 17985 841 18021 842
rect 18093 841 18129 842
rect 18195 875 18232 876
rect 18195 874 18233 875
rect 18195 866 18259 874
rect 18195 846 18204 866
rect 18224 852 18259 866
rect 18279 852 18282 872
rect 18224 847 18282 852
rect 18224 846 18259 847
rect 17138 813 17185 826
rect 14523 788 14531 810
rect 14555 788 14563 810
rect 17478 807 17519 832
rect 17664 807 17701 838
rect 17882 816 17919 838
rect 18195 834 18259 846
rect 17877 807 17919 816
rect 18299 808 18326 986
rect 17478 795 17523 807
rect 14523 780 14563 788
rect 101 698 506 725
rect 542 698 545 725
rect 4465 711 4870 738
rect 4906 711 4909 738
rect 8842 723 9247 750
rect 9283 723 9286 750
rect 13206 736 13611 763
rect 13647 736 13650 763
rect 17474 737 17523 795
rect 17664 781 17726 807
rect 17877 806 17962 807
rect 18158 806 18326 808
rect 17877 780 18326 806
rect 17877 737 17916 780
rect 18158 779 18326 780
rect 18789 784 18829 1008
rect 18955 1007 19123 1008
rect 19187 1040 19220 1373
rect 19825 1372 19852 1550
rect 19892 1512 19956 1524
rect 20232 1520 20269 1552
rect 20295 1551 20486 1573
rect 20621 1571 20730 1591
rect 20750 1571 20759 1591
rect 20621 1564 20759 1571
rect 20817 1591 20965 1600
rect 20817 1571 20826 1591
rect 20846 1571 20936 1591
rect 20956 1571 20965 1591
rect 20621 1562 20717 1564
rect 20817 1561 20965 1571
rect 21024 1591 21061 1601
rect 21024 1571 21032 1591
rect 21052 1571 21061 1591
rect 20873 1560 20909 1561
rect 20450 1549 20486 1551
rect 20450 1520 20487 1549
rect 19892 1511 19927 1512
rect 19869 1506 19927 1511
rect 19869 1486 19872 1506
rect 19892 1492 19927 1506
rect 19947 1492 19956 1512
rect 19892 1484 19956 1492
rect 19918 1483 19956 1484
rect 19919 1482 19956 1483
rect 20022 1516 20058 1517
rect 20130 1516 20166 1517
rect 20022 1508 20166 1516
rect 20022 1488 20030 1508
rect 20050 1507 20138 1508
rect 20050 1488 20085 1507
rect 20106 1488 20138 1507
rect 20158 1488 20166 1508
rect 20022 1482 20166 1488
rect 20232 1512 20270 1520
rect 20348 1516 20384 1517
rect 20232 1492 20241 1512
rect 20261 1492 20270 1512
rect 20232 1483 20270 1492
rect 20299 1508 20384 1516
rect 20299 1488 20356 1508
rect 20376 1488 20384 1508
rect 20232 1482 20269 1483
rect 20299 1482 20384 1488
rect 20450 1512 20488 1520
rect 20450 1492 20459 1512
rect 20479 1492 20488 1512
rect 20721 1501 20758 1502
rect 21024 1501 21061 1571
rect 21096 1600 21127 1651
rect 21423 1646 21468 1652
rect 21423 1628 21441 1646
rect 21459 1628 21468 1646
rect 22929 1646 22938 1666
rect 22958 1646 22966 1666
rect 22929 1636 22966 1646
rect 23025 1666 23112 1676
rect 23025 1646 23034 1666
rect 23054 1646 23112 1666
rect 23025 1637 23112 1646
rect 23025 1636 23062 1637
rect 21423 1618 21468 1628
rect 21146 1600 21183 1601
rect 21096 1591 21183 1600
rect 21096 1571 21154 1591
rect 21174 1571 21183 1591
rect 21096 1561 21183 1571
rect 21242 1591 21279 1601
rect 21242 1571 21250 1591
rect 21270 1571 21279 1591
rect 21423 1576 21466 1618
rect 21850 1607 21902 1609
rect 21329 1574 21466 1576
rect 21096 1560 21127 1561
rect 21242 1501 21279 1571
rect 20720 1500 21061 1501
rect 20450 1483 20488 1492
rect 20645 1495 21061 1500
rect 20450 1482 20487 1483
rect 19911 1454 20001 1460
rect 19911 1434 19927 1454
rect 19947 1452 20001 1454
rect 19947 1434 19972 1452
rect 19911 1432 19972 1434
rect 19992 1432 20001 1452
rect 19911 1426 20001 1432
rect 19924 1372 19961 1373
rect 20020 1372 20057 1373
rect 20076 1372 20112 1482
rect 20299 1461 20330 1482
rect 20645 1475 20648 1495
rect 20668 1475 21061 1495
rect 21245 1485 21279 1501
rect 21323 1553 21466 1574
rect 21848 1603 22281 1607
rect 21848 1597 22287 1603
rect 21848 1579 21869 1597
rect 21887 1579 22287 1597
rect 23081 1586 23112 1637
rect 23147 1666 23184 1736
rect 23450 1735 23487 1736
rect 23299 1676 23335 1677
rect 23147 1646 23156 1666
rect 23176 1646 23184 1666
rect 23147 1636 23184 1646
rect 23243 1666 23391 1676
rect 23491 1673 23587 1675
rect 23243 1646 23252 1666
rect 23272 1646 23362 1666
rect 23382 1646 23391 1666
rect 23243 1637 23391 1646
rect 23449 1666 23587 1673
rect 23449 1646 23458 1666
rect 23478 1646 23587 1666
rect 23449 1637 23587 1646
rect 23243 1636 23280 1637
rect 22973 1583 23014 1584
rect 21848 1561 22287 1579
rect 21021 1466 21061 1475
rect 21323 1466 21350 1553
rect 21423 1527 21466 1553
rect 21423 1509 21436 1527
rect 21454 1509 21466 1527
rect 21423 1498 21466 1509
rect 20295 1460 20330 1461
rect 20173 1450 20330 1460
rect 20173 1430 20190 1450
rect 20210 1430 20330 1450
rect 20173 1423 20330 1430
rect 20397 1453 20546 1461
rect 20397 1433 20408 1453
rect 20428 1433 20467 1453
rect 20487 1433 20546 1453
rect 21021 1449 21350 1466
rect 21021 1448 21061 1449
rect 20397 1426 20546 1433
rect 21418 1437 21458 1440
rect 21418 1431 21461 1437
rect 21043 1428 21461 1431
rect 20397 1425 20438 1426
rect 20131 1372 20168 1373
rect 19824 1363 19962 1372
rect 19824 1343 19933 1363
rect 19953 1343 19962 1363
rect 19824 1336 19962 1343
rect 20020 1363 20168 1372
rect 20020 1343 20029 1363
rect 20049 1343 20139 1363
rect 20159 1343 20168 1363
rect 19824 1334 19920 1336
rect 20020 1333 20168 1343
rect 20227 1363 20264 1373
rect 20227 1343 20235 1363
rect 20255 1343 20264 1363
rect 20076 1332 20112 1333
rect 19924 1273 19961 1274
rect 20227 1273 20264 1343
rect 20299 1372 20330 1423
rect 21043 1410 21434 1428
rect 21452 1410 21461 1428
rect 21043 1408 21461 1410
rect 21043 1400 21070 1408
rect 21311 1405 21461 1408
rect 20623 1394 20791 1395
rect 21042 1394 21070 1400
rect 20623 1378 21070 1394
rect 21418 1400 21461 1405
rect 20349 1372 20386 1373
rect 20299 1363 20386 1372
rect 20299 1343 20357 1363
rect 20377 1343 20386 1363
rect 20299 1333 20386 1343
rect 20445 1363 20482 1373
rect 20445 1343 20453 1363
rect 20473 1343 20482 1363
rect 20299 1332 20330 1333
rect 19923 1272 20264 1273
rect 20445 1272 20482 1343
rect 19848 1267 20264 1272
rect 19848 1247 19851 1267
rect 19871 1247 20264 1267
rect 20295 1248 20482 1272
rect 20623 1368 21067 1378
rect 20623 1366 20791 1368
rect 20623 1188 20650 1366
rect 20690 1328 20754 1340
rect 21030 1336 21067 1368
rect 21093 1367 21284 1389
rect 21248 1365 21284 1367
rect 21248 1336 21285 1365
rect 21418 1344 21458 1400
rect 20690 1327 20725 1328
rect 20667 1322 20725 1327
rect 20667 1302 20670 1322
rect 20690 1308 20725 1322
rect 20745 1308 20754 1328
rect 20690 1300 20754 1308
rect 20716 1299 20754 1300
rect 20717 1298 20754 1299
rect 20820 1332 20856 1333
rect 20928 1332 20964 1333
rect 20820 1324 20964 1332
rect 20820 1304 20828 1324
rect 20848 1304 20883 1324
rect 20903 1304 20936 1324
rect 20956 1304 20964 1324
rect 20820 1298 20964 1304
rect 21030 1328 21068 1336
rect 21146 1332 21182 1333
rect 21030 1308 21039 1328
rect 21059 1308 21068 1328
rect 21030 1299 21068 1308
rect 21097 1324 21182 1332
rect 21097 1304 21154 1324
rect 21174 1304 21182 1324
rect 21030 1298 21067 1299
rect 21097 1298 21182 1304
rect 21248 1328 21286 1336
rect 21248 1308 21257 1328
rect 21277 1308 21286 1328
rect 21418 1326 21430 1344
rect 21448 1326 21458 1344
rect 21850 1372 21902 1561
rect 22248 1536 22287 1561
rect 22865 1576 23014 1583
rect 22865 1556 22924 1576
rect 22944 1556 22983 1576
rect 23003 1556 23014 1576
rect 22865 1548 23014 1556
rect 23081 1579 23238 1586
rect 23081 1559 23201 1579
rect 23221 1559 23238 1579
rect 23081 1549 23238 1559
rect 23081 1548 23116 1549
rect 22032 1511 22219 1535
rect 22248 1516 22643 1536
rect 22663 1516 22666 1536
rect 23081 1527 23112 1548
rect 23299 1527 23335 1637
rect 23354 1636 23391 1637
rect 23450 1636 23487 1637
rect 23410 1577 23500 1583
rect 23410 1557 23419 1577
rect 23439 1575 23500 1577
rect 23439 1557 23464 1575
rect 23410 1555 23464 1557
rect 23484 1555 23500 1575
rect 23410 1549 23500 1555
rect 22924 1526 22961 1527
rect 22248 1511 22666 1516
rect 22923 1517 22961 1526
rect 22032 1440 22069 1511
rect 22248 1510 22591 1511
rect 22248 1507 22287 1510
rect 22553 1509 22590 1510
rect 22184 1450 22215 1451
rect 22032 1420 22041 1440
rect 22061 1420 22069 1440
rect 22032 1410 22069 1420
rect 22128 1440 22215 1450
rect 22128 1420 22137 1440
rect 22157 1420 22215 1440
rect 22128 1411 22215 1420
rect 22128 1410 22165 1411
rect 21850 1354 21866 1372
rect 21884 1354 21902 1372
rect 22184 1360 22215 1411
rect 22250 1440 22287 1507
rect 22923 1497 22932 1517
rect 22952 1497 22961 1517
rect 22923 1489 22961 1497
rect 23027 1521 23112 1527
rect 23142 1526 23179 1527
rect 23027 1501 23035 1521
rect 23055 1501 23112 1521
rect 23027 1493 23112 1501
rect 23141 1517 23179 1526
rect 23141 1497 23150 1517
rect 23170 1497 23179 1517
rect 23027 1492 23063 1493
rect 23141 1489 23179 1497
rect 23245 1521 23389 1527
rect 23245 1501 23253 1521
rect 23273 1516 23361 1521
rect 23273 1501 23309 1516
rect 23245 1499 23309 1501
rect 23328 1501 23361 1516
rect 23381 1501 23389 1521
rect 23328 1499 23389 1501
rect 23245 1493 23389 1499
rect 23245 1492 23281 1493
rect 23353 1492 23389 1493
rect 23455 1526 23492 1527
rect 23455 1525 23493 1526
rect 23455 1517 23519 1525
rect 23455 1497 23464 1517
rect 23484 1503 23519 1517
rect 23539 1503 23542 1523
rect 23484 1498 23542 1503
rect 23484 1497 23519 1498
rect 22924 1460 22961 1489
rect 22925 1458 22961 1460
rect 22402 1450 22438 1451
rect 22250 1420 22259 1440
rect 22279 1420 22287 1440
rect 22250 1410 22287 1420
rect 22346 1440 22494 1450
rect 22594 1447 22690 1449
rect 22346 1420 22355 1440
rect 22375 1420 22465 1440
rect 22485 1420 22494 1440
rect 22346 1411 22494 1420
rect 22552 1440 22690 1447
rect 22552 1420 22561 1440
rect 22581 1420 22690 1440
rect 22925 1436 23116 1458
rect 23142 1457 23179 1489
rect 23455 1485 23519 1497
rect 23559 1459 23586 1637
rect 23418 1457 23586 1459
rect 23142 1443 23586 1457
rect 24189 1591 24357 1592
rect 24483 1591 24523 1815
rect 24986 1819 25154 1820
rect 25389 1819 25429 1852
rect 25785 1819 25832 1852
rect 26236 1850 26277 1875
rect 26422 1850 26459 1881
rect 26640 1850 26677 1881
rect 26953 1877 27017 1889
rect 27057 1851 27084 2029
rect 26236 1823 26285 1850
rect 26421 1824 26470 1850
rect 26639 1849 26720 1850
rect 26916 1849 27084 1851
rect 26639 1824 27084 1849
rect 26640 1823 27084 1824
rect 24986 1818 25430 1819
rect 24986 1793 25431 1818
rect 24986 1791 25154 1793
rect 25350 1792 25431 1793
rect 25600 1792 25649 1818
rect 25785 1792 25834 1819
rect 24986 1613 25013 1791
rect 25053 1753 25117 1765
rect 25393 1761 25430 1792
rect 25611 1761 25648 1792
rect 25793 1767 25834 1792
rect 26238 1790 26285 1823
rect 26641 1790 26681 1823
rect 26916 1822 27084 1823
rect 27547 1827 27587 2051
rect 27713 2050 27881 2051
rect 28484 2185 28928 2199
rect 28484 2183 28652 2185
rect 28484 2005 28511 2183
rect 28551 2145 28615 2157
rect 28891 2153 28928 2185
rect 28954 2184 29145 2206
rect 29380 2202 29489 2222
rect 29509 2202 29518 2222
rect 29380 2195 29518 2202
rect 29576 2222 29724 2231
rect 29576 2202 29585 2222
rect 29605 2202 29695 2222
rect 29715 2202 29724 2222
rect 29380 2193 29476 2195
rect 29576 2192 29724 2202
rect 29783 2222 29820 2232
rect 29783 2202 29791 2222
rect 29811 2202 29820 2222
rect 29632 2191 29668 2192
rect 29109 2182 29145 2184
rect 29109 2153 29146 2182
rect 28551 2144 28586 2145
rect 28528 2139 28586 2144
rect 28528 2119 28531 2139
rect 28551 2125 28586 2139
rect 28606 2125 28615 2145
rect 28551 2117 28615 2125
rect 28577 2116 28615 2117
rect 28578 2115 28615 2116
rect 28681 2149 28717 2150
rect 28789 2149 28825 2150
rect 28681 2141 28825 2149
rect 28681 2121 28689 2141
rect 28709 2139 28797 2141
rect 28709 2121 28742 2139
rect 28681 2120 28742 2121
rect 28763 2121 28797 2139
rect 28817 2121 28825 2141
rect 28763 2120 28825 2121
rect 28681 2115 28825 2120
rect 28891 2145 28929 2153
rect 29007 2149 29043 2150
rect 28891 2125 28900 2145
rect 28920 2125 28929 2145
rect 28891 2116 28929 2125
rect 28958 2141 29043 2149
rect 28958 2121 29015 2141
rect 29035 2121 29043 2141
rect 28891 2115 28928 2116
rect 28958 2115 29043 2121
rect 29109 2145 29147 2153
rect 29109 2125 29118 2145
rect 29138 2125 29147 2145
rect 29783 2135 29820 2202
rect 29855 2231 29886 2282
rect 30168 2270 30186 2288
rect 30204 2270 30220 2288
rect 29905 2231 29942 2232
rect 29855 2222 29942 2231
rect 29855 2202 29913 2222
rect 29933 2202 29942 2222
rect 29855 2192 29942 2202
rect 30001 2222 30038 2232
rect 30001 2202 30009 2222
rect 30029 2202 30038 2222
rect 29855 2191 29886 2192
rect 29480 2132 29517 2133
rect 29783 2132 29822 2135
rect 29479 2131 29822 2132
rect 30001 2131 30038 2202
rect 29109 2116 29147 2125
rect 29404 2126 29822 2131
rect 29109 2115 29146 2116
rect 28570 2087 28660 2093
rect 28570 2067 28586 2087
rect 28606 2085 28660 2087
rect 28606 2067 28631 2085
rect 28570 2065 28631 2067
rect 28651 2065 28660 2085
rect 28570 2059 28660 2065
rect 28583 2005 28620 2006
rect 28679 2005 28716 2006
rect 28735 2005 28771 2115
rect 28958 2094 28989 2115
rect 29404 2106 29407 2126
rect 29427 2106 29822 2126
rect 29851 2107 30038 2131
rect 28954 2093 28989 2094
rect 28832 2083 28989 2093
rect 28832 2063 28849 2083
rect 28869 2063 28989 2083
rect 28832 2056 28989 2063
rect 29056 2086 29205 2094
rect 29056 2066 29067 2086
rect 29087 2066 29126 2086
rect 29146 2066 29205 2086
rect 29056 2059 29205 2066
rect 29783 2081 29822 2106
rect 30168 2081 30220 2270
rect 30612 2298 30622 2316
rect 30640 2298 30652 2316
rect 30784 2314 30793 2334
rect 30813 2314 30822 2334
rect 30784 2306 30822 2314
rect 30888 2338 30973 2344
rect 31003 2343 31040 2344
rect 30888 2318 30896 2338
rect 30916 2318 30973 2338
rect 30888 2310 30973 2318
rect 31002 2334 31040 2343
rect 31002 2314 31011 2334
rect 31031 2314 31040 2334
rect 30888 2309 30924 2310
rect 31002 2306 31040 2314
rect 31106 2338 31250 2344
rect 31106 2318 31114 2338
rect 31134 2318 31167 2338
rect 31187 2318 31222 2338
rect 31242 2318 31250 2338
rect 31106 2310 31250 2318
rect 31106 2309 31142 2310
rect 31214 2309 31250 2310
rect 31316 2343 31353 2344
rect 31316 2342 31354 2343
rect 31316 2334 31380 2342
rect 31316 2314 31325 2334
rect 31345 2320 31380 2334
rect 31400 2320 31403 2340
rect 31345 2315 31403 2320
rect 31345 2314 31380 2315
rect 30612 2242 30652 2298
rect 30785 2277 30822 2306
rect 30786 2275 30822 2277
rect 30786 2253 30977 2275
rect 31003 2274 31040 2306
rect 31316 2302 31380 2314
rect 31420 2276 31447 2454
rect 31279 2274 31447 2276
rect 31003 2264 31447 2274
rect 31588 2370 31775 2394
rect 31806 2375 32199 2395
rect 32219 2375 32222 2395
rect 31806 2370 32222 2375
rect 31588 2299 31625 2370
rect 31806 2369 32147 2370
rect 31740 2309 31771 2310
rect 31588 2279 31597 2299
rect 31617 2279 31625 2299
rect 31588 2269 31625 2279
rect 31684 2299 31771 2309
rect 31684 2279 31693 2299
rect 31713 2279 31771 2299
rect 31684 2270 31771 2279
rect 31684 2269 31721 2270
rect 30609 2237 30652 2242
rect 31000 2248 31447 2264
rect 31000 2242 31028 2248
rect 31279 2247 31447 2248
rect 30609 2234 30759 2237
rect 31000 2234 31027 2242
rect 30609 2232 31027 2234
rect 30609 2214 30618 2232
rect 30636 2214 31027 2232
rect 31740 2219 31771 2270
rect 31806 2299 31843 2369
rect 32109 2368 32146 2369
rect 32347 2311 32380 2470
rect 31958 2309 31994 2310
rect 31806 2279 31815 2299
rect 31835 2279 31843 2299
rect 31806 2269 31843 2279
rect 31902 2299 32050 2309
rect 32150 2306 32246 2308
rect 31902 2279 31911 2299
rect 31931 2279 32021 2299
rect 32041 2279 32050 2299
rect 31902 2270 32050 2279
rect 32108 2299 32246 2306
rect 32108 2279 32117 2299
rect 32137 2279 32246 2299
rect 32347 2307 32383 2311
rect 32347 2289 32356 2307
rect 32378 2289 32383 2307
rect 32347 2283 32383 2289
rect 32108 2270 32246 2279
rect 31902 2269 31939 2270
rect 31632 2216 31673 2217
rect 30609 2211 31027 2214
rect 30609 2205 30652 2211
rect 30612 2202 30652 2205
rect 31524 2209 31673 2216
rect 31009 2193 31049 2194
rect 30720 2176 31049 2193
rect 31524 2189 31583 2209
rect 31603 2189 31642 2209
rect 31662 2189 31673 2209
rect 31524 2181 31673 2189
rect 31740 2212 31897 2219
rect 31740 2192 31860 2212
rect 31880 2192 31897 2212
rect 31740 2182 31897 2192
rect 31740 2181 31775 2182
rect 30604 2133 30647 2144
rect 30604 2115 30616 2133
rect 30634 2115 30647 2133
rect 30604 2089 30647 2115
rect 30720 2089 30747 2176
rect 31009 2167 31049 2176
rect 29783 2063 30222 2081
rect 29056 2058 29097 2059
rect 28790 2005 28827 2006
rect 28483 1996 28621 2005
rect 28483 1976 28592 1996
rect 28612 1976 28621 1996
rect 28483 1969 28621 1976
rect 28679 1996 28827 2005
rect 28679 1976 28688 1996
rect 28708 1976 28798 1996
rect 28818 1976 28827 1996
rect 28483 1967 28579 1969
rect 28679 1966 28827 1976
rect 28886 1996 28923 2006
rect 28886 1976 28894 1996
rect 28914 1976 28923 1996
rect 28735 1965 28771 1966
rect 28583 1906 28620 1907
rect 28886 1906 28923 1976
rect 28958 2005 28989 2056
rect 29783 2045 30183 2063
rect 30201 2045 30222 2063
rect 29783 2039 30222 2045
rect 29789 2035 30222 2039
rect 30604 2068 30747 2089
rect 30791 2141 30825 2157
rect 31009 2147 31402 2167
rect 31422 2147 31425 2167
rect 31740 2160 31771 2181
rect 31958 2160 31994 2270
rect 32013 2269 32050 2270
rect 32109 2269 32146 2270
rect 32069 2210 32159 2216
rect 32069 2190 32078 2210
rect 32098 2208 32159 2210
rect 32098 2190 32123 2208
rect 32069 2188 32123 2190
rect 32143 2188 32159 2208
rect 32069 2182 32159 2188
rect 31583 2159 31620 2160
rect 31009 2142 31425 2147
rect 31582 2150 31620 2159
rect 31009 2141 31350 2142
rect 30791 2071 30828 2141
rect 30943 2081 30974 2082
rect 30604 2066 30741 2068
rect 30168 2033 30220 2035
rect 30604 2024 30647 2066
rect 30791 2051 30800 2071
rect 30820 2051 30828 2071
rect 30791 2041 30828 2051
rect 30887 2071 30974 2081
rect 30887 2051 30896 2071
rect 30916 2051 30974 2071
rect 30887 2042 30974 2051
rect 30887 2041 30924 2042
rect 30602 2014 30647 2024
rect 29008 2005 29045 2006
rect 28958 1996 29045 2005
rect 28958 1976 29016 1996
rect 29036 1976 29045 1996
rect 28958 1966 29045 1976
rect 29104 1996 29141 2006
rect 29104 1976 29112 1996
rect 29132 1976 29141 1996
rect 30602 1996 30611 2014
rect 30629 1996 30647 2014
rect 30602 1990 30647 1996
rect 30943 1991 30974 2042
rect 31009 2071 31046 2141
rect 31312 2140 31349 2141
rect 31582 2130 31591 2150
rect 31611 2130 31620 2150
rect 31582 2122 31620 2130
rect 31686 2154 31771 2160
rect 31801 2159 31838 2160
rect 31686 2134 31694 2154
rect 31714 2134 31771 2154
rect 31686 2126 31771 2134
rect 31800 2150 31838 2159
rect 31800 2130 31809 2150
rect 31829 2130 31838 2150
rect 31686 2125 31722 2126
rect 31800 2122 31838 2130
rect 31904 2154 32048 2160
rect 31904 2134 31912 2154
rect 31932 2135 31964 2154
rect 31985 2135 32020 2154
rect 31932 2134 32020 2135
rect 32040 2134 32048 2154
rect 31904 2126 32048 2134
rect 31904 2125 31940 2126
rect 32012 2125 32048 2126
rect 32114 2159 32151 2160
rect 32114 2158 32152 2159
rect 32114 2150 32178 2158
rect 32114 2130 32123 2150
rect 32143 2136 32178 2150
rect 32198 2136 32201 2156
rect 32143 2131 32201 2136
rect 32143 2130 32178 2131
rect 31583 2093 31620 2122
rect 31584 2091 31620 2093
rect 31161 2081 31197 2082
rect 31009 2051 31018 2071
rect 31038 2051 31046 2071
rect 31009 2041 31046 2051
rect 31105 2071 31253 2081
rect 31353 2078 31449 2080
rect 31105 2051 31114 2071
rect 31134 2051 31224 2071
rect 31244 2051 31253 2071
rect 31105 2042 31253 2051
rect 31311 2071 31449 2078
rect 31311 2051 31320 2071
rect 31340 2051 31449 2071
rect 31584 2069 31775 2091
rect 31801 2090 31838 2122
rect 32114 2118 32178 2130
rect 32218 2092 32245 2270
rect 32850 2269 32883 2602
rect 32947 2634 33115 2635
rect 33241 2634 33281 2858
rect 33744 2862 33912 2863
rect 34148 2862 34189 2896
rect 34546 2875 34593 2896
rect 33744 2852 34189 2862
rect 34261 2860 34404 2861
rect 33744 2836 34188 2852
rect 33744 2834 33912 2836
rect 34108 2835 34188 2836
rect 34261 2835 34406 2860
rect 34548 2835 34593 2875
rect 33744 2656 33771 2834
rect 33811 2796 33875 2808
rect 34151 2804 34188 2835
rect 34369 2804 34406 2835
rect 34551 2828 34593 2835
rect 33811 2795 33846 2796
rect 33788 2790 33846 2795
rect 33788 2770 33791 2790
rect 33811 2776 33846 2790
rect 33866 2776 33875 2796
rect 33811 2768 33875 2776
rect 33837 2767 33875 2768
rect 33838 2766 33875 2767
rect 33941 2800 33977 2801
rect 34049 2800 34085 2801
rect 33941 2792 34085 2800
rect 33941 2772 33949 2792
rect 33969 2788 34057 2792
rect 33969 2772 34013 2788
rect 33941 2768 34013 2772
rect 34033 2772 34057 2788
rect 34077 2772 34085 2792
rect 34033 2768 34085 2772
rect 33941 2766 34085 2768
rect 34151 2796 34189 2804
rect 34267 2800 34303 2801
rect 34151 2776 34160 2796
rect 34180 2776 34189 2796
rect 34151 2767 34189 2776
rect 34218 2792 34303 2800
rect 34218 2772 34275 2792
rect 34295 2772 34303 2792
rect 34151 2766 34188 2767
rect 34218 2766 34303 2772
rect 34369 2796 34407 2804
rect 34369 2776 34378 2796
rect 34398 2776 34407 2796
rect 34369 2767 34407 2776
rect 34551 2801 34594 2828
rect 34551 2783 34565 2801
rect 34583 2783 34594 2801
rect 34551 2775 34594 2783
rect 34556 2773 34594 2775
rect 34369 2766 34406 2767
rect 33830 2738 33920 2744
rect 33830 2718 33846 2738
rect 33866 2736 33920 2738
rect 33866 2718 33891 2736
rect 33830 2716 33891 2718
rect 33911 2716 33920 2736
rect 33830 2710 33920 2716
rect 33843 2656 33880 2657
rect 33939 2656 33976 2657
rect 33995 2656 34031 2766
rect 34218 2745 34249 2766
rect 34214 2744 34249 2745
rect 34092 2734 34249 2744
rect 34092 2714 34109 2734
rect 34129 2714 34249 2734
rect 34092 2707 34249 2714
rect 34316 2737 34465 2745
rect 34316 2717 34327 2737
rect 34347 2717 34386 2737
rect 34406 2717 34465 2737
rect 34316 2710 34465 2717
rect 34316 2709 34357 2710
rect 34553 2708 34590 2711
rect 34050 2656 34087 2657
rect 33743 2647 33881 2656
rect 32947 2608 33391 2634
rect 32947 2606 33115 2608
rect 32947 2428 32974 2606
rect 33014 2568 33078 2580
rect 33354 2576 33391 2608
rect 33417 2607 33608 2629
rect 33743 2627 33852 2647
rect 33872 2627 33881 2647
rect 33743 2620 33881 2627
rect 33939 2647 34087 2656
rect 33939 2627 33948 2647
rect 33968 2627 34058 2647
rect 34078 2627 34087 2647
rect 33743 2618 33839 2620
rect 33939 2617 34087 2627
rect 34146 2647 34183 2657
rect 34146 2627 34154 2647
rect 34174 2627 34183 2647
rect 33995 2616 34031 2617
rect 33572 2605 33608 2607
rect 33572 2576 33609 2605
rect 33014 2567 33049 2568
rect 32991 2562 33049 2567
rect 32991 2542 32994 2562
rect 33014 2548 33049 2562
rect 33069 2548 33078 2568
rect 33014 2542 33078 2548
rect 32991 2540 33078 2542
rect 32991 2536 33018 2540
rect 33040 2539 33078 2540
rect 33041 2538 33078 2539
rect 33144 2572 33180 2573
rect 33252 2572 33288 2573
rect 33144 2565 33288 2572
rect 33144 2564 33206 2565
rect 33144 2544 33152 2564
rect 33172 2547 33206 2564
rect 33225 2564 33288 2565
rect 33225 2547 33260 2564
rect 33172 2544 33260 2547
rect 33280 2544 33288 2564
rect 33144 2538 33288 2544
rect 33354 2568 33392 2576
rect 33470 2572 33506 2573
rect 33354 2548 33363 2568
rect 33383 2548 33392 2568
rect 33354 2539 33392 2548
rect 33421 2564 33506 2572
rect 33421 2544 33478 2564
rect 33498 2544 33506 2564
rect 33354 2538 33391 2539
rect 33421 2538 33506 2544
rect 33572 2568 33610 2576
rect 33572 2548 33581 2568
rect 33601 2548 33610 2568
rect 33843 2557 33880 2558
rect 34146 2557 34183 2627
rect 34218 2656 34249 2707
rect 34545 2702 34590 2708
rect 34545 2684 34563 2702
rect 34581 2684 34590 2702
rect 34545 2674 34590 2684
rect 34268 2656 34305 2657
rect 34218 2647 34305 2656
rect 34218 2627 34276 2647
rect 34296 2627 34305 2647
rect 34218 2617 34305 2627
rect 34364 2647 34401 2657
rect 34364 2627 34372 2647
rect 34392 2627 34401 2647
rect 34545 2632 34588 2674
rect 34451 2630 34588 2632
rect 34218 2616 34249 2617
rect 34364 2557 34401 2627
rect 33842 2556 34183 2557
rect 33572 2539 33610 2548
rect 33767 2551 34183 2556
rect 33572 2538 33609 2539
rect 33033 2510 33123 2516
rect 33033 2490 33049 2510
rect 33069 2508 33123 2510
rect 33069 2490 33094 2508
rect 33033 2488 33094 2490
rect 33114 2488 33123 2508
rect 33033 2482 33123 2488
rect 33046 2428 33083 2429
rect 33142 2428 33179 2429
rect 33198 2428 33234 2538
rect 33421 2517 33452 2538
rect 33767 2531 33770 2551
rect 33790 2531 34183 2551
rect 34367 2541 34401 2557
rect 34445 2609 34588 2630
rect 34143 2522 34183 2531
rect 34445 2522 34472 2609
rect 34545 2583 34588 2609
rect 34545 2565 34558 2583
rect 34576 2565 34588 2583
rect 34545 2554 34588 2565
rect 33417 2516 33452 2517
rect 33295 2506 33452 2516
rect 33295 2486 33312 2506
rect 33332 2486 33452 2506
rect 33295 2479 33452 2486
rect 33519 2509 33665 2517
rect 33519 2489 33530 2509
rect 33550 2489 33589 2509
rect 33609 2489 33665 2509
rect 34143 2505 34472 2522
rect 34143 2504 34183 2505
rect 33519 2482 33665 2489
rect 34540 2493 34580 2496
rect 34540 2487 34583 2493
rect 34165 2484 34583 2487
rect 33519 2481 33560 2482
rect 33253 2428 33290 2429
rect 32946 2419 33084 2428
rect 32946 2399 33055 2419
rect 33075 2399 33084 2419
rect 32946 2392 33084 2399
rect 33142 2419 33290 2428
rect 33142 2399 33151 2419
rect 33171 2399 33261 2419
rect 33281 2399 33290 2419
rect 32946 2390 33042 2392
rect 33142 2389 33290 2399
rect 33349 2419 33386 2429
rect 33349 2399 33357 2419
rect 33377 2399 33386 2419
rect 33198 2388 33234 2389
rect 33046 2329 33083 2330
rect 33349 2329 33386 2399
rect 33421 2428 33452 2479
rect 34165 2466 34556 2484
rect 34574 2466 34583 2484
rect 34165 2464 34583 2466
rect 34165 2456 34192 2464
rect 34433 2461 34583 2464
rect 33745 2450 33913 2451
rect 34164 2450 34192 2456
rect 33745 2434 34192 2450
rect 34540 2456 34583 2461
rect 33471 2428 33508 2429
rect 33421 2419 33508 2428
rect 33421 2399 33479 2419
rect 33499 2399 33508 2419
rect 33421 2389 33508 2399
rect 33567 2419 33604 2429
rect 33567 2399 33575 2419
rect 33595 2399 33604 2419
rect 33421 2388 33452 2389
rect 33045 2328 33386 2329
rect 33567 2328 33604 2399
rect 32970 2323 33386 2328
rect 32970 2303 32973 2323
rect 32993 2303 33386 2323
rect 33417 2304 33604 2328
rect 33745 2424 34189 2434
rect 33745 2422 33913 2424
rect 32845 2224 32887 2269
rect 33745 2244 33772 2422
rect 33812 2384 33876 2396
rect 34152 2392 34189 2424
rect 34215 2423 34406 2445
rect 34370 2421 34406 2423
rect 34370 2392 34407 2421
rect 34540 2400 34580 2456
rect 33812 2383 33847 2384
rect 33789 2378 33847 2383
rect 33789 2358 33792 2378
rect 33812 2364 33847 2378
rect 33867 2364 33876 2384
rect 33812 2356 33876 2364
rect 33838 2355 33876 2356
rect 33839 2354 33876 2355
rect 33942 2388 33978 2389
rect 34050 2388 34086 2389
rect 33942 2380 34086 2388
rect 33942 2360 33950 2380
rect 33970 2360 34005 2380
rect 34025 2360 34058 2380
rect 34078 2360 34086 2380
rect 33942 2354 34086 2360
rect 34152 2384 34190 2392
rect 34268 2388 34304 2389
rect 34152 2364 34161 2384
rect 34181 2364 34190 2384
rect 34152 2355 34190 2364
rect 34219 2380 34304 2388
rect 34219 2360 34276 2380
rect 34296 2360 34304 2380
rect 34152 2354 34189 2355
rect 34219 2354 34304 2360
rect 34370 2384 34408 2392
rect 34370 2364 34379 2384
rect 34399 2364 34408 2384
rect 34540 2382 34552 2400
rect 34570 2382 34580 2400
rect 34540 2372 34580 2382
rect 34370 2355 34408 2364
rect 34370 2354 34407 2355
rect 33831 2326 33921 2332
rect 33831 2306 33847 2326
rect 33867 2324 33921 2326
rect 33867 2306 33892 2324
rect 33831 2304 33892 2306
rect 33912 2304 33921 2324
rect 33831 2298 33921 2304
rect 33844 2244 33881 2245
rect 33940 2244 33977 2245
rect 33996 2244 34032 2354
rect 34219 2333 34250 2354
rect 34215 2332 34250 2333
rect 34093 2322 34250 2332
rect 34093 2302 34110 2322
rect 34130 2302 34250 2322
rect 34093 2295 34250 2302
rect 34317 2325 34466 2333
rect 34317 2305 34328 2325
rect 34348 2305 34387 2325
rect 34407 2305 34466 2325
rect 34317 2298 34466 2305
rect 34532 2301 34584 2319
rect 34317 2297 34358 2298
rect 34051 2244 34088 2245
rect 33744 2235 33882 2244
rect 33216 2224 33249 2226
rect 32845 2212 33292 2224
rect 32077 2090 32245 2092
rect 31801 2064 32245 2090
rect 31311 2042 31449 2051
rect 31105 2041 31142 2042
rect 30602 1987 30639 1990
rect 30835 1988 30876 1989
rect 28958 1965 28989 1966
rect 28582 1905 28923 1906
rect 29104 1905 29141 1976
rect 30727 1981 30876 1988
rect 30171 1968 30208 1973
rect 30162 1964 30209 1968
rect 30162 1946 30181 1964
rect 30199 1946 30209 1964
rect 30727 1961 30786 1981
rect 30806 1961 30845 1981
rect 30865 1961 30876 1981
rect 30727 1953 30876 1961
rect 30943 1984 31100 1991
rect 30943 1964 31063 1984
rect 31083 1964 31100 1984
rect 30943 1954 31100 1964
rect 30943 1953 30978 1954
rect 28507 1900 28923 1905
rect 28507 1880 28510 1900
rect 28530 1880 28923 1900
rect 28954 1881 29141 1905
rect 29766 1903 29806 1908
rect 30162 1903 30209 1946
rect 30943 1932 30974 1953
rect 31161 1932 31197 2042
rect 31216 2041 31253 2042
rect 31312 2041 31349 2042
rect 31272 1982 31362 1988
rect 31272 1962 31281 1982
rect 31301 1980 31362 1982
rect 31301 1962 31326 1980
rect 31272 1960 31326 1962
rect 31346 1960 31362 1980
rect 31272 1954 31362 1960
rect 30786 1931 30823 1932
rect 29766 1864 30209 1903
rect 30599 1923 30636 1925
rect 30599 1915 30641 1923
rect 30599 1897 30609 1915
rect 30627 1897 30641 1915
rect 30599 1888 30641 1897
rect 30785 1922 30823 1931
rect 30785 1902 30794 1922
rect 30814 1902 30823 1922
rect 30785 1894 30823 1902
rect 30889 1926 30974 1932
rect 31004 1931 31041 1932
rect 30889 1906 30897 1926
rect 30917 1906 30974 1926
rect 30889 1898 30974 1906
rect 31003 1922 31041 1931
rect 31003 1902 31012 1922
rect 31032 1902 31041 1922
rect 30889 1897 30925 1898
rect 31003 1894 31041 1902
rect 31107 1930 31251 1932
rect 31107 1926 31159 1930
rect 31107 1906 31115 1926
rect 31135 1910 31159 1926
rect 31179 1926 31251 1930
rect 31179 1910 31223 1926
rect 31135 1906 31223 1910
rect 31243 1906 31251 1926
rect 31107 1898 31251 1906
rect 31107 1897 31143 1898
rect 31215 1897 31251 1898
rect 31317 1931 31354 1932
rect 31317 1930 31355 1931
rect 31317 1922 31381 1930
rect 31317 1902 31326 1922
rect 31346 1908 31381 1922
rect 31401 1908 31404 1928
rect 31346 1903 31404 1908
rect 31346 1902 31381 1903
rect 27547 1805 27555 1827
rect 27579 1805 27587 1827
rect 27547 1797 27587 1805
rect 28860 1849 28900 1857
rect 28860 1827 28868 1849
rect 28892 1827 28900 1849
rect 25053 1752 25088 1753
rect 25030 1747 25088 1752
rect 25030 1727 25033 1747
rect 25053 1733 25088 1747
rect 25108 1733 25117 1753
rect 25053 1725 25117 1733
rect 25079 1724 25117 1725
rect 25080 1723 25117 1724
rect 25183 1757 25219 1758
rect 25291 1757 25327 1758
rect 25183 1749 25327 1757
rect 25183 1729 25191 1749
rect 25211 1745 25299 1749
rect 25211 1729 25255 1745
rect 25183 1725 25255 1729
rect 25275 1729 25299 1745
rect 25319 1729 25327 1749
rect 25275 1725 25327 1729
rect 25183 1723 25327 1725
rect 25393 1753 25431 1761
rect 25509 1757 25545 1758
rect 25393 1733 25402 1753
rect 25422 1733 25431 1753
rect 25393 1724 25431 1733
rect 25460 1749 25545 1757
rect 25460 1729 25517 1749
rect 25537 1729 25545 1749
rect 25393 1723 25430 1724
rect 25460 1723 25545 1729
rect 25611 1753 25649 1761
rect 25611 1733 25620 1753
rect 25640 1733 25649 1753
rect 25611 1724 25649 1733
rect 25793 1758 25835 1767
rect 25793 1740 25807 1758
rect 25825 1740 25835 1758
rect 25793 1732 25835 1740
rect 25798 1730 25835 1732
rect 26238 1751 26681 1790
rect 25611 1723 25648 1724
rect 25072 1695 25162 1701
rect 25072 1675 25088 1695
rect 25108 1693 25162 1695
rect 25108 1675 25133 1693
rect 25072 1673 25133 1675
rect 25153 1673 25162 1693
rect 25072 1667 25162 1673
rect 25085 1613 25122 1614
rect 25181 1613 25218 1614
rect 25237 1613 25273 1723
rect 25460 1702 25491 1723
rect 26238 1708 26285 1751
rect 26641 1746 26681 1751
rect 27306 1749 27493 1773
rect 27524 1754 27917 1774
rect 27937 1754 27940 1774
rect 27524 1749 27940 1754
rect 25456 1701 25491 1702
rect 25334 1691 25491 1701
rect 25334 1671 25351 1691
rect 25371 1671 25491 1691
rect 25334 1664 25491 1671
rect 25558 1694 25707 1702
rect 25558 1674 25569 1694
rect 25589 1674 25628 1694
rect 25648 1674 25707 1694
rect 26238 1690 26248 1708
rect 26266 1690 26285 1708
rect 26238 1686 26285 1690
rect 26239 1681 26276 1686
rect 25558 1667 25707 1674
rect 27306 1678 27343 1749
rect 27524 1748 27865 1749
rect 27458 1688 27489 1689
rect 25558 1666 25599 1667
rect 25795 1665 25832 1668
rect 25292 1613 25329 1614
rect 24985 1604 25123 1613
rect 24189 1565 24633 1591
rect 24189 1563 24357 1565
rect 23142 1431 23589 1443
rect 23185 1429 23218 1431
rect 22552 1411 22690 1420
rect 22346 1410 22383 1411
rect 22076 1357 22117 1358
rect 21850 1336 21902 1354
rect 21968 1350 22117 1357
rect 21418 1316 21458 1326
rect 21968 1330 22027 1350
rect 22047 1330 22086 1350
rect 22106 1330 22117 1350
rect 21968 1322 22117 1330
rect 22184 1353 22341 1360
rect 22184 1333 22304 1353
rect 22324 1333 22341 1353
rect 22184 1323 22341 1333
rect 22184 1322 22219 1323
rect 21248 1299 21286 1308
rect 22184 1301 22215 1322
rect 22402 1301 22438 1411
rect 22457 1410 22494 1411
rect 22553 1410 22590 1411
rect 22513 1351 22603 1357
rect 22513 1331 22522 1351
rect 22542 1349 22603 1351
rect 22542 1331 22567 1349
rect 22513 1329 22567 1331
rect 22587 1329 22603 1349
rect 22513 1323 22603 1329
rect 22027 1300 22064 1301
rect 21248 1298 21285 1299
rect 20709 1270 20799 1276
rect 20709 1250 20725 1270
rect 20745 1268 20799 1270
rect 20745 1250 20770 1268
rect 20709 1248 20770 1250
rect 20790 1248 20799 1268
rect 20709 1242 20799 1248
rect 20722 1188 20759 1189
rect 20818 1188 20855 1189
rect 20874 1188 20910 1298
rect 21097 1277 21128 1298
rect 22026 1291 22064 1300
rect 21093 1276 21128 1277
rect 20971 1266 21128 1276
rect 20971 1246 20988 1266
rect 21008 1246 21128 1266
rect 20971 1239 21128 1246
rect 21195 1269 21344 1277
rect 21195 1249 21206 1269
rect 21226 1249 21265 1269
rect 21285 1249 21344 1269
rect 21854 1273 21894 1283
rect 21195 1242 21344 1249
rect 21410 1245 21462 1263
rect 21195 1241 21236 1242
rect 20929 1188 20966 1189
rect 20622 1179 20760 1188
rect 20622 1159 20731 1179
rect 20751 1159 20760 1179
rect 20622 1152 20760 1159
rect 20818 1179 20966 1188
rect 20818 1159 20827 1179
rect 20847 1159 20937 1179
rect 20957 1159 20966 1179
rect 20622 1150 20718 1152
rect 20818 1149 20966 1159
rect 21025 1179 21062 1189
rect 21025 1159 21033 1179
rect 21053 1159 21062 1179
rect 20874 1148 20910 1149
rect 21025 1092 21062 1159
rect 21097 1188 21128 1239
rect 21410 1227 21428 1245
rect 21446 1227 21462 1245
rect 21147 1188 21184 1189
rect 21097 1179 21184 1188
rect 21097 1159 21155 1179
rect 21175 1159 21184 1179
rect 21097 1149 21184 1159
rect 21243 1179 21280 1189
rect 21243 1159 21251 1179
rect 21271 1159 21280 1179
rect 21097 1148 21128 1149
rect 20722 1089 20759 1090
rect 21025 1089 21064 1092
rect 20721 1088 21064 1089
rect 21243 1088 21280 1159
rect 20646 1083 21064 1088
rect 20646 1063 20649 1083
rect 20669 1063 21064 1083
rect 21093 1064 21280 1088
rect 19187 1032 19224 1040
rect 19187 1013 19195 1032
rect 19216 1013 19224 1032
rect 19187 1007 19224 1013
rect 21025 1038 21064 1063
rect 21410 1038 21462 1227
rect 21854 1255 21864 1273
rect 21882 1255 21894 1273
rect 22026 1271 22035 1291
rect 22055 1271 22064 1291
rect 22026 1263 22064 1271
rect 22130 1295 22215 1301
rect 22245 1300 22282 1301
rect 22130 1275 22138 1295
rect 22158 1275 22215 1295
rect 22130 1267 22215 1275
rect 22244 1291 22282 1300
rect 22244 1271 22253 1291
rect 22273 1271 22282 1291
rect 22130 1266 22166 1267
rect 22244 1263 22282 1271
rect 22348 1295 22492 1301
rect 22348 1275 22356 1295
rect 22376 1275 22409 1295
rect 22429 1275 22464 1295
rect 22484 1275 22492 1295
rect 22348 1267 22492 1275
rect 22348 1266 22384 1267
rect 22456 1266 22492 1267
rect 22558 1300 22595 1301
rect 22558 1299 22596 1300
rect 22558 1291 22622 1299
rect 22558 1271 22567 1291
rect 22587 1277 22622 1291
rect 22642 1277 22645 1297
rect 22587 1272 22645 1277
rect 22587 1271 22622 1272
rect 21854 1199 21894 1255
rect 22027 1234 22064 1263
rect 22028 1232 22064 1234
rect 22028 1210 22219 1232
rect 22245 1231 22282 1263
rect 22558 1259 22622 1271
rect 22662 1233 22689 1411
rect 23547 1386 23589 1431
rect 22521 1231 22689 1233
rect 22245 1221 22689 1231
rect 22830 1327 23017 1351
rect 23048 1332 23441 1352
rect 23461 1332 23464 1352
rect 23048 1327 23464 1332
rect 22830 1256 22867 1327
rect 23048 1326 23389 1327
rect 22982 1266 23013 1267
rect 22830 1236 22839 1256
rect 22859 1236 22867 1256
rect 22830 1226 22867 1236
rect 22926 1256 23013 1266
rect 22926 1236 22935 1256
rect 22955 1236 23013 1256
rect 22926 1227 23013 1236
rect 22926 1226 22963 1227
rect 21851 1194 21894 1199
rect 22242 1205 22689 1221
rect 22242 1199 22270 1205
rect 22521 1204 22689 1205
rect 21851 1191 22001 1194
rect 22242 1191 22269 1199
rect 21851 1189 22269 1191
rect 21851 1171 21860 1189
rect 21878 1171 22269 1189
rect 22982 1176 23013 1227
rect 23048 1256 23085 1326
rect 23351 1325 23388 1326
rect 23200 1266 23236 1267
rect 23048 1236 23057 1256
rect 23077 1236 23085 1256
rect 23048 1226 23085 1236
rect 23144 1256 23292 1266
rect 23392 1263 23488 1265
rect 23144 1236 23153 1256
rect 23173 1236 23263 1256
rect 23283 1236 23292 1256
rect 23144 1227 23292 1236
rect 23350 1256 23488 1263
rect 23350 1236 23359 1256
rect 23379 1236 23488 1256
rect 23350 1227 23488 1236
rect 23144 1226 23181 1227
rect 22874 1173 22915 1174
rect 21851 1168 22269 1171
rect 21851 1162 21894 1168
rect 21854 1159 21894 1162
rect 22769 1166 22915 1173
rect 22251 1150 22291 1151
rect 21962 1133 22291 1150
rect 22769 1146 22825 1166
rect 22845 1146 22884 1166
rect 22904 1146 22915 1166
rect 22769 1138 22915 1146
rect 22982 1169 23139 1176
rect 22982 1149 23102 1169
rect 23122 1149 23139 1169
rect 22982 1139 23139 1149
rect 22982 1138 23017 1139
rect 21846 1090 21889 1101
rect 21846 1072 21858 1090
rect 21876 1072 21889 1090
rect 21846 1046 21889 1072
rect 21962 1046 21989 1133
rect 22251 1124 22291 1133
rect 21025 1020 21464 1038
rect 21025 1002 21425 1020
rect 21443 1002 21464 1020
rect 21025 996 21464 1002
rect 21031 992 21464 996
rect 21846 1025 21989 1046
rect 22033 1098 22067 1114
rect 22251 1104 22644 1124
rect 22664 1104 22667 1124
rect 22982 1117 23013 1138
rect 23200 1117 23236 1227
rect 23255 1226 23292 1227
rect 23351 1226 23388 1227
rect 23311 1167 23401 1173
rect 23311 1147 23320 1167
rect 23340 1165 23401 1167
rect 23340 1147 23365 1165
rect 23311 1145 23365 1147
rect 23385 1145 23401 1165
rect 23311 1139 23401 1145
rect 22825 1116 22862 1117
rect 22251 1099 22667 1104
rect 22824 1107 22862 1116
rect 22251 1098 22592 1099
rect 22033 1028 22070 1098
rect 22185 1038 22216 1039
rect 21846 1023 21983 1025
rect 21410 990 21462 992
rect 21846 981 21889 1023
rect 22033 1008 22042 1028
rect 22062 1008 22070 1028
rect 22033 998 22070 1008
rect 22129 1028 22216 1038
rect 22129 1008 22138 1028
rect 22158 1008 22216 1028
rect 22129 999 22216 1008
rect 22129 998 22166 999
rect 21844 971 21889 981
rect 21844 953 21853 971
rect 21871 953 21889 971
rect 21844 947 21889 953
rect 22185 948 22216 999
rect 22251 1028 22288 1098
rect 22554 1097 22591 1098
rect 22824 1087 22833 1107
rect 22853 1087 22862 1107
rect 22824 1079 22862 1087
rect 22928 1111 23013 1117
rect 23043 1116 23080 1117
rect 22928 1091 22936 1111
rect 22956 1091 23013 1111
rect 22928 1083 23013 1091
rect 23042 1107 23080 1116
rect 23042 1087 23051 1107
rect 23071 1087 23080 1107
rect 22928 1082 22964 1083
rect 23042 1079 23080 1087
rect 23146 1111 23290 1117
rect 23146 1091 23154 1111
rect 23174 1108 23262 1111
rect 23174 1091 23209 1108
rect 23146 1090 23209 1091
rect 23228 1091 23262 1108
rect 23282 1091 23290 1111
rect 23228 1090 23290 1091
rect 23146 1083 23290 1090
rect 23146 1082 23182 1083
rect 23254 1082 23290 1083
rect 23356 1116 23393 1117
rect 23356 1115 23394 1116
rect 23416 1115 23443 1119
rect 23356 1113 23443 1115
rect 23356 1107 23420 1113
rect 23356 1087 23365 1107
rect 23385 1093 23420 1107
rect 23440 1093 23443 1113
rect 23385 1088 23443 1093
rect 23385 1087 23420 1088
rect 22825 1050 22862 1079
rect 22826 1048 22862 1050
rect 22403 1038 22439 1039
rect 22251 1008 22260 1028
rect 22280 1008 22288 1028
rect 22251 998 22288 1008
rect 22347 1028 22495 1038
rect 22595 1035 22691 1037
rect 22347 1008 22356 1028
rect 22376 1008 22466 1028
rect 22486 1008 22495 1028
rect 22347 999 22495 1008
rect 22553 1028 22691 1035
rect 22553 1008 22562 1028
rect 22582 1008 22691 1028
rect 22826 1026 23017 1048
rect 23043 1047 23080 1079
rect 23356 1075 23420 1087
rect 23460 1049 23487 1227
rect 23319 1047 23487 1049
rect 23043 1021 23487 1047
rect 22553 999 22691 1008
rect 22347 998 22384 999
rect 21844 944 21881 947
rect 22077 945 22118 946
rect 21969 938 22118 945
rect 21413 925 21450 930
rect 21404 921 21451 925
rect 21404 903 21423 921
rect 21441 903 21451 921
rect 21969 918 22028 938
rect 22048 918 22087 938
rect 22107 918 22118 938
rect 21969 910 22118 918
rect 22185 941 22342 948
rect 22185 921 22305 941
rect 22325 921 22342 941
rect 22185 911 22342 921
rect 22185 910 22220 911
rect 21404 840 21451 903
rect 22185 889 22216 910
rect 22403 889 22439 999
rect 22458 998 22495 999
rect 22554 998 22591 999
rect 22514 939 22604 945
rect 22514 919 22523 939
rect 22543 937 22604 939
rect 22543 919 22568 937
rect 22514 917 22568 919
rect 22588 917 22604 937
rect 22514 911 22604 917
rect 22028 888 22065 889
rect 21841 880 21878 882
rect 21841 872 21883 880
rect 21841 854 21851 872
rect 21869 854 21883 872
rect 21841 845 21883 854
rect 22027 879 22065 888
rect 22027 859 22036 879
rect 22056 859 22065 879
rect 22027 851 22065 859
rect 22131 883 22216 889
rect 22246 888 22283 889
rect 22131 863 22139 883
rect 22159 863 22216 883
rect 22131 855 22216 863
rect 22245 879 22283 888
rect 22245 859 22254 879
rect 22274 859 22283 879
rect 22131 854 22167 855
rect 22245 851 22283 859
rect 22349 887 22493 889
rect 22349 883 22401 887
rect 22349 863 22357 883
rect 22377 867 22401 883
rect 22421 883 22493 887
rect 22421 867 22465 883
rect 22377 863 22465 867
rect 22485 863 22493 883
rect 22349 855 22493 863
rect 22349 854 22385 855
rect 22457 854 22493 855
rect 22559 888 22596 889
rect 22559 887 22597 888
rect 22559 879 22623 887
rect 22559 859 22568 879
rect 22588 865 22623 879
rect 22643 865 22646 885
rect 22588 860 22646 865
rect 22588 859 22623 860
rect 21404 825 21454 840
rect 21404 800 21418 825
rect 21450 800 21454 825
rect 21842 820 21883 845
rect 22028 820 22065 851
rect 22246 829 22283 851
rect 22559 847 22623 859
rect 22241 820 22283 829
rect 22663 821 22690 999
rect 21842 808 21887 820
rect 21404 787 21451 800
rect 18789 762 18797 784
rect 18821 762 18829 784
rect 18789 754 18829 762
rect 21838 750 21887 808
rect 22028 794 22090 820
rect 22241 819 22326 820
rect 22522 819 22690 821
rect 22241 793 22690 819
rect 22241 750 22280 793
rect 22522 792 22690 793
rect 23153 797 23193 1021
rect 23319 1020 23487 1021
rect 23551 1053 23584 1386
rect 24189 1385 24216 1563
rect 24256 1525 24320 1537
rect 24596 1533 24633 1565
rect 24659 1564 24850 1586
rect 24985 1584 25094 1604
rect 25114 1584 25123 1604
rect 24985 1577 25123 1584
rect 25181 1604 25329 1613
rect 25181 1584 25190 1604
rect 25210 1584 25300 1604
rect 25320 1584 25329 1604
rect 24985 1575 25081 1577
rect 25181 1574 25329 1584
rect 25388 1604 25425 1614
rect 25388 1584 25396 1604
rect 25416 1584 25425 1604
rect 25237 1573 25273 1574
rect 24814 1562 24850 1564
rect 24814 1533 24851 1562
rect 24256 1524 24291 1525
rect 24233 1519 24291 1524
rect 24233 1499 24236 1519
rect 24256 1505 24291 1519
rect 24311 1505 24320 1525
rect 24256 1497 24320 1505
rect 24282 1496 24320 1497
rect 24283 1495 24320 1496
rect 24386 1529 24422 1530
rect 24494 1529 24530 1530
rect 24386 1521 24530 1529
rect 24386 1501 24394 1521
rect 24414 1520 24502 1521
rect 24414 1501 24449 1520
rect 24470 1501 24502 1520
rect 24522 1501 24530 1521
rect 24386 1495 24530 1501
rect 24596 1525 24634 1533
rect 24712 1529 24748 1530
rect 24596 1505 24605 1525
rect 24625 1505 24634 1525
rect 24596 1496 24634 1505
rect 24663 1521 24748 1529
rect 24663 1501 24720 1521
rect 24740 1501 24748 1521
rect 24596 1495 24633 1496
rect 24663 1495 24748 1501
rect 24814 1525 24852 1533
rect 24814 1505 24823 1525
rect 24843 1505 24852 1525
rect 25085 1514 25122 1515
rect 25388 1514 25425 1584
rect 25460 1613 25491 1664
rect 25787 1659 25832 1665
rect 25787 1641 25805 1659
rect 25823 1641 25832 1659
rect 27306 1658 27315 1678
rect 27335 1658 27343 1678
rect 27306 1648 27343 1658
rect 27402 1678 27489 1688
rect 27402 1658 27411 1678
rect 27431 1658 27489 1678
rect 27402 1649 27489 1658
rect 27402 1648 27439 1649
rect 25787 1631 25832 1641
rect 25510 1613 25547 1614
rect 25460 1604 25547 1613
rect 25460 1584 25518 1604
rect 25538 1584 25547 1604
rect 25460 1574 25547 1584
rect 25606 1604 25643 1614
rect 25606 1584 25614 1604
rect 25634 1584 25643 1604
rect 25787 1589 25830 1631
rect 26227 1619 26279 1621
rect 25693 1587 25830 1589
rect 25460 1573 25491 1574
rect 25606 1514 25643 1584
rect 25084 1513 25425 1514
rect 24814 1496 24852 1505
rect 25009 1508 25425 1513
rect 24814 1495 24851 1496
rect 24275 1467 24365 1473
rect 24275 1447 24291 1467
rect 24311 1465 24365 1467
rect 24311 1447 24336 1465
rect 24275 1445 24336 1447
rect 24356 1445 24365 1465
rect 24275 1439 24365 1445
rect 24288 1385 24325 1386
rect 24384 1385 24421 1386
rect 24440 1385 24476 1495
rect 24663 1474 24694 1495
rect 25009 1488 25012 1508
rect 25032 1488 25425 1508
rect 25609 1498 25643 1514
rect 25687 1566 25830 1587
rect 26225 1615 26658 1619
rect 26225 1609 26664 1615
rect 26225 1591 26246 1609
rect 26264 1591 26664 1609
rect 27458 1598 27489 1649
rect 27524 1678 27561 1748
rect 27827 1747 27864 1748
rect 27676 1688 27712 1689
rect 27524 1658 27533 1678
rect 27553 1658 27561 1678
rect 27524 1648 27561 1658
rect 27620 1678 27768 1688
rect 27868 1685 27964 1687
rect 27620 1658 27629 1678
rect 27649 1658 27739 1678
rect 27759 1658 27768 1678
rect 27620 1649 27768 1658
rect 27826 1678 27964 1685
rect 27826 1658 27835 1678
rect 27855 1658 27964 1678
rect 27826 1649 27964 1658
rect 27620 1648 27657 1649
rect 27350 1595 27391 1596
rect 26225 1573 26664 1591
rect 25385 1479 25425 1488
rect 25687 1479 25714 1566
rect 25787 1540 25830 1566
rect 25787 1522 25800 1540
rect 25818 1522 25830 1540
rect 25787 1511 25830 1522
rect 24659 1473 24694 1474
rect 24537 1463 24694 1473
rect 24537 1443 24554 1463
rect 24574 1443 24694 1463
rect 24537 1436 24694 1443
rect 24761 1466 24910 1474
rect 24761 1446 24772 1466
rect 24792 1446 24831 1466
rect 24851 1446 24910 1466
rect 25385 1462 25714 1479
rect 25385 1461 25425 1462
rect 24761 1439 24910 1446
rect 25782 1450 25822 1453
rect 25782 1444 25825 1450
rect 25407 1441 25825 1444
rect 24761 1438 24802 1439
rect 24495 1385 24532 1386
rect 24188 1376 24326 1385
rect 24188 1356 24297 1376
rect 24317 1356 24326 1376
rect 24188 1349 24326 1356
rect 24384 1376 24532 1385
rect 24384 1356 24393 1376
rect 24413 1356 24503 1376
rect 24523 1356 24532 1376
rect 24188 1347 24284 1349
rect 24384 1346 24532 1356
rect 24591 1376 24628 1386
rect 24591 1356 24599 1376
rect 24619 1356 24628 1376
rect 24440 1345 24476 1346
rect 24288 1286 24325 1287
rect 24591 1286 24628 1356
rect 24663 1385 24694 1436
rect 25407 1423 25798 1441
rect 25816 1423 25825 1441
rect 25407 1421 25825 1423
rect 25407 1413 25434 1421
rect 25675 1418 25825 1421
rect 24987 1407 25155 1408
rect 25406 1407 25434 1413
rect 24987 1391 25434 1407
rect 25782 1413 25825 1418
rect 24713 1385 24750 1386
rect 24663 1376 24750 1385
rect 24663 1356 24721 1376
rect 24741 1356 24750 1376
rect 24663 1346 24750 1356
rect 24809 1376 24846 1386
rect 24809 1356 24817 1376
rect 24837 1356 24846 1376
rect 24663 1345 24694 1346
rect 24287 1285 24628 1286
rect 24809 1285 24846 1356
rect 24212 1280 24628 1285
rect 24212 1260 24215 1280
rect 24235 1260 24628 1280
rect 24659 1261 24846 1285
rect 24987 1381 25431 1391
rect 24987 1379 25155 1381
rect 24987 1201 25014 1379
rect 25054 1341 25118 1353
rect 25394 1349 25431 1381
rect 25457 1380 25648 1402
rect 25612 1378 25648 1380
rect 25612 1349 25649 1378
rect 25782 1357 25822 1413
rect 25054 1340 25089 1341
rect 25031 1335 25089 1340
rect 25031 1315 25034 1335
rect 25054 1321 25089 1335
rect 25109 1321 25118 1341
rect 25054 1313 25118 1321
rect 25080 1312 25118 1313
rect 25081 1311 25118 1312
rect 25184 1345 25220 1346
rect 25292 1345 25328 1346
rect 25184 1337 25328 1345
rect 25184 1317 25192 1337
rect 25212 1317 25247 1337
rect 25267 1317 25300 1337
rect 25320 1317 25328 1337
rect 25184 1311 25328 1317
rect 25394 1341 25432 1349
rect 25510 1345 25546 1346
rect 25394 1321 25403 1341
rect 25423 1321 25432 1341
rect 25394 1312 25432 1321
rect 25461 1337 25546 1345
rect 25461 1317 25518 1337
rect 25538 1317 25546 1337
rect 25394 1311 25431 1312
rect 25461 1311 25546 1317
rect 25612 1341 25650 1349
rect 25612 1321 25621 1341
rect 25641 1321 25650 1341
rect 25782 1339 25794 1357
rect 25812 1339 25822 1357
rect 26227 1384 26279 1573
rect 26625 1548 26664 1573
rect 27242 1588 27391 1595
rect 27242 1568 27301 1588
rect 27321 1568 27360 1588
rect 27380 1568 27391 1588
rect 27242 1560 27391 1568
rect 27458 1591 27615 1598
rect 27458 1571 27578 1591
rect 27598 1571 27615 1591
rect 27458 1561 27615 1571
rect 27458 1560 27493 1561
rect 26409 1523 26596 1547
rect 26625 1528 27020 1548
rect 27040 1528 27043 1548
rect 27458 1539 27489 1560
rect 27676 1539 27712 1649
rect 27731 1648 27768 1649
rect 27827 1648 27864 1649
rect 27787 1589 27877 1595
rect 27787 1569 27796 1589
rect 27816 1587 27877 1589
rect 27816 1569 27841 1587
rect 27787 1567 27841 1569
rect 27861 1567 27877 1587
rect 27787 1561 27877 1567
rect 27301 1538 27338 1539
rect 26625 1523 27043 1528
rect 27300 1529 27338 1538
rect 26409 1452 26446 1523
rect 26625 1522 26968 1523
rect 26625 1519 26664 1522
rect 26930 1521 26967 1522
rect 26561 1462 26592 1463
rect 26409 1432 26418 1452
rect 26438 1432 26446 1452
rect 26409 1422 26446 1432
rect 26505 1452 26592 1462
rect 26505 1432 26514 1452
rect 26534 1432 26592 1452
rect 26505 1423 26592 1432
rect 26505 1422 26542 1423
rect 26227 1366 26243 1384
rect 26261 1366 26279 1384
rect 26561 1372 26592 1423
rect 26627 1452 26664 1519
rect 27300 1509 27309 1529
rect 27329 1509 27338 1529
rect 27300 1501 27338 1509
rect 27404 1533 27489 1539
rect 27519 1538 27556 1539
rect 27404 1513 27412 1533
rect 27432 1513 27489 1533
rect 27404 1505 27489 1513
rect 27518 1529 27556 1538
rect 27518 1509 27527 1529
rect 27547 1509 27556 1529
rect 27404 1504 27440 1505
rect 27518 1501 27556 1509
rect 27622 1533 27766 1539
rect 27622 1513 27630 1533
rect 27650 1528 27738 1533
rect 27650 1513 27686 1528
rect 27622 1511 27686 1513
rect 27705 1513 27738 1528
rect 27758 1513 27766 1533
rect 27705 1511 27766 1513
rect 27622 1505 27766 1511
rect 27622 1504 27658 1505
rect 27730 1504 27766 1505
rect 27832 1538 27869 1539
rect 27832 1537 27870 1538
rect 27832 1529 27896 1537
rect 27832 1509 27841 1529
rect 27861 1515 27896 1529
rect 27916 1515 27919 1535
rect 27861 1510 27919 1515
rect 27861 1509 27896 1510
rect 27301 1472 27338 1501
rect 27302 1470 27338 1472
rect 26779 1462 26815 1463
rect 26627 1432 26636 1452
rect 26656 1432 26664 1452
rect 26627 1422 26664 1432
rect 26723 1452 26871 1462
rect 26971 1459 27067 1461
rect 26723 1432 26732 1452
rect 26752 1432 26842 1452
rect 26862 1432 26871 1452
rect 26723 1423 26871 1432
rect 26929 1452 27067 1459
rect 26929 1432 26938 1452
rect 26958 1432 27067 1452
rect 27302 1448 27493 1470
rect 27519 1469 27556 1501
rect 27832 1497 27896 1509
rect 27936 1471 27963 1649
rect 27795 1469 27963 1471
rect 27519 1455 27963 1469
rect 28566 1603 28734 1604
rect 28860 1603 28900 1827
rect 29363 1831 29531 1832
rect 29766 1831 29806 1864
rect 30162 1831 30209 1864
rect 30600 1863 30641 1888
rect 30786 1863 30823 1894
rect 31004 1863 31041 1894
rect 31317 1890 31381 1902
rect 31421 1864 31448 2042
rect 30600 1836 30649 1863
rect 30785 1837 30834 1863
rect 31003 1862 31084 1863
rect 31280 1862 31448 1864
rect 31003 1837 31448 1862
rect 31004 1836 31448 1837
rect 29363 1830 29807 1831
rect 29363 1805 29808 1830
rect 29363 1803 29531 1805
rect 29727 1804 29808 1805
rect 29977 1804 30026 1830
rect 30162 1804 30211 1831
rect 29363 1625 29390 1803
rect 29430 1765 29494 1777
rect 29770 1773 29807 1804
rect 29988 1773 30025 1804
rect 30170 1779 30211 1804
rect 30602 1803 30649 1836
rect 31005 1803 31045 1836
rect 31280 1835 31448 1836
rect 31911 1840 31951 2064
rect 32077 2063 32245 2064
rect 32848 2198 33292 2212
rect 32848 2196 33016 2198
rect 32848 2018 32875 2196
rect 32915 2158 32979 2170
rect 33255 2166 33292 2198
rect 33318 2197 33509 2219
rect 33744 2215 33853 2235
rect 33873 2215 33882 2235
rect 33744 2208 33882 2215
rect 33940 2235 34088 2244
rect 33940 2215 33949 2235
rect 33969 2215 34059 2235
rect 34079 2215 34088 2235
rect 33744 2206 33840 2208
rect 33940 2205 34088 2215
rect 34147 2235 34184 2245
rect 34147 2215 34155 2235
rect 34175 2215 34184 2235
rect 33996 2204 34032 2205
rect 33473 2195 33509 2197
rect 33473 2166 33510 2195
rect 32915 2157 32950 2158
rect 32892 2152 32950 2157
rect 32892 2132 32895 2152
rect 32915 2138 32950 2152
rect 32970 2138 32979 2158
rect 32915 2130 32979 2138
rect 32941 2129 32979 2130
rect 32942 2128 32979 2129
rect 33045 2162 33081 2163
rect 33153 2162 33189 2163
rect 33045 2154 33189 2162
rect 33045 2134 33053 2154
rect 33073 2152 33161 2154
rect 33073 2134 33106 2152
rect 33045 2133 33106 2134
rect 33127 2134 33161 2152
rect 33181 2134 33189 2154
rect 33127 2133 33189 2134
rect 33045 2128 33189 2133
rect 33255 2158 33293 2166
rect 33371 2162 33407 2163
rect 33255 2138 33264 2158
rect 33284 2138 33293 2158
rect 33255 2129 33293 2138
rect 33322 2154 33407 2162
rect 33322 2134 33379 2154
rect 33399 2134 33407 2154
rect 33255 2128 33292 2129
rect 33322 2128 33407 2134
rect 33473 2158 33511 2166
rect 33473 2138 33482 2158
rect 33502 2138 33511 2158
rect 34147 2148 34184 2215
rect 34219 2244 34250 2295
rect 34532 2283 34550 2301
rect 34568 2283 34584 2301
rect 34269 2244 34306 2245
rect 34219 2235 34306 2244
rect 34219 2215 34277 2235
rect 34297 2215 34306 2235
rect 34219 2205 34306 2215
rect 34365 2235 34402 2245
rect 34365 2215 34373 2235
rect 34393 2215 34402 2235
rect 34219 2204 34250 2205
rect 33844 2145 33881 2146
rect 34147 2145 34186 2148
rect 33843 2144 34186 2145
rect 34365 2144 34402 2215
rect 33473 2129 33511 2138
rect 33768 2139 34186 2144
rect 33473 2128 33510 2129
rect 32934 2100 33024 2106
rect 32934 2080 32950 2100
rect 32970 2098 33024 2100
rect 32970 2080 32995 2098
rect 32934 2078 32995 2080
rect 33015 2078 33024 2098
rect 32934 2072 33024 2078
rect 32947 2018 32984 2019
rect 33043 2018 33080 2019
rect 33099 2018 33135 2128
rect 33322 2107 33353 2128
rect 33768 2119 33771 2139
rect 33791 2119 34186 2139
rect 34215 2120 34402 2144
rect 33318 2106 33353 2107
rect 33196 2096 33353 2106
rect 33196 2076 33213 2096
rect 33233 2076 33353 2096
rect 33196 2069 33353 2076
rect 33420 2099 33569 2107
rect 33420 2079 33431 2099
rect 33451 2079 33490 2099
rect 33510 2079 33569 2099
rect 33420 2072 33569 2079
rect 34147 2094 34186 2119
rect 34532 2094 34584 2283
rect 34147 2076 34586 2094
rect 33420 2071 33461 2072
rect 33154 2018 33191 2019
rect 32847 2009 32985 2018
rect 32847 1989 32956 2009
rect 32976 1989 32985 2009
rect 32847 1982 32985 1989
rect 33043 2009 33191 2018
rect 33043 1989 33052 2009
rect 33072 1989 33162 2009
rect 33182 1989 33191 2009
rect 32847 1980 32943 1982
rect 33043 1979 33191 1989
rect 33250 2009 33287 2019
rect 33250 1989 33258 2009
rect 33278 1989 33287 2009
rect 33099 1978 33135 1979
rect 32947 1919 32984 1920
rect 33250 1919 33287 1989
rect 33322 2018 33353 2069
rect 34147 2058 34547 2076
rect 34565 2058 34586 2076
rect 34147 2052 34586 2058
rect 34153 2048 34586 2052
rect 34532 2046 34584 2048
rect 33372 2018 33409 2019
rect 33322 2009 33409 2018
rect 33322 1989 33380 2009
rect 33400 1989 33409 2009
rect 33322 1979 33409 1989
rect 33468 2009 33505 2019
rect 33468 1989 33476 2009
rect 33496 1989 33505 2009
rect 33322 1978 33353 1979
rect 32946 1918 33287 1919
rect 33468 1918 33505 1989
rect 34535 1981 34572 1986
rect 34526 1977 34573 1981
rect 34526 1959 34545 1977
rect 34563 1959 34573 1977
rect 32871 1913 33287 1918
rect 32871 1893 32874 1913
rect 32894 1893 33287 1913
rect 33318 1894 33505 1918
rect 34130 1916 34170 1921
rect 34526 1916 34573 1959
rect 34130 1877 34573 1916
rect 31911 1818 31919 1840
rect 31943 1818 31951 1840
rect 31911 1810 31951 1818
rect 33224 1862 33264 1870
rect 33224 1840 33232 1862
rect 33256 1840 33264 1862
rect 29430 1764 29465 1765
rect 29407 1759 29465 1764
rect 29407 1739 29410 1759
rect 29430 1745 29465 1759
rect 29485 1745 29494 1765
rect 29430 1737 29494 1745
rect 29456 1736 29494 1737
rect 29457 1735 29494 1736
rect 29560 1769 29596 1770
rect 29668 1769 29704 1770
rect 29560 1761 29704 1769
rect 29560 1741 29568 1761
rect 29588 1757 29676 1761
rect 29588 1741 29632 1757
rect 29560 1737 29632 1741
rect 29652 1741 29676 1757
rect 29696 1741 29704 1761
rect 29652 1737 29704 1741
rect 29560 1735 29704 1737
rect 29770 1765 29808 1773
rect 29886 1769 29922 1770
rect 29770 1745 29779 1765
rect 29799 1745 29808 1765
rect 29770 1736 29808 1745
rect 29837 1761 29922 1769
rect 29837 1741 29894 1761
rect 29914 1741 29922 1761
rect 29770 1735 29807 1736
rect 29837 1735 29922 1741
rect 29988 1765 30026 1773
rect 29988 1745 29997 1765
rect 30017 1745 30026 1765
rect 29988 1736 30026 1745
rect 30170 1770 30212 1779
rect 30170 1752 30184 1770
rect 30202 1752 30212 1770
rect 30170 1744 30212 1752
rect 30175 1742 30212 1744
rect 30602 1764 31045 1803
rect 29988 1735 30025 1736
rect 29449 1707 29539 1713
rect 29449 1687 29465 1707
rect 29485 1705 29539 1707
rect 29485 1687 29510 1705
rect 29449 1685 29510 1687
rect 29530 1685 29539 1705
rect 29449 1679 29539 1685
rect 29462 1625 29499 1626
rect 29558 1625 29595 1626
rect 29614 1625 29650 1735
rect 29837 1714 29868 1735
rect 30602 1721 30649 1764
rect 31005 1759 31045 1764
rect 31670 1762 31857 1786
rect 31888 1767 32281 1787
rect 32301 1767 32304 1787
rect 31888 1762 32304 1767
rect 29833 1713 29868 1714
rect 29711 1703 29868 1713
rect 29711 1683 29728 1703
rect 29748 1683 29868 1703
rect 29711 1676 29868 1683
rect 29935 1706 30084 1714
rect 29935 1686 29946 1706
rect 29966 1686 30005 1706
rect 30025 1686 30084 1706
rect 30602 1703 30612 1721
rect 30630 1703 30649 1721
rect 30602 1699 30649 1703
rect 30603 1694 30640 1699
rect 29935 1679 30084 1686
rect 31670 1691 31707 1762
rect 31888 1761 32229 1762
rect 31822 1701 31853 1702
rect 29935 1678 29976 1679
rect 30172 1677 30209 1680
rect 29669 1625 29706 1626
rect 29362 1616 29500 1625
rect 28566 1577 29010 1603
rect 28566 1575 28734 1577
rect 27519 1443 27966 1455
rect 27562 1441 27595 1443
rect 26929 1423 27067 1432
rect 26723 1422 26760 1423
rect 26453 1369 26494 1370
rect 26227 1348 26279 1366
rect 26345 1362 26494 1369
rect 25782 1329 25822 1339
rect 26345 1342 26404 1362
rect 26424 1342 26463 1362
rect 26483 1342 26494 1362
rect 26345 1334 26494 1342
rect 26561 1365 26718 1372
rect 26561 1345 26681 1365
rect 26701 1345 26718 1365
rect 26561 1335 26718 1345
rect 26561 1334 26596 1335
rect 25612 1312 25650 1321
rect 26561 1313 26592 1334
rect 26779 1313 26815 1423
rect 26834 1422 26871 1423
rect 26930 1422 26967 1423
rect 26890 1363 26980 1369
rect 26890 1343 26899 1363
rect 26919 1361 26980 1363
rect 26919 1343 26944 1361
rect 26890 1341 26944 1343
rect 26964 1341 26980 1361
rect 26890 1335 26980 1341
rect 26404 1312 26441 1313
rect 25612 1311 25649 1312
rect 25073 1283 25163 1289
rect 25073 1263 25089 1283
rect 25109 1281 25163 1283
rect 25109 1263 25134 1281
rect 25073 1261 25134 1263
rect 25154 1261 25163 1281
rect 25073 1255 25163 1261
rect 25086 1201 25123 1202
rect 25182 1201 25219 1202
rect 25238 1201 25274 1311
rect 25461 1290 25492 1311
rect 26403 1303 26441 1312
rect 25457 1289 25492 1290
rect 25335 1279 25492 1289
rect 25335 1259 25352 1279
rect 25372 1259 25492 1279
rect 25335 1252 25492 1259
rect 25559 1282 25708 1290
rect 25559 1262 25570 1282
rect 25590 1262 25629 1282
rect 25649 1262 25708 1282
rect 26231 1285 26271 1295
rect 25559 1255 25708 1262
rect 25774 1258 25826 1276
rect 25559 1254 25600 1255
rect 25293 1201 25330 1202
rect 24986 1192 25124 1201
rect 24986 1172 25095 1192
rect 25115 1172 25124 1192
rect 24986 1165 25124 1172
rect 25182 1192 25330 1201
rect 25182 1172 25191 1192
rect 25211 1172 25301 1192
rect 25321 1172 25330 1192
rect 24986 1163 25082 1165
rect 25182 1162 25330 1172
rect 25389 1192 25426 1202
rect 25389 1172 25397 1192
rect 25417 1172 25426 1192
rect 25238 1161 25274 1162
rect 25389 1105 25426 1172
rect 25461 1201 25492 1252
rect 25774 1240 25792 1258
rect 25810 1240 25826 1258
rect 25511 1201 25548 1202
rect 25461 1192 25548 1201
rect 25461 1172 25519 1192
rect 25539 1172 25548 1192
rect 25461 1162 25548 1172
rect 25607 1192 25644 1202
rect 25607 1172 25615 1192
rect 25635 1172 25644 1192
rect 25461 1161 25492 1162
rect 25086 1102 25123 1103
rect 25389 1102 25428 1105
rect 25085 1101 25428 1102
rect 25607 1101 25644 1172
rect 25010 1096 25428 1101
rect 25010 1076 25013 1096
rect 25033 1076 25428 1096
rect 25457 1077 25644 1101
rect 23551 1045 23588 1053
rect 23551 1026 23559 1045
rect 23580 1026 23588 1045
rect 23551 1020 23588 1026
rect 25389 1051 25428 1076
rect 25774 1051 25826 1240
rect 26231 1267 26241 1285
rect 26259 1267 26271 1285
rect 26403 1283 26412 1303
rect 26432 1283 26441 1303
rect 26403 1275 26441 1283
rect 26507 1307 26592 1313
rect 26622 1312 26659 1313
rect 26507 1287 26515 1307
rect 26535 1287 26592 1307
rect 26507 1279 26592 1287
rect 26621 1303 26659 1312
rect 26621 1283 26630 1303
rect 26650 1283 26659 1303
rect 26507 1278 26543 1279
rect 26621 1275 26659 1283
rect 26725 1307 26869 1313
rect 26725 1287 26733 1307
rect 26753 1287 26786 1307
rect 26806 1287 26841 1307
rect 26861 1287 26869 1307
rect 26725 1279 26869 1287
rect 26725 1278 26761 1279
rect 26833 1278 26869 1279
rect 26935 1312 26972 1313
rect 26935 1311 26973 1312
rect 26935 1303 26999 1311
rect 26935 1283 26944 1303
rect 26964 1289 26999 1303
rect 27019 1289 27022 1309
rect 26964 1284 27022 1289
rect 26964 1283 26999 1284
rect 26231 1211 26271 1267
rect 26404 1246 26441 1275
rect 26405 1244 26441 1246
rect 26405 1222 26596 1244
rect 26622 1243 26659 1275
rect 26935 1271 26999 1283
rect 27039 1245 27066 1423
rect 27924 1398 27966 1443
rect 26898 1243 27066 1245
rect 26622 1233 27066 1243
rect 27207 1339 27394 1363
rect 27425 1344 27818 1364
rect 27838 1344 27841 1364
rect 27425 1339 27841 1344
rect 27207 1268 27244 1339
rect 27425 1338 27766 1339
rect 27359 1278 27390 1279
rect 27207 1248 27216 1268
rect 27236 1248 27244 1268
rect 27207 1238 27244 1248
rect 27303 1268 27390 1278
rect 27303 1248 27312 1268
rect 27332 1248 27390 1268
rect 27303 1239 27390 1248
rect 27303 1238 27340 1239
rect 26228 1206 26271 1211
rect 26619 1217 27066 1233
rect 26619 1211 26647 1217
rect 26898 1216 27066 1217
rect 26228 1203 26378 1206
rect 26619 1203 26646 1211
rect 26228 1201 26646 1203
rect 26228 1183 26237 1201
rect 26255 1183 26646 1201
rect 27359 1188 27390 1239
rect 27425 1268 27462 1338
rect 27728 1337 27765 1338
rect 27577 1278 27613 1279
rect 27425 1248 27434 1268
rect 27454 1248 27462 1268
rect 27425 1238 27462 1248
rect 27521 1268 27669 1278
rect 27769 1275 27865 1277
rect 27521 1248 27530 1268
rect 27550 1248 27640 1268
rect 27660 1248 27669 1268
rect 27521 1239 27669 1248
rect 27727 1268 27865 1275
rect 27727 1248 27736 1268
rect 27756 1248 27865 1268
rect 27727 1239 27865 1248
rect 27521 1238 27558 1239
rect 27251 1185 27292 1186
rect 26228 1180 26646 1183
rect 26228 1174 26271 1180
rect 26231 1171 26271 1174
rect 27146 1178 27292 1185
rect 26628 1162 26668 1163
rect 26339 1145 26668 1162
rect 27146 1158 27202 1178
rect 27222 1158 27261 1178
rect 27281 1158 27292 1178
rect 27146 1150 27292 1158
rect 27359 1181 27516 1188
rect 27359 1161 27479 1181
rect 27499 1161 27516 1181
rect 27359 1151 27516 1161
rect 27359 1150 27394 1151
rect 26223 1102 26266 1113
rect 26223 1084 26235 1102
rect 26253 1084 26266 1102
rect 26223 1058 26266 1084
rect 26339 1058 26366 1145
rect 26628 1136 26668 1145
rect 25389 1033 25828 1051
rect 25389 1015 25789 1033
rect 25807 1015 25828 1033
rect 25389 1009 25828 1015
rect 25395 1005 25828 1009
rect 26223 1037 26366 1058
rect 26410 1110 26444 1126
rect 26628 1116 27021 1136
rect 27041 1116 27044 1136
rect 27359 1129 27390 1150
rect 27577 1129 27613 1239
rect 27632 1238 27669 1239
rect 27728 1238 27765 1239
rect 27688 1179 27778 1185
rect 27688 1159 27697 1179
rect 27717 1177 27778 1179
rect 27717 1159 27742 1177
rect 27688 1157 27742 1159
rect 27762 1157 27778 1177
rect 27688 1151 27778 1157
rect 27202 1128 27239 1129
rect 26628 1111 27044 1116
rect 27201 1119 27239 1128
rect 26628 1110 26969 1111
rect 26410 1040 26447 1110
rect 26562 1050 26593 1051
rect 26223 1035 26360 1037
rect 25774 1003 25826 1005
rect 26223 993 26266 1035
rect 26410 1020 26419 1040
rect 26439 1020 26447 1040
rect 26410 1010 26447 1020
rect 26506 1040 26593 1050
rect 26506 1020 26515 1040
rect 26535 1020 26593 1040
rect 26506 1011 26593 1020
rect 26506 1010 26543 1011
rect 26221 983 26266 993
rect 26221 965 26230 983
rect 26248 965 26266 983
rect 26221 959 26266 965
rect 26562 960 26593 1011
rect 26628 1040 26665 1110
rect 26931 1109 26968 1110
rect 27201 1099 27210 1119
rect 27230 1099 27239 1119
rect 27201 1091 27239 1099
rect 27305 1123 27390 1129
rect 27420 1128 27457 1129
rect 27305 1103 27313 1123
rect 27333 1103 27390 1123
rect 27305 1095 27390 1103
rect 27419 1119 27457 1128
rect 27419 1099 27428 1119
rect 27448 1099 27457 1119
rect 27305 1094 27341 1095
rect 27419 1091 27457 1099
rect 27523 1123 27667 1129
rect 27523 1103 27531 1123
rect 27551 1120 27639 1123
rect 27551 1103 27586 1120
rect 27523 1102 27586 1103
rect 27605 1103 27639 1120
rect 27659 1103 27667 1123
rect 27605 1102 27667 1103
rect 27523 1095 27667 1102
rect 27523 1094 27559 1095
rect 27631 1094 27667 1095
rect 27733 1128 27770 1129
rect 27733 1127 27771 1128
rect 27793 1127 27820 1131
rect 27733 1125 27820 1127
rect 27733 1119 27797 1125
rect 27733 1099 27742 1119
rect 27762 1105 27797 1119
rect 27817 1105 27820 1125
rect 27762 1100 27820 1105
rect 27762 1099 27797 1100
rect 27202 1062 27239 1091
rect 27203 1060 27239 1062
rect 26780 1050 26816 1051
rect 26628 1020 26637 1040
rect 26657 1020 26665 1040
rect 26628 1010 26665 1020
rect 26724 1040 26872 1050
rect 26972 1047 27068 1049
rect 26724 1020 26733 1040
rect 26753 1020 26843 1040
rect 26863 1020 26872 1040
rect 26724 1011 26872 1020
rect 26930 1040 27068 1047
rect 26930 1020 26939 1040
rect 26959 1020 27068 1040
rect 27203 1038 27394 1060
rect 27420 1059 27457 1091
rect 27733 1087 27797 1099
rect 27837 1061 27864 1239
rect 27696 1059 27864 1061
rect 27420 1033 27864 1059
rect 26930 1011 27068 1020
rect 26724 1010 26761 1011
rect 26221 956 26258 959
rect 26454 957 26495 958
rect 26346 950 26495 957
rect 25777 938 25814 943
rect 25768 934 25815 938
rect 25768 916 25787 934
rect 25805 916 25815 934
rect 26346 930 26405 950
rect 26425 930 26464 950
rect 26484 930 26495 950
rect 26346 922 26495 930
rect 26562 953 26719 960
rect 26562 933 26682 953
rect 26702 933 26719 953
rect 26562 923 26719 933
rect 26562 922 26597 923
rect 25768 853 25815 916
rect 26562 901 26593 922
rect 26780 901 26816 1011
rect 26835 1010 26872 1011
rect 26931 1010 26968 1011
rect 26891 951 26981 957
rect 26891 931 26900 951
rect 26920 949 26981 951
rect 26920 931 26945 949
rect 26891 929 26945 931
rect 26965 929 26981 949
rect 26891 923 26981 929
rect 26405 900 26442 901
rect 26218 892 26255 894
rect 26218 884 26260 892
rect 26218 866 26228 884
rect 26246 866 26260 884
rect 26218 857 26260 866
rect 26404 891 26442 900
rect 26404 871 26413 891
rect 26433 871 26442 891
rect 26404 863 26442 871
rect 26508 895 26593 901
rect 26623 900 26660 901
rect 26508 875 26516 895
rect 26536 875 26593 895
rect 26508 867 26593 875
rect 26622 891 26660 900
rect 26622 871 26631 891
rect 26651 871 26660 891
rect 26508 866 26544 867
rect 26622 863 26660 871
rect 26726 899 26870 901
rect 26726 895 26778 899
rect 26726 875 26734 895
rect 26754 879 26778 895
rect 26798 895 26870 899
rect 26798 879 26842 895
rect 26754 875 26842 879
rect 26862 875 26870 895
rect 26726 867 26870 875
rect 26726 866 26762 867
rect 26834 866 26870 867
rect 26936 900 26973 901
rect 26936 899 26974 900
rect 26936 891 27000 899
rect 26936 871 26945 891
rect 26965 877 27000 891
rect 27020 877 27023 897
rect 26965 872 27023 877
rect 26965 871 27000 872
rect 25768 838 25818 853
rect 25768 813 25782 838
rect 25814 813 25818 838
rect 26219 832 26260 857
rect 26405 832 26442 863
rect 26623 841 26660 863
rect 26936 859 27000 871
rect 26618 832 26660 841
rect 27040 833 27067 1011
rect 26219 820 26264 832
rect 25768 800 25815 813
rect 23153 775 23161 797
rect 23185 775 23193 797
rect 23153 767 23193 775
rect 26215 762 26264 820
rect 26405 806 26467 832
rect 26618 831 26703 832
rect 26899 831 27067 833
rect 26618 805 27067 831
rect 26618 762 26657 805
rect 26899 804 27067 805
rect 27530 809 27570 1033
rect 27696 1032 27864 1033
rect 27928 1065 27961 1398
rect 28566 1397 28593 1575
rect 28633 1537 28697 1549
rect 28973 1545 29010 1577
rect 29036 1576 29227 1598
rect 29362 1596 29471 1616
rect 29491 1596 29500 1616
rect 29362 1589 29500 1596
rect 29558 1616 29706 1625
rect 29558 1596 29567 1616
rect 29587 1596 29677 1616
rect 29697 1596 29706 1616
rect 29362 1587 29458 1589
rect 29558 1586 29706 1596
rect 29765 1616 29802 1626
rect 29765 1596 29773 1616
rect 29793 1596 29802 1616
rect 29614 1585 29650 1586
rect 29191 1574 29227 1576
rect 29191 1545 29228 1574
rect 28633 1536 28668 1537
rect 28610 1531 28668 1536
rect 28610 1511 28613 1531
rect 28633 1517 28668 1531
rect 28688 1517 28697 1537
rect 28633 1509 28697 1517
rect 28659 1508 28697 1509
rect 28660 1507 28697 1508
rect 28763 1541 28799 1542
rect 28871 1541 28907 1542
rect 28763 1533 28907 1541
rect 28763 1513 28771 1533
rect 28791 1532 28879 1533
rect 28791 1513 28826 1532
rect 28847 1513 28879 1532
rect 28899 1513 28907 1533
rect 28763 1507 28907 1513
rect 28973 1537 29011 1545
rect 29089 1541 29125 1542
rect 28973 1517 28982 1537
rect 29002 1517 29011 1537
rect 28973 1508 29011 1517
rect 29040 1533 29125 1541
rect 29040 1513 29097 1533
rect 29117 1513 29125 1533
rect 28973 1507 29010 1508
rect 29040 1507 29125 1513
rect 29191 1537 29229 1545
rect 29191 1517 29200 1537
rect 29220 1517 29229 1537
rect 29462 1526 29499 1527
rect 29765 1526 29802 1596
rect 29837 1625 29868 1676
rect 30164 1671 30209 1677
rect 30164 1653 30182 1671
rect 30200 1653 30209 1671
rect 31670 1671 31679 1691
rect 31699 1671 31707 1691
rect 31670 1661 31707 1671
rect 31766 1691 31853 1701
rect 31766 1671 31775 1691
rect 31795 1671 31853 1691
rect 31766 1662 31853 1671
rect 31766 1661 31803 1662
rect 30164 1643 30209 1653
rect 29887 1625 29924 1626
rect 29837 1616 29924 1625
rect 29837 1596 29895 1616
rect 29915 1596 29924 1616
rect 29837 1586 29924 1596
rect 29983 1616 30020 1626
rect 29983 1596 29991 1616
rect 30011 1596 30020 1616
rect 30164 1601 30207 1643
rect 30591 1632 30643 1634
rect 30070 1599 30207 1601
rect 29837 1585 29868 1586
rect 29983 1526 30020 1596
rect 29461 1525 29802 1526
rect 29191 1508 29229 1517
rect 29386 1520 29802 1525
rect 29191 1507 29228 1508
rect 28652 1479 28742 1485
rect 28652 1459 28668 1479
rect 28688 1477 28742 1479
rect 28688 1459 28713 1477
rect 28652 1457 28713 1459
rect 28733 1457 28742 1477
rect 28652 1451 28742 1457
rect 28665 1397 28702 1398
rect 28761 1397 28798 1398
rect 28817 1397 28853 1507
rect 29040 1486 29071 1507
rect 29386 1500 29389 1520
rect 29409 1500 29802 1520
rect 29986 1510 30020 1526
rect 30064 1578 30207 1599
rect 30589 1628 31022 1632
rect 30589 1622 31028 1628
rect 30589 1604 30610 1622
rect 30628 1604 31028 1622
rect 31822 1611 31853 1662
rect 31888 1691 31925 1761
rect 32191 1760 32228 1761
rect 32040 1701 32076 1702
rect 31888 1671 31897 1691
rect 31917 1671 31925 1691
rect 31888 1661 31925 1671
rect 31984 1691 32132 1701
rect 32232 1698 32328 1700
rect 31984 1671 31993 1691
rect 32013 1671 32103 1691
rect 32123 1671 32132 1691
rect 31984 1662 32132 1671
rect 32190 1691 32328 1698
rect 32190 1671 32199 1691
rect 32219 1671 32328 1691
rect 32190 1662 32328 1671
rect 31984 1661 32021 1662
rect 31714 1608 31755 1609
rect 30589 1586 31028 1604
rect 29762 1491 29802 1500
rect 30064 1491 30091 1578
rect 30164 1552 30207 1578
rect 30164 1534 30177 1552
rect 30195 1534 30207 1552
rect 30164 1523 30207 1534
rect 29036 1485 29071 1486
rect 28914 1475 29071 1485
rect 28914 1455 28931 1475
rect 28951 1455 29071 1475
rect 28914 1448 29071 1455
rect 29138 1478 29287 1486
rect 29138 1458 29149 1478
rect 29169 1458 29208 1478
rect 29228 1458 29287 1478
rect 29762 1474 30091 1491
rect 29762 1473 29802 1474
rect 29138 1451 29287 1458
rect 30159 1462 30199 1465
rect 30159 1456 30202 1462
rect 29784 1453 30202 1456
rect 29138 1450 29179 1451
rect 28872 1397 28909 1398
rect 28565 1388 28703 1397
rect 28565 1368 28674 1388
rect 28694 1368 28703 1388
rect 28565 1361 28703 1368
rect 28761 1388 28909 1397
rect 28761 1368 28770 1388
rect 28790 1368 28880 1388
rect 28900 1368 28909 1388
rect 28565 1359 28661 1361
rect 28761 1358 28909 1368
rect 28968 1388 29005 1398
rect 28968 1368 28976 1388
rect 28996 1368 29005 1388
rect 28817 1357 28853 1358
rect 28665 1298 28702 1299
rect 28968 1298 29005 1368
rect 29040 1397 29071 1448
rect 29784 1435 30175 1453
rect 30193 1435 30202 1453
rect 29784 1433 30202 1435
rect 29784 1425 29811 1433
rect 30052 1430 30202 1433
rect 29364 1419 29532 1420
rect 29783 1419 29811 1425
rect 29364 1403 29811 1419
rect 30159 1425 30202 1430
rect 29090 1397 29127 1398
rect 29040 1388 29127 1397
rect 29040 1368 29098 1388
rect 29118 1368 29127 1388
rect 29040 1358 29127 1368
rect 29186 1388 29223 1398
rect 29186 1368 29194 1388
rect 29214 1368 29223 1388
rect 29040 1357 29071 1358
rect 28664 1297 29005 1298
rect 29186 1297 29223 1368
rect 28589 1292 29005 1297
rect 28589 1272 28592 1292
rect 28612 1272 29005 1292
rect 29036 1273 29223 1297
rect 29364 1393 29808 1403
rect 29364 1391 29532 1393
rect 29364 1213 29391 1391
rect 29431 1353 29495 1365
rect 29771 1361 29808 1393
rect 29834 1392 30025 1414
rect 29989 1390 30025 1392
rect 29989 1361 30026 1390
rect 30159 1369 30199 1425
rect 29431 1352 29466 1353
rect 29408 1347 29466 1352
rect 29408 1327 29411 1347
rect 29431 1333 29466 1347
rect 29486 1333 29495 1353
rect 29431 1325 29495 1333
rect 29457 1324 29495 1325
rect 29458 1323 29495 1324
rect 29561 1357 29597 1358
rect 29669 1357 29705 1358
rect 29561 1349 29705 1357
rect 29561 1329 29569 1349
rect 29589 1329 29624 1349
rect 29644 1329 29677 1349
rect 29697 1329 29705 1349
rect 29561 1323 29705 1329
rect 29771 1353 29809 1361
rect 29887 1357 29923 1358
rect 29771 1333 29780 1353
rect 29800 1333 29809 1353
rect 29771 1324 29809 1333
rect 29838 1349 29923 1357
rect 29838 1329 29895 1349
rect 29915 1329 29923 1349
rect 29771 1323 29808 1324
rect 29838 1323 29923 1329
rect 29989 1353 30027 1361
rect 29989 1333 29998 1353
rect 30018 1333 30027 1353
rect 30159 1351 30171 1369
rect 30189 1351 30199 1369
rect 30591 1397 30643 1586
rect 30989 1561 31028 1586
rect 31606 1601 31755 1608
rect 31606 1581 31665 1601
rect 31685 1581 31724 1601
rect 31744 1581 31755 1601
rect 31606 1573 31755 1581
rect 31822 1604 31979 1611
rect 31822 1584 31942 1604
rect 31962 1584 31979 1604
rect 31822 1574 31979 1584
rect 31822 1573 31857 1574
rect 30773 1536 30960 1560
rect 30989 1541 31384 1561
rect 31404 1541 31407 1561
rect 31822 1552 31853 1573
rect 32040 1552 32076 1662
rect 32095 1661 32132 1662
rect 32191 1661 32228 1662
rect 32151 1602 32241 1608
rect 32151 1582 32160 1602
rect 32180 1600 32241 1602
rect 32180 1582 32205 1600
rect 32151 1580 32205 1582
rect 32225 1580 32241 1600
rect 32151 1574 32241 1580
rect 31665 1551 31702 1552
rect 30989 1536 31407 1541
rect 31664 1542 31702 1551
rect 30773 1465 30810 1536
rect 30989 1535 31332 1536
rect 30989 1532 31028 1535
rect 31294 1534 31331 1535
rect 30925 1475 30956 1476
rect 30773 1445 30782 1465
rect 30802 1445 30810 1465
rect 30773 1435 30810 1445
rect 30869 1465 30956 1475
rect 30869 1445 30878 1465
rect 30898 1445 30956 1465
rect 30869 1436 30956 1445
rect 30869 1435 30906 1436
rect 30591 1379 30607 1397
rect 30625 1379 30643 1397
rect 30925 1385 30956 1436
rect 30991 1465 31028 1532
rect 31664 1522 31673 1542
rect 31693 1522 31702 1542
rect 31664 1514 31702 1522
rect 31768 1546 31853 1552
rect 31883 1551 31920 1552
rect 31768 1526 31776 1546
rect 31796 1526 31853 1546
rect 31768 1518 31853 1526
rect 31882 1542 31920 1551
rect 31882 1522 31891 1542
rect 31911 1522 31920 1542
rect 31768 1517 31804 1518
rect 31882 1514 31920 1522
rect 31986 1546 32130 1552
rect 31986 1526 31994 1546
rect 32014 1541 32102 1546
rect 32014 1526 32050 1541
rect 31986 1524 32050 1526
rect 32069 1526 32102 1541
rect 32122 1526 32130 1546
rect 32069 1524 32130 1526
rect 31986 1518 32130 1524
rect 31986 1517 32022 1518
rect 32094 1517 32130 1518
rect 32196 1551 32233 1552
rect 32196 1550 32234 1551
rect 32196 1542 32260 1550
rect 32196 1522 32205 1542
rect 32225 1528 32260 1542
rect 32280 1528 32283 1548
rect 32225 1523 32283 1528
rect 32225 1522 32260 1523
rect 31665 1485 31702 1514
rect 31666 1483 31702 1485
rect 31143 1475 31179 1476
rect 30991 1445 31000 1465
rect 31020 1445 31028 1465
rect 30991 1435 31028 1445
rect 31087 1465 31235 1475
rect 31335 1472 31431 1474
rect 31087 1445 31096 1465
rect 31116 1445 31206 1465
rect 31226 1445 31235 1465
rect 31087 1436 31235 1445
rect 31293 1465 31431 1472
rect 31293 1445 31302 1465
rect 31322 1445 31431 1465
rect 31666 1461 31857 1483
rect 31883 1482 31920 1514
rect 32196 1510 32260 1522
rect 32300 1484 32327 1662
rect 32159 1482 32327 1484
rect 31883 1468 32327 1482
rect 32930 1616 33098 1617
rect 33224 1616 33264 1840
rect 33727 1844 33895 1845
rect 34130 1844 34170 1877
rect 34526 1844 34573 1877
rect 33727 1843 34171 1844
rect 33727 1818 34172 1843
rect 33727 1816 33895 1818
rect 34091 1817 34172 1818
rect 34341 1817 34390 1843
rect 34526 1817 34575 1844
rect 33727 1638 33754 1816
rect 33794 1778 33858 1790
rect 34134 1786 34171 1817
rect 34352 1786 34389 1817
rect 34534 1792 34575 1817
rect 33794 1777 33829 1778
rect 33771 1772 33829 1777
rect 33771 1752 33774 1772
rect 33794 1758 33829 1772
rect 33849 1758 33858 1778
rect 33794 1750 33858 1758
rect 33820 1749 33858 1750
rect 33821 1748 33858 1749
rect 33924 1782 33960 1783
rect 34032 1782 34068 1783
rect 33924 1774 34068 1782
rect 33924 1754 33932 1774
rect 33952 1770 34040 1774
rect 33952 1754 33996 1770
rect 33924 1750 33996 1754
rect 34016 1754 34040 1770
rect 34060 1754 34068 1774
rect 34016 1750 34068 1754
rect 33924 1748 34068 1750
rect 34134 1778 34172 1786
rect 34250 1782 34286 1783
rect 34134 1758 34143 1778
rect 34163 1758 34172 1778
rect 34134 1749 34172 1758
rect 34201 1774 34286 1782
rect 34201 1754 34258 1774
rect 34278 1754 34286 1774
rect 34134 1748 34171 1749
rect 34201 1748 34286 1754
rect 34352 1778 34390 1786
rect 34352 1758 34361 1778
rect 34381 1758 34390 1778
rect 34352 1749 34390 1758
rect 34534 1783 34576 1792
rect 34534 1765 34548 1783
rect 34566 1765 34576 1783
rect 34534 1757 34576 1765
rect 34539 1755 34576 1757
rect 34352 1748 34389 1749
rect 33813 1720 33903 1726
rect 33813 1700 33829 1720
rect 33849 1718 33903 1720
rect 33849 1700 33874 1718
rect 33813 1698 33874 1700
rect 33894 1698 33903 1718
rect 33813 1692 33903 1698
rect 33826 1638 33863 1639
rect 33922 1638 33959 1639
rect 33978 1638 34014 1748
rect 34201 1727 34232 1748
rect 34197 1726 34232 1727
rect 34075 1716 34232 1726
rect 34075 1696 34092 1716
rect 34112 1696 34232 1716
rect 34075 1689 34232 1696
rect 34299 1719 34448 1727
rect 34299 1699 34310 1719
rect 34330 1699 34369 1719
rect 34389 1699 34448 1719
rect 34299 1692 34448 1699
rect 34299 1691 34340 1692
rect 34536 1690 34573 1693
rect 34033 1638 34070 1639
rect 33726 1629 33864 1638
rect 32930 1590 33374 1616
rect 32930 1588 33098 1590
rect 31883 1456 32330 1468
rect 31926 1454 31959 1456
rect 31293 1436 31431 1445
rect 31087 1435 31124 1436
rect 30817 1382 30858 1383
rect 30591 1361 30643 1379
rect 30709 1375 30858 1382
rect 30159 1341 30199 1351
rect 30709 1355 30768 1375
rect 30788 1355 30827 1375
rect 30847 1355 30858 1375
rect 30709 1347 30858 1355
rect 30925 1378 31082 1385
rect 30925 1358 31045 1378
rect 31065 1358 31082 1378
rect 30925 1348 31082 1358
rect 30925 1347 30960 1348
rect 29989 1324 30027 1333
rect 30925 1326 30956 1347
rect 31143 1326 31179 1436
rect 31198 1435 31235 1436
rect 31294 1435 31331 1436
rect 31254 1376 31344 1382
rect 31254 1356 31263 1376
rect 31283 1374 31344 1376
rect 31283 1356 31308 1374
rect 31254 1354 31308 1356
rect 31328 1354 31344 1374
rect 31254 1348 31344 1354
rect 30768 1325 30805 1326
rect 29989 1323 30026 1324
rect 29450 1295 29540 1301
rect 29450 1275 29466 1295
rect 29486 1293 29540 1295
rect 29486 1275 29511 1293
rect 29450 1273 29511 1275
rect 29531 1273 29540 1293
rect 29450 1267 29540 1273
rect 29463 1213 29500 1214
rect 29559 1213 29596 1214
rect 29615 1213 29651 1323
rect 29838 1302 29869 1323
rect 30767 1316 30805 1325
rect 29834 1301 29869 1302
rect 29712 1291 29869 1301
rect 29712 1271 29729 1291
rect 29749 1271 29869 1291
rect 29712 1264 29869 1271
rect 29936 1294 30085 1302
rect 29936 1274 29947 1294
rect 29967 1274 30006 1294
rect 30026 1274 30085 1294
rect 30595 1298 30635 1308
rect 29936 1267 30085 1274
rect 30151 1270 30203 1288
rect 29936 1266 29977 1267
rect 29670 1213 29707 1214
rect 29363 1204 29501 1213
rect 29363 1184 29472 1204
rect 29492 1184 29501 1204
rect 29363 1177 29501 1184
rect 29559 1204 29707 1213
rect 29559 1184 29568 1204
rect 29588 1184 29678 1204
rect 29698 1184 29707 1204
rect 29363 1175 29459 1177
rect 29559 1174 29707 1184
rect 29766 1204 29803 1214
rect 29766 1184 29774 1204
rect 29794 1184 29803 1204
rect 29615 1173 29651 1174
rect 29766 1117 29803 1184
rect 29838 1213 29869 1264
rect 30151 1252 30169 1270
rect 30187 1252 30203 1270
rect 29888 1213 29925 1214
rect 29838 1204 29925 1213
rect 29838 1184 29896 1204
rect 29916 1184 29925 1204
rect 29838 1174 29925 1184
rect 29984 1204 30021 1214
rect 29984 1184 29992 1204
rect 30012 1184 30021 1204
rect 29838 1173 29869 1174
rect 29463 1114 29500 1115
rect 29766 1114 29805 1117
rect 29462 1113 29805 1114
rect 29984 1113 30021 1184
rect 29387 1108 29805 1113
rect 29387 1088 29390 1108
rect 29410 1088 29805 1108
rect 29834 1089 30021 1113
rect 27928 1057 27965 1065
rect 27928 1038 27936 1057
rect 27957 1038 27965 1057
rect 27928 1032 27965 1038
rect 29766 1063 29805 1088
rect 30151 1063 30203 1252
rect 30595 1280 30605 1298
rect 30623 1280 30635 1298
rect 30767 1296 30776 1316
rect 30796 1296 30805 1316
rect 30767 1288 30805 1296
rect 30871 1320 30956 1326
rect 30986 1325 31023 1326
rect 30871 1300 30879 1320
rect 30899 1300 30956 1320
rect 30871 1292 30956 1300
rect 30985 1316 31023 1325
rect 30985 1296 30994 1316
rect 31014 1296 31023 1316
rect 30871 1291 30907 1292
rect 30985 1288 31023 1296
rect 31089 1320 31233 1326
rect 31089 1300 31097 1320
rect 31117 1300 31150 1320
rect 31170 1300 31205 1320
rect 31225 1300 31233 1320
rect 31089 1292 31233 1300
rect 31089 1291 31125 1292
rect 31197 1291 31233 1292
rect 31299 1325 31336 1326
rect 31299 1324 31337 1325
rect 31299 1316 31363 1324
rect 31299 1296 31308 1316
rect 31328 1302 31363 1316
rect 31383 1302 31386 1322
rect 31328 1297 31386 1302
rect 31328 1296 31363 1297
rect 30595 1224 30635 1280
rect 30768 1259 30805 1288
rect 30769 1257 30805 1259
rect 30769 1235 30960 1257
rect 30986 1256 31023 1288
rect 31299 1284 31363 1296
rect 31403 1258 31430 1436
rect 32288 1411 32330 1456
rect 31262 1256 31430 1258
rect 30986 1246 31430 1256
rect 31571 1352 31758 1376
rect 31789 1357 32182 1377
rect 32202 1357 32205 1377
rect 31789 1352 32205 1357
rect 31571 1281 31608 1352
rect 31789 1351 32130 1352
rect 31723 1291 31754 1292
rect 31571 1261 31580 1281
rect 31600 1261 31608 1281
rect 31571 1251 31608 1261
rect 31667 1281 31754 1291
rect 31667 1261 31676 1281
rect 31696 1261 31754 1281
rect 31667 1252 31754 1261
rect 31667 1251 31704 1252
rect 30592 1219 30635 1224
rect 30983 1230 31430 1246
rect 30983 1224 31011 1230
rect 31262 1229 31430 1230
rect 30592 1216 30742 1219
rect 30983 1216 31010 1224
rect 30592 1214 31010 1216
rect 30592 1196 30601 1214
rect 30619 1196 31010 1214
rect 31723 1201 31754 1252
rect 31789 1281 31826 1351
rect 32092 1350 32129 1351
rect 31941 1291 31977 1292
rect 31789 1261 31798 1281
rect 31818 1261 31826 1281
rect 31789 1251 31826 1261
rect 31885 1281 32033 1291
rect 32133 1288 32229 1290
rect 31885 1261 31894 1281
rect 31914 1261 32004 1281
rect 32024 1261 32033 1281
rect 31885 1252 32033 1261
rect 32091 1281 32229 1288
rect 32091 1261 32100 1281
rect 32120 1261 32229 1281
rect 32091 1252 32229 1261
rect 31885 1251 31922 1252
rect 31615 1198 31656 1199
rect 30592 1193 31010 1196
rect 30592 1187 30635 1193
rect 30595 1184 30635 1187
rect 31510 1191 31656 1198
rect 30992 1175 31032 1176
rect 30703 1158 31032 1175
rect 31510 1171 31566 1191
rect 31586 1171 31625 1191
rect 31645 1171 31656 1191
rect 31510 1163 31656 1171
rect 31723 1194 31880 1201
rect 31723 1174 31843 1194
rect 31863 1174 31880 1194
rect 31723 1164 31880 1174
rect 31723 1163 31758 1164
rect 30587 1115 30630 1126
rect 30587 1097 30599 1115
rect 30617 1097 30630 1115
rect 30587 1071 30630 1097
rect 30703 1071 30730 1158
rect 30992 1149 31032 1158
rect 29766 1045 30205 1063
rect 29766 1027 30166 1045
rect 30184 1027 30205 1045
rect 29766 1021 30205 1027
rect 29772 1017 30205 1021
rect 30587 1050 30730 1071
rect 30774 1123 30808 1139
rect 30992 1129 31385 1149
rect 31405 1129 31408 1149
rect 31723 1142 31754 1163
rect 31941 1142 31977 1252
rect 31996 1251 32033 1252
rect 32092 1251 32129 1252
rect 32052 1192 32142 1198
rect 32052 1172 32061 1192
rect 32081 1190 32142 1192
rect 32081 1172 32106 1190
rect 32052 1170 32106 1172
rect 32126 1170 32142 1190
rect 32052 1164 32142 1170
rect 31566 1141 31603 1142
rect 30992 1124 31408 1129
rect 31565 1132 31603 1141
rect 30992 1123 31333 1124
rect 30774 1053 30811 1123
rect 30926 1063 30957 1064
rect 30587 1048 30724 1050
rect 30151 1015 30203 1017
rect 30587 1006 30630 1048
rect 30774 1033 30783 1053
rect 30803 1033 30811 1053
rect 30774 1023 30811 1033
rect 30870 1053 30957 1063
rect 30870 1033 30879 1053
rect 30899 1033 30957 1053
rect 30870 1024 30957 1033
rect 30870 1023 30907 1024
rect 30585 996 30630 1006
rect 30585 978 30594 996
rect 30612 978 30630 996
rect 30585 972 30630 978
rect 30926 973 30957 1024
rect 30992 1053 31029 1123
rect 31295 1122 31332 1123
rect 31565 1112 31574 1132
rect 31594 1112 31603 1132
rect 31565 1104 31603 1112
rect 31669 1136 31754 1142
rect 31784 1141 31821 1142
rect 31669 1116 31677 1136
rect 31697 1116 31754 1136
rect 31669 1108 31754 1116
rect 31783 1132 31821 1141
rect 31783 1112 31792 1132
rect 31812 1112 31821 1132
rect 31669 1107 31705 1108
rect 31783 1104 31821 1112
rect 31887 1136 32031 1142
rect 31887 1116 31895 1136
rect 31915 1133 32003 1136
rect 31915 1116 31950 1133
rect 31887 1115 31950 1116
rect 31969 1116 32003 1133
rect 32023 1116 32031 1136
rect 31969 1115 32031 1116
rect 31887 1108 32031 1115
rect 31887 1107 31923 1108
rect 31995 1107 32031 1108
rect 32097 1141 32134 1142
rect 32097 1140 32135 1141
rect 32157 1140 32184 1144
rect 32097 1138 32184 1140
rect 32097 1132 32161 1138
rect 32097 1112 32106 1132
rect 32126 1118 32161 1132
rect 32181 1118 32184 1138
rect 32126 1113 32184 1118
rect 32126 1112 32161 1113
rect 31566 1075 31603 1104
rect 31567 1073 31603 1075
rect 31144 1063 31180 1064
rect 30992 1033 31001 1053
rect 31021 1033 31029 1053
rect 30992 1023 31029 1033
rect 31088 1053 31236 1063
rect 31336 1060 31432 1062
rect 31088 1033 31097 1053
rect 31117 1033 31207 1053
rect 31227 1033 31236 1053
rect 31088 1024 31236 1033
rect 31294 1053 31432 1060
rect 31294 1033 31303 1053
rect 31323 1033 31432 1053
rect 31567 1051 31758 1073
rect 31784 1072 31821 1104
rect 32097 1100 32161 1112
rect 32201 1074 32228 1252
rect 32060 1072 32228 1074
rect 31784 1046 32228 1072
rect 31294 1024 31432 1033
rect 31088 1023 31125 1024
rect 30585 969 30622 972
rect 30818 970 30859 971
rect 30710 963 30859 970
rect 30154 950 30191 955
rect 30145 946 30192 950
rect 30145 928 30164 946
rect 30182 928 30192 946
rect 30710 943 30769 963
rect 30789 943 30828 963
rect 30848 943 30859 963
rect 30710 935 30859 943
rect 30926 966 31083 973
rect 30926 946 31046 966
rect 31066 946 31083 966
rect 30926 936 31083 946
rect 30926 935 30961 936
rect 30145 865 30192 928
rect 30926 914 30957 935
rect 31144 914 31180 1024
rect 31199 1023 31236 1024
rect 31295 1023 31332 1024
rect 31255 964 31345 970
rect 31255 944 31264 964
rect 31284 962 31345 964
rect 31284 944 31309 962
rect 31255 942 31309 944
rect 31329 942 31345 962
rect 31255 936 31345 942
rect 30769 913 30806 914
rect 30582 905 30619 907
rect 30582 897 30624 905
rect 30582 879 30592 897
rect 30610 879 30624 897
rect 30582 870 30624 879
rect 30768 904 30806 913
rect 30768 884 30777 904
rect 30797 884 30806 904
rect 30768 876 30806 884
rect 30872 908 30957 914
rect 30987 913 31024 914
rect 30872 888 30880 908
rect 30900 888 30957 908
rect 30872 880 30957 888
rect 30986 904 31024 913
rect 30986 884 30995 904
rect 31015 884 31024 904
rect 30872 879 30908 880
rect 30986 876 31024 884
rect 31090 912 31234 914
rect 31090 908 31142 912
rect 31090 888 31098 908
rect 31118 892 31142 908
rect 31162 908 31234 912
rect 31162 892 31206 908
rect 31118 888 31206 892
rect 31226 888 31234 908
rect 31090 880 31234 888
rect 31090 879 31126 880
rect 31198 879 31234 880
rect 31300 913 31337 914
rect 31300 912 31338 913
rect 31300 904 31364 912
rect 31300 884 31309 904
rect 31329 890 31364 904
rect 31384 890 31387 910
rect 31329 885 31387 890
rect 31329 884 31364 885
rect 30145 850 30195 865
rect 30145 825 30159 850
rect 30191 825 30195 850
rect 30583 845 30624 870
rect 30769 845 30806 876
rect 30987 854 31024 876
rect 31300 872 31364 884
rect 30982 845 31024 854
rect 31404 846 31431 1024
rect 30583 833 30628 845
rect 30145 812 30192 825
rect 27530 787 27538 809
rect 27562 787 27570 809
rect 27530 779 27570 787
rect 30579 775 30628 833
rect 30769 819 30831 845
rect 30982 844 31067 845
rect 31263 844 31431 846
rect 30982 818 31431 844
rect 30982 775 31021 818
rect 31263 817 31431 818
rect 31894 822 31934 1046
rect 32060 1045 32228 1046
rect 32292 1078 32325 1411
rect 32930 1410 32957 1588
rect 32997 1550 33061 1562
rect 33337 1558 33374 1590
rect 33400 1589 33591 1611
rect 33726 1609 33835 1629
rect 33855 1609 33864 1629
rect 33726 1602 33864 1609
rect 33922 1629 34070 1638
rect 33922 1609 33931 1629
rect 33951 1609 34041 1629
rect 34061 1609 34070 1629
rect 33726 1600 33822 1602
rect 33922 1599 34070 1609
rect 34129 1629 34166 1639
rect 34129 1609 34137 1629
rect 34157 1609 34166 1629
rect 33978 1598 34014 1599
rect 33555 1587 33591 1589
rect 33555 1558 33592 1587
rect 32997 1549 33032 1550
rect 32974 1544 33032 1549
rect 32974 1524 32977 1544
rect 32997 1530 33032 1544
rect 33052 1530 33061 1550
rect 32997 1522 33061 1530
rect 33023 1521 33061 1522
rect 33024 1520 33061 1521
rect 33127 1554 33163 1555
rect 33235 1554 33271 1555
rect 33127 1546 33271 1554
rect 33127 1526 33135 1546
rect 33155 1545 33243 1546
rect 33155 1526 33190 1545
rect 33211 1526 33243 1545
rect 33263 1526 33271 1546
rect 33127 1520 33271 1526
rect 33337 1550 33375 1558
rect 33453 1554 33489 1555
rect 33337 1530 33346 1550
rect 33366 1530 33375 1550
rect 33337 1521 33375 1530
rect 33404 1546 33489 1554
rect 33404 1526 33461 1546
rect 33481 1526 33489 1546
rect 33337 1520 33374 1521
rect 33404 1520 33489 1526
rect 33555 1550 33593 1558
rect 33555 1530 33564 1550
rect 33584 1530 33593 1550
rect 33826 1539 33863 1540
rect 34129 1539 34166 1609
rect 34201 1638 34232 1689
rect 34528 1684 34573 1690
rect 34528 1666 34546 1684
rect 34564 1666 34573 1684
rect 34528 1656 34573 1666
rect 34251 1638 34288 1639
rect 34201 1629 34288 1638
rect 34201 1609 34259 1629
rect 34279 1609 34288 1629
rect 34201 1599 34288 1609
rect 34347 1629 34384 1639
rect 34347 1609 34355 1629
rect 34375 1609 34384 1629
rect 34528 1614 34571 1656
rect 34434 1612 34571 1614
rect 34201 1598 34232 1599
rect 34347 1539 34384 1609
rect 33825 1538 34166 1539
rect 33555 1521 33593 1530
rect 33750 1533 34166 1538
rect 33555 1520 33592 1521
rect 33016 1492 33106 1498
rect 33016 1472 33032 1492
rect 33052 1490 33106 1492
rect 33052 1472 33077 1490
rect 33016 1470 33077 1472
rect 33097 1470 33106 1490
rect 33016 1464 33106 1470
rect 33029 1410 33066 1411
rect 33125 1410 33162 1411
rect 33181 1410 33217 1520
rect 33404 1499 33435 1520
rect 33750 1513 33753 1533
rect 33773 1513 34166 1533
rect 34350 1523 34384 1539
rect 34428 1591 34571 1612
rect 34126 1504 34166 1513
rect 34428 1504 34455 1591
rect 34528 1565 34571 1591
rect 34528 1547 34541 1565
rect 34559 1547 34571 1565
rect 34528 1536 34571 1547
rect 33400 1498 33435 1499
rect 33278 1488 33435 1498
rect 33278 1468 33295 1488
rect 33315 1468 33435 1488
rect 33278 1461 33435 1468
rect 33502 1491 33651 1499
rect 33502 1471 33513 1491
rect 33533 1471 33572 1491
rect 33592 1471 33651 1491
rect 34126 1487 34455 1504
rect 34126 1486 34166 1487
rect 33502 1464 33651 1471
rect 34523 1475 34563 1478
rect 34523 1469 34566 1475
rect 34148 1466 34566 1469
rect 33502 1463 33543 1464
rect 33236 1410 33273 1411
rect 32929 1401 33067 1410
rect 32929 1381 33038 1401
rect 33058 1381 33067 1401
rect 32929 1374 33067 1381
rect 33125 1401 33273 1410
rect 33125 1381 33134 1401
rect 33154 1381 33244 1401
rect 33264 1381 33273 1401
rect 32929 1372 33025 1374
rect 33125 1371 33273 1381
rect 33332 1401 33369 1411
rect 33332 1381 33340 1401
rect 33360 1381 33369 1401
rect 33181 1370 33217 1371
rect 33029 1311 33066 1312
rect 33332 1311 33369 1381
rect 33404 1410 33435 1461
rect 34148 1448 34539 1466
rect 34557 1448 34566 1466
rect 34148 1446 34566 1448
rect 34148 1438 34175 1446
rect 34416 1443 34566 1446
rect 33728 1432 33896 1433
rect 34147 1432 34175 1438
rect 33728 1416 34175 1432
rect 34523 1438 34566 1443
rect 33454 1410 33491 1411
rect 33404 1401 33491 1410
rect 33404 1381 33462 1401
rect 33482 1381 33491 1401
rect 33404 1371 33491 1381
rect 33550 1401 33587 1411
rect 33550 1381 33558 1401
rect 33578 1381 33587 1401
rect 33404 1370 33435 1371
rect 33028 1310 33369 1311
rect 33550 1310 33587 1381
rect 32953 1305 33369 1310
rect 32953 1285 32956 1305
rect 32976 1285 33369 1305
rect 33400 1286 33587 1310
rect 33728 1406 34172 1416
rect 33728 1404 33896 1406
rect 33728 1226 33755 1404
rect 33795 1366 33859 1378
rect 34135 1374 34172 1406
rect 34198 1405 34389 1427
rect 34353 1403 34389 1405
rect 34353 1374 34390 1403
rect 34523 1382 34563 1438
rect 33795 1365 33830 1366
rect 33772 1360 33830 1365
rect 33772 1340 33775 1360
rect 33795 1346 33830 1360
rect 33850 1346 33859 1366
rect 33795 1338 33859 1346
rect 33821 1337 33859 1338
rect 33822 1336 33859 1337
rect 33925 1370 33961 1371
rect 34033 1370 34069 1371
rect 33925 1362 34069 1370
rect 33925 1342 33933 1362
rect 33953 1342 33988 1362
rect 34008 1342 34041 1362
rect 34061 1342 34069 1362
rect 33925 1336 34069 1342
rect 34135 1366 34173 1374
rect 34251 1370 34287 1371
rect 34135 1346 34144 1366
rect 34164 1346 34173 1366
rect 34135 1337 34173 1346
rect 34202 1362 34287 1370
rect 34202 1342 34259 1362
rect 34279 1342 34287 1362
rect 34135 1336 34172 1337
rect 34202 1336 34287 1342
rect 34353 1366 34391 1374
rect 34353 1346 34362 1366
rect 34382 1346 34391 1366
rect 34523 1364 34535 1382
rect 34553 1364 34563 1382
rect 34523 1354 34563 1364
rect 34353 1337 34391 1346
rect 34353 1336 34390 1337
rect 33814 1308 33904 1314
rect 33814 1288 33830 1308
rect 33850 1306 33904 1308
rect 33850 1288 33875 1306
rect 33814 1286 33875 1288
rect 33895 1286 33904 1306
rect 33814 1280 33904 1286
rect 33827 1226 33864 1227
rect 33923 1226 33960 1227
rect 33979 1226 34015 1336
rect 34202 1315 34233 1336
rect 34198 1314 34233 1315
rect 34076 1304 34233 1314
rect 34076 1284 34093 1304
rect 34113 1284 34233 1304
rect 34076 1277 34233 1284
rect 34300 1307 34449 1315
rect 34300 1287 34311 1307
rect 34331 1287 34370 1307
rect 34390 1287 34449 1307
rect 34300 1280 34449 1287
rect 34515 1283 34567 1301
rect 34300 1279 34341 1280
rect 34034 1226 34071 1227
rect 33727 1217 33865 1226
rect 33727 1197 33836 1217
rect 33856 1197 33865 1217
rect 33727 1190 33865 1197
rect 33923 1217 34071 1226
rect 33923 1197 33932 1217
rect 33952 1197 34042 1217
rect 34062 1197 34071 1217
rect 33727 1188 33823 1190
rect 33923 1187 34071 1197
rect 34130 1217 34167 1227
rect 34130 1197 34138 1217
rect 34158 1197 34167 1217
rect 33979 1186 34015 1187
rect 34130 1130 34167 1197
rect 34202 1226 34233 1277
rect 34515 1265 34533 1283
rect 34551 1265 34567 1283
rect 34252 1226 34289 1227
rect 34202 1217 34289 1226
rect 34202 1197 34260 1217
rect 34280 1197 34289 1217
rect 34202 1187 34289 1197
rect 34348 1217 34385 1227
rect 34348 1197 34356 1217
rect 34376 1197 34385 1217
rect 34202 1186 34233 1187
rect 33827 1127 33864 1128
rect 34130 1127 34169 1130
rect 33826 1126 34169 1127
rect 34348 1126 34385 1197
rect 33751 1121 34169 1126
rect 33751 1101 33754 1121
rect 33774 1101 34169 1121
rect 34198 1102 34385 1126
rect 32292 1070 32329 1078
rect 32292 1051 32300 1070
rect 32321 1051 32329 1070
rect 32292 1045 32329 1051
rect 34130 1076 34169 1101
rect 34515 1076 34567 1265
rect 34130 1058 34569 1076
rect 34130 1040 34530 1058
rect 34548 1040 34569 1058
rect 34130 1034 34569 1040
rect 34136 1030 34569 1034
rect 34515 1028 34567 1030
rect 34518 963 34555 968
rect 34509 959 34556 963
rect 34509 941 34528 959
rect 34546 941 34556 959
rect 34509 878 34556 941
rect 34509 863 34559 878
rect 34509 838 34523 863
rect 34555 838 34559 863
rect 34509 825 34556 838
rect 31894 800 31902 822
rect 31926 800 31934 822
rect 31894 792 31934 800
rect 13206 732 13650 736
rect 13206 731 13632 732
rect 8842 719 9286 723
rect 8842 718 9268 719
rect 4465 707 4909 711
rect 17472 710 17877 737
rect 17913 710 17916 737
rect 21836 723 22241 750
rect 22277 723 22280 750
rect 26213 735 26618 762
rect 26654 735 26657 762
rect 30577 748 30982 775
rect 31018 748 31021 775
rect 30577 744 31021 748
rect 30577 743 31003 744
rect 26213 731 26657 735
rect 26213 730 26639 731
rect 21836 719 22280 723
rect 21836 718 22262 719
rect 4465 706 4891 707
rect 17472 706 17916 710
rect 17472 705 17898 706
rect 101 694 545 698
rect 101 693 527 694
rect 32336 573 32401 574
rect 14965 561 15030 562
rect 10601 548 10666 549
rect 6224 536 6289 537
rect 1860 523 1925 524
rect 1511 498 1698 522
rect 1729 502 2122 523
rect 2143 502 2145 523
rect 1729 498 2145 502
rect 5875 511 6062 535
rect 6093 515 6486 536
rect 6507 515 6509 536
rect 6093 511 6509 515
rect 10252 523 10439 547
rect 10470 527 10863 548
rect 10884 527 10886 548
rect 10470 523 10886 527
rect 14616 536 14803 560
rect 14834 540 15227 561
rect 15248 540 15250 561
rect 27972 560 28037 561
rect 23595 548 23660 549
rect 14834 536 15250 540
rect 1511 427 1548 498
rect 1729 497 2070 498
rect 1663 437 1694 438
rect 1511 407 1520 427
rect 1540 407 1548 427
rect 1511 397 1548 407
rect 1607 427 1694 437
rect 1607 407 1616 427
rect 1636 407 1694 427
rect 1607 398 1694 407
rect 1607 397 1644 398
rect 1663 347 1694 398
rect 1729 427 1766 497
rect 2032 496 2069 497
rect 4349 449 4414 450
rect 1881 437 1917 438
rect 1729 407 1738 427
rect 1758 407 1766 427
rect 1729 397 1766 407
rect 1825 427 1973 437
rect 2073 434 2234 436
rect 1825 407 1834 427
rect 1854 407 1944 427
rect 1964 407 1973 427
rect 1825 398 1973 407
rect 2031 429 2234 434
rect 2031 427 2204 429
rect 2031 407 2040 427
rect 2060 409 2204 427
rect 2224 409 2234 429
rect 2060 407 2234 409
rect 2031 400 2234 407
rect 4000 424 4187 448
rect 4218 428 4611 449
rect 4632 428 4634 449
rect 4218 424 4634 428
rect 5875 440 5912 511
rect 6093 510 6434 511
rect 6027 450 6058 451
rect 2031 398 2169 400
rect 1825 397 1862 398
rect 1555 344 1596 345
rect 1447 337 1596 344
rect 1447 317 1506 337
rect 1526 317 1565 337
rect 1585 317 1596 337
rect 1447 309 1596 317
rect 1663 340 1820 347
rect 1663 320 1783 340
rect 1803 320 1820 340
rect 1663 310 1820 320
rect 1663 309 1698 310
rect 1663 288 1694 309
rect 1881 288 1917 398
rect 1936 397 1973 398
rect 2032 397 2069 398
rect 1992 338 2082 344
rect 1992 318 2001 338
rect 2021 336 2082 338
rect 2021 318 2046 336
rect 1992 316 2046 318
rect 2066 316 2082 336
rect 1992 310 2082 316
rect 1506 287 1543 288
rect 1505 278 1543 287
rect 1505 258 1514 278
rect 1534 258 1543 278
rect 1505 250 1543 258
rect 1609 282 1694 288
rect 1724 287 1761 288
rect 1609 262 1617 282
rect 1637 262 1694 282
rect 1609 254 1694 262
rect 1723 278 1761 287
rect 1723 258 1732 278
rect 1752 258 1761 278
rect 1609 253 1645 254
rect 1723 250 1761 258
rect 1827 283 1971 288
rect 1827 282 1888 283
rect 1827 262 1835 282
rect 1855 262 1888 282
rect 1827 259 1888 262
rect 1911 282 1971 283
rect 1911 262 1943 282
rect 1963 262 1971 282
rect 1911 259 1971 262
rect 1827 254 1971 259
rect 1827 253 1863 254
rect 1935 253 1971 254
rect 2037 287 2074 288
rect 2037 286 2075 287
rect 2037 278 2101 286
rect 2037 258 2046 278
rect 2066 264 2101 278
rect 2121 264 2124 284
rect 2066 259 2124 264
rect 2066 258 2101 259
rect 1506 221 1543 250
rect 1507 219 1543 221
rect 1507 197 1698 219
rect 1724 218 1761 250
rect 2037 246 2101 258
rect 2141 220 2168 398
rect 4000 353 4037 424
rect 4218 423 4559 424
rect 4152 363 4183 364
rect 4000 333 4009 353
rect 4029 333 4037 353
rect 4000 323 4037 333
rect 4096 353 4183 363
rect 4096 333 4105 353
rect 4125 333 4183 353
rect 4096 324 4183 333
rect 4096 323 4133 324
rect 4152 273 4183 324
rect 4218 353 4255 423
rect 4521 422 4558 423
rect 5875 420 5884 440
rect 5904 420 5912 440
rect 5875 410 5912 420
rect 5971 440 6058 450
rect 5971 420 5980 440
rect 6000 420 6058 440
rect 5971 411 6058 420
rect 5971 410 6008 411
rect 4370 363 4406 364
rect 4218 333 4227 353
rect 4247 333 4255 353
rect 4218 323 4255 333
rect 4314 353 4462 363
rect 4562 360 4684 362
rect 4314 333 4323 353
rect 4343 333 4433 353
rect 4453 333 4462 353
rect 4314 324 4462 333
rect 4520 358 4684 360
rect 6027 360 6058 411
rect 6093 440 6130 510
rect 6396 509 6433 510
rect 8797 473 8862 474
rect 6245 450 6281 451
rect 6093 420 6102 440
rect 6122 420 6130 440
rect 6093 410 6130 420
rect 6189 440 6337 450
rect 6437 447 6598 449
rect 6189 420 6198 440
rect 6218 420 6308 440
rect 6328 420 6337 440
rect 6189 411 6337 420
rect 6395 442 6598 447
rect 6395 440 6568 442
rect 6395 420 6404 440
rect 6424 422 6568 440
rect 6588 422 6598 442
rect 6424 420 6598 422
rect 6395 413 6598 420
rect 8448 448 8635 472
rect 8666 452 9059 473
rect 9080 452 9082 473
rect 8666 448 9082 452
rect 10252 452 10289 523
rect 10470 522 10811 523
rect 10404 462 10435 463
rect 6395 411 6533 413
rect 6189 410 6226 411
rect 4520 355 4723 358
rect 5919 357 5960 358
rect 4520 353 4693 355
rect 4520 333 4529 353
rect 4549 335 4693 353
rect 4713 335 4723 355
rect 4549 333 4723 335
rect 4520 326 4723 333
rect 5811 350 5960 357
rect 5811 330 5870 350
rect 5890 330 5929 350
rect 5949 330 5960 350
rect 4520 324 4658 326
rect 4314 323 4351 324
rect 4044 270 4085 271
rect 3936 263 4085 270
rect 3936 243 3995 263
rect 4015 243 4054 263
rect 4074 243 4085 263
rect 3936 235 4085 243
rect 4152 266 4309 273
rect 4152 246 4272 266
rect 4292 246 4309 266
rect 4152 236 4309 246
rect 4152 235 4187 236
rect 2000 218 2168 220
rect 1724 192 2168 218
rect 4152 214 4183 235
rect 4370 214 4406 324
rect 4425 323 4462 324
rect 4521 323 4558 324
rect 4481 264 4571 270
rect 4481 244 4490 264
rect 4510 262 4571 264
rect 4510 244 4535 262
rect 4481 242 4535 244
rect 4555 242 4571 262
rect 4481 236 4571 242
rect 3995 213 4032 214
rect 1834 189 1874 192
rect 2000 191 2168 192
rect 3994 204 4032 213
rect 3994 184 4003 204
rect 4023 184 4032 204
rect 3994 176 4032 184
rect 4098 208 4183 214
rect 4213 213 4250 214
rect 4098 188 4106 208
rect 4126 188 4183 208
rect 4098 180 4183 188
rect 4212 204 4250 213
rect 4212 184 4221 204
rect 4241 184 4250 204
rect 4098 179 4134 180
rect 4212 176 4250 184
rect 4316 208 4460 214
rect 4316 188 4324 208
rect 4344 205 4432 208
rect 4344 188 4380 205
rect 4316 184 4380 188
rect 4397 188 4432 205
rect 4452 188 4460 208
rect 4397 184 4460 188
rect 4316 180 4460 184
rect 4316 179 4352 180
rect 4424 179 4460 180
rect 4526 213 4563 214
rect 4526 212 4564 213
rect 4526 204 4590 212
rect 4526 184 4535 204
rect 4555 190 4590 204
rect 4610 190 4613 210
rect 4555 185 4613 190
rect 4555 184 4590 185
rect 3995 147 4032 176
rect 3996 145 4032 147
rect 3996 123 4187 145
rect 4213 144 4250 176
rect 4526 172 4590 184
rect 4630 146 4657 324
rect 5811 322 5960 330
rect 6027 353 6184 360
rect 6027 333 6147 353
rect 6167 333 6184 353
rect 6027 323 6184 333
rect 6027 322 6062 323
rect 6027 301 6058 322
rect 6245 301 6281 411
rect 6300 410 6337 411
rect 6396 410 6433 411
rect 6356 351 6446 357
rect 6356 331 6365 351
rect 6385 349 6446 351
rect 6385 331 6410 349
rect 6356 329 6410 331
rect 6430 329 6446 349
rect 6356 323 6446 329
rect 5870 300 5907 301
rect 5869 291 5907 300
rect 5869 271 5878 291
rect 5898 271 5907 291
rect 5869 263 5907 271
rect 5973 295 6058 301
rect 6088 300 6125 301
rect 5973 275 5981 295
rect 6001 275 6058 295
rect 5973 267 6058 275
rect 6087 291 6125 300
rect 6087 271 6096 291
rect 6116 271 6125 291
rect 5973 266 6009 267
rect 6087 263 6125 271
rect 6191 297 6335 301
rect 6191 295 6255 297
rect 6191 275 6199 295
rect 6219 275 6255 295
rect 6191 273 6255 275
rect 6278 295 6335 297
rect 6278 275 6307 295
rect 6327 275 6335 295
rect 6278 273 6335 275
rect 6191 267 6335 273
rect 6191 266 6227 267
rect 6299 266 6335 267
rect 6401 300 6438 301
rect 6401 299 6439 300
rect 6401 291 6465 299
rect 6401 271 6410 291
rect 6430 277 6465 291
rect 6485 277 6488 297
rect 6430 272 6488 277
rect 6430 271 6465 272
rect 5870 234 5907 263
rect 5871 232 5907 234
rect 5871 210 6062 232
rect 6088 231 6125 263
rect 6401 259 6465 271
rect 6505 233 6532 411
rect 8448 377 8485 448
rect 8666 447 9007 448
rect 8600 387 8631 388
rect 8448 357 8457 377
rect 8477 357 8485 377
rect 8448 347 8485 357
rect 8544 377 8631 387
rect 8544 357 8553 377
rect 8573 357 8631 377
rect 8544 348 8631 357
rect 8544 347 8581 348
rect 8600 297 8631 348
rect 8666 377 8703 447
rect 8969 446 9006 447
rect 10252 432 10261 452
rect 10281 432 10289 452
rect 10252 422 10289 432
rect 10348 452 10435 462
rect 10348 432 10357 452
rect 10377 432 10435 452
rect 10348 423 10435 432
rect 10348 422 10385 423
rect 8818 387 8854 388
rect 8666 357 8675 377
rect 8695 357 8703 377
rect 8666 347 8703 357
rect 8762 377 8910 387
rect 9010 384 9132 386
rect 8762 357 8771 377
rect 8791 357 8881 377
rect 8901 357 8910 377
rect 8762 348 8910 357
rect 8968 382 9132 384
rect 8968 379 9171 382
rect 8968 377 9141 379
rect 8968 357 8977 377
rect 8997 359 9141 377
rect 9161 359 9171 379
rect 10404 372 10435 423
rect 10470 452 10507 522
rect 10773 521 10810 522
rect 13090 474 13155 475
rect 10622 462 10658 463
rect 10470 432 10479 452
rect 10499 432 10507 452
rect 10470 422 10507 432
rect 10566 452 10714 462
rect 10814 459 10975 461
rect 10566 432 10575 452
rect 10595 432 10685 452
rect 10705 432 10714 452
rect 10566 423 10714 432
rect 10772 454 10975 459
rect 10772 452 10945 454
rect 10772 432 10781 452
rect 10801 434 10945 452
rect 10965 434 10975 454
rect 10801 432 10975 434
rect 10772 425 10975 432
rect 12741 449 12928 473
rect 12959 453 13352 474
rect 13373 453 13375 474
rect 12959 449 13375 453
rect 14616 465 14653 536
rect 14834 535 15175 536
rect 19231 535 19296 536
rect 14768 475 14799 476
rect 10772 423 10910 425
rect 10566 422 10603 423
rect 10296 369 10337 370
rect 8997 357 9171 359
rect 8968 350 9171 357
rect 10188 362 10337 369
rect 8968 348 9106 350
rect 8762 347 8799 348
rect 8492 294 8533 295
rect 8379 287 8533 294
rect 8379 267 8443 287
rect 8463 267 8502 287
rect 8522 267 8533 287
rect 8379 260 8533 267
rect 8384 259 8533 260
rect 8600 290 8757 297
rect 8600 270 8720 290
rect 8740 270 8757 290
rect 8600 260 8757 270
rect 8600 259 8635 260
rect 8600 238 8631 259
rect 8818 238 8854 348
rect 8873 347 8910 348
rect 8969 347 9006 348
rect 8929 288 9019 294
rect 8929 268 8938 288
rect 8958 286 9019 288
rect 8958 268 8983 286
rect 8929 266 8983 268
rect 9003 266 9019 286
rect 8929 260 9019 266
rect 8443 237 8480 238
rect 6364 231 6532 233
rect 6088 205 6532 231
rect 6198 202 6238 205
rect 6364 204 6532 205
rect 8442 228 8480 237
rect 8442 208 8451 228
rect 8471 208 8480 228
rect 8442 200 8480 208
rect 8546 232 8631 238
rect 8661 237 8698 238
rect 8546 212 8554 232
rect 8574 212 8631 232
rect 8546 204 8631 212
rect 8660 228 8698 237
rect 8660 208 8669 228
rect 8689 208 8698 228
rect 8546 203 8582 204
rect 8660 200 8698 208
rect 8764 232 8908 238
rect 8764 212 8772 232
rect 8792 227 8880 232
rect 8792 212 8819 227
rect 8764 209 8819 212
rect 8840 212 8880 227
rect 8900 212 8908 232
rect 8840 209 8908 212
rect 8764 204 8908 209
rect 8764 203 8800 204
rect 8872 203 8908 204
rect 8974 237 9011 238
rect 8974 236 9012 237
rect 8974 228 9038 236
rect 8974 208 8983 228
rect 9003 214 9038 228
rect 9058 214 9061 234
rect 9003 209 9061 214
rect 9003 208 9038 209
rect 8443 171 8480 200
rect 8444 169 8480 171
rect 8444 147 8635 169
rect 8661 168 8698 200
rect 8974 196 9038 208
rect 9078 170 9105 348
rect 10188 342 10247 362
rect 10267 342 10306 362
rect 10326 342 10337 362
rect 10188 334 10337 342
rect 10404 365 10561 372
rect 10404 345 10524 365
rect 10544 345 10561 365
rect 10404 335 10561 345
rect 10404 334 10439 335
rect 10404 313 10435 334
rect 10622 313 10658 423
rect 10677 422 10714 423
rect 10773 422 10810 423
rect 10733 363 10823 369
rect 10733 343 10742 363
rect 10762 361 10823 363
rect 10762 343 10787 361
rect 10733 341 10787 343
rect 10807 341 10823 361
rect 10733 335 10823 341
rect 10247 312 10284 313
rect 10246 303 10284 312
rect 10246 283 10255 303
rect 10275 283 10284 303
rect 10246 275 10284 283
rect 10350 307 10435 313
rect 10465 312 10502 313
rect 10350 287 10358 307
rect 10378 287 10435 307
rect 10350 279 10435 287
rect 10464 303 10502 312
rect 10464 283 10473 303
rect 10493 283 10502 303
rect 10350 278 10386 279
rect 10464 275 10502 283
rect 10568 308 10712 313
rect 10568 307 10629 308
rect 10568 287 10576 307
rect 10596 287 10629 307
rect 10568 284 10629 287
rect 10652 307 10712 308
rect 10652 287 10684 307
rect 10704 287 10712 307
rect 10652 284 10712 287
rect 10568 279 10712 284
rect 10568 278 10604 279
rect 10676 278 10712 279
rect 10778 312 10815 313
rect 10778 311 10816 312
rect 10778 303 10842 311
rect 10778 283 10787 303
rect 10807 289 10842 303
rect 10862 289 10865 309
rect 10807 284 10865 289
rect 10807 283 10842 284
rect 10247 246 10284 275
rect 10248 244 10284 246
rect 10248 222 10439 244
rect 10465 243 10502 275
rect 10778 271 10842 283
rect 10882 245 10909 423
rect 12741 378 12778 449
rect 12959 448 13300 449
rect 12893 388 12924 389
rect 12741 358 12750 378
rect 12770 358 12778 378
rect 12741 348 12778 358
rect 12837 378 12924 388
rect 12837 358 12846 378
rect 12866 358 12924 378
rect 12837 349 12924 358
rect 12837 348 12874 349
rect 12893 298 12924 349
rect 12959 378 12996 448
rect 13262 447 13299 448
rect 14616 445 14625 465
rect 14645 445 14653 465
rect 14616 435 14653 445
rect 14712 465 14799 475
rect 14712 445 14721 465
rect 14741 445 14799 465
rect 14712 436 14799 445
rect 14712 435 14749 436
rect 13111 388 13147 389
rect 12959 358 12968 378
rect 12988 358 12996 378
rect 12959 348 12996 358
rect 13055 378 13203 388
rect 13303 385 13425 387
rect 13055 358 13064 378
rect 13084 358 13174 378
rect 13194 358 13203 378
rect 13055 349 13203 358
rect 13261 383 13425 385
rect 14768 385 14799 436
rect 14834 465 14871 535
rect 15137 534 15174 535
rect 18882 510 19069 534
rect 19100 514 19493 535
rect 19514 514 19516 535
rect 19100 510 19516 514
rect 23246 523 23433 547
rect 23464 527 23857 548
rect 23878 527 23880 548
rect 23464 523 23880 527
rect 27623 535 27810 559
rect 27841 539 28234 560
rect 28255 539 28257 560
rect 27841 535 28257 539
rect 31987 548 32174 572
rect 32205 552 32598 573
rect 32619 552 32621 573
rect 32205 548 32621 552
rect 14986 475 15022 476
rect 14834 445 14843 465
rect 14863 445 14871 465
rect 14834 435 14871 445
rect 14930 465 15078 475
rect 15178 472 15339 474
rect 14930 445 14939 465
rect 14959 445 15049 465
rect 15069 445 15078 465
rect 14930 436 15078 445
rect 15136 467 15339 472
rect 15136 465 15309 467
rect 15136 445 15145 465
rect 15165 447 15309 465
rect 15329 447 15339 467
rect 15165 445 15339 447
rect 15136 438 15339 445
rect 18882 439 18919 510
rect 19100 509 19441 510
rect 19034 449 19065 450
rect 15136 436 15274 438
rect 14930 435 14967 436
rect 13261 380 13464 383
rect 14660 382 14701 383
rect 13261 378 13434 380
rect 13261 358 13270 378
rect 13290 360 13434 378
rect 13454 360 13464 380
rect 13290 358 13464 360
rect 13261 351 13464 358
rect 14552 375 14701 382
rect 14552 355 14611 375
rect 14631 355 14670 375
rect 14690 355 14701 375
rect 13261 349 13399 351
rect 13055 348 13092 349
rect 12785 295 12826 296
rect 12677 288 12826 295
rect 12677 268 12736 288
rect 12756 268 12795 288
rect 12815 268 12826 288
rect 12677 260 12826 268
rect 12893 291 13050 298
rect 12893 271 13013 291
rect 13033 271 13050 291
rect 12893 261 13050 271
rect 12893 260 12928 261
rect 10741 243 10909 245
rect 10465 217 10909 243
rect 12893 239 12924 260
rect 13111 239 13147 349
rect 13166 348 13203 349
rect 13262 348 13299 349
rect 13222 289 13312 295
rect 13222 269 13231 289
rect 13251 287 13312 289
rect 13251 269 13276 287
rect 13222 267 13276 269
rect 13296 267 13312 287
rect 13222 261 13312 267
rect 12736 238 12773 239
rect 10575 214 10615 217
rect 10741 216 10909 217
rect 12735 229 12773 238
rect 12735 209 12744 229
rect 12764 209 12773 229
rect 12735 201 12773 209
rect 12839 233 12924 239
rect 12954 238 12991 239
rect 12839 213 12847 233
rect 12867 213 12924 233
rect 12839 205 12924 213
rect 12953 229 12991 238
rect 12953 209 12962 229
rect 12982 209 12991 229
rect 12839 204 12875 205
rect 12953 201 12991 209
rect 13057 233 13201 239
rect 13057 213 13065 233
rect 13085 213 13117 233
rect 13057 211 13117 213
rect 13138 213 13173 233
rect 13193 213 13201 233
rect 13138 211 13201 213
rect 13057 205 13201 211
rect 13057 204 13093 205
rect 13165 204 13201 205
rect 13267 238 13304 239
rect 13267 237 13305 238
rect 13267 229 13331 237
rect 13267 209 13276 229
rect 13296 215 13331 229
rect 13351 215 13354 235
rect 13296 210 13354 215
rect 13296 209 13331 210
rect 12736 172 12773 201
rect 8937 168 9105 170
rect 4489 144 4657 146
rect 4213 118 4657 144
rect 8661 142 9105 168
rect 12737 170 12773 172
rect 12737 148 12928 170
rect 12954 169 12991 201
rect 13267 197 13331 209
rect 13371 171 13398 349
rect 14552 347 14701 355
rect 14768 378 14925 385
rect 14768 358 14888 378
rect 14908 358 14925 378
rect 14768 348 14925 358
rect 14768 347 14803 348
rect 14768 326 14799 347
rect 14986 326 15022 436
rect 15041 435 15078 436
rect 15137 435 15174 436
rect 15097 376 15187 382
rect 15097 356 15106 376
rect 15126 374 15187 376
rect 15126 356 15151 374
rect 15097 354 15151 356
rect 15171 354 15187 374
rect 15097 348 15187 354
rect 14611 325 14648 326
rect 14610 316 14648 325
rect 14610 296 14619 316
rect 14639 296 14648 316
rect 14610 288 14648 296
rect 14714 320 14799 326
rect 14829 325 14866 326
rect 14714 300 14722 320
rect 14742 300 14799 320
rect 14714 292 14799 300
rect 14828 316 14866 325
rect 14828 296 14837 316
rect 14857 296 14866 316
rect 14714 291 14750 292
rect 14828 288 14866 296
rect 14932 322 15076 326
rect 14932 320 14996 322
rect 14932 300 14940 320
rect 14960 300 14996 320
rect 14932 298 14996 300
rect 15019 320 15076 322
rect 15019 300 15048 320
rect 15068 300 15076 320
rect 15019 298 15076 300
rect 14932 292 15076 298
rect 14932 291 14968 292
rect 15040 291 15076 292
rect 15142 325 15179 326
rect 15142 324 15180 325
rect 15142 316 15206 324
rect 15142 296 15151 316
rect 15171 302 15206 316
rect 15226 302 15229 322
rect 15171 297 15229 302
rect 15171 296 15206 297
rect 14611 259 14648 288
rect 14612 257 14648 259
rect 14612 235 14803 257
rect 14829 256 14866 288
rect 15142 284 15206 296
rect 15246 258 15273 436
rect 18882 419 18891 439
rect 18911 419 18919 439
rect 17287 410 17352 411
rect 16938 385 17125 409
rect 17156 389 17549 410
rect 17570 389 17572 410
rect 18882 409 18919 419
rect 18978 439 19065 449
rect 18978 419 18987 439
rect 19007 419 19065 439
rect 18978 410 19065 419
rect 18978 409 19015 410
rect 17156 385 17572 389
rect 16938 314 16975 385
rect 17156 384 17497 385
rect 17090 324 17121 325
rect 16938 294 16947 314
rect 16967 294 16975 314
rect 16938 284 16975 294
rect 17034 314 17121 324
rect 17034 294 17043 314
rect 17063 294 17121 314
rect 17034 285 17121 294
rect 17034 284 17071 285
rect 15105 256 15273 258
rect 14829 230 15273 256
rect 17090 234 17121 285
rect 17156 314 17193 384
rect 17459 383 17496 384
rect 19034 359 19065 410
rect 19100 439 19137 509
rect 19403 508 19440 509
rect 21720 461 21785 462
rect 19252 449 19288 450
rect 19100 419 19109 439
rect 19129 419 19137 439
rect 19100 409 19137 419
rect 19196 439 19344 449
rect 19444 446 19605 448
rect 19196 419 19205 439
rect 19225 419 19315 439
rect 19335 419 19344 439
rect 19196 410 19344 419
rect 19402 441 19605 446
rect 19402 439 19575 441
rect 19402 419 19411 439
rect 19431 421 19575 439
rect 19595 421 19605 441
rect 19431 419 19605 421
rect 19402 412 19605 419
rect 21371 436 21558 460
rect 21589 440 21982 461
rect 22003 440 22005 461
rect 21589 436 22005 440
rect 23246 452 23283 523
rect 23464 522 23805 523
rect 23398 462 23429 463
rect 19402 410 19540 412
rect 19196 409 19233 410
rect 18926 356 18967 357
rect 18818 349 18967 356
rect 18818 329 18877 349
rect 18897 329 18936 349
rect 18956 329 18967 349
rect 17308 324 17344 325
rect 17156 294 17165 314
rect 17185 294 17193 314
rect 17156 284 17193 294
rect 17252 314 17400 324
rect 17500 321 17622 323
rect 18818 321 18967 329
rect 19034 352 19191 359
rect 19034 332 19154 352
rect 19174 332 19191 352
rect 19034 322 19191 332
rect 19034 321 19069 322
rect 17252 294 17261 314
rect 17281 294 17371 314
rect 17391 294 17400 314
rect 17252 285 17400 294
rect 17458 319 17622 321
rect 17458 316 17661 319
rect 17458 314 17631 316
rect 17458 294 17467 314
rect 17487 296 17631 314
rect 17651 296 17661 316
rect 19034 300 19065 321
rect 19252 300 19288 410
rect 19307 409 19344 410
rect 19403 409 19440 410
rect 19363 350 19453 356
rect 19363 330 19372 350
rect 19392 348 19453 350
rect 19392 330 19417 348
rect 19363 328 19417 330
rect 19437 328 19453 348
rect 19363 322 19453 328
rect 18877 299 18914 300
rect 17487 294 17661 296
rect 17458 287 17661 294
rect 18876 290 18914 299
rect 17458 285 17596 287
rect 17252 284 17289 285
rect 16982 231 17023 232
rect 14939 227 14979 230
rect 15105 229 15273 230
rect 16869 224 17023 231
rect 16869 204 16933 224
rect 16953 204 16992 224
rect 17012 204 17023 224
rect 16869 197 17023 204
rect 16874 196 17023 197
rect 17090 227 17247 234
rect 17090 207 17210 227
rect 17230 207 17247 227
rect 17090 197 17247 207
rect 17090 196 17125 197
rect 17090 175 17121 196
rect 17308 175 17344 285
rect 17363 284 17400 285
rect 17459 284 17496 285
rect 17419 225 17509 231
rect 17419 205 17428 225
rect 17448 223 17509 225
rect 17448 205 17473 223
rect 17419 203 17473 205
rect 17493 203 17509 223
rect 17419 197 17509 203
rect 16933 174 16970 175
rect 13230 169 13398 171
rect 12954 143 13398 169
rect 8771 139 8811 142
rect 8937 141 9105 142
rect 13064 140 13104 143
rect 13230 142 13398 143
rect 16932 165 16970 174
rect 16932 145 16941 165
rect 16961 145 16970 165
rect 16932 137 16970 145
rect 17036 169 17121 175
rect 17151 174 17188 175
rect 17036 149 17044 169
rect 17064 149 17121 169
rect 17036 141 17121 149
rect 17150 165 17188 174
rect 17150 145 17159 165
rect 17179 145 17188 165
rect 17036 140 17072 141
rect 17150 137 17188 145
rect 17254 169 17398 175
rect 17254 149 17262 169
rect 17282 149 17370 169
rect 17390 149 17398 169
rect 17254 141 17398 149
rect 17254 140 17290 141
rect 17362 140 17398 141
rect 17464 174 17501 175
rect 17464 173 17502 174
rect 17464 165 17528 173
rect 17464 145 17473 165
rect 17493 151 17528 165
rect 17548 151 17551 171
rect 17493 146 17551 151
rect 17493 145 17528 146
rect 4323 115 4363 118
rect 4489 117 4657 118
rect 16933 108 16970 137
rect 16934 106 16970 108
rect 16934 84 17125 106
rect 17151 105 17188 137
rect 17464 133 17528 145
rect 17568 107 17595 285
rect 18876 270 18885 290
rect 18905 270 18914 290
rect 18876 262 18914 270
rect 18980 294 19065 300
rect 19095 299 19132 300
rect 18980 274 18988 294
rect 19008 274 19065 294
rect 18980 266 19065 274
rect 19094 290 19132 299
rect 19094 270 19103 290
rect 19123 270 19132 290
rect 18980 265 19016 266
rect 19094 262 19132 270
rect 19198 295 19342 300
rect 19198 294 19259 295
rect 19198 274 19206 294
rect 19226 274 19259 294
rect 19198 271 19259 274
rect 19282 294 19342 295
rect 19282 274 19314 294
rect 19334 274 19342 294
rect 19282 271 19342 274
rect 19198 266 19342 271
rect 19198 265 19234 266
rect 19306 265 19342 266
rect 19408 299 19445 300
rect 19408 298 19446 299
rect 19408 290 19472 298
rect 19408 270 19417 290
rect 19437 276 19472 290
rect 19492 276 19495 296
rect 19437 271 19495 276
rect 19437 270 19472 271
rect 18877 233 18914 262
rect 18878 231 18914 233
rect 18878 209 19069 231
rect 19095 230 19132 262
rect 19408 258 19472 270
rect 19512 232 19539 410
rect 21371 365 21408 436
rect 21589 435 21930 436
rect 21523 375 21554 376
rect 21371 345 21380 365
rect 21400 345 21408 365
rect 21371 335 21408 345
rect 21467 365 21554 375
rect 21467 345 21476 365
rect 21496 345 21554 365
rect 21467 336 21554 345
rect 21467 335 21504 336
rect 21523 285 21554 336
rect 21589 365 21626 435
rect 21892 434 21929 435
rect 23246 432 23255 452
rect 23275 432 23283 452
rect 23246 422 23283 432
rect 23342 452 23429 462
rect 23342 432 23351 452
rect 23371 432 23429 452
rect 23342 423 23429 432
rect 23342 422 23379 423
rect 21741 375 21777 376
rect 21589 345 21598 365
rect 21618 345 21626 365
rect 21589 335 21626 345
rect 21685 365 21833 375
rect 21933 372 22055 374
rect 21685 345 21694 365
rect 21714 345 21804 365
rect 21824 345 21833 365
rect 21685 336 21833 345
rect 21891 370 22055 372
rect 23398 372 23429 423
rect 23464 452 23501 522
rect 23767 521 23804 522
rect 26168 485 26233 486
rect 23616 462 23652 463
rect 23464 432 23473 452
rect 23493 432 23501 452
rect 23464 422 23501 432
rect 23560 452 23708 462
rect 23808 459 23969 461
rect 23560 432 23569 452
rect 23589 432 23679 452
rect 23699 432 23708 452
rect 23560 423 23708 432
rect 23766 454 23969 459
rect 23766 452 23939 454
rect 23766 432 23775 452
rect 23795 434 23939 452
rect 23959 434 23969 454
rect 23795 432 23969 434
rect 23766 425 23969 432
rect 25819 460 26006 484
rect 26037 464 26430 485
rect 26451 464 26453 485
rect 26037 460 26453 464
rect 27623 464 27660 535
rect 27841 534 28182 535
rect 27775 474 27806 475
rect 23766 423 23904 425
rect 23560 422 23597 423
rect 21891 367 22094 370
rect 23290 369 23331 370
rect 21891 365 22064 367
rect 21891 345 21900 365
rect 21920 347 22064 365
rect 22084 347 22094 367
rect 21920 345 22094 347
rect 21891 338 22094 345
rect 23182 362 23331 369
rect 23182 342 23241 362
rect 23261 342 23300 362
rect 23320 342 23331 362
rect 21891 336 22029 338
rect 21685 335 21722 336
rect 21415 282 21456 283
rect 21307 275 21456 282
rect 21307 255 21366 275
rect 21386 255 21425 275
rect 21445 255 21456 275
rect 21307 247 21456 255
rect 21523 278 21680 285
rect 21523 258 21643 278
rect 21663 258 21680 278
rect 21523 248 21680 258
rect 21523 247 21558 248
rect 19371 230 19539 232
rect 19095 204 19539 230
rect 21523 226 21554 247
rect 21741 226 21777 336
rect 21796 335 21833 336
rect 21892 335 21929 336
rect 21852 276 21942 282
rect 21852 256 21861 276
rect 21881 274 21942 276
rect 21881 256 21906 274
rect 21852 254 21906 256
rect 21926 254 21942 274
rect 21852 248 21942 254
rect 21366 225 21403 226
rect 19205 201 19245 204
rect 19371 203 19539 204
rect 21365 216 21403 225
rect 21365 196 21374 216
rect 21394 196 21403 216
rect 21365 188 21403 196
rect 21469 220 21554 226
rect 21584 225 21621 226
rect 21469 200 21477 220
rect 21497 200 21554 220
rect 21469 192 21554 200
rect 21583 216 21621 225
rect 21583 196 21592 216
rect 21612 196 21621 216
rect 21469 191 21505 192
rect 21583 188 21621 196
rect 21687 220 21831 226
rect 21687 200 21695 220
rect 21715 217 21803 220
rect 21715 200 21751 217
rect 21687 196 21751 200
rect 21768 200 21803 217
rect 21823 200 21831 220
rect 21768 196 21831 200
rect 21687 192 21831 196
rect 21687 191 21723 192
rect 21795 191 21831 192
rect 21897 225 21934 226
rect 21897 224 21935 225
rect 21897 216 21961 224
rect 21897 196 21906 216
rect 21926 202 21961 216
rect 21981 202 21984 222
rect 21926 197 21984 202
rect 21926 196 21961 197
rect 21366 159 21403 188
rect 21367 157 21403 159
rect 21367 135 21558 157
rect 21584 156 21621 188
rect 21897 184 21961 196
rect 22001 158 22028 336
rect 23182 334 23331 342
rect 23398 365 23555 372
rect 23398 345 23518 365
rect 23538 345 23555 365
rect 23398 335 23555 345
rect 23398 334 23433 335
rect 23398 313 23429 334
rect 23616 313 23652 423
rect 23671 422 23708 423
rect 23767 422 23804 423
rect 23727 363 23817 369
rect 23727 343 23736 363
rect 23756 361 23817 363
rect 23756 343 23781 361
rect 23727 341 23781 343
rect 23801 341 23817 361
rect 23727 335 23817 341
rect 23241 312 23278 313
rect 23240 303 23278 312
rect 23240 283 23249 303
rect 23269 283 23278 303
rect 23240 275 23278 283
rect 23344 307 23429 313
rect 23459 312 23496 313
rect 23344 287 23352 307
rect 23372 287 23429 307
rect 23344 279 23429 287
rect 23458 303 23496 312
rect 23458 283 23467 303
rect 23487 283 23496 303
rect 23344 278 23380 279
rect 23458 275 23496 283
rect 23562 309 23706 313
rect 23562 307 23626 309
rect 23562 287 23570 307
rect 23590 287 23626 307
rect 23562 285 23626 287
rect 23649 307 23706 309
rect 23649 287 23678 307
rect 23698 287 23706 307
rect 23649 285 23706 287
rect 23562 279 23706 285
rect 23562 278 23598 279
rect 23670 278 23706 279
rect 23772 312 23809 313
rect 23772 311 23810 312
rect 23772 303 23836 311
rect 23772 283 23781 303
rect 23801 289 23836 303
rect 23856 289 23859 309
rect 23801 284 23859 289
rect 23801 283 23836 284
rect 23241 246 23278 275
rect 23242 244 23278 246
rect 23242 222 23433 244
rect 23459 243 23496 275
rect 23772 271 23836 283
rect 23876 245 23903 423
rect 25819 389 25856 460
rect 26037 459 26378 460
rect 25971 399 26002 400
rect 25819 369 25828 389
rect 25848 369 25856 389
rect 25819 359 25856 369
rect 25915 389 26002 399
rect 25915 369 25924 389
rect 25944 369 26002 389
rect 25915 360 26002 369
rect 25915 359 25952 360
rect 25971 309 26002 360
rect 26037 389 26074 459
rect 26340 458 26377 459
rect 27623 444 27632 464
rect 27652 444 27660 464
rect 27623 434 27660 444
rect 27719 464 27806 474
rect 27719 444 27728 464
rect 27748 444 27806 464
rect 27719 435 27806 444
rect 27719 434 27756 435
rect 26189 399 26225 400
rect 26037 369 26046 389
rect 26066 369 26074 389
rect 26037 359 26074 369
rect 26133 389 26281 399
rect 26381 396 26503 398
rect 26133 369 26142 389
rect 26162 369 26252 389
rect 26272 369 26281 389
rect 26133 360 26281 369
rect 26339 394 26503 396
rect 26339 391 26542 394
rect 26339 389 26512 391
rect 26339 369 26348 389
rect 26368 371 26512 389
rect 26532 371 26542 391
rect 27775 384 27806 435
rect 27841 464 27878 534
rect 28144 533 28181 534
rect 30461 486 30526 487
rect 27993 474 28029 475
rect 27841 444 27850 464
rect 27870 444 27878 464
rect 27841 434 27878 444
rect 27937 464 28085 474
rect 28185 471 28346 473
rect 27937 444 27946 464
rect 27966 444 28056 464
rect 28076 444 28085 464
rect 27937 435 28085 444
rect 28143 466 28346 471
rect 28143 464 28316 466
rect 28143 444 28152 464
rect 28172 446 28316 464
rect 28336 446 28346 466
rect 28172 444 28346 446
rect 28143 437 28346 444
rect 30112 461 30299 485
rect 30330 465 30723 486
rect 30744 465 30746 486
rect 30330 461 30746 465
rect 31987 477 32024 548
rect 32205 547 32546 548
rect 32139 487 32170 488
rect 28143 435 28281 437
rect 27937 434 27974 435
rect 27667 381 27708 382
rect 26368 369 26542 371
rect 26339 362 26542 369
rect 27559 374 27708 381
rect 26339 360 26477 362
rect 26133 359 26170 360
rect 25863 306 25904 307
rect 25750 299 25904 306
rect 25750 279 25814 299
rect 25834 279 25873 299
rect 25893 279 25904 299
rect 25750 272 25904 279
rect 25755 271 25904 272
rect 25971 302 26128 309
rect 25971 282 26091 302
rect 26111 282 26128 302
rect 25971 272 26128 282
rect 25971 271 26006 272
rect 25971 250 26002 271
rect 26189 250 26225 360
rect 26244 359 26281 360
rect 26340 359 26377 360
rect 26300 300 26390 306
rect 26300 280 26309 300
rect 26329 298 26390 300
rect 26329 280 26354 298
rect 26300 278 26354 280
rect 26374 278 26390 298
rect 26300 272 26390 278
rect 25814 249 25851 250
rect 23735 243 23903 245
rect 23459 217 23903 243
rect 23569 214 23609 217
rect 23735 216 23903 217
rect 25813 240 25851 249
rect 25813 220 25822 240
rect 25842 220 25851 240
rect 25813 212 25851 220
rect 25917 244 26002 250
rect 26032 249 26069 250
rect 25917 224 25925 244
rect 25945 224 26002 244
rect 25917 216 26002 224
rect 26031 240 26069 249
rect 26031 220 26040 240
rect 26060 220 26069 240
rect 25917 215 25953 216
rect 26031 212 26069 220
rect 26135 244 26279 250
rect 26135 224 26143 244
rect 26163 242 26251 244
rect 26163 224 26195 242
rect 26135 221 26195 224
rect 26218 224 26251 242
rect 26271 224 26279 244
rect 26218 221 26279 224
rect 26135 216 26279 221
rect 26135 215 26171 216
rect 26243 215 26279 216
rect 26345 249 26382 250
rect 26345 248 26383 249
rect 26345 240 26409 248
rect 26345 220 26354 240
rect 26374 226 26409 240
rect 26429 226 26432 246
rect 26374 221 26432 226
rect 26374 220 26409 221
rect 25814 183 25851 212
rect 25815 181 25851 183
rect 25815 159 26006 181
rect 26032 180 26069 212
rect 26345 208 26409 220
rect 26449 182 26476 360
rect 27559 354 27618 374
rect 27638 354 27677 374
rect 27697 354 27708 374
rect 27559 346 27708 354
rect 27775 377 27932 384
rect 27775 357 27895 377
rect 27915 357 27932 377
rect 27775 347 27932 357
rect 27775 346 27810 347
rect 27775 325 27806 346
rect 27993 325 28029 435
rect 28048 434 28085 435
rect 28144 434 28181 435
rect 28104 375 28194 381
rect 28104 355 28113 375
rect 28133 373 28194 375
rect 28133 355 28158 373
rect 28104 353 28158 355
rect 28178 353 28194 373
rect 28104 347 28194 353
rect 27618 324 27655 325
rect 27617 315 27655 324
rect 27617 295 27626 315
rect 27646 295 27655 315
rect 27617 287 27655 295
rect 27721 319 27806 325
rect 27836 324 27873 325
rect 27721 299 27729 319
rect 27749 299 27806 319
rect 27721 291 27806 299
rect 27835 315 27873 324
rect 27835 295 27844 315
rect 27864 295 27873 315
rect 27721 290 27757 291
rect 27835 287 27873 295
rect 27939 320 28083 325
rect 27939 319 28000 320
rect 27939 299 27947 319
rect 27967 299 28000 319
rect 27939 296 28000 299
rect 28023 319 28083 320
rect 28023 299 28055 319
rect 28075 299 28083 319
rect 28023 296 28083 299
rect 27939 291 28083 296
rect 27939 290 27975 291
rect 28047 290 28083 291
rect 28149 324 28186 325
rect 28149 323 28187 324
rect 28149 315 28213 323
rect 28149 295 28158 315
rect 28178 301 28213 315
rect 28233 301 28236 321
rect 28178 296 28236 301
rect 28178 295 28213 296
rect 27618 258 27655 287
rect 27619 256 27655 258
rect 27619 234 27810 256
rect 27836 255 27873 287
rect 28149 283 28213 295
rect 28253 257 28280 435
rect 30112 390 30149 461
rect 30330 460 30671 461
rect 30264 400 30295 401
rect 30112 370 30121 390
rect 30141 370 30149 390
rect 30112 360 30149 370
rect 30208 390 30295 400
rect 30208 370 30217 390
rect 30237 370 30295 390
rect 30208 361 30295 370
rect 30208 360 30245 361
rect 30264 310 30295 361
rect 30330 390 30367 460
rect 30633 459 30670 460
rect 31987 457 31996 477
rect 32016 457 32024 477
rect 31987 447 32024 457
rect 32083 477 32170 487
rect 32083 457 32092 477
rect 32112 457 32170 477
rect 32083 448 32170 457
rect 32083 447 32120 448
rect 30482 400 30518 401
rect 30330 370 30339 390
rect 30359 370 30367 390
rect 30330 360 30367 370
rect 30426 390 30574 400
rect 30674 397 30796 399
rect 30426 370 30435 390
rect 30455 370 30545 390
rect 30565 370 30574 390
rect 30426 361 30574 370
rect 30632 395 30796 397
rect 32139 397 32170 448
rect 32205 477 32242 547
rect 32508 546 32545 547
rect 32357 487 32393 488
rect 32205 457 32214 477
rect 32234 457 32242 477
rect 32205 447 32242 457
rect 32301 477 32449 487
rect 32549 484 32710 486
rect 32301 457 32310 477
rect 32330 457 32420 477
rect 32440 457 32449 477
rect 32301 448 32449 457
rect 32507 479 32710 484
rect 32507 477 32680 479
rect 32507 457 32516 477
rect 32536 459 32680 477
rect 32700 459 32710 479
rect 32536 457 32710 459
rect 32507 450 32710 457
rect 32507 448 32645 450
rect 32301 447 32338 448
rect 30632 392 30835 395
rect 32031 394 32072 395
rect 30632 390 30805 392
rect 30632 370 30641 390
rect 30661 372 30805 390
rect 30825 372 30835 392
rect 30661 370 30835 372
rect 30632 363 30835 370
rect 31923 387 32072 394
rect 31923 367 31982 387
rect 32002 367 32041 387
rect 32061 367 32072 387
rect 30632 361 30770 363
rect 30426 360 30463 361
rect 30156 307 30197 308
rect 30048 300 30197 307
rect 30048 280 30107 300
rect 30127 280 30166 300
rect 30186 280 30197 300
rect 30048 272 30197 280
rect 30264 303 30421 310
rect 30264 283 30384 303
rect 30404 283 30421 303
rect 30264 273 30421 283
rect 30264 272 30299 273
rect 28112 255 28280 257
rect 27836 229 28280 255
rect 30264 251 30295 272
rect 30482 251 30518 361
rect 30537 360 30574 361
rect 30633 360 30670 361
rect 30593 301 30683 307
rect 30593 281 30602 301
rect 30622 299 30683 301
rect 30622 281 30647 299
rect 30593 279 30647 281
rect 30667 279 30683 299
rect 30593 273 30683 279
rect 30107 250 30144 251
rect 27946 226 27986 229
rect 28112 228 28280 229
rect 30106 241 30144 250
rect 30106 221 30115 241
rect 30135 221 30144 241
rect 30106 213 30144 221
rect 30210 245 30295 251
rect 30325 250 30362 251
rect 30210 225 30218 245
rect 30238 225 30295 245
rect 30210 217 30295 225
rect 30324 241 30362 250
rect 30324 221 30333 241
rect 30353 221 30362 241
rect 30210 216 30246 217
rect 30324 213 30362 221
rect 30428 245 30572 251
rect 30428 225 30436 245
rect 30456 225 30488 245
rect 30428 223 30488 225
rect 30509 225 30544 245
rect 30564 225 30572 245
rect 30509 223 30572 225
rect 30428 217 30572 223
rect 30428 216 30464 217
rect 30536 216 30572 217
rect 30638 250 30675 251
rect 30638 249 30676 250
rect 30638 241 30702 249
rect 30638 221 30647 241
rect 30667 227 30702 241
rect 30722 227 30725 247
rect 30667 222 30725 227
rect 30667 221 30702 222
rect 30107 184 30144 213
rect 26308 180 26476 182
rect 21860 156 22028 158
rect 21584 130 22028 156
rect 26032 154 26476 180
rect 30108 182 30144 184
rect 30108 160 30299 182
rect 30325 181 30362 213
rect 30638 209 30702 221
rect 30742 183 30769 361
rect 31923 359 32072 367
rect 32139 390 32296 397
rect 32139 370 32259 390
rect 32279 370 32296 390
rect 32139 360 32296 370
rect 32139 359 32174 360
rect 32139 338 32170 359
rect 32357 338 32393 448
rect 32412 447 32449 448
rect 32508 447 32545 448
rect 32468 388 32558 394
rect 32468 368 32477 388
rect 32497 386 32558 388
rect 32497 368 32522 386
rect 32468 366 32522 368
rect 32542 366 32558 386
rect 32468 360 32558 366
rect 31982 337 32019 338
rect 31981 328 32019 337
rect 31981 308 31990 328
rect 32010 308 32019 328
rect 31981 300 32019 308
rect 32085 332 32170 338
rect 32200 337 32237 338
rect 32085 312 32093 332
rect 32113 312 32170 332
rect 32085 304 32170 312
rect 32199 328 32237 337
rect 32199 308 32208 328
rect 32228 308 32237 328
rect 32085 303 32121 304
rect 32199 300 32237 308
rect 32303 334 32447 338
rect 32303 332 32367 334
rect 32303 312 32311 332
rect 32331 312 32367 332
rect 32303 310 32367 312
rect 32390 332 32447 334
rect 32390 312 32419 332
rect 32439 312 32447 332
rect 32390 310 32447 312
rect 32303 304 32447 310
rect 32303 303 32339 304
rect 32411 303 32447 304
rect 32513 337 32550 338
rect 32513 336 32551 337
rect 32513 328 32577 336
rect 32513 308 32522 328
rect 32542 314 32577 328
rect 32597 314 32600 334
rect 32542 309 32600 314
rect 32542 308 32577 309
rect 31982 271 32019 300
rect 31983 269 32019 271
rect 31983 247 32174 269
rect 32200 268 32237 300
rect 32513 296 32577 308
rect 32617 270 32644 448
rect 32476 268 32644 270
rect 32200 242 32644 268
rect 32310 239 32350 242
rect 32476 241 32644 242
rect 30601 181 30769 183
rect 30325 155 30769 181
rect 26142 151 26182 154
rect 26308 153 26476 154
rect 30435 152 30475 155
rect 30601 154 30769 155
rect 21694 127 21734 130
rect 21860 129 22028 130
rect 17427 105 17595 107
rect 17151 79 17595 105
rect 17261 76 17301 79
rect 17427 78 17595 79
<< viali >>
rect 2883 8916 2907 8938
rect 2488 8668 2509 8687
rect 1035 8617 1055 8637
rect 419 8431 439 8451
rect 959 8430 979 8450
rect 801 8376 821 8396
rect 1014 8378 1034 8398
rect 1833 8433 1853 8453
rect 1217 8247 1237 8267
rect 1036 8205 1056 8225
rect 1757 8246 1777 8266
rect 1598 8193 1619 8212
rect 1812 8194 1832 8214
rect 7247 8929 7271 8951
rect 3425 8828 3445 8848
rect 3647 8826 3667 8846
rect 3480 8776 3500 8796
rect 4020 8775 4040 8795
rect 2628 8600 2648 8620
rect 2840 8605 2859 8623
rect 2683 8548 2703 8568
rect 3404 8589 3424 8609
rect 3223 8547 3243 8567
rect 2607 8361 2627 8381
rect 3426 8416 3446 8436
rect 3639 8418 3659 8438
rect 6852 8681 6873 8700
rect 5399 8630 5419 8650
rect 4783 8444 4803 8464
rect 5323 8443 5343 8463
rect 3481 8364 3501 8384
rect 4021 8363 4041 8383
rect 420 8019 440 8039
rect 960 8018 980 8038
rect 793 7968 813 7988
rect 1015 7966 1035 7986
rect 2529 8190 2549 8210
rect 2740 8197 2759 8214
rect 2584 8138 2604 8158
rect 3405 8177 3425 8197
rect 3124 8137 3144 8157
rect 5165 8389 5185 8409
rect 5378 8391 5398 8411
rect 6197 8446 6217 8466
rect 5581 8260 5601 8280
rect 5400 8218 5420 8238
rect 6121 8259 6141 8279
rect 5962 8206 5983 8225
rect 6176 8207 6196 8227
rect 7789 8841 7809 8861
rect 8011 8839 8031 8859
rect 11624 8941 11648 8963
rect 7844 8789 7864 8809
rect 8384 8788 8404 8808
rect 6992 8613 7012 8633
rect 7204 8618 7223 8636
rect 7047 8561 7067 8581
rect 7768 8602 7788 8622
rect 7587 8560 7607 8580
rect 6971 8374 6991 8394
rect 7790 8429 7810 8449
rect 8003 8431 8023 8451
rect 11229 8693 11250 8712
rect 9776 8642 9796 8662
rect 9160 8456 9180 8476
rect 9700 8455 9720 8475
rect 7845 8377 7865 8397
rect 8385 8376 8405 8396
rect 4784 8032 4804 8052
rect 2508 7951 2528 7971
rect 5324 8031 5344 8051
rect 5157 7981 5177 8001
rect 5379 7979 5399 7999
rect 1553 7876 1577 7898
rect 2866 7898 2890 7920
rect 1915 7825 1935 7845
rect 1299 7639 1319 7659
rect 1018 7599 1038 7619
rect 1839 7638 1859 7658
rect 1682 7586 1703 7605
rect 1894 7586 1914 7606
rect 6893 8203 6913 8223
rect 7104 8210 7123 8227
rect 6948 8151 6968 8171
rect 7769 8190 7789 8210
rect 7488 8150 7508 8170
rect 9542 8401 9562 8421
rect 9755 8403 9775 8423
rect 10574 8458 10594 8478
rect 9958 8272 9978 8292
rect 9777 8230 9797 8250
rect 10498 8271 10518 8291
rect 10339 8218 10360 8237
rect 10553 8219 10573 8239
rect 15988 8954 16012 8976
rect 12166 8853 12186 8873
rect 12388 8851 12408 8871
rect 12221 8801 12241 8821
rect 12761 8800 12781 8820
rect 11369 8625 11389 8645
rect 11581 8630 11600 8648
rect 11424 8573 11444 8593
rect 12145 8614 12165 8634
rect 11964 8572 11984 8592
rect 11348 8386 11368 8406
rect 12167 8441 12187 8461
rect 12380 8443 12400 8463
rect 15593 8706 15614 8725
rect 14140 8655 14160 8675
rect 13524 8469 13544 8489
rect 14064 8468 14084 8488
rect 12222 8389 12242 8409
rect 12762 8388 12782 8408
rect 9161 8044 9181 8064
rect 6872 7964 6892 7984
rect 9701 8043 9721 8063
rect 9534 7993 9554 8013
rect 9756 7991 9776 8011
rect 5917 7889 5941 7911
rect 7230 7911 7254 7933
rect 3408 7810 3428 7830
rect 3630 7808 3650 7828
rect 3463 7758 3483 7778
rect 6279 7838 6299 7858
rect 4003 7757 4023 7777
rect 402 7413 422 7433
rect 942 7412 962 7432
rect 784 7358 804 7378
rect 997 7360 1017 7380
rect 1816 7415 1836 7435
rect 1200 7229 1220 7249
rect 1019 7187 1039 7207
rect 1740 7228 1760 7248
rect 1584 7173 1603 7191
rect 1795 7176 1815 7196
rect 403 7001 423 7021
rect 943 7000 963 7020
rect 776 6950 796 6970
rect 998 6948 1018 6968
rect 2611 7582 2631 7602
rect 2824 7584 2845 7603
rect 2666 7530 2686 7550
rect 3387 7571 3407 7591
rect 3206 7529 3226 7549
rect 2431 7431 2453 7449
rect 2590 7343 2610 7363
rect 3409 7398 3429 7418
rect 3622 7400 3642 7420
rect 5663 7652 5683 7672
rect 5382 7612 5402 7632
rect 6203 7651 6223 7671
rect 6046 7599 6067 7618
rect 6258 7599 6278 7619
rect 11270 8215 11290 8235
rect 11481 8222 11500 8239
rect 11325 8163 11345 8183
rect 12146 8202 12166 8222
rect 11865 8162 11885 8182
rect 13906 8414 13926 8434
rect 14119 8416 14139 8436
rect 14938 8471 14958 8491
rect 14322 8285 14342 8305
rect 14141 8243 14161 8263
rect 14862 8284 14882 8304
rect 14703 8231 14724 8250
rect 14917 8232 14937 8252
rect 20254 8928 20278 8950
rect 16530 8866 16550 8886
rect 16752 8864 16772 8884
rect 16585 8814 16605 8834
rect 17125 8813 17145 8833
rect 15733 8638 15753 8658
rect 15945 8643 15964 8661
rect 15788 8586 15808 8606
rect 16509 8627 16529 8647
rect 16328 8585 16348 8605
rect 15712 8399 15732 8419
rect 16531 8454 16551 8474
rect 16744 8456 16764 8476
rect 19859 8680 19880 8699
rect 18406 8629 18426 8649
rect 16586 8402 16606 8422
rect 17790 8443 17810 8463
rect 17126 8401 17146 8421
rect 18330 8442 18350 8462
rect 13525 8057 13545 8077
rect 11249 7976 11269 7996
rect 14065 8056 14085 8076
rect 13898 8006 13918 8026
rect 14120 8004 14140 8024
rect 10294 7901 10318 7923
rect 11607 7923 11631 7945
rect 7772 7823 7792 7843
rect 7994 7821 8014 7841
rect 7827 7771 7847 7791
rect 10656 7850 10676 7870
rect 8367 7770 8387 7790
rect 4766 7426 4786 7446
rect 5306 7425 5326 7445
rect 3464 7346 3484 7366
rect 4004 7345 4024 7365
rect 2232 7235 2256 7257
rect 1934 7109 1955 7128
rect 1536 6858 1560 6880
rect 1961 6805 1981 6825
rect 1345 6619 1365 6639
rect 998 6581 1018 6601
rect 1885 6618 1905 6638
rect 1729 6565 1747 6583
rect 1940 6566 1960 6586
rect 382 6395 402 6415
rect 922 6394 942 6414
rect 764 6340 784 6360
rect 977 6342 997 6362
rect 1796 6397 1816 6417
rect 1180 6211 1200 6231
rect 999 6169 1019 6189
rect 1720 6210 1740 6230
rect 1561 6157 1582 6176
rect 1775 6158 1795 6178
rect 383 5983 403 6003
rect 923 5982 943 6002
rect 756 5932 776 5952
rect 978 5930 998 5950
rect 1516 5840 1540 5862
rect 1878 5789 1898 5809
rect 1262 5603 1282 5623
rect 981 5563 1001 5583
rect 1802 5602 1822 5622
rect 1647 5546 1666 5563
rect 1857 5550 1877 5570
rect 365 5377 385 5397
rect 905 5376 925 5396
rect 747 5322 767 5342
rect 960 5324 980 5344
rect 1959 5479 1981 5497
rect 1779 5379 1799 5399
rect 1163 5193 1183 5213
rect 982 5151 1002 5171
rect 1703 5192 1723 5212
rect 1547 5137 1566 5155
rect 1758 5140 1778 5160
rect 366 4965 386 4985
rect 906 4964 926 4984
rect 739 4914 759 4934
rect 961 4912 981 4932
rect 2446 7174 2466 7194
rect 2657 7172 2680 7194
rect 2501 7122 2521 7142
rect 3388 7159 3408 7179
rect 3041 7121 3061 7141
rect 5148 7371 5168 7391
rect 5361 7373 5381 7393
rect 6180 7428 6200 7448
rect 5564 7242 5584 7262
rect 5383 7200 5403 7220
rect 6104 7241 6124 7261
rect 5948 7186 5967 7204
rect 6159 7189 6179 7209
rect 2425 6935 2445 6955
rect 4767 7014 4787 7034
rect 5307 7013 5327 7033
rect 5140 6963 5160 6983
rect 5362 6961 5382 6981
rect 2846 6880 2870 6902
rect 2451 6632 2472 6651
rect 6975 7595 6995 7615
rect 7188 7597 7209 7616
rect 7030 7543 7050 7563
rect 7751 7584 7771 7604
rect 7570 7542 7590 7562
rect 6795 7444 6817 7462
rect 6954 7356 6974 7376
rect 7773 7411 7793 7431
rect 7986 7413 8006 7433
rect 10040 7664 10060 7684
rect 9759 7624 9779 7644
rect 10580 7663 10600 7683
rect 10423 7611 10444 7630
rect 10635 7611 10655 7631
rect 15634 8228 15654 8248
rect 15845 8235 15864 8252
rect 15689 8176 15709 8196
rect 16510 8215 16530 8235
rect 16229 8175 16249 8195
rect 18172 8388 18192 8408
rect 18385 8390 18405 8410
rect 19204 8445 19224 8465
rect 18588 8259 18608 8279
rect 18407 8217 18427 8237
rect 19128 8258 19148 8278
rect 18969 8205 18990 8224
rect 19183 8206 19203 8226
rect 24618 8941 24642 8963
rect 20796 8840 20816 8860
rect 21018 8838 21038 8858
rect 20851 8788 20871 8808
rect 21391 8787 21411 8807
rect 19999 8612 20019 8632
rect 20211 8617 20230 8635
rect 20054 8560 20074 8580
rect 20775 8601 20795 8621
rect 20594 8559 20614 8579
rect 19978 8373 19998 8393
rect 20797 8428 20817 8448
rect 21010 8430 21030 8450
rect 24223 8693 24244 8712
rect 22770 8642 22790 8662
rect 22154 8456 22174 8476
rect 22694 8455 22714 8475
rect 20852 8376 20872 8396
rect 21392 8375 21412 8395
rect 15613 7989 15633 8009
rect 17791 8031 17811 8051
rect 18331 8030 18351 8050
rect 14658 7914 14682 7936
rect 15971 7936 15995 7958
rect 12149 7835 12169 7855
rect 12371 7833 12391 7853
rect 12204 7783 12224 7803
rect 15020 7863 15040 7883
rect 12744 7782 12764 7802
rect 9143 7438 9163 7458
rect 9683 7437 9703 7457
rect 7828 7359 7848 7379
rect 8368 7358 8388 7378
rect 6596 7248 6620 7270
rect 6298 7122 6319 7141
rect 5900 6871 5924 6893
rect 3388 6792 3408 6812
rect 3610 6790 3630 6810
rect 3443 6740 3463 6760
rect 3983 6739 4003 6759
rect 6325 6818 6345 6838
rect 2591 6564 2611 6584
rect 2803 6569 2822 6587
rect 2646 6512 2666 6532
rect 3367 6553 3387 6573
rect 3186 6511 3206 6531
rect 2570 6325 2590 6345
rect 3389 6380 3409 6400
rect 3602 6382 3622 6402
rect 5709 6632 5729 6652
rect 5362 6594 5382 6614
rect 6249 6631 6269 6651
rect 6093 6578 6111 6596
rect 6304 6579 6324 6599
rect 4746 6408 4766 6428
rect 5286 6407 5306 6427
rect 3444 6328 3464 6348
rect 3984 6327 4004 6347
rect 2492 6154 2512 6174
rect 2703 6155 2724 6174
rect 2547 6102 2567 6122
rect 3368 6141 3388 6161
rect 3087 6101 3107 6121
rect 5128 6353 5148 6373
rect 5341 6355 5361 6375
rect 6160 6410 6180 6430
rect 5544 6224 5564 6244
rect 5363 6182 5383 6202
rect 6084 6223 6104 6243
rect 5925 6170 5946 6189
rect 6139 6171 6159 6191
rect 4747 5996 4767 6016
rect 2471 5915 2491 5935
rect 5287 5995 5307 6015
rect 5120 5945 5140 5965
rect 5342 5943 5362 5963
rect 2829 5862 2853 5884
rect 5880 5853 5904 5875
rect 3371 5774 3391 5794
rect 3593 5772 3613 5792
rect 3426 5722 3446 5742
rect 6242 5802 6262 5822
rect 3966 5721 3986 5741
rect 2574 5546 2594 5566
rect 2787 5548 2808 5567
rect 2629 5494 2649 5514
rect 3350 5535 3370 5555
rect 3169 5493 3189 5513
rect 2553 5307 2573 5327
rect 3372 5362 3392 5382
rect 3585 5364 3605 5384
rect 5626 5616 5646 5636
rect 5345 5576 5365 5596
rect 6166 5615 6186 5635
rect 6011 5559 6030 5576
rect 6221 5563 6241 5583
rect 4729 5390 4749 5410
rect 5269 5389 5289 5409
rect 3427 5310 3447 5330
rect 3967 5309 3987 5329
rect 1897 5073 1918 5092
rect 2270 5140 2290 5160
rect 2482 5139 2508 5165
rect 2325 5088 2345 5108
rect 3351 5123 3371 5143
rect 2865 5087 2885 5107
rect 5111 5335 5131 5355
rect 5324 5337 5344 5357
rect 6323 5492 6345 5510
rect 6143 5392 6163 5412
rect 5527 5206 5547 5226
rect 5346 5164 5366 5184
rect 6067 5205 6087 5225
rect 5911 5150 5930 5168
rect 6122 5153 6142 5173
rect 2249 4901 2269 4921
rect 4730 4978 4750 4998
rect 5270 4977 5290 4997
rect 5103 4927 5123 4947
rect 5325 4925 5345 4945
rect 1499 4822 1523 4844
rect 2810 4844 2834 4866
rect 2064 4767 2084 4787
rect 1448 4581 1468 4601
rect 962 4545 982 4565
rect 1988 4580 2008 4600
rect 1826 4517 1849 4540
rect 2043 4528 2063 4548
rect 2415 4596 2436 4615
rect 346 4359 366 4379
rect 886 4358 906 4378
rect 728 4304 748 4324
rect 941 4306 961 4326
rect 1760 4361 1780 4381
rect 1144 4175 1164 4195
rect 963 4133 983 4153
rect 1684 4174 1704 4194
rect 1525 4121 1546 4140
rect 1739 4122 1759 4142
rect 347 3947 367 3967
rect 887 3946 907 3966
rect 720 3896 740 3916
rect 942 3894 962 3914
rect 1480 3804 1504 3826
rect 1842 3753 1862 3773
rect 1226 3567 1246 3587
rect 945 3527 965 3547
rect 1766 3566 1786 3586
rect 1609 3514 1630 3533
rect 1821 3514 1841 3534
rect 329 3341 349 3361
rect 869 3340 889 3360
rect 711 3286 731 3306
rect 924 3288 944 3308
rect 1743 3343 1763 3363
rect 1127 3157 1147 3177
rect 946 3115 966 3135
rect 1667 3156 1687 3176
rect 1511 3101 1530 3119
rect 1722 3104 1742 3124
rect 330 2929 350 2949
rect 870 2928 890 2948
rect 703 2878 723 2898
rect 925 2876 945 2896
rect 1861 3037 1882 3056
rect 1463 2786 1487 2808
rect 1888 2733 1908 2753
rect 1272 2547 1292 2567
rect 925 2509 945 2529
rect 1812 2546 1832 2566
rect 1653 2494 1676 2516
rect 1867 2494 1887 2514
rect 6810 7187 6830 7207
rect 7021 7185 7044 7207
rect 6865 7135 6885 7155
rect 7752 7172 7772 7192
rect 7405 7134 7425 7154
rect 9525 7383 9545 7403
rect 9738 7385 9758 7405
rect 10557 7440 10577 7460
rect 9941 7254 9961 7274
rect 9760 7212 9780 7232
rect 10481 7253 10501 7273
rect 10325 7198 10344 7216
rect 10536 7201 10556 7221
rect 6789 6948 6809 6968
rect 9144 7026 9164 7046
rect 9684 7025 9704 7045
rect 9517 6975 9537 6995
rect 9739 6973 9759 6993
rect 7210 6893 7234 6915
rect 6815 6645 6836 6664
rect 11352 7607 11372 7627
rect 11565 7609 11586 7628
rect 11407 7555 11427 7575
rect 12128 7596 12148 7616
rect 11947 7554 11967 7574
rect 11172 7456 11194 7474
rect 11331 7368 11351 7388
rect 12150 7423 12170 7443
rect 12363 7425 12383 7445
rect 14404 7677 14424 7697
rect 14123 7637 14143 7657
rect 14944 7676 14964 7696
rect 14787 7624 14808 7643
rect 14999 7624 15019 7644
rect 18164 7980 18184 8000
rect 18386 7978 18406 7998
rect 16513 7848 16533 7868
rect 16735 7846 16755 7866
rect 19900 8202 19920 8222
rect 20111 8209 20130 8226
rect 19955 8150 19975 8170
rect 20776 8189 20796 8209
rect 20495 8149 20515 8169
rect 22536 8401 22556 8421
rect 22749 8403 22769 8423
rect 23568 8458 23588 8478
rect 22952 8272 22972 8292
rect 22771 8230 22791 8250
rect 23492 8271 23512 8291
rect 23333 8218 23354 8237
rect 23547 8219 23567 8239
rect 25160 8853 25180 8873
rect 25382 8851 25402 8871
rect 28995 8953 29019 8975
rect 25215 8801 25235 8821
rect 25755 8800 25775 8820
rect 24363 8625 24383 8645
rect 24575 8630 24594 8648
rect 24418 8573 24438 8593
rect 25139 8614 25159 8634
rect 24958 8572 24978 8592
rect 24342 8386 24362 8406
rect 25161 8441 25181 8461
rect 25374 8443 25394 8463
rect 28600 8705 28621 8724
rect 27147 8654 27167 8674
rect 26531 8468 26551 8488
rect 27071 8467 27091 8487
rect 25216 8389 25236 8409
rect 25756 8388 25776 8408
rect 22155 8044 22175 8064
rect 19879 7963 19899 7983
rect 22695 8043 22715 8063
rect 22528 7993 22548 8013
rect 22750 7991 22770 8011
rect 18924 7888 18948 7910
rect 20237 7910 20261 7932
rect 16568 7796 16588 7816
rect 17108 7795 17128 7815
rect 19286 7837 19306 7857
rect 13507 7451 13527 7471
rect 14047 7450 14067 7470
rect 12205 7371 12225 7391
rect 12745 7370 12765 7390
rect 10973 7260 10997 7282
rect 10675 7134 10696 7153
rect 10277 6883 10301 6905
rect 7752 6805 7772 6825
rect 7974 6803 7994 6823
rect 7807 6753 7827 6773
rect 8347 6752 8367 6772
rect 10702 6830 10722 6850
rect 6955 6577 6975 6597
rect 7167 6582 7186 6600
rect 7010 6525 7030 6545
rect 7731 6566 7751 6586
rect 7550 6524 7570 6544
rect 6934 6338 6954 6358
rect 7753 6393 7773 6413
rect 7966 6395 7986 6415
rect 10086 6644 10106 6664
rect 9739 6606 9759 6626
rect 10626 6643 10646 6663
rect 10470 6590 10488 6608
rect 10681 6591 10701 6611
rect 9123 6420 9143 6440
rect 9663 6419 9683 6439
rect 7808 6341 7828 6361
rect 8348 6340 8368 6360
rect 6856 6167 6876 6187
rect 7067 6168 7088 6187
rect 6911 6115 6931 6135
rect 7732 6154 7752 6174
rect 7451 6114 7471 6134
rect 9505 6365 9525 6385
rect 9718 6367 9738 6387
rect 10537 6422 10557 6442
rect 9921 6236 9941 6256
rect 9740 6194 9760 6214
rect 10461 6235 10481 6255
rect 10302 6182 10323 6201
rect 10516 6183 10536 6203
rect 9124 6008 9144 6028
rect 6835 5928 6855 5948
rect 9664 6007 9684 6027
rect 9497 5957 9517 5977
rect 9719 5955 9739 5975
rect 7193 5875 7217 5897
rect 10257 5865 10281 5887
rect 7735 5787 7755 5807
rect 7957 5785 7977 5805
rect 7790 5735 7810 5755
rect 10619 5814 10639 5834
rect 8330 5734 8350 5754
rect 6938 5559 6958 5579
rect 7151 5561 7172 5580
rect 6993 5507 7013 5527
rect 7714 5548 7734 5568
rect 7533 5506 7553 5526
rect 6917 5320 6937 5340
rect 7736 5375 7756 5395
rect 7949 5377 7969 5397
rect 10003 5628 10023 5648
rect 9722 5588 9742 5608
rect 10543 5627 10563 5647
rect 10388 5571 10407 5588
rect 10598 5575 10618 5595
rect 9106 5402 9126 5422
rect 9646 5401 9666 5421
rect 7791 5323 7811 5343
rect 8331 5322 8351 5342
rect 6261 5086 6282 5105
rect 6634 5153 6654 5173
rect 6846 5152 6872 5178
rect 6689 5101 6709 5121
rect 7715 5136 7735 5156
rect 7229 5100 7249 5120
rect 9488 5347 9508 5367
rect 9701 5349 9721 5369
rect 10700 5504 10722 5522
rect 10520 5404 10540 5424
rect 9904 5218 9924 5238
rect 9723 5176 9743 5196
rect 10444 5217 10464 5237
rect 10288 5162 10307 5180
rect 10499 5165 10519 5185
rect 6613 4914 6633 4934
rect 9107 4990 9127 5010
rect 9647 4989 9667 5009
rect 9480 4939 9500 4959
rect 9702 4937 9722 4957
rect 5863 4835 5887 4857
rect 7174 4857 7198 4879
rect 3352 4756 3372 4776
rect 3574 4754 3594 4774
rect 3407 4704 3427 4724
rect 3947 4703 3967 4723
rect 6428 4780 6448 4800
rect 2555 4528 2575 4548
rect 2767 4533 2786 4551
rect 2610 4476 2630 4496
rect 3331 4517 3351 4537
rect 3150 4475 3170 4495
rect 2534 4289 2554 4309
rect 2352 4191 2374 4209
rect 3353 4344 3373 4364
rect 3566 4346 3586 4366
rect 5812 4594 5832 4614
rect 5326 4558 5346 4578
rect 6352 4593 6372 4613
rect 6190 4530 6213 4553
rect 6407 4541 6427 4561
rect 6779 4609 6800 4628
rect 4710 4372 4730 4392
rect 5250 4371 5270 4391
rect 3408 4292 3428 4312
rect 3948 4291 3968 4311
rect 2456 4118 2476 4138
rect 2667 4125 2686 4142
rect 2511 4066 2531 4086
rect 3332 4105 3352 4125
rect 3051 4065 3071 4085
rect 5092 4317 5112 4337
rect 5305 4319 5325 4339
rect 6124 4374 6144 4394
rect 5508 4188 5528 4208
rect 5327 4146 5347 4166
rect 6048 4187 6068 4207
rect 5889 4134 5910 4153
rect 6103 4135 6123 4155
rect 4711 3960 4731 3980
rect 2435 3879 2455 3899
rect 5251 3959 5271 3979
rect 5084 3909 5104 3929
rect 5306 3907 5326 3927
rect 2793 3826 2817 3848
rect 5844 3817 5868 3839
rect 3335 3738 3355 3758
rect 3557 3736 3577 3756
rect 3390 3686 3410 3706
rect 6206 3766 6226 3786
rect 3930 3685 3950 3705
rect 2538 3510 2558 3530
rect 2751 3512 2772 3531
rect 2593 3458 2613 3478
rect 3314 3499 3334 3519
rect 3133 3457 3153 3477
rect 2517 3271 2537 3291
rect 3336 3326 3356 3346
rect 3549 3328 3569 3348
rect 5590 3580 5610 3600
rect 5309 3540 5329 3560
rect 6130 3579 6150 3599
rect 5973 3527 5994 3546
rect 6185 3527 6205 3547
rect 4693 3354 4713 3374
rect 5233 3353 5253 3373
rect 3391 3274 3411 3294
rect 3931 3273 3951 3293
rect 2373 3102 2393 3122
rect 2586 3105 2604 3123
rect 2428 3050 2448 3070
rect 3315 3087 3335 3107
rect 2968 3049 2988 3069
rect 5075 3299 5095 3319
rect 5288 3301 5308 3321
rect 6107 3356 6127 3376
rect 5491 3170 5511 3190
rect 5310 3128 5330 3148
rect 6031 3169 6051 3189
rect 5875 3114 5894 3132
rect 6086 3117 6106 3137
rect 2352 2863 2372 2883
rect 4694 2942 4714 2962
rect 5234 2941 5254 2961
rect 5067 2891 5087 2911
rect 5289 2889 5309 2909
rect 2773 2808 2797 2830
rect 2378 2560 2399 2579
rect 2077 2431 2101 2453
rect 309 2323 329 2343
rect 849 2322 869 2342
rect 691 2268 711 2288
rect 904 2270 924 2290
rect 1723 2325 1743 2345
rect 1880 2239 1902 2257
rect 1107 2139 1127 2159
rect 926 2097 946 2117
rect 1647 2138 1667 2158
rect 1488 2085 1509 2104
rect 1702 2086 1722 2106
rect 6225 3050 6246 3069
rect 5827 2799 5851 2821
rect 3315 2720 3335 2740
rect 3537 2718 3557 2738
rect 3370 2668 3390 2688
rect 3910 2667 3930 2687
rect 6252 2746 6272 2766
rect 2518 2492 2538 2512
rect 2730 2497 2749 2515
rect 2573 2440 2593 2460
rect 3294 2481 3314 2501
rect 3113 2439 3133 2459
rect 2497 2253 2517 2273
rect 3316 2308 3336 2328
rect 3529 2310 3549 2330
rect 5636 2560 5656 2580
rect 5289 2522 5309 2542
rect 6176 2559 6196 2579
rect 6017 2507 6040 2529
rect 6231 2507 6251 2527
rect 11187 7199 11207 7219
rect 11398 7197 11421 7219
rect 11242 7147 11262 7167
rect 12129 7184 12149 7204
rect 11782 7146 11802 7166
rect 13889 7396 13909 7416
rect 14102 7398 14122 7418
rect 14921 7453 14941 7473
rect 14305 7267 14325 7287
rect 14124 7225 14144 7245
rect 14845 7266 14865 7286
rect 14689 7211 14708 7229
rect 14900 7214 14920 7234
rect 11166 6960 11186 6980
rect 13508 7039 13528 7059
rect 14048 7038 14068 7058
rect 13881 6988 13901 7008
rect 14103 6986 14123 7006
rect 11587 6905 11611 6927
rect 11192 6657 11213 6676
rect 15716 7620 15736 7640
rect 15929 7622 15950 7641
rect 15771 7568 15791 7588
rect 16492 7609 16512 7629
rect 16311 7567 16331 7587
rect 15536 7469 15558 7487
rect 15695 7381 15715 7401
rect 16514 7436 16534 7456
rect 16727 7438 16747 7458
rect 18670 7651 18690 7671
rect 18389 7611 18409 7631
rect 19210 7650 19230 7670
rect 19053 7598 19074 7617
rect 19265 7598 19285 7618
rect 24264 8215 24284 8235
rect 24475 8222 24494 8239
rect 24319 8163 24339 8183
rect 25140 8202 25160 8222
rect 24859 8162 24879 8182
rect 26913 8413 26933 8433
rect 27126 8415 27146 8435
rect 27945 8470 27965 8490
rect 27329 8284 27349 8304
rect 27148 8242 27168 8262
rect 27869 8283 27889 8303
rect 27710 8230 27731 8249
rect 27924 8231 27944 8251
rect 33359 8966 33383 8988
rect 29537 8865 29557 8885
rect 29759 8863 29779 8883
rect 29592 8813 29612 8833
rect 30132 8812 30152 8832
rect 28740 8637 28760 8657
rect 28952 8642 28971 8660
rect 28795 8585 28815 8605
rect 29516 8626 29536 8646
rect 29335 8584 29355 8604
rect 28719 8398 28739 8418
rect 29538 8453 29558 8473
rect 29751 8455 29771 8475
rect 32964 8718 32985 8737
rect 31511 8667 31531 8687
rect 30895 8481 30915 8501
rect 31435 8480 31455 8500
rect 29593 8401 29613 8421
rect 30133 8400 30153 8420
rect 26532 8056 26552 8076
rect 24243 7976 24263 7996
rect 27072 8055 27092 8075
rect 26905 8005 26925 8025
rect 27127 8003 27147 8023
rect 23288 7901 23312 7923
rect 24601 7923 24625 7945
rect 20779 7822 20799 7842
rect 21001 7820 21021 7840
rect 20834 7770 20854 7790
rect 23650 7850 23670 7870
rect 21374 7769 21394 7789
rect 16569 7384 16589 7404
rect 17773 7425 17793 7445
rect 17109 7383 17129 7403
rect 18313 7424 18333 7444
rect 15337 7273 15361 7295
rect 15039 7147 15060 7166
rect 14641 6896 14665 6918
rect 12129 6817 12149 6837
rect 12351 6815 12371 6835
rect 12184 6765 12204 6785
rect 12724 6764 12744 6784
rect 15066 6843 15086 6863
rect 11332 6589 11352 6609
rect 11544 6594 11563 6612
rect 11387 6537 11407 6557
rect 12108 6578 12128 6598
rect 11927 6536 11947 6556
rect 11311 6350 11331 6370
rect 12130 6405 12150 6425
rect 12343 6407 12363 6427
rect 14450 6657 14470 6677
rect 14103 6619 14123 6639
rect 14990 6656 15010 6676
rect 14834 6603 14852 6621
rect 15045 6604 15065 6624
rect 13487 6433 13507 6453
rect 14027 6432 14047 6452
rect 12185 6353 12205 6373
rect 12725 6352 12745 6372
rect 11233 6179 11253 6199
rect 11444 6180 11465 6199
rect 11288 6127 11308 6147
rect 12109 6166 12129 6186
rect 11828 6126 11848 6146
rect 13869 6378 13889 6398
rect 14082 6380 14102 6400
rect 14901 6435 14921 6455
rect 14285 6249 14305 6269
rect 14104 6207 14124 6227
rect 14825 6248 14845 6268
rect 14666 6195 14687 6214
rect 14880 6196 14900 6216
rect 13488 6021 13508 6041
rect 11212 5940 11232 5960
rect 14028 6020 14048 6040
rect 13861 5970 13881 5990
rect 14083 5968 14103 5988
rect 11570 5887 11594 5909
rect 14621 5878 14645 5900
rect 12112 5799 12132 5819
rect 12334 5797 12354 5817
rect 12167 5747 12187 5767
rect 14983 5827 15003 5847
rect 12707 5746 12727 5766
rect 11315 5571 11335 5591
rect 11528 5573 11549 5592
rect 11370 5519 11390 5539
rect 12091 5560 12111 5580
rect 11910 5518 11930 5538
rect 11294 5332 11314 5352
rect 12113 5387 12133 5407
rect 12326 5389 12346 5409
rect 14367 5641 14387 5661
rect 14086 5601 14106 5621
rect 14907 5640 14927 5660
rect 14752 5584 14771 5601
rect 14962 5588 14982 5608
rect 13470 5415 13490 5435
rect 14010 5414 14030 5434
rect 12168 5335 12188 5355
rect 12708 5334 12728 5354
rect 10638 5098 10659 5117
rect 11011 5165 11031 5185
rect 11223 5164 11249 5190
rect 11066 5113 11086 5133
rect 12092 5148 12112 5168
rect 11606 5112 11626 5132
rect 13852 5360 13872 5380
rect 14065 5362 14085 5382
rect 15064 5517 15086 5535
rect 14884 5417 14904 5437
rect 14268 5231 14288 5251
rect 14087 5189 14107 5209
rect 14808 5230 14828 5250
rect 14652 5175 14671 5193
rect 14863 5178 14883 5198
rect 10990 4926 11010 4946
rect 13471 5003 13491 5023
rect 14011 5002 14031 5022
rect 13844 4952 13864 4972
rect 14066 4950 14086 4970
rect 10240 4847 10264 4869
rect 11551 4869 11575 4891
rect 7716 4769 7736 4789
rect 7938 4767 7958 4787
rect 7771 4717 7791 4737
rect 8311 4716 8331 4736
rect 10805 4792 10825 4812
rect 6919 4541 6939 4561
rect 7131 4546 7150 4564
rect 6974 4489 6994 4509
rect 7695 4530 7715 4550
rect 7514 4488 7534 4508
rect 6898 4302 6918 4322
rect 6716 4204 6738 4222
rect 7717 4357 7737 4377
rect 7930 4359 7950 4379
rect 10189 4606 10209 4626
rect 9703 4570 9723 4590
rect 10729 4605 10749 4625
rect 10567 4542 10590 4565
rect 10784 4553 10804 4573
rect 11156 4621 11177 4640
rect 9087 4384 9107 4404
rect 9627 4383 9647 4403
rect 7772 4305 7792 4325
rect 8312 4304 8332 4324
rect 6820 4131 6840 4151
rect 7031 4138 7050 4155
rect 6875 4079 6895 4099
rect 7696 4118 7716 4138
rect 7415 4078 7435 4098
rect 9469 4329 9489 4349
rect 9682 4331 9702 4351
rect 10501 4386 10521 4406
rect 9885 4200 9905 4220
rect 9704 4158 9724 4178
rect 10425 4199 10445 4219
rect 10266 4146 10287 4165
rect 10480 4147 10500 4167
rect 9088 3972 9108 3992
rect 6799 3892 6819 3912
rect 9628 3971 9648 3991
rect 9461 3921 9481 3941
rect 9683 3919 9703 3939
rect 7157 3839 7181 3861
rect 10221 3829 10245 3851
rect 7699 3751 7719 3771
rect 7921 3749 7941 3769
rect 7754 3699 7774 3719
rect 10583 3778 10603 3798
rect 8294 3698 8314 3718
rect 6902 3523 6922 3543
rect 7115 3525 7136 3544
rect 6957 3471 6977 3491
rect 7678 3512 7698 3532
rect 7497 3470 7517 3490
rect 6881 3284 6901 3304
rect 7700 3339 7720 3359
rect 7913 3341 7933 3361
rect 9967 3592 9987 3612
rect 9686 3552 9706 3572
rect 10507 3591 10527 3611
rect 10350 3539 10371 3558
rect 10562 3539 10582 3559
rect 9070 3366 9090 3386
rect 9610 3365 9630 3385
rect 7755 3287 7775 3307
rect 8295 3286 8315 3306
rect 6737 3115 6757 3135
rect 6950 3118 6968 3136
rect 6792 3063 6812 3083
rect 7679 3100 7699 3120
rect 7332 3062 7352 3082
rect 9452 3311 9472 3331
rect 9665 3313 9685 3333
rect 10484 3368 10504 3388
rect 9868 3182 9888 3202
rect 9687 3140 9707 3160
rect 10408 3181 10428 3201
rect 10252 3126 10271 3144
rect 10463 3129 10483 3149
rect 6716 2876 6736 2896
rect 9071 2954 9091 2974
rect 9611 2953 9631 2973
rect 9444 2903 9464 2923
rect 9666 2901 9686 2921
rect 7137 2821 7161 2843
rect 6742 2573 6763 2592
rect 6441 2444 6465 2466
rect 4673 2336 4693 2356
rect 5213 2335 5233 2355
rect 3371 2256 3391 2276
rect 3911 2255 3931 2275
rect 310 1911 330 1931
rect 850 1910 870 1930
rect 683 1860 703 1880
rect 905 1858 925 1878
rect 2419 2082 2439 2102
rect 2630 2083 2651 2102
rect 2474 2030 2494 2050
rect 3295 2069 3315 2089
rect 3014 2029 3034 2049
rect 5055 2281 5075 2301
rect 5268 2283 5288 2303
rect 6087 2338 6107 2358
rect 6244 2252 6266 2270
rect 5471 2152 5491 2172
rect 5290 2110 5310 2130
rect 6011 2151 6031 2171
rect 5852 2098 5873 2117
rect 6066 2099 6086 2119
rect 10602 3062 10623 3081
rect 10204 2811 10228 2833
rect 7679 2733 7699 2753
rect 7901 2731 7921 2751
rect 7734 2681 7754 2701
rect 8274 2680 8294 2700
rect 10629 2758 10649 2778
rect 6882 2505 6902 2525
rect 7094 2510 7113 2528
rect 6937 2453 6957 2473
rect 7658 2494 7678 2514
rect 7477 2452 7497 2472
rect 6861 2266 6881 2286
rect 7680 2321 7700 2341
rect 7893 2323 7913 2343
rect 10013 2572 10033 2592
rect 9666 2534 9686 2554
rect 10553 2571 10573 2591
rect 10394 2519 10417 2541
rect 10608 2519 10628 2539
rect 15551 7212 15571 7232
rect 15762 7210 15785 7232
rect 15606 7160 15626 7180
rect 16493 7197 16513 7217
rect 16146 7159 16166 7179
rect 18155 7370 18175 7390
rect 18368 7372 18388 7392
rect 19187 7427 19207 7447
rect 18571 7241 18591 7261
rect 18390 7199 18410 7219
rect 19111 7240 19131 7260
rect 15530 6973 15550 6993
rect 18955 7185 18974 7203
rect 19166 7188 19186 7208
rect 17774 7013 17794 7033
rect 18314 7012 18334 7032
rect 15951 6918 15975 6940
rect 15556 6670 15577 6689
rect 18147 6962 18167 6982
rect 18369 6960 18389 6980
rect 16493 6830 16513 6850
rect 16715 6828 16735 6848
rect 19982 7594 20002 7614
rect 20195 7596 20216 7615
rect 20037 7542 20057 7562
rect 20758 7583 20778 7603
rect 20577 7541 20597 7561
rect 19802 7443 19824 7461
rect 19961 7355 19981 7375
rect 20780 7410 20800 7430
rect 20993 7412 21013 7432
rect 23034 7664 23054 7684
rect 22753 7624 22773 7644
rect 23574 7663 23594 7683
rect 23417 7611 23438 7630
rect 23629 7611 23649 7631
rect 28641 8227 28661 8247
rect 28852 8234 28871 8251
rect 28696 8175 28716 8195
rect 29517 8214 29537 8234
rect 29236 8174 29256 8194
rect 31277 8426 31297 8446
rect 31490 8428 31510 8448
rect 32309 8483 32329 8503
rect 31693 8297 31713 8317
rect 31512 8255 31532 8275
rect 32233 8296 32253 8316
rect 32074 8243 32095 8262
rect 32288 8244 32308 8264
rect 33901 8878 33921 8898
rect 34123 8876 34143 8896
rect 33956 8826 33976 8846
rect 34496 8825 34516 8845
rect 33104 8650 33124 8670
rect 33316 8655 33335 8673
rect 33159 8598 33179 8618
rect 33880 8639 33900 8659
rect 33699 8597 33719 8617
rect 33083 8411 33103 8431
rect 33902 8466 33922 8486
rect 34115 8468 34135 8488
rect 33957 8414 33977 8434
rect 34497 8413 34517 8433
rect 30896 8069 30916 8089
rect 28620 7988 28640 8008
rect 31436 8068 31456 8088
rect 31269 8018 31289 8038
rect 31491 8016 31511 8036
rect 27665 7913 27689 7935
rect 28978 7935 29002 7957
rect 25143 7835 25163 7855
rect 25365 7833 25385 7853
rect 25198 7783 25218 7803
rect 28027 7862 28047 7882
rect 25738 7782 25758 7802
rect 22137 7438 22157 7458
rect 22677 7437 22697 7457
rect 20835 7358 20855 7378
rect 21375 7357 21395 7377
rect 19603 7247 19627 7269
rect 19305 7121 19326 7140
rect 18907 6870 18931 6892
rect 16548 6778 16568 6798
rect 17088 6777 17108 6797
rect 15696 6602 15716 6622
rect 15908 6607 15927 6625
rect 19332 6817 19352 6837
rect 15751 6550 15771 6570
rect 16472 6591 16492 6611
rect 16291 6549 16311 6569
rect 15675 6363 15695 6383
rect 16494 6418 16514 6438
rect 16707 6420 16727 6440
rect 18716 6631 18736 6651
rect 18369 6593 18389 6613
rect 19256 6630 19276 6650
rect 19100 6577 19118 6595
rect 19311 6578 19331 6598
rect 16549 6366 16569 6386
rect 17753 6407 17773 6427
rect 17089 6365 17109 6385
rect 18293 6406 18313 6426
rect 15597 6192 15617 6212
rect 15808 6193 15829 6212
rect 15652 6140 15672 6160
rect 16473 6179 16493 6199
rect 16192 6139 16212 6159
rect 18135 6352 18155 6372
rect 18348 6354 18368 6374
rect 19167 6409 19187 6429
rect 18551 6223 18571 6243
rect 18370 6181 18390 6201
rect 19091 6222 19111 6242
rect 18932 6169 18953 6188
rect 19146 6170 19166 6190
rect 15576 5953 15596 5973
rect 17754 5995 17774 6015
rect 18294 5994 18314 6014
rect 15934 5900 15958 5922
rect 18127 5944 18147 5964
rect 18349 5942 18369 5962
rect 16476 5812 16496 5832
rect 16698 5810 16718 5830
rect 18887 5852 18911 5874
rect 16531 5760 16551 5780
rect 17071 5759 17091 5779
rect 19249 5801 19269 5821
rect 15679 5584 15699 5604
rect 15892 5586 15913 5605
rect 15734 5532 15754 5552
rect 16455 5573 16475 5593
rect 16274 5531 16294 5551
rect 15658 5345 15678 5365
rect 16477 5400 16497 5420
rect 16690 5402 16710 5422
rect 18633 5615 18653 5635
rect 18352 5575 18372 5595
rect 19173 5614 19193 5634
rect 19018 5558 19037 5575
rect 19228 5562 19248 5582
rect 16532 5348 16552 5368
rect 17736 5389 17756 5409
rect 17072 5347 17092 5367
rect 18276 5388 18296 5408
rect 15002 5111 15023 5130
rect 15375 5178 15395 5198
rect 15587 5177 15613 5203
rect 15430 5126 15450 5146
rect 16456 5161 16476 5181
rect 15970 5125 15990 5145
rect 18118 5334 18138 5354
rect 18331 5336 18351 5356
rect 19330 5491 19352 5509
rect 19150 5391 19170 5411
rect 18534 5205 18554 5225
rect 18353 5163 18373 5183
rect 19074 5204 19094 5224
rect 15354 4939 15374 4959
rect 18918 5149 18937 5167
rect 19129 5152 19149 5172
rect 17737 4977 17757 4997
rect 18277 4976 18297 4996
rect 14604 4860 14628 4882
rect 15915 4882 15939 4904
rect 18110 4926 18130 4946
rect 18332 4924 18352 4944
rect 12093 4781 12113 4801
rect 12315 4779 12335 4799
rect 12148 4729 12168 4749
rect 12688 4728 12708 4748
rect 15169 4805 15189 4825
rect 11296 4553 11316 4573
rect 11508 4558 11527 4576
rect 11351 4501 11371 4521
rect 12072 4542 12092 4562
rect 11891 4500 11911 4520
rect 11275 4314 11295 4334
rect 11093 4216 11115 4234
rect 12094 4369 12114 4389
rect 12307 4371 12327 4391
rect 14553 4619 14573 4639
rect 14067 4583 14087 4603
rect 15093 4618 15113 4638
rect 14931 4555 14954 4578
rect 15148 4566 15168 4586
rect 15520 4634 15541 4653
rect 13451 4397 13471 4417
rect 13991 4396 14011 4416
rect 12149 4317 12169 4337
rect 12689 4316 12709 4336
rect 11197 4143 11217 4163
rect 11408 4150 11427 4167
rect 11252 4091 11272 4111
rect 12073 4130 12093 4150
rect 11792 4090 11812 4110
rect 13833 4342 13853 4362
rect 14046 4344 14066 4364
rect 14865 4399 14885 4419
rect 14249 4213 14269 4233
rect 14068 4171 14088 4191
rect 14789 4212 14809 4232
rect 14630 4159 14651 4178
rect 14844 4160 14864 4180
rect 13452 3985 13472 4005
rect 11176 3904 11196 3924
rect 13992 3984 14012 4004
rect 13825 3934 13845 3954
rect 14047 3932 14067 3952
rect 11534 3851 11558 3873
rect 14585 3842 14609 3864
rect 12076 3763 12096 3783
rect 12298 3761 12318 3781
rect 12131 3711 12151 3731
rect 14947 3791 14967 3811
rect 12671 3710 12691 3730
rect 11279 3535 11299 3555
rect 11492 3537 11513 3556
rect 11334 3483 11354 3503
rect 12055 3524 12075 3544
rect 11874 3482 11894 3502
rect 11258 3296 11278 3316
rect 12077 3351 12097 3371
rect 12290 3353 12310 3373
rect 14331 3605 14351 3625
rect 14050 3565 14070 3585
rect 14871 3604 14891 3624
rect 14714 3552 14735 3571
rect 14926 3552 14946 3572
rect 13434 3379 13454 3399
rect 13974 3378 13994 3398
rect 12132 3299 12152 3319
rect 12672 3298 12692 3318
rect 11114 3127 11134 3147
rect 11327 3130 11345 3148
rect 11169 3075 11189 3095
rect 12056 3112 12076 3132
rect 11709 3074 11729 3094
rect 13816 3324 13836 3344
rect 14029 3326 14049 3346
rect 14848 3381 14868 3401
rect 14232 3195 14252 3215
rect 14051 3153 14071 3173
rect 14772 3194 14792 3214
rect 14616 3139 14635 3157
rect 14827 3142 14847 3162
rect 11093 2888 11113 2908
rect 13435 2967 13455 2987
rect 13975 2966 13995 2986
rect 13808 2916 13828 2936
rect 14030 2914 14050 2934
rect 11514 2833 11538 2855
rect 11119 2585 11140 2604
rect 10818 2456 10842 2478
rect 9050 2348 9070 2368
rect 9590 2347 9610 2367
rect 7735 2269 7755 2289
rect 8275 2268 8295 2288
rect 4674 1924 4694 1944
rect 2398 1843 2418 1863
rect 5214 1923 5234 1943
rect 5047 1873 5067 1893
rect 5269 1871 5289 1891
rect 1443 1768 1467 1790
rect 2756 1790 2780 1812
rect 1805 1717 1825 1737
rect 1189 1531 1209 1551
rect 908 1491 928 1511
rect 1729 1530 1749 1550
rect 1574 1474 1593 1491
rect 1784 1478 1804 1498
rect 6783 2095 6803 2115
rect 6994 2096 7015 2115
rect 6838 2043 6858 2063
rect 7659 2082 7679 2102
rect 7378 2042 7398 2062
rect 9432 2293 9452 2313
rect 9645 2295 9665 2315
rect 10464 2350 10484 2370
rect 10621 2264 10643 2282
rect 9848 2164 9868 2184
rect 9667 2122 9687 2142
rect 10388 2163 10408 2183
rect 10229 2110 10250 2129
rect 10443 2111 10463 2131
rect 14966 3075 14987 3094
rect 14568 2824 14592 2846
rect 12056 2745 12076 2765
rect 12278 2743 12298 2763
rect 12111 2693 12131 2713
rect 12651 2692 12671 2712
rect 14993 2771 15013 2791
rect 11259 2517 11279 2537
rect 11471 2522 11490 2540
rect 11314 2465 11334 2485
rect 12035 2506 12055 2526
rect 11854 2464 11874 2484
rect 11238 2278 11258 2298
rect 12057 2333 12077 2353
rect 12270 2335 12290 2355
rect 14377 2585 14397 2605
rect 14030 2547 14050 2567
rect 14917 2584 14937 2604
rect 14758 2532 14781 2554
rect 14972 2532 14992 2552
rect 19817 7186 19837 7206
rect 20028 7184 20051 7206
rect 19872 7134 19892 7154
rect 20759 7171 20779 7191
rect 20412 7133 20432 7153
rect 22519 7383 22539 7403
rect 22732 7385 22752 7405
rect 23551 7440 23571 7460
rect 22935 7254 22955 7274
rect 22754 7212 22774 7232
rect 23475 7253 23495 7273
rect 23319 7198 23338 7216
rect 23530 7201 23550 7221
rect 19796 6947 19816 6967
rect 22138 7026 22158 7046
rect 22678 7025 22698 7045
rect 22511 6975 22531 6995
rect 22733 6973 22753 6993
rect 20217 6892 20241 6914
rect 19822 6644 19843 6663
rect 24346 7607 24366 7627
rect 24559 7609 24580 7628
rect 24401 7555 24421 7575
rect 25122 7596 25142 7616
rect 24941 7554 24961 7574
rect 24166 7456 24188 7474
rect 24325 7368 24345 7388
rect 25144 7423 25164 7443
rect 25357 7425 25377 7445
rect 27411 7676 27431 7696
rect 27130 7636 27150 7656
rect 27951 7675 27971 7695
rect 27794 7623 27815 7642
rect 28006 7623 28026 7643
rect 33005 8240 33025 8260
rect 33216 8247 33235 8264
rect 33060 8188 33080 8208
rect 33881 8227 33901 8247
rect 33600 8187 33620 8207
rect 32984 8001 33004 8021
rect 32029 7926 32053 7948
rect 33342 7948 33366 7970
rect 29520 7847 29540 7867
rect 29742 7845 29762 7865
rect 29575 7795 29595 7815
rect 32391 7875 32411 7895
rect 30115 7794 30135 7814
rect 26514 7450 26534 7470
rect 27054 7449 27074 7469
rect 25199 7371 25219 7391
rect 25739 7370 25759 7390
rect 23967 7260 23991 7282
rect 23669 7134 23690 7153
rect 23271 6883 23295 6905
rect 20759 6804 20779 6824
rect 20981 6802 21001 6822
rect 20814 6752 20834 6772
rect 21354 6751 21374 6771
rect 23696 6830 23716 6850
rect 19962 6576 19982 6596
rect 20174 6581 20193 6599
rect 20017 6524 20037 6544
rect 20738 6565 20758 6585
rect 20557 6523 20577 6543
rect 19941 6337 19961 6357
rect 20760 6392 20780 6412
rect 20973 6394 20993 6414
rect 23080 6644 23100 6664
rect 22733 6606 22753 6626
rect 23620 6643 23640 6663
rect 23464 6590 23482 6608
rect 23675 6591 23695 6611
rect 22117 6420 22137 6440
rect 22657 6419 22677 6439
rect 20815 6340 20835 6360
rect 21355 6339 21375 6359
rect 19863 6166 19883 6186
rect 20074 6167 20095 6186
rect 19918 6114 19938 6134
rect 20739 6153 20759 6173
rect 20458 6113 20478 6133
rect 22499 6365 22519 6385
rect 22712 6367 22732 6387
rect 23531 6422 23551 6442
rect 22915 6236 22935 6256
rect 22734 6194 22754 6214
rect 23455 6235 23475 6255
rect 23296 6182 23317 6201
rect 23510 6183 23530 6203
rect 22118 6008 22138 6028
rect 19842 5927 19862 5947
rect 22658 6007 22678 6027
rect 22491 5957 22511 5977
rect 22713 5955 22733 5975
rect 20200 5874 20224 5896
rect 23251 5865 23275 5887
rect 20742 5786 20762 5806
rect 20964 5784 20984 5804
rect 20797 5734 20817 5754
rect 23613 5814 23633 5834
rect 21337 5733 21357 5753
rect 19945 5558 19965 5578
rect 20158 5560 20179 5579
rect 20000 5506 20020 5526
rect 20721 5547 20741 5567
rect 20540 5505 20560 5525
rect 19924 5319 19944 5339
rect 20743 5374 20763 5394
rect 20956 5376 20976 5396
rect 22997 5628 23017 5648
rect 22716 5588 22736 5608
rect 23537 5627 23557 5647
rect 23382 5571 23401 5588
rect 23592 5575 23612 5595
rect 22100 5402 22120 5422
rect 22640 5401 22660 5421
rect 20798 5322 20818 5342
rect 21338 5321 21358 5341
rect 19268 5085 19289 5104
rect 19641 5152 19661 5172
rect 19853 5151 19879 5177
rect 19696 5100 19716 5120
rect 20722 5135 20742 5155
rect 20236 5099 20256 5119
rect 22482 5347 22502 5367
rect 22695 5349 22715 5369
rect 23694 5504 23716 5522
rect 23514 5404 23534 5424
rect 22898 5218 22918 5238
rect 22717 5176 22737 5196
rect 23438 5217 23458 5237
rect 23282 5162 23301 5180
rect 23493 5165 23513 5185
rect 19620 4913 19640 4933
rect 22101 4990 22121 5010
rect 22641 4989 22661 5009
rect 22474 4939 22494 4959
rect 22696 4937 22716 4957
rect 16457 4794 16477 4814
rect 16679 4792 16699 4812
rect 18870 4834 18894 4856
rect 20181 4856 20205 4878
rect 16512 4742 16532 4762
rect 17052 4741 17072 4761
rect 15660 4566 15680 4586
rect 15872 4571 15891 4589
rect 19435 4779 19455 4799
rect 15715 4514 15735 4534
rect 16436 4555 16456 4575
rect 16255 4513 16275 4533
rect 15639 4327 15659 4347
rect 15457 4229 15479 4247
rect 16458 4382 16478 4402
rect 16671 4384 16691 4404
rect 18819 4593 18839 4613
rect 18333 4557 18353 4577
rect 19359 4592 19379 4612
rect 19197 4529 19220 4552
rect 19414 4540 19434 4560
rect 19786 4608 19807 4627
rect 16513 4330 16533 4350
rect 17717 4371 17737 4391
rect 17053 4329 17073 4349
rect 18257 4370 18277 4390
rect 15561 4156 15581 4176
rect 15772 4163 15791 4180
rect 15616 4104 15636 4124
rect 16437 4143 16457 4163
rect 16156 4103 16176 4123
rect 18099 4316 18119 4336
rect 18312 4318 18332 4338
rect 19131 4373 19151 4393
rect 18515 4187 18535 4207
rect 18334 4145 18354 4165
rect 19055 4186 19075 4206
rect 18896 4133 18917 4152
rect 19110 4134 19130 4154
rect 15540 3917 15560 3937
rect 17718 3959 17738 3979
rect 18258 3958 18278 3978
rect 15898 3864 15922 3886
rect 18091 3908 18111 3928
rect 18313 3906 18333 3926
rect 16440 3776 16460 3796
rect 16662 3774 16682 3794
rect 18851 3816 18875 3838
rect 16495 3724 16515 3744
rect 17035 3723 17055 3743
rect 19213 3765 19233 3785
rect 15643 3548 15663 3568
rect 15856 3550 15877 3569
rect 15698 3496 15718 3516
rect 16419 3537 16439 3557
rect 16238 3495 16258 3515
rect 15622 3309 15642 3329
rect 16441 3364 16461 3384
rect 16654 3366 16674 3386
rect 18597 3579 18617 3599
rect 18316 3539 18336 3559
rect 19137 3578 19157 3598
rect 18980 3526 19001 3545
rect 19192 3526 19212 3546
rect 16496 3312 16516 3332
rect 17700 3353 17720 3373
rect 17036 3311 17056 3331
rect 18240 3352 18260 3372
rect 15478 3140 15498 3160
rect 15691 3143 15709 3161
rect 15533 3088 15553 3108
rect 16420 3125 16440 3145
rect 16073 3087 16093 3107
rect 18082 3298 18102 3318
rect 18295 3300 18315 3320
rect 19114 3355 19134 3375
rect 18498 3169 18518 3189
rect 18317 3127 18337 3147
rect 19038 3168 19058 3188
rect 15457 2901 15477 2921
rect 18882 3113 18901 3131
rect 19093 3116 19113 3136
rect 17701 2941 17721 2961
rect 18241 2940 18261 2960
rect 15878 2846 15902 2868
rect 15483 2598 15504 2617
rect 15182 2469 15206 2491
rect 13414 2361 13434 2381
rect 13954 2360 13974 2380
rect 12112 2281 12132 2301
rect 12652 2280 12672 2300
rect 9051 1936 9071 1956
rect 6762 1856 6782 1876
rect 9591 1935 9611 1955
rect 9424 1885 9444 1905
rect 9646 1883 9666 1903
rect 5807 1781 5831 1803
rect 7120 1803 7144 1825
rect 3298 1702 3318 1722
rect 3520 1700 3540 1720
rect 3353 1650 3373 1670
rect 6169 1730 6189 1750
rect 3893 1649 3913 1669
rect 292 1305 312 1325
rect 832 1304 852 1324
rect 674 1250 694 1270
rect 887 1252 907 1272
rect 1706 1307 1726 1327
rect 1090 1121 1110 1141
rect 909 1079 929 1099
rect 1630 1120 1650 1140
rect 1474 1065 1493 1083
rect 1685 1068 1705 1088
rect 293 893 313 913
rect 833 892 853 912
rect 666 842 686 862
rect 888 840 908 860
rect 2501 1474 2521 1494
rect 2714 1476 2735 1495
rect 2556 1422 2576 1442
rect 3277 1463 3297 1483
rect 3096 1421 3116 1441
rect 2480 1235 2500 1255
rect 3299 1290 3319 1310
rect 3512 1292 3532 1312
rect 5553 1544 5573 1564
rect 5272 1504 5292 1524
rect 6093 1543 6113 1563
rect 5938 1487 5957 1504
rect 6148 1491 6168 1511
rect 11160 2107 11180 2127
rect 11371 2108 11392 2127
rect 11215 2055 11235 2075
rect 12036 2094 12056 2114
rect 11755 2054 11775 2074
rect 13796 2306 13816 2326
rect 14009 2308 14029 2328
rect 14828 2363 14848 2383
rect 14985 2277 15007 2295
rect 14212 2177 14232 2197
rect 14031 2135 14051 2155
rect 14752 2176 14772 2196
rect 14593 2123 14614 2142
rect 14807 2124 14827 2144
rect 18074 2890 18094 2910
rect 18296 2888 18316 2908
rect 16420 2758 16440 2778
rect 16642 2756 16662 2776
rect 19232 3049 19253 3068
rect 18834 2798 18858 2820
rect 16475 2706 16495 2726
rect 17015 2705 17035 2725
rect 15623 2530 15643 2550
rect 15835 2535 15854 2553
rect 19259 2745 19279 2765
rect 15678 2478 15698 2498
rect 16399 2519 16419 2539
rect 16218 2477 16238 2497
rect 15602 2291 15622 2311
rect 16421 2346 16441 2366
rect 16634 2348 16654 2368
rect 18643 2559 18663 2579
rect 18296 2521 18316 2541
rect 19183 2558 19203 2578
rect 19024 2506 19047 2528
rect 19238 2506 19258 2526
rect 24181 7199 24201 7219
rect 24392 7197 24415 7219
rect 24236 7147 24256 7167
rect 25123 7184 25143 7204
rect 24776 7146 24796 7166
rect 26896 7395 26916 7415
rect 27109 7397 27129 7417
rect 27928 7452 27948 7472
rect 27312 7266 27332 7286
rect 27131 7224 27151 7244
rect 27852 7265 27872 7285
rect 27696 7210 27715 7228
rect 27907 7213 27927 7233
rect 24160 6960 24180 6980
rect 26515 7038 26535 7058
rect 27055 7037 27075 7057
rect 26888 6987 26908 7007
rect 27110 6985 27130 7005
rect 24581 6905 24605 6927
rect 24186 6657 24207 6676
rect 28723 7619 28743 7639
rect 28936 7621 28957 7640
rect 28778 7567 28798 7587
rect 29499 7608 29519 7628
rect 29318 7566 29338 7586
rect 28543 7468 28565 7486
rect 28702 7380 28722 7400
rect 29521 7435 29541 7455
rect 29734 7437 29754 7457
rect 31775 7689 31795 7709
rect 31494 7649 31514 7669
rect 32315 7688 32335 7708
rect 32158 7636 32179 7655
rect 32370 7636 32390 7656
rect 33884 7860 33904 7880
rect 34106 7858 34126 7878
rect 33939 7808 33959 7828
rect 34479 7807 34499 7827
rect 30878 7463 30898 7483
rect 31418 7462 31438 7482
rect 29576 7383 29596 7403
rect 30116 7382 30136 7402
rect 28344 7272 28368 7294
rect 28046 7146 28067 7165
rect 27648 6895 27672 6917
rect 25123 6817 25143 6837
rect 25345 6815 25365 6835
rect 25178 6765 25198 6785
rect 25718 6764 25738 6784
rect 28073 6842 28093 6862
rect 24326 6589 24346 6609
rect 24538 6594 24557 6612
rect 24381 6537 24401 6557
rect 25102 6578 25122 6598
rect 24921 6536 24941 6556
rect 24305 6350 24325 6370
rect 25124 6405 25144 6425
rect 25337 6407 25357 6427
rect 27457 6656 27477 6676
rect 27110 6618 27130 6638
rect 27997 6655 28017 6675
rect 27841 6602 27859 6620
rect 28052 6603 28072 6623
rect 26494 6432 26514 6452
rect 27034 6431 27054 6451
rect 25179 6353 25199 6373
rect 25719 6352 25739 6372
rect 24227 6179 24247 6199
rect 24438 6180 24459 6199
rect 24282 6127 24302 6147
rect 25103 6166 25123 6186
rect 24822 6126 24842 6146
rect 26876 6377 26896 6397
rect 27089 6379 27109 6399
rect 27908 6434 27928 6454
rect 27292 6248 27312 6268
rect 27111 6206 27131 6226
rect 27832 6247 27852 6267
rect 27673 6194 27694 6213
rect 27887 6195 27907 6215
rect 26495 6020 26515 6040
rect 24206 5940 24226 5960
rect 27035 6019 27055 6039
rect 26868 5969 26888 5989
rect 27090 5967 27110 5987
rect 24564 5887 24588 5909
rect 27628 5877 27652 5899
rect 25106 5799 25126 5819
rect 25328 5797 25348 5817
rect 25161 5747 25181 5767
rect 27990 5826 28010 5846
rect 25701 5746 25721 5766
rect 24309 5571 24329 5591
rect 24522 5573 24543 5592
rect 24364 5519 24384 5539
rect 25085 5560 25105 5580
rect 24904 5518 24924 5538
rect 24288 5332 24308 5352
rect 25107 5387 25127 5407
rect 25320 5389 25340 5409
rect 27374 5640 27394 5660
rect 27093 5600 27113 5620
rect 27914 5639 27934 5659
rect 27759 5583 27778 5600
rect 27969 5587 27989 5607
rect 26477 5414 26497 5434
rect 27017 5413 27037 5433
rect 25162 5335 25182 5355
rect 25702 5334 25722 5354
rect 23632 5098 23653 5117
rect 24005 5165 24025 5185
rect 24217 5164 24243 5190
rect 24060 5113 24080 5133
rect 25086 5148 25106 5168
rect 24600 5112 24620 5132
rect 26859 5359 26879 5379
rect 27072 5361 27092 5381
rect 28071 5516 28093 5534
rect 27891 5416 27911 5436
rect 27275 5230 27295 5250
rect 27094 5188 27114 5208
rect 27815 5229 27835 5249
rect 27659 5174 27678 5192
rect 27870 5177 27890 5197
rect 23984 4926 24004 4946
rect 26478 5002 26498 5022
rect 27018 5001 27038 5021
rect 26851 4951 26871 4971
rect 27073 4949 27093 4969
rect 23234 4847 23258 4869
rect 24545 4869 24569 4891
rect 20723 4768 20743 4788
rect 20945 4766 20965 4786
rect 20778 4716 20798 4736
rect 21318 4715 21338 4735
rect 23799 4792 23819 4812
rect 19926 4540 19946 4560
rect 20138 4545 20157 4563
rect 19981 4488 20001 4508
rect 20702 4529 20722 4549
rect 20521 4487 20541 4507
rect 19905 4301 19925 4321
rect 19723 4203 19745 4221
rect 20724 4356 20744 4376
rect 20937 4358 20957 4378
rect 23183 4606 23203 4626
rect 22697 4570 22717 4590
rect 23723 4605 23743 4625
rect 23561 4542 23584 4565
rect 23778 4553 23798 4573
rect 24150 4621 24171 4640
rect 22081 4384 22101 4404
rect 22621 4383 22641 4403
rect 20779 4304 20799 4324
rect 21319 4303 21339 4323
rect 19827 4130 19847 4150
rect 20038 4137 20057 4154
rect 19882 4078 19902 4098
rect 20703 4117 20723 4137
rect 20422 4077 20442 4097
rect 22463 4329 22483 4349
rect 22676 4331 22696 4351
rect 23495 4386 23515 4406
rect 22879 4200 22899 4220
rect 22698 4158 22718 4178
rect 23419 4199 23439 4219
rect 23260 4146 23281 4165
rect 23474 4147 23494 4167
rect 22082 3972 22102 3992
rect 19806 3891 19826 3911
rect 22622 3971 22642 3991
rect 22455 3921 22475 3941
rect 22677 3919 22697 3939
rect 20164 3838 20188 3860
rect 23215 3829 23239 3851
rect 20706 3750 20726 3770
rect 20928 3748 20948 3768
rect 20761 3698 20781 3718
rect 23577 3778 23597 3798
rect 21301 3697 21321 3717
rect 19909 3522 19929 3542
rect 20122 3524 20143 3543
rect 19964 3470 19984 3490
rect 20685 3511 20705 3531
rect 20504 3469 20524 3489
rect 19888 3283 19908 3303
rect 20707 3338 20727 3358
rect 20920 3340 20940 3360
rect 22961 3592 22981 3612
rect 22680 3552 22700 3572
rect 23501 3591 23521 3611
rect 23344 3539 23365 3558
rect 23556 3539 23576 3559
rect 22064 3366 22084 3386
rect 22604 3365 22624 3385
rect 20762 3286 20782 3306
rect 21302 3285 21322 3305
rect 19744 3114 19764 3134
rect 19957 3117 19975 3135
rect 19799 3062 19819 3082
rect 20686 3099 20706 3119
rect 20339 3061 20359 3081
rect 22446 3311 22466 3331
rect 22659 3313 22679 3333
rect 23478 3368 23498 3388
rect 22862 3182 22882 3202
rect 22681 3140 22701 3160
rect 23402 3181 23422 3201
rect 23246 3126 23265 3144
rect 23457 3129 23477 3149
rect 19723 2875 19743 2895
rect 22065 2954 22085 2974
rect 22605 2953 22625 2973
rect 22438 2903 22458 2923
rect 22660 2901 22680 2921
rect 20144 2820 20168 2842
rect 19749 2572 19770 2591
rect 19448 2443 19472 2465
rect 16476 2294 16496 2314
rect 17680 2335 17700 2355
rect 17016 2293 17036 2313
rect 18220 2334 18240 2354
rect 13415 1949 13435 1969
rect 11139 1868 11159 1888
rect 13955 1948 13975 1968
rect 13788 1898 13808 1918
rect 14010 1896 14030 1916
rect 10184 1793 10208 1815
rect 11497 1815 11521 1837
rect 7662 1715 7682 1735
rect 7884 1713 7904 1733
rect 7717 1663 7737 1683
rect 10546 1742 10566 1762
rect 8257 1662 8277 1682
rect 4656 1318 4676 1338
rect 5196 1317 5216 1337
rect 3354 1238 3374 1258
rect 3894 1237 3914 1257
rect 3278 1051 3298 1071
rect 1824 1001 1845 1020
rect 5038 1263 5058 1283
rect 5251 1265 5271 1285
rect 6070 1320 6090 1340
rect 5454 1134 5474 1154
rect 5273 1092 5293 1112
rect 5994 1133 6014 1153
rect 5838 1078 5857 1096
rect 6049 1081 6069 1101
rect 4657 906 4677 926
rect 5197 905 5217 925
rect 5030 855 5050 875
rect 5252 853 5272 873
rect 4047 788 4079 813
rect 1426 750 1450 772
rect 6865 1487 6885 1507
rect 7078 1489 7099 1508
rect 6920 1435 6940 1455
rect 7641 1476 7661 1496
rect 7460 1434 7480 1454
rect 6844 1248 6864 1268
rect 7663 1303 7683 1323
rect 7876 1305 7896 1325
rect 9930 1556 9950 1576
rect 9649 1516 9669 1536
rect 10470 1555 10490 1575
rect 10315 1499 10334 1516
rect 10525 1503 10545 1523
rect 15524 2120 15544 2140
rect 15735 2121 15756 2140
rect 15579 2068 15599 2088
rect 16400 2107 16420 2127
rect 16119 2067 16139 2087
rect 18062 2280 18082 2300
rect 18275 2282 18295 2302
rect 19094 2337 19114 2357
rect 19251 2251 19273 2269
rect 18478 2151 18498 2171
rect 18297 2109 18317 2129
rect 19018 2150 19038 2170
rect 18859 2097 18880 2116
rect 19073 2098 19093 2118
rect 23596 3062 23617 3081
rect 23198 2811 23222 2833
rect 20686 2732 20706 2752
rect 20908 2730 20928 2750
rect 20741 2680 20761 2700
rect 21281 2679 21301 2699
rect 23623 2758 23643 2778
rect 19889 2504 19909 2524
rect 20101 2509 20120 2527
rect 19944 2452 19964 2472
rect 20665 2493 20685 2513
rect 20484 2451 20504 2471
rect 19868 2265 19888 2285
rect 20687 2320 20707 2340
rect 20900 2322 20920 2342
rect 23007 2572 23027 2592
rect 22660 2534 22680 2554
rect 23547 2571 23567 2591
rect 23388 2519 23411 2541
rect 23602 2519 23622 2539
rect 28558 7211 28578 7231
rect 28769 7209 28792 7231
rect 28613 7159 28633 7179
rect 29500 7196 29520 7216
rect 29153 7158 29173 7178
rect 31260 7408 31280 7428
rect 31473 7410 31493 7430
rect 32292 7465 32312 7485
rect 31676 7279 31696 7299
rect 31495 7237 31515 7257
rect 32216 7278 32236 7298
rect 32060 7223 32079 7241
rect 32271 7226 32291 7246
rect 28537 6972 28557 6992
rect 30879 7051 30899 7071
rect 31419 7050 31439 7070
rect 31252 7000 31272 7020
rect 31474 6998 31494 7018
rect 28958 6917 28982 6939
rect 28563 6669 28584 6688
rect 33087 7632 33107 7652
rect 33300 7634 33321 7653
rect 33142 7580 33162 7600
rect 33863 7621 33883 7641
rect 33682 7579 33702 7599
rect 32907 7481 32929 7499
rect 33066 7393 33086 7413
rect 33885 7448 33905 7468
rect 34098 7450 34118 7470
rect 33940 7396 33960 7416
rect 34480 7395 34500 7415
rect 32708 7285 32732 7307
rect 32410 7159 32431 7178
rect 32012 6908 32036 6930
rect 29500 6829 29520 6849
rect 29722 6827 29742 6847
rect 29555 6777 29575 6797
rect 30095 6776 30115 6796
rect 32437 6855 32457 6875
rect 28703 6601 28723 6621
rect 28915 6606 28934 6624
rect 28758 6549 28778 6569
rect 29479 6590 29499 6610
rect 29298 6548 29318 6568
rect 28682 6362 28702 6382
rect 29501 6417 29521 6437
rect 29714 6419 29734 6439
rect 31821 6669 31841 6689
rect 31474 6631 31494 6651
rect 32361 6668 32381 6688
rect 32205 6615 32223 6633
rect 32416 6616 32436 6636
rect 30858 6445 30878 6465
rect 31398 6444 31418 6464
rect 29556 6365 29576 6385
rect 30096 6364 30116 6384
rect 28604 6191 28624 6211
rect 28815 6192 28836 6211
rect 28659 6139 28679 6159
rect 29480 6178 29500 6198
rect 29199 6138 29219 6158
rect 31240 6390 31260 6410
rect 31453 6392 31473 6412
rect 32272 6447 32292 6467
rect 31656 6261 31676 6281
rect 31475 6219 31495 6239
rect 32196 6260 32216 6280
rect 32037 6207 32058 6226
rect 32251 6208 32271 6228
rect 30859 6033 30879 6053
rect 28583 5952 28603 5972
rect 31399 6032 31419 6052
rect 31232 5982 31252 6002
rect 31454 5980 31474 6000
rect 28941 5899 28965 5921
rect 31992 5890 32016 5912
rect 29483 5811 29503 5831
rect 29705 5809 29725 5829
rect 29538 5759 29558 5779
rect 32354 5839 32374 5859
rect 30078 5758 30098 5778
rect 28686 5583 28706 5603
rect 28899 5585 28920 5604
rect 28741 5531 28761 5551
rect 29462 5572 29482 5592
rect 29281 5530 29301 5550
rect 28665 5344 28685 5364
rect 29484 5399 29504 5419
rect 29697 5401 29717 5421
rect 31738 5653 31758 5673
rect 31457 5613 31477 5633
rect 32278 5652 32298 5672
rect 32123 5596 32142 5613
rect 32333 5600 32353 5620
rect 30841 5427 30861 5447
rect 31381 5426 31401 5446
rect 29539 5347 29559 5367
rect 30079 5346 30099 5366
rect 28009 5110 28030 5129
rect 28382 5177 28402 5197
rect 28594 5176 28620 5202
rect 28437 5125 28457 5145
rect 29463 5160 29483 5180
rect 28977 5124 28997 5144
rect 31223 5372 31243 5392
rect 31436 5374 31456 5394
rect 32435 5529 32457 5547
rect 32255 5429 32275 5449
rect 31639 5243 31659 5263
rect 31458 5201 31478 5221
rect 32179 5242 32199 5262
rect 32023 5187 32042 5205
rect 32234 5190 32254 5210
rect 28361 4938 28381 4958
rect 30842 5015 30862 5035
rect 31382 5014 31402 5034
rect 31215 4964 31235 4984
rect 31437 4962 31457 4982
rect 27611 4859 27635 4881
rect 28922 4881 28946 4903
rect 25087 4781 25107 4801
rect 25309 4779 25329 4799
rect 25142 4729 25162 4749
rect 25682 4728 25702 4748
rect 28176 4804 28196 4824
rect 24290 4553 24310 4573
rect 24502 4558 24521 4576
rect 24345 4501 24365 4521
rect 25066 4542 25086 4562
rect 24885 4500 24905 4520
rect 24269 4314 24289 4334
rect 24087 4216 24109 4234
rect 25088 4369 25108 4389
rect 25301 4371 25321 4391
rect 27560 4618 27580 4638
rect 27074 4582 27094 4602
rect 28100 4617 28120 4637
rect 27938 4554 27961 4577
rect 28155 4565 28175 4585
rect 28527 4633 28548 4652
rect 26458 4396 26478 4416
rect 26998 4395 27018 4415
rect 25143 4317 25163 4337
rect 25683 4316 25703 4336
rect 24191 4143 24211 4163
rect 24402 4150 24421 4167
rect 24246 4091 24266 4111
rect 25067 4130 25087 4150
rect 24786 4090 24806 4110
rect 26840 4341 26860 4361
rect 27053 4343 27073 4363
rect 27872 4398 27892 4418
rect 27256 4212 27276 4232
rect 27075 4170 27095 4190
rect 27796 4211 27816 4231
rect 27637 4158 27658 4177
rect 27851 4159 27871 4179
rect 26459 3984 26479 4004
rect 24170 3904 24190 3924
rect 26999 3983 27019 4003
rect 26832 3933 26852 3953
rect 27054 3931 27074 3951
rect 24528 3851 24552 3873
rect 27592 3841 27616 3863
rect 25070 3763 25090 3783
rect 25292 3761 25312 3781
rect 25125 3711 25145 3731
rect 27954 3790 27974 3810
rect 25665 3710 25685 3730
rect 24273 3535 24293 3555
rect 24486 3537 24507 3556
rect 24328 3483 24348 3503
rect 25049 3524 25069 3544
rect 24868 3482 24888 3502
rect 24252 3296 24272 3316
rect 25071 3351 25091 3371
rect 25284 3353 25304 3373
rect 27338 3604 27358 3624
rect 27057 3564 27077 3584
rect 27878 3603 27898 3623
rect 27721 3551 27742 3570
rect 27933 3551 27953 3571
rect 26441 3378 26461 3398
rect 26981 3377 27001 3397
rect 25126 3299 25146 3319
rect 25666 3298 25686 3318
rect 24108 3127 24128 3147
rect 24321 3130 24339 3148
rect 24163 3075 24183 3095
rect 25050 3112 25070 3132
rect 24703 3074 24723 3094
rect 26823 3323 26843 3343
rect 27036 3325 27056 3345
rect 27855 3380 27875 3400
rect 27239 3194 27259 3214
rect 27058 3152 27078 3172
rect 27779 3193 27799 3213
rect 27623 3138 27642 3156
rect 27834 3141 27854 3161
rect 24087 2888 24107 2908
rect 26442 2966 26462 2986
rect 26982 2965 27002 2985
rect 26815 2915 26835 2935
rect 27037 2913 27057 2933
rect 24508 2833 24532 2855
rect 24113 2585 24134 2604
rect 23812 2456 23836 2478
rect 22044 2348 22064 2368
rect 22584 2347 22604 2367
rect 20742 2268 20762 2288
rect 21282 2267 21302 2287
rect 15503 1881 15523 1901
rect 17681 1923 17701 1943
rect 18221 1922 18241 1942
rect 14548 1806 14572 1828
rect 15861 1828 15885 1850
rect 12039 1727 12059 1747
rect 12261 1725 12281 1745
rect 12094 1675 12114 1695
rect 14910 1755 14930 1775
rect 12634 1674 12654 1694
rect 9033 1330 9053 1350
rect 9573 1329 9593 1349
rect 7718 1251 7738 1271
rect 8258 1250 8278 1270
rect 7642 1064 7662 1084
rect 6188 1014 6209 1033
rect 9415 1275 9435 1295
rect 9628 1277 9648 1297
rect 10447 1332 10467 1352
rect 9831 1146 9851 1166
rect 9650 1104 9670 1124
rect 10371 1145 10391 1165
rect 10215 1090 10234 1108
rect 10426 1093 10446 1113
rect 9034 918 9054 938
rect 9574 917 9594 937
rect 9407 867 9427 887
rect 9629 865 9649 885
rect 8411 801 8443 826
rect 5790 763 5814 785
rect 11242 1499 11262 1519
rect 11455 1501 11476 1520
rect 11297 1447 11317 1467
rect 12018 1488 12038 1508
rect 11837 1446 11857 1466
rect 11221 1260 11241 1280
rect 12040 1315 12060 1335
rect 12253 1317 12273 1337
rect 14294 1569 14314 1589
rect 14013 1529 14033 1549
rect 14834 1568 14854 1588
rect 14679 1512 14698 1529
rect 14889 1516 14909 1536
rect 18054 1872 18074 1892
rect 18276 1870 18296 1890
rect 16403 1740 16423 1760
rect 16625 1738 16645 1758
rect 19790 2094 19810 2114
rect 20001 2095 20022 2114
rect 19845 2042 19865 2062
rect 20666 2081 20686 2101
rect 20385 2041 20405 2061
rect 22426 2293 22446 2313
rect 22639 2295 22659 2315
rect 23458 2350 23478 2370
rect 23615 2264 23637 2282
rect 22842 2164 22862 2184
rect 22661 2122 22681 2142
rect 23382 2163 23402 2183
rect 23223 2110 23244 2129
rect 23437 2111 23457 2131
rect 27973 3074 27994 3093
rect 27575 2823 27599 2845
rect 25050 2745 25070 2765
rect 25272 2743 25292 2763
rect 25105 2693 25125 2713
rect 25645 2692 25665 2712
rect 28000 2770 28020 2790
rect 24253 2517 24273 2537
rect 24465 2522 24484 2540
rect 24308 2465 24328 2485
rect 25029 2506 25049 2526
rect 24848 2464 24868 2484
rect 24232 2278 24252 2298
rect 25051 2333 25071 2353
rect 25264 2335 25284 2355
rect 27384 2584 27404 2604
rect 27037 2546 27057 2566
rect 27924 2583 27944 2603
rect 27765 2531 27788 2553
rect 27979 2531 27999 2551
rect 32922 7224 32942 7244
rect 33133 7222 33156 7244
rect 32977 7172 32997 7192
rect 33864 7209 33884 7229
rect 33517 7171 33537 7191
rect 32901 6985 32921 7005
rect 33322 6930 33346 6952
rect 32927 6682 32948 6701
rect 33864 6842 33884 6862
rect 34086 6840 34106 6860
rect 33919 6790 33939 6810
rect 34459 6789 34479 6809
rect 33067 6614 33087 6634
rect 33279 6619 33298 6637
rect 33122 6562 33142 6582
rect 33843 6603 33863 6623
rect 33662 6561 33682 6581
rect 33046 6375 33066 6395
rect 33865 6430 33885 6450
rect 34078 6432 34098 6452
rect 33920 6378 33940 6398
rect 34460 6377 34480 6397
rect 32968 6204 32988 6224
rect 33179 6205 33200 6224
rect 33023 6152 33043 6172
rect 33844 6191 33864 6211
rect 33563 6151 33583 6171
rect 32947 5965 32967 5985
rect 33305 5912 33329 5934
rect 33847 5824 33867 5844
rect 34069 5822 34089 5842
rect 33902 5772 33922 5792
rect 34442 5771 34462 5791
rect 33050 5596 33070 5616
rect 33263 5598 33284 5617
rect 33105 5544 33125 5564
rect 33826 5585 33846 5605
rect 33645 5543 33665 5563
rect 33029 5357 33049 5377
rect 33848 5412 33868 5432
rect 34061 5414 34081 5434
rect 33903 5360 33923 5380
rect 34443 5359 34463 5379
rect 32373 5123 32394 5142
rect 32746 5190 32766 5210
rect 32958 5189 32984 5215
rect 32801 5138 32821 5158
rect 33827 5173 33847 5193
rect 33341 5137 33361 5157
rect 32725 4951 32745 4971
rect 31975 4872 31999 4894
rect 33286 4894 33310 4916
rect 29464 4793 29484 4813
rect 29686 4791 29706 4811
rect 29519 4741 29539 4761
rect 30059 4740 30079 4760
rect 32540 4817 32560 4837
rect 28667 4565 28687 4585
rect 28879 4570 28898 4588
rect 28722 4513 28742 4533
rect 29443 4554 29463 4574
rect 29262 4512 29282 4532
rect 28646 4326 28666 4346
rect 28464 4228 28486 4246
rect 29465 4381 29485 4401
rect 29678 4383 29698 4403
rect 31924 4631 31944 4651
rect 31438 4595 31458 4615
rect 32464 4630 32484 4650
rect 32302 4567 32325 4590
rect 32519 4578 32539 4598
rect 32891 4646 32912 4665
rect 30822 4409 30842 4429
rect 31362 4408 31382 4428
rect 29520 4329 29540 4349
rect 30060 4328 30080 4348
rect 28568 4155 28588 4175
rect 28779 4162 28798 4179
rect 28623 4103 28643 4123
rect 29444 4142 29464 4162
rect 29163 4102 29183 4122
rect 31204 4354 31224 4374
rect 31417 4356 31437 4376
rect 32236 4411 32256 4431
rect 31620 4225 31640 4245
rect 31439 4183 31459 4203
rect 32160 4224 32180 4244
rect 32001 4171 32022 4190
rect 32215 4172 32235 4192
rect 30823 3997 30843 4017
rect 28547 3916 28567 3936
rect 31363 3996 31383 4016
rect 31196 3946 31216 3966
rect 31418 3944 31438 3964
rect 28905 3863 28929 3885
rect 31956 3854 31980 3876
rect 29447 3775 29467 3795
rect 29669 3773 29689 3793
rect 29502 3723 29522 3743
rect 32318 3803 32338 3823
rect 30042 3722 30062 3742
rect 28650 3547 28670 3567
rect 28863 3549 28884 3568
rect 28705 3495 28725 3515
rect 29426 3536 29446 3556
rect 29245 3494 29265 3514
rect 28629 3308 28649 3328
rect 29448 3363 29468 3383
rect 29661 3365 29681 3385
rect 31702 3617 31722 3637
rect 31421 3577 31441 3597
rect 32242 3616 32262 3636
rect 32085 3564 32106 3583
rect 32297 3564 32317 3584
rect 30805 3391 30825 3411
rect 31345 3390 31365 3410
rect 29503 3311 29523 3331
rect 30043 3310 30063 3330
rect 28485 3139 28505 3159
rect 28698 3142 28716 3160
rect 28540 3087 28560 3107
rect 29427 3124 29447 3144
rect 29080 3086 29100 3106
rect 31187 3336 31207 3356
rect 31400 3338 31420 3358
rect 32219 3393 32239 3413
rect 31603 3207 31623 3227
rect 31422 3165 31442 3185
rect 32143 3206 32163 3226
rect 31987 3151 32006 3169
rect 32198 3154 32218 3174
rect 28464 2900 28484 2920
rect 30806 2979 30826 2999
rect 31346 2978 31366 2998
rect 31179 2928 31199 2948
rect 31401 2926 31421 2946
rect 28885 2845 28909 2867
rect 28490 2597 28511 2616
rect 28189 2468 28213 2490
rect 26421 2360 26441 2380
rect 26961 2359 26981 2379
rect 25106 2281 25126 2301
rect 25646 2280 25666 2300
rect 22045 1936 22065 1956
rect 19769 1855 19789 1875
rect 22585 1935 22605 1955
rect 22418 1885 22438 1905
rect 22640 1883 22660 1903
rect 18814 1780 18838 1802
rect 20127 1802 20151 1824
rect 16458 1688 16478 1708
rect 16998 1687 17018 1707
rect 19176 1729 19196 1749
rect 13397 1343 13417 1363
rect 13937 1342 13957 1362
rect 12095 1263 12115 1283
rect 12635 1262 12655 1282
rect 12019 1076 12039 1096
rect 10565 1026 10586 1045
rect 13779 1288 13799 1308
rect 13992 1290 14012 1310
rect 14811 1345 14831 1365
rect 14195 1159 14215 1179
rect 14014 1117 14034 1137
rect 14735 1158 14755 1178
rect 14579 1103 14598 1121
rect 14790 1106 14810 1126
rect 13398 931 13418 951
rect 13938 930 13958 950
rect 13771 880 13791 900
rect 13993 878 14013 898
rect 12788 813 12820 838
rect 10167 775 10191 797
rect 15606 1512 15626 1532
rect 15819 1514 15840 1533
rect 15661 1460 15681 1480
rect 16382 1501 16402 1521
rect 16201 1459 16221 1479
rect 15585 1273 15605 1293
rect 16404 1328 16424 1348
rect 16617 1330 16637 1350
rect 18560 1543 18580 1563
rect 18279 1503 18299 1523
rect 19100 1542 19120 1562
rect 18945 1486 18964 1503
rect 19155 1490 19175 1510
rect 24154 2107 24174 2127
rect 24365 2108 24386 2127
rect 24209 2055 24229 2075
rect 25030 2094 25050 2114
rect 24749 2054 24769 2074
rect 26803 2305 26823 2325
rect 27016 2307 27036 2327
rect 27835 2362 27855 2382
rect 27992 2276 28014 2294
rect 27219 2176 27239 2196
rect 27038 2134 27058 2154
rect 27759 2175 27779 2195
rect 27600 2122 27621 2141
rect 27814 2123 27834 2143
rect 32337 3087 32358 3106
rect 31939 2836 31963 2858
rect 29427 2757 29447 2777
rect 29649 2755 29669 2775
rect 29482 2705 29502 2725
rect 30022 2704 30042 2724
rect 32364 2783 32384 2803
rect 28630 2529 28650 2549
rect 28842 2534 28861 2552
rect 28685 2477 28705 2497
rect 29406 2518 29426 2538
rect 29225 2476 29245 2496
rect 28609 2290 28629 2310
rect 29428 2345 29448 2365
rect 29641 2347 29661 2367
rect 31748 2597 31768 2617
rect 31401 2559 31421 2579
rect 32288 2596 32308 2616
rect 32129 2544 32152 2566
rect 32343 2544 32363 2564
rect 33828 4806 33848 4826
rect 34050 4804 34070 4824
rect 33883 4754 33903 4774
rect 34423 4753 34443 4773
rect 33031 4578 33051 4598
rect 33243 4583 33262 4601
rect 33086 4526 33106 4546
rect 33807 4567 33827 4587
rect 33626 4525 33646 4545
rect 33010 4339 33030 4359
rect 32828 4241 32850 4259
rect 33829 4394 33849 4414
rect 34042 4396 34062 4416
rect 33884 4342 33904 4362
rect 34424 4341 34444 4361
rect 32932 4168 32952 4188
rect 33143 4175 33162 4192
rect 32987 4116 33007 4136
rect 33808 4155 33828 4175
rect 33527 4115 33547 4135
rect 32911 3929 32931 3949
rect 33269 3876 33293 3898
rect 33811 3788 33831 3808
rect 34033 3786 34053 3806
rect 33866 3736 33886 3756
rect 34406 3735 34426 3755
rect 33014 3560 33034 3580
rect 33227 3562 33248 3581
rect 33069 3508 33089 3528
rect 33790 3549 33810 3569
rect 33609 3507 33629 3527
rect 32993 3321 33013 3341
rect 33812 3376 33832 3396
rect 34025 3378 34045 3398
rect 33867 3324 33887 3344
rect 34407 3323 34427 3343
rect 32849 3152 32869 3172
rect 33062 3155 33080 3173
rect 32904 3100 32924 3120
rect 33791 3137 33811 3157
rect 33444 3099 33464 3119
rect 32828 2913 32848 2933
rect 33249 2858 33273 2880
rect 32854 2610 32875 2629
rect 32553 2481 32577 2503
rect 30785 2373 30805 2393
rect 31325 2372 31345 2392
rect 29483 2293 29503 2313
rect 30023 2292 30043 2312
rect 26422 1948 26442 1968
rect 24133 1868 24153 1888
rect 26962 1947 26982 1967
rect 26795 1897 26815 1917
rect 27017 1895 27037 1915
rect 23178 1793 23202 1815
rect 24491 1815 24515 1837
rect 20669 1714 20689 1734
rect 20891 1712 20911 1732
rect 20724 1662 20744 1682
rect 23540 1742 23560 1762
rect 21264 1661 21284 1681
rect 16459 1276 16479 1296
rect 17663 1317 17683 1337
rect 16999 1275 17019 1295
rect 18203 1316 18223 1336
rect 16383 1089 16403 1109
rect 14929 1039 14950 1058
rect 18045 1262 18065 1282
rect 18258 1264 18278 1284
rect 19077 1319 19097 1339
rect 18461 1133 18481 1153
rect 18280 1091 18300 1111
rect 19001 1132 19021 1152
rect 18845 1077 18864 1095
rect 19056 1080 19076 1100
rect 17664 905 17684 925
rect 18204 904 18224 924
rect 17152 826 17184 851
rect 18037 854 18057 874
rect 18259 852 18279 872
rect 14531 788 14555 810
rect 506 698 542 725
rect 4870 711 4906 738
rect 9247 723 9283 750
rect 13611 736 13647 763
rect 19872 1486 19892 1506
rect 20085 1488 20106 1507
rect 19927 1434 19947 1454
rect 20648 1475 20668 1495
rect 20467 1433 20487 1453
rect 19851 1247 19871 1267
rect 20670 1302 20690 1322
rect 20883 1304 20903 1324
rect 22924 1556 22944 1576
rect 22643 1516 22663 1536
rect 23464 1555 23484 1575
rect 23309 1499 23328 1516
rect 23519 1503 23539 1523
rect 28531 2119 28551 2139
rect 28742 2120 28763 2139
rect 28586 2067 28606 2087
rect 29407 2106 29427 2126
rect 29126 2066 29146 2086
rect 31167 2318 31187 2338
rect 31380 2320 31400 2340
rect 32199 2375 32219 2395
rect 32356 2289 32378 2307
rect 31583 2189 31603 2209
rect 31402 2147 31422 2167
rect 32123 2188 32143 2208
rect 31964 2135 31985 2154
rect 32178 2136 32198 2156
rect 33791 2770 33811 2790
rect 34013 2768 34033 2788
rect 33846 2718 33866 2738
rect 34386 2717 34406 2737
rect 32994 2542 33014 2562
rect 33206 2547 33225 2565
rect 33049 2490 33069 2510
rect 33770 2531 33790 2551
rect 33589 2489 33609 2509
rect 32973 2303 32993 2323
rect 33792 2358 33812 2378
rect 34005 2360 34025 2380
rect 33847 2306 33867 2326
rect 34387 2305 34407 2325
rect 30786 1961 30806 1981
rect 28510 1880 28530 1900
rect 31326 1960 31346 1980
rect 31159 1910 31179 1930
rect 31381 1908 31401 1928
rect 27555 1805 27579 1827
rect 28868 1827 28892 1849
rect 25033 1727 25053 1747
rect 25255 1725 25275 1745
rect 25088 1675 25108 1695
rect 27917 1754 27937 1774
rect 25628 1674 25648 1694
rect 22027 1330 22047 1350
rect 22567 1329 22587 1349
rect 20725 1250 20745 1270
rect 21265 1249 21285 1269
rect 20649 1063 20669 1083
rect 19195 1013 19216 1032
rect 22409 1275 22429 1295
rect 22622 1277 22642 1297
rect 23441 1332 23461 1352
rect 22825 1146 22845 1166
rect 22644 1104 22664 1124
rect 23365 1145 23385 1165
rect 23209 1090 23228 1108
rect 23420 1093 23440 1113
rect 22028 918 22048 938
rect 22568 917 22588 937
rect 22401 867 22421 887
rect 22623 865 22643 885
rect 21418 800 21450 825
rect 18797 762 18821 784
rect 24236 1499 24256 1519
rect 24449 1501 24470 1520
rect 24291 1447 24311 1467
rect 25012 1488 25032 1508
rect 24831 1446 24851 1466
rect 24215 1260 24235 1280
rect 25034 1315 25054 1335
rect 25247 1317 25267 1337
rect 27301 1568 27321 1588
rect 27020 1528 27040 1548
rect 27841 1567 27861 1587
rect 27686 1511 27705 1528
rect 27896 1515 27916 1535
rect 32895 2132 32915 2152
rect 33106 2133 33127 2152
rect 32950 2080 32970 2100
rect 33771 2119 33791 2139
rect 33490 2079 33510 2099
rect 32874 1893 32894 1913
rect 31919 1818 31943 1840
rect 33232 1840 33256 1862
rect 29410 1739 29430 1759
rect 29632 1737 29652 1757
rect 29465 1687 29485 1707
rect 32281 1767 32301 1787
rect 30005 1686 30025 1706
rect 26404 1342 26424 1362
rect 26944 1341 26964 1361
rect 25089 1263 25109 1283
rect 25629 1262 25649 1282
rect 25013 1076 25033 1096
rect 23559 1026 23580 1045
rect 26786 1287 26806 1307
rect 26999 1289 27019 1309
rect 27818 1344 27838 1364
rect 27202 1158 27222 1178
rect 27021 1116 27041 1136
rect 27742 1157 27762 1177
rect 27586 1102 27605 1120
rect 27797 1105 27817 1125
rect 26405 930 26425 950
rect 26945 929 26965 949
rect 26778 879 26798 899
rect 27000 877 27020 897
rect 25782 813 25814 838
rect 23161 775 23185 797
rect 28613 1511 28633 1531
rect 28826 1513 28847 1532
rect 28668 1459 28688 1479
rect 29389 1500 29409 1520
rect 29208 1458 29228 1478
rect 28592 1272 28612 1292
rect 29411 1327 29431 1347
rect 29624 1329 29644 1349
rect 31665 1581 31685 1601
rect 31384 1541 31404 1561
rect 32205 1580 32225 1600
rect 32050 1524 32069 1541
rect 32260 1528 32280 1548
rect 33774 1752 33794 1772
rect 33996 1750 34016 1770
rect 33829 1700 33849 1720
rect 34369 1699 34389 1719
rect 30768 1355 30788 1375
rect 31308 1354 31328 1374
rect 29466 1275 29486 1295
rect 30006 1274 30026 1294
rect 29390 1088 29410 1108
rect 27936 1038 27957 1057
rect 31150 1300 31170 1320
rect 31363 1302 31383 1322
rect 32182 1357 32202 1377
rect 31566 1171 31586 1191
rect 31385 1129 31405 1149
rect 32106 1170 32126 1190
rect 31950 1115 31969 1133
rect 32161 1118 32181 1138
rect 30769 943 30789 963
rect 31309 942 31329 962
rect 31142 892 31162 912
rect 31364 890 31384 910
rect 30159 825 30191 850
rect 27538 787 27562 809
rect 32977 1524 32997 1544
rect 33190 1526 33211 1545
rect 33032 1472 33052 1492
rect 33753 1513 33773 1533
rect 33572 1471 33592 1491
rect 32956 1285 32976 1305
rect 33775 1340 33795 1360
rect 33988 1342 34008 1362
rect 33830 1288 33850 1308
rect 34370 1287 34390 1307
rect 33754 1101 33774 1121
rect 32300 1051 32321 1070
rect 34523 838 34555 863
rect 31902 800 31926 822
rect 17877 710 17913 737
rect 22241 723 22277 750
rect 26618 735 26654 762
rect 30982 748 31018 775
rect 2122 502 2143 523
rect 6486 515 6507 536
rect 10863 527 10884 548
rect 15227 540 15248 561
rect 2204 409 2224 429
rect 4611 428 4632 449
rect 1506 317 1526 337
rect 2046 316 2066 336
rect 1888 259 1911 283
rect 2101 264 2121 284
rect 6568 422 6588 442
rect 9059 452 9080 473
rect 4693 335 4713 355
rect 5870 330 5890 350
rect 3995 243 4015 263
rect 4535 242 4555 262
rect 4380 184 4397 205
rect 4590 190 4610 210
rect 6410 329 6430 349
rect 6255 273 6278 297
rect 6465 277 6485 297
rect 9141 359 9161 379
rect 10945 434 10965 454
rect 13352 453 13373 474
rect 8443 267 8463 287
rect 8983 266 9003 286
rect 8819 209 8840 227
rect 9038 214 9058 234
rect 10247 342 10267 362
rect 10787 341 10807 361
rect 10629 284 10652 308
rect 10842 289 10862 309
rect 19493 514 19514 535
rect 23857 527 23878 548
rect 28234 539 28255 560
rect 32598 552 32619 573
rect 15309 447 15329 467
rect 13434 360 13454 380
rect 14611 355 14631 375
rect 12736 268 12756 288
rect 13276 267 13296 287
rect 13117 211 13138 233
rect 13331 215 13351 235
rect 15151 354 15171 374
rect 14996 298 15019 322
rect 15206 302 15226 322
rect 17549 389 17570 410
rect 19575 421 19595 441
rect 21982 440 22003 461
rect 18877 329 18897 349
rect 17631 296 17651 316
rect 19417 328 19437 348
rect 16933 204 16953 224
rect 17473 203 17493 223
rect 17528 151 17548 171
rect 19259 271 19282 295
rect 19472 276 19492 296
rect 23939 434 23959 454
rect 26430 464 26451 485
rect 22064 347 22084 367
rect 23241 342 23261 362
rect 21366 255 21386 275
rect 21906 254 21926 274
rect 21751 196 21768 217
rect 21961 202 21981 222
rect 23781 341 23801 361
rect 23626 285 23649 309
rect 23836 289 23856 309
rect 26512 371 26532 391
rect 28316 446 28336 466
rect 30723 465 30744 486
rect 25814 279 25834 299
rect 26354 278 26374 298
rect 26195 221 26218 242
rect 26409 226 26429 246
rect 27618 354 27638 374
rect 28158 353 28178 373
rect 28000 296 28023 320
rect 28213 301 28233 321
rect 32680 459 32700 479
rect 30805 372 30825 392
rect 31982 367 32002 387
rect 30107 280 30127 300
rect 30647 279 30667 299
rect 30488 223 30509 245
rect 30702 227 30722 247
rect 32522 366 32542 386
rect 32367 310 32390 334
rect 32577 314 32597 334
<< metal1 >>
rect 33863 8996 34149 8997
rect 33348 8988 34151 8996
rect 16492 8984 16778 8985
rect 15977 8976 16780 8984
rect 29499 8983 29785 8984
rect 12128 8971 12414 8972
rect 11613 8963 12416 8971
rect 7751 8959 8037 8960
rect 7236 8951 8039 8959
rect 3387 8946 3673 8947
rect 2872 8938 3675 8946
rect 2872 8921 2883 8938
rect 2873 8916 2883 8921
rect 2907 8921 3675 8938
rect 7236 8934 7247 8951
rect 2907 8916 2912 8921
rect 2873 8903 2912 8916
rect 3417 8855 3452 8856
rect 3396 8848 3452 8855
rect 3396 8828 3425 8848
rect 3445 8828 3452 8848
rect 3396 8823 3452 8828
rect 3636 8846 3675 8921
rect 7237 8929 7247 8934
rect 7271 8934 8039 8951
rect 11613 8946 11624 8963
rect 7271 8929 7276 8934
rect 7237 8916 7276 8929
rect 7781 8868 7816 8869
rect 3636 8826 3647 8846
rect 3667 8826 3675 8846
rect 2480 8687 2862 8692
rect 2480 8668 2488 8687
rect 2509 8668 2862 8687
rect 2480 8660 2862 8668
rect 1031 8642 1063 8643
rect 1028 8637 1063 8642
rect 1028 8617 1035 8637
rect 1055 8617 1063 8637
rect 2833 8630 2862 8660
rect 2620 8627 2655 8628
rect 1028 8609 1063 8617
rect 410 8451 995 8459
rect 410 8431 419 8451
rect 439 8450 995 8451
rect 439 8431 959 8450
rect 410 8430 959 8431
rect 979 8430 995 8450
rect 410 8424 995 8430
rect 1029 8403 1063 8609
rect 2599 8620 2655 8627
rect 2599 8600 2628 8620
rect 2648 8600 2655 8620
rect 2599 8595 2655 8600
rect 2832 8623 2866 8630
rect 2832 8605 2840 8623
rect 2859 8605 2866 8623
rect 2832 8597 2866 8605
rect 3396 8617 3430 8823
rect 3636 8822 3675 8826
rect 7760 8861 7816 8868
rect 7760 8841 7789 8861
rect 7809 8841 7816 8861
rect 7760 8836 7816 8841
rect 8000 8859 8039 8934
rect 11614 8941 11624 8946
rect 11648 8946 12416 8963
rect 15977 8959 15988 8976
rect 11648 8941 11653 8946
rect 11614 8928 11653 8941
rect 12158 8880 12193 8881
rect 8000 8839 8011 8859
rect 8031 8839 8039 8859
rect 3464 8796 4049 8802
rect 3464 8776 3480 8796
rect 3500 8795 4049 8796
rect 3500 8776 4020 8795
rect 3464 8775 4020 8776
rect 4040 8775 4049 8795
rect 3464 8767 4049 8775
rect 6844 8700 7226 8705
rect 6844 8681 6852 8700
rect 6873 8681 7226 8700
rect 6844 8673 7226 8681
rect 5395 8655 5427 8656
rect 5392 8650 5427 8655
rect 5392 8630 5399 8650
rect 5419 8630 5427 8650
rect 7197 8643 7226 8673
rect 6984 8640 7019 8641
rect 5392 8622 5427 8630
rect 3396 8609 3431 8617
rect 793 8396 828 8403
rect 793 8376 801 8396
rect 821 8376 828 8396
rect 793 8303 828 8376
rect 1007 8398 1063 8403
rect 1007 8378 1014 8398
rect 1034 8378 1063 8398
rect 1007 8371 1063 8378
rect 1098 8505 1128 8507
rect 1827 8505 1860 8506
rect 1098 8479 1861 8505
rect 1007 8370 1042 8371
rect 1098 8304 1128 8479
rect 1827 8458 1861 8479
rect 1826 8453 1861 8458
rect 1826 8433 1833 8453
rect 1853 8433 1861 8453
rect 1826 8425 1861 8433
rect 1093 8303 1128 8304
rect 792 8276 1128 8303
rect 1098 8275 1128 8276
rect 1208 8267 1793 8275
rect 1208 8247 1217 8267
rect 1237 8266 1793 8267
rect 1237 8247 1757 8266
rect 1208 8246 1757 8247
rect 1777 8246 1793 8266
rect 1208 8240 1793 8246
rect 1032 8230 1064 8231
rect 1029 8225 1064 8230
rect 1029 8205 1036 8225
rect 1056 8205 1064 8225
rect 1827 8219 1861 8425
rect 2599 8389 2633 8595
rect 3396 8589 3404 8609
rect 3424 8589 3431 8609
rect 3396 8584 3431 8589
rect 3396 8583 3428 8584
rect 2667 8568 3252 8574
rect 2667 8548 2683 8568
rect 2703 8567 3252 8568
rect 2703 8548 3223 8567
rect 2667 8547 3223 8548
rect 3243 8547 3252 8567
rect 2667 8539 3252 8547
rect 3332 8538 3362 8539
rect 3332 8511 3668 8538
rect 3332 8510 3367 8511
rect 2599 8381 2634 8389
rect 2599 8361 2607 8381
rect 2627 8361 2634 8381
rect 2599 8356 2634 8361
rect 2599 8335 2633 8356
rect 3332 8335 3362 8510
rect 3418 8443 3453 8444
rect 2599 8309 3362 8335
rect 2600 8308 2633 8309
rect 3332 8307 3362 8309
rect 3397 8436 3453 8443
rect 3397 8416 3426 8436
rect 3446 8416 3453 8436
rect 3397 8411 3453 8416
rect 3632 8438 3667 8511
rect 3632 8418 3639 8438
rect 3659 8418 3667 8438
rect 4774 8464 5359 8472
rect 4774 8444 4783 8464
rect 4803 8463 5359 8464
rect 4803 8444 5323 8463
rect 4774 8443 5323 8444
rect 5343 8443 5359 8463
rect 4774 8437 5359 8443
rect 3632 8411 3667 8418
rect 5393 8416 5427 8622
rect 6963 8633 7019 8640
rect 6963 8613 6992 8633
rect 7012 8613 7019 8633
rect 6963 8608 7019 8613
rect 7196 8636 7230 8643
rect 7196 8618 7204 8636
rect 7223 8618 7230 8636
rect 7196 8610 7230 8618
rect 7760 8630 7794 8836
rect 8000 8835 8039 8839
rect 12137 8873 12193 8880
rect 12137 8853 12166 8873
rect 12186 8853 12193 8873
rect 12137 8848 12193 8853
rect 12377 8871 12416 8946
rect 15978 8954 15988 8959
rect 16012 8959 16780 8976
rect 28984 8975 29787 8983
rect 25122 8971 25408 8972
rect 24607 8963 25410 8971
rect 16012 8954 16017 8959
rect 15978 8941 16017 8954
rect 16522 8893 16557 8894
rect 12377 8851 12388 8871
rect 12408 8851 12416 8871
rect 7828 8809 8413 8815
rect 7828 8789 7844 8809
rect 7864 8808 8413 8809
rect 7864 8789 8384 8808
rect 7828 8788 8384 8789
rect 8404 8788 8413 8808
rect 7828 8780 8413 8788
rect 11221 8712 11603 8717
rect 11221 8693 11229 8712
rect 11250 8693 11603 8712
rect 11221 8685 11603 8693
rect 9772 8667 9804 8668
rect 9769 8662 9804 8667
rect 9769 8642 9776 8662
rect 9796 8642 9804 8662
rect 11574 8655 11603 8685
rect 11361 8652 11396 8653
rect 9769 8634 9804 8642
rect 7760 8622 7795 8630
rect 1029 8197 1064 8205
rect 411 8039 996 8047
rect 411 8019 420 8039
rect 440 8038 996 8039
rect 440 8019 960 8038
rect 411 8018 960 8019
rect 980 8018 996 8038
rect 411 8012 996 8018
rect 785 7988 824 7992
rect 1030 7991 1064 8197
rect 1593 8212 1628 8218
rect 1593 8193 1598 8212
rect 1619 8193 1628 8212
rect 1593 8184 1628 8193
rect 1805 8214 1861 8219
rect 1805 8194 1812 8214
rect 1832 8194 1861 8214
rect 1805 8187 1861 8194
rect 2428 8258 2762 8286
rect 1805 8186 1840 8187
rect 1597 8116 1626 8184
rect 1597 8082 1943 8116
rect 785 7968 793 7988
rect 813 7968 824 7988
rect 785 7893 824 7968
rect 1008 7986 1064 7991
rect 1008 7966 1015 7986
rect 1035 7966 1064 7986
rect 1008 7959 1064 7966
rect 1008 7958 1043 7959
rect 1548 7898 1587 7911
rect 1548 7893 1553 7898
rect 785 7876 1553 7893
rect 1577 7893 1587 7898
rect 1577 7876 1588 7893
rect 785 7868 1588 7876
rect 787 7867 1073 7868
rect 1904 7845 1943 8082
rect 1904 7833 1915 7845
rect 1908 7825 1915 7833
rect 1935 7825 1943 7845
rect 1908 7817 1943 7825
rect 1290 7659 1875 7667
rect 1290 7639 1299 7659
rect 1319 7658 1875 7659
rect 1319 7639 1839 7658
rect 1290 7638 1839 7639
rect 1859 7638 1875 7658
rect 1290 7632 1875 7638
rect 1014 7624 1046 7625
rect 1011 7619 1046 7624
rect 1011 7599 1018 7619
rect 1038 7599 1046 7619
rect 1909 7611 1943 7817
rect 1011 7591 1046 7599
rect 393 7433 978 7441
rect 393 7413 402 7433
rect 422 7432 978 7433
rect 422 7413 942 7432
rect 393 7412 942 7413
rect 962 7412 978 7432
rect 393 7406 978 7412
rect 1012 7385 1046 7591
rect 1677 7605 1708 7611
rect 1677 7586 1682 7605
rect 1703 7586 1708 7605
rect 1677 7544 1708 7586
rect 1887 7606 1943 7611
rect 1887 7586 1894 7606
rect 1914 7586 1943 7606
rect 1887 7579 1943 7586
rect 1887 7578 1922 7579
rect 1677 7516 2016 7544
rect 776 7378 811 7385
rect 776 7358 784 7378
rect 804 7358 811 7378
rect 776 7285 811 7358
rect 990 7380 1046 7385
rect 990 7360 997 7380
rect 1017 7360 1046 7380
rect 990 7353 1046 7360
rect 1081 7487 1111 7489
rect 1810 7487 1843 7488
rect 1081 7461 1844 7487
rect 990 7352 1025 7353
rect 1081 7286 1111 7461
rect 1810 7440 1844 7461
rect 1809 7435 1844 7440
rect 1809 7415 1816 7435
rect 1836 7415 1844 7435
rect 1809 7407 1844 7415
rect 1076 7285 1111 7286
rect 775 7258 1111 7285
rect 1081 7257 1111 7258
rect 1191 7249 1776 7257
rect 1191 7229 1200 7249
rect 1220 7248 1776 7249
rect 1220 7229 1740 7248
rect 1191 7228 1740 7229
rect 1760 7228 1776 7248
rect 1191 7222 1776 7228
rect 1015 7212 1047 7213
rect 1012 7207 1047 7212
rect 1012 7187 1019 7207
rect 1039 7187 1047 7207
rect 1810 7201 1844 7407
rect 1012 7179 1047 7187
rect 394 7021 979 7029
rect 394 7001 403 7021
rect 423 7020 979 7021
rect 423 7001 943 7020
rect 394 7000 943 7001
rect 963 7000 979 7020
rect 394 6994 979 7000
rect 768 6970 807 6974
rect 1013 6973 1047 7179
rect 1577 7191 1611 7199
rect 1577 7173 1584 7191
rect 1603 7173 1611 7191
rect 1577 7166 1611 7173
rect 1788 7196 1844 7201
rect 1788 7176 1795 7196
rect 1815 7176 1844 7196
rect 1788 7169 1844 7176
rect 1788 7168 1823 7169
rect 1581 7136 1610 7166
rect 1581 7128 1963 7136
rect 1581 7109 1934 7128
rect 1955 7109 1963 7128
rect 1581 7104 1963 7109
rect 768 6950 776 6970
rect 796 6950 807 6970
rect 768 6875 807 6950
rect 991 6968 1047 6973
rect 991 6948 998 6968
rect 1018 6948 1047 6968
rect 991 6941 1047 6948
rect 991 6940 1026 6941
rect 1531 6880 1570 6893
rect 1531 6875 1536 6880
rect 768 6858 1536 6875
rect 1560 6875 1570 6880
rect 1560 6858 1571 6875
rect 768 6850 1571 6858
rect 770 6849 1056 6850
rect 1987 6831 2016 7516
rect 2428 7449 2460 8258
rect 2736 8223 2762 8258
rect 2521 8217 2556 8218
rect 2500 8210 2556 8217
rect 2500 8190 2529 8210
rect 2549 8190 2556 8210
rect 2500 8185 2556 8190
rect 2732 8214 2768 8223
rect 2732 8197 2740 8214
rect 2759 8197 2768 8214
rect 2732 8188 2768 8197
rect 3397 8205 3431 8411
rect 5157 8409 5192 8416
rect 3465 8384 4050 8390
rect 3465 8364 3481 8384
rect 3501 8383 4050 8384
rect 3501 8364 4021 8383
rect 3465 8363 4021 8364
rect 4041 8363 4050 8383
rect 3465 8355 4050 8363
rect 5157 8389 5165 8409
rect 5185 8389 5192 8409
rect 5157 8316 5192 8389
rect 5371 8411 5427 8416
rect 5371 8391 5378 8411
rect 5398 8391 5427 8411
rect 5371 8384 5427 8391
rect 5462 8518 5492 8520
rect 6191 8518 6224 8519
rect 5462 8492 6225 8518
rect 5371 8383 5406 8384
rect 5462 8317 5492 8492
rect 6191 8471 6225 8492
rect 6190 8466 6225 8471
rect 6190 8446 6197 8466
rect 6217 8446 6225 8466
rect 6190 8438 6225 8446
rect 5457 8316 5492 8317
rect 5156 8289 5492 8316
rect 5462 8288 5492 8289
rect 5572 8280 6157 8288
rect 5572 8260 5581 8280
rect 5601 8279 6157 8280
rect 5601 8260 6121 8279
rect 5572 8259 6121 8260
rect 6141 8259 6157 8279
rect 5572 8253 6157 8259
rect 5396 8243 5428 8244
rect 5393 8238 5428 8243
rect 5393 8218 5400 8238
rect 5420 8218 5428 8238
rect 6191 8232 6225 8438
rect 6963 8402 6997 8608
rect 7760 8602 7768 8622
rect 7788 8602 7795 8622
rect 7760 8597 7795 8602
rect 7760 8596 7792 8597
rect 7031 8581 7616 8587
rect 7031 8561 7047 8581
rect 7067 8580 7616 8581
rect 7067 8561 7587 8580
rect 7031 8560 7587 8561
rect 7607 8560 7616 8580
rect 7031 8552 7616 8560
rect 7696 8551 7726 8552
rect 7696 8524 8032 8551
rect 7696 8523 7731 8524
rect 6963 8394 6998 8402
rect 6963 8374 6971 8394
rect 6991 8374 6998 8394
rect 6963 8369 6998 8374
rect 6963 8348 6997 8369
rect 7696 8348 7726 8523
rect 7782 8456 7817 8457
rect 6963 8322 7726 8348
rect 6964 8321 6997 8322
rect 7696 8320 7726 8322
rect 7761 8449 7817 8456
rect 7761 8429 7790 8449
rect 7810 8429 7817 8449
rect 7761 8424 7817 8429
rect 7996 8451 8031 8524
rect 7996 8431 8003 8451
rect 8023 8431 8031 8451
rect 9151 8476 9736 8484
rect 9151 8456 9160 8476
rect 9180 8475 9736 8476
rect 9180 8456 9700 8475
rect 9151 8455 9700 8456
rect 9720 8455 9736 8475
rect 9151 8449 9736 8455
rect 7996 8424 8031 8431
rect 9770 8428 9804 8634
rect 11340 8645 11396 8652
rect 11340 8625 11369 8645
rect 11389 8625 11396 8645
rect 11340 8620 11396 8625
rect 11573 8648 11607 8655
rect 11573 8630 11581 8648
rect 11600 8630 11607 8648
rect 11573 8622 11607 8630
rect 12137 8642 12171 8848
rect 12377 8847 12416 8851
rect 16501 8886 16557 8893
rect 16501 8866 16530 8886
rect 16550 8866 16557 8886
rect 16501 8861 16557 8866
rect 16741 8884 16780 8959
rect 20758 8958 21044 8959
rect 20243 8950 21046 8958
rect 20243 8933 20254 8950
rect 20244 8928 20254 8933
rect 20278 8933 21046 8950
rect 24607 8946 24618 8963
rect 20278 8928 20283 8933
rect 20244 8915 20283 8928
rect 16741 8864 16752 8884
rect 16772 8864 16780 8884
rect 20788 8867 20823 8868
rect 12205 8821 12790 8827
rect 12205 8801 12221 8821
rect 12241 8820 12790 8821
rect 12241 8801 12761 8820
rect 12205 8800 12761 8801
rect 12781 8800 12790 8820
rect 12205 8792 12790 8800
rect 15585 8725 15967 8730
rect 15585 8706 15593 8725
rect 15614 8706 15967 8725
rect 15585 8698 15967 8706
rect 14136 8680 14168 8681
rect 14133 8675 14168 8680
rect 14133 8655 14140 8675
rect 14160 8655 14168 8675
rect 15938 8668 15967 8698
rect 15725 8665 15760 8666
rect 14133 8647 14168 8655
rect 12137 8634 12172 8642
rect 5393 8210 5428 8218
rect 3397 8197 3432 8205
rect 2500 7979 2534 8185
rect 3397 8177 3405 8197
rect 3425 8177 3432 8197
rect 3397 8172 3432 8177
rect 3397 8171 3429 8172
rect 2568 8158 3153 8164
rect 2568 8138 2584 8158
rect 2604 8157 3153 8158
rect 2604 8138 3124 8157
rect 2568 8137 3124 8138
rect 3144 8137 3153 8157
rect 2568 8129 3153 8137
rect 4775 8052 5360 8060
rect 4775 8032 4784 8052
rect 4804 8051 5360 8052
rect 4804 8032 5324 8051
rect 4775 8031 5324 8032
rect 5344 8031 5360 8051
rect 4775 8025 5360 8031
rect 5149 8001 5188 8005
rect 5394 8004 5428 8210
rect 5957 8225 5992 8231
rect 5957 8206 5962 8225
rect 5983 8206 5992 8225
rect 5957 8197 5992 8206
rect 6169 8227 6225 8232
rect 6169 8207 6176 8227
rect 6196 8207 6225 8227
rect 6169 8200 6225 8207
rect 6792 8271 7126 8299
rect 6169 8199 6204 8200
rect 5961 8129 5990 8197
rect 5961 8095 6307 8129
rect 5149 7981 5157 8001
rect 5177 7981 5188 8001
rect 2500 7971 2535 7979
rect 2500 7951 2508 7971
rect 2528 7963 2535 7971
rect 2528 7951 2539 7963
rect 2500 7714 2539 7951
rect 3370 7928 3656 7929
rect 2855 7920 3658 7928
rect 2855 7903 2866 7920
rect 2856 7898 2866 7903
rect 2890 7903 3658 7920
rect 2890 7898 2895 7903
rect 2856 7885 2895 7898
rect 3400 7837 3435 7838
rect 3379 7830 3435 7837
rect 3379 7810 3408 7830
rect 3428 7810 3435 7830
rect 3379 7805 3435 7810
rect 3619 7828 3658 7903
rect 5149 7906 5188 7981
rect 5372 7999 5428 8004
rect 5372 7979 5379 7999
rect 5399 7979 5428 7999
rect 5372 7972 5428 7979
rect 5372 7971 5407 7972
rect 5912 7911 5951 7924
rect 5912 7906 5917 7911
rect 5149 7889 5917 7906
rect 5941 7906 5951 7911
rect 5941 7889 5952 7906
rect 5149 7881 5952 7889
rect 5151 7880 5437 7881
rect 6268 7858 6307 8095
rect 6268 7846 6279 7858
rect 6272 7838 6279 7846
rect 6299 7838 6307 7858
rect 6272 7830 6307 7838
rect 3619 7808 3630 7828
rect 3650 7808 3658 7828
rect 2500 7680 2846 7714
rect 2817 7612 2846 7680
rect 2603 7609 2638 7610
rect 2428 7431 2431 7449
rect 2453 7431 2460 7449
rect 2428 7419 2460 7431
rect 2582 7602 2638 7609
rect 2582 7582 2611 7602
rect 2631 7582 2638 7602
rect 2582 7577 2638 7582
rect 2815 7603 2850 7612
rect 2815 7584 2824 7603
rect 2845 7584 2850 7603
rect 2815 7578 2850 7584
rect 3379 7599 3413 7805
rect 3619 7804 3658 7808
rect 3447 7778 4032 7784
rect 3447 7758 3463 7778
rect 3483 7777 4032 7778
rect 3483 7758 4003 7777
rect 3447 7757 4003 7758
rect 4023 7757 4032 7777
rect 3447 7749 4032 7757
rect 5654 7672 6239 7680
rect 5654 7652 5663 7672
rect 5683 7671 6239 7672
rect 5683 7652 6203 7671
rect 5654 7651 6203 7652
rect 6223 7651 6239 7671
rect 5654 7645 6239 7651
rect 5378 7637 5410 7638
rect 5375 7632 5410 7637
rect 5375 7612 5382 7632
rect 5402 7612 5410 7632
rect 6273 7624 6307 7830
rect 5375 7604 5410 7612
rect 3379 7591 3414 7599
rect 2582 7371 2616 7577
rect 3379 7571 3387 7591
rect 3407 7571 3414 7591
rect 3379 7566 3414 7571
rect 3379 7565 3411 7566
rect 2650 7550 3235 7556
rect 2650 7530 2666 7550
rect 2686 7549 3235 7550
rect 2686 7530 3206 7549
rect 2650 7529 3206 7530
rect 3226 7529 3235 7549
rect 2650 7521 3235 7529
rect 3315 7520 3345 7521
rect 3315 7493 3651 7520
rect 3315 7492 3350 7493
rect 2582 7363 2617 7371
rect 2582 7343 2590 7363
rect 2610 7343 2617 7363
rect 2582 7338 2617 7343
rect 2582 7317 2616 7338
rect 3315 7317 3345 7492
rect 3401 7425 3436 7426
rect 2582 7291 3345 7317
rect 2583 7290 2616 7291
rect 3315 7289 3345 7291
rect 3380 7418 3436 7425
rect 3380 7398 3409 7418
rect 3429 7398 3436 7418
rect 3380 7393 3436 7398
rect 3615 7420 3650 7493
rect 3615 7400 3622 7420
rect 3642 7400 3650 7420
rect 4757 7446 5342 7454
rect 4757 7426 4766 7446
rect 4786 7445 5342 7446
rect 4786 7426 5306 7445
rect 4757 7425 5306 7426
rect 5326 7425 5342 7445
rect 4757 7419 5342 7425
rect 3615 7393 3650 7400
rect 5376 7398 5410 7604
rect 6041 7618 6072 7624
rect 6041 7599 6046 7618
rect 6067 7599 6072 7618
rect 6041 7557 6072 7599
rect 6251 7619 6307 7624
rect 6251 7599 6258 7619
rect 6278 7599 6307 7619
rect 6251 7592 6307 7599
rect 6251 7591 6286 7592
rect 6041 7529 6380 7557
rect 2220 7257 2683 7265
rect 2220 7235 2232 7257
rect 2256 7235 2683 7257
rect 2220 7234 2683 7235
rect 2222 7222 2261 7234
rect 2656 7203 2683 7234
rect 2438 7201 2473 7202
rect 2417 7194 2473 7201
rect 2417 7174 2446 7194
rect 2466 7174 2473 7194
rect 2417 7169 2473 7174
rect 2652 7194 2685 7203
rect 2652 7172 2657 7194
rect 2680 7172 2685 7194
rect 2417 6963 2451 7169
rect 2652 7166 2685 7172
rect 3380 7187 3414 7393
rect 5140 7391 5175 7398
rect 3448 7366 4033 7372
rect 3448 7346 3464 7366
rect 3484 7365 4033 7366
rect 3484 7346 4004 7365
rect 3448 7345 4004 7346
rect 4024 7345 4033 7365
rect 3448 7337 4033 7345
rect 5140 7371 5148 7391
rect 5168 7371 5175 7391
rect 5140 7298 5175 7371
rect 5354 7393 5410 7398
rect 5354 7373 5361 7393
rect 5381 7373 5410 7393
rect 5354 7366 5410 7373
rect 5445 7500 5475 7502
rect 6174 7500 6207 7501
rect 5445 7474 6208 7500
rect 5354 7365 5389 7366
rect 5445 7299 5475 7474
rect 6174 7453 6208 7474
rect 6173 7448 6208 7453
rect 6173 7428 6180 7448
rect 6200 7428 6208 7448
rect 6173 7420 6208 7428
rect 5440 7298 5475 7299
rect 5139 7271 5475 7298
rect 5445 7270 5475 7271
rect 5555 7262 6140 7270
rect 5555 7242 5564 7262
rect 5584 7261 6140 7262
rect 5584 7242 6104 7261
rect 5555 7241 6104 7242
rect 6124 7241 6140 7261
rect 5555 7235 6140 7241
rect 5379 7225 5411 7226
rect 5376 7220 5411 7225
rect 5376 7200 5383 7220
rect 5403 7200 5411 7220
rect 6174 7214 6208 7420
rect 5376 7192 5411 7200
rect 3380 7179 3415 7187
rect 3380 7159 3388 7179
rect 3408 7159 3415 7179
rect 3380 7154 3415 7159
rect 3380 7153 3412 7154
rect 2485 7142 3070 7148
rect 2485 7122 2501 7142
rect 2521 7141 3070 7142
rect 2521 7122 3041 7141
rect 2485 7121 3041 7122
rect 3061 7121 3070 7141
rect 2485 7113 3070 7121
rect 4758 7034 5343 7042
rect 4758 7014 4767 7034
rect 4787 7033 5343 7034
rect 4787 7014 5307 7033
rect 4758 7013 5307 7014
rect 5327 7013 5343 7033
rect 4758 7007 5343 7013
rect 5132 6983 5171 6987
rect 5377 6986 5411 7192
rect 5941 7204 5975 7212
rect 5941 7186 5948 7204
rect 5967 7186 5975 7204
rect 5941 7179 5975 7186
rect 6152 7209 6208 7214
rect 6152 7189 6159 7209
rect 6179 7189 6208 7209
rect 6152 7182 6208 7189
rect 6152 7181 6187 7182
rect 5945 7149 5974 7179
rect 5945 7141 6327 7149
rect 5945 7122 6298 7141
rect 6319 7122 6327 7141
rect 5945 7117 6327 7122
rect 5132 6963 5140 6983
rect 5160 6963 5171 6983
rect 2417 6962 2452 6963
rect 2385 6955 2452 6962
rect 2385 6935 2425 6955
rect 2445 6935 2452 6955
rect 2385 6932 2452 6935
rect 2385 6929 2450 6932
rect 1956 6828 2021 6831
rect 1954 6825 2021 6828
rect 1954 6805 1961 6825
rect 1981 6805 2021 6825
rect 1954 6798 2021 6805
rect 1954 6797 1989 6798
rect 1336 6639 1921 6647
rect 1336 6619 1345 6639
rect 1365 6638 1921 6639
rect 1365 6619 1885 6638
rect 1336 6618 1885 6619
rect 1905 6618 1921 6638
rect 1336 6612 1921 6618
rect 994 6606 1026 6607
rect 991 6601 1026 6606
rect 991 6581 998 6601
rect 1018 6581 1026 6601
rect 991 6573 1026 6581
rect 373 6415 958 6423
rect 373 6395 382 6415
rect 402 6414 958 6415
rect 402 6395 922 6414
rect 373 6394 922 6395
rect 942 6394 958 6414
rect 373 6388 958 6394
rect 992 6367 1026 6573
rect 1719 6583 1760 6594
rect 1955 6591 1989 6797
rect 1719 6565 1729 6583
rect 1747 6565 1760 6583
rect 1719 6557 1760 6565
rect 1933 6586 1989 6591
rect 1933 6566 1940 6586
rect 1960 6566 1989 6586
rect 1933 6559 1989 6566
rect 1933 6558 1968 6559
rect 1728 6527 1754 6557
rect 1728 6526 2066 6527
rect 1728 6490 2082 6526
rect 756 6360 791 6367
rect 756 6340 764 6360
rect 784 6340 791 6360
rect 756 6267 791 6340
rect 970 6362 1026 6367
rect 970 6342 977 6362
rect 997 6342 1026 6362
rect 970 6335 1026 6342
rect 1061 6469 1091 6471
rect 1790 6469 1823 6470
rect 1061 6443 1824 6469
rect 970 6334 1005 6335
rect 1061 6268 1091 6443
rect 1790 6422 1824 6443
rect 1789 6417 1824 6422
rect 1789 6397 1796 6417
rect 1816 6397 1824 6417
rect 1789 6389 1824 6397
rect 1056 6267 1091 6268
rect 755 6240 1091 6267
rect 1061 6239 1091 6240
rect 1171 6231 1756 6239
rect 1171 6211 1180 6231
rect 1200 6230 1756 6231
rect 1200 6211 1720 6230
rect 1171 6210 1720 6211
rect 1740 6210 1756 6230
rect 1171 6204 1756 6210
rect 995 6194 1027 6195
rect 992 6189 1027 6194
rect 992 6169 999 6189
rect 1019 6169 1027 6189
rect 1790 6183 1824 6389
rect 992 6161 1027 6169
rect 374 6003 959 6011
rect 374 5983 383 6003
rect 403 6002 959 6003
rect 403 5983 923 6002
rect 374 5982 923 5983
rect 943 5982 959 6002
rect 374 5976 959 5982
rect 748 5952 787 5956
rect 993 5955 1027 6161
rect 1556 6176 1591 6182
rect 1556 6157 1561 6176
rect 1582 6157 1591 6176
rect 1556 6148 1591 6157
rect 1768 6178 1824 6183
rect 1768 6158 1775 6178
rect 1795 6158 1824 6178
rect 1768 6151 1824 6158
rect 1768 6150 1803 6151
rect 1560 6080 1589 6148
rect 1560 6046 1906 6080
rect 748 5932 756 5952
rect 776 5932 787 5952
rect 748 5857 787 5932
rect 971 5950 1027 5955
rect 971 5930 978 5950
rect 998 5930 1027 5950
rect 971 5923 1027 5930
rect 971 5922 1006 5923
rect 1511 5862 1550 5875
rect 1511 5857 1516 5862
rect 748 5840 1516 5857
rect 1540 5857 1550 5862
rect 1540 5840 1551 5857
rect 748 5832 1551 5840
rect 750 5831 1036 5832
rect 1867 5809 1906 6046
rect 1867 5797 1878 5809
rect 1871 5789 1878 5797
rect 1898 5789 1906 5809
rect 1871 5781 1906 5789
rect 1253 5623 1838 5631
rect 1253 5603 1262 5623
rect 1282 5622 1838 5623
rect 1282 5603 1802 5622
rect 1253 5602 1802 5603
rect 1822 5602 1838 5622
rect 1253 5596 1838 5602
rect 977 5588 1009 5589
rect 974 5583 1009 5588
rect 974 5563 981 5583
rect 1001 5563 1009 5583
rect 1872 5575 1906 5781
rect 974 5555 1009 5563
rect 356 5397 941 5405
rect 356 5377 365 5397
rect 385 5396 941 5397
rect 385 5377 905 5396
rect 356 5376 905 5377
rect 925 5376 941 5396
rect 356 5370 941 5376
rect 975 5349 1009 5555
rect 1638 5563 1674 5572
rect 1638 5546 1647 5563
rect 1666 5546 1674 5563
rect 1638 5537 1674 5546
rect 1850 5570 1906 5575
rect 1850 5550 1857 5570
rect 1877 5550 1906 5570
rect 1850 5543 1906 5550
rect 1850 5542 1885 5543
rect 1644 5502 1670 5537
rect 1952 5502 1984 5503
rect 1644 5497 1984 5502
rect 1644 5479 1959 5497
rect 1981 5479 1984 5497
rect 1644 5474 1984 5479
rect 1952 5473 1984 5474
rect 739 5342 774 5349
rect 739 5322 747 5342
rect 767 5322 774 5342
rect 739 5249 774 5322
rect 953 5344 1009 5349
rect 953 5324 960 5344
rect 980 5324 1009 5344
rect 953 5317 1009 5324
rect 1044 5451 1074 5453
rect 1773 5451 1806 5452
rect 1044 5425 1807 5451
rect 953 5316 988 5317
rect 1044 5250 1074 5425
rect 1773 5404 1807 5425
rect 1772 5399 1807 5404
rect 1772 5379 1779 5399
rect 1799 5379 1807 5399
rect 1772 5371 1807 5379
rect 1039 5249 1074 5250
rect 738 5222 1074 5249
rect 1044 5221 1074 5222
rect 1154 5213 1739 5221
rect 1154 5193 1163 5213
rect 1183 5212 1739 5213
rect 1183 5193 1703 5212
rect 1154 5192 1703 5193
rect 1723 5192 1739 5212
rect 1154 5186 1739 5192
rect 978 5176 1010 5177
rect 975 5171 1010 5176
rect 975 5151 982 5171
rect 1002 5151 1010 5171
rect 1773 5165 1807 5371
rect 975 5143 1010 5151
rect 357 4985 942 4993
rect 357 4965 366 4985
rect 386 4984 942 4985
rect 386 4965 906 4984
rect 357 4964 906 4965
rect 926 4964 942 4984
rect 357 4958 942 4964
rect 731 4934 770 4938
rect 976 4937 1010 5143
rect 1540 5155 1574 5163
rect 1540 5137 1547 5155
rect 1566 5137 1574 5155
rect 1540 5130 1574 5137
rect 1751 5160 1807 5165
rect 1751 5140 1758 5160
rect 1778 5140 1807 5160
rect 1751 5133 1807 5140
rect 1751 5132 1786 5133
rect 1544 5100 1573 5130
rect 1544 5092 1926 5100
rect 1544 5073 1897 5092
rect 1918 5073 1926 5092
rect 1544 5068 1926 5073
rect 731 4914 739 4934
rect 759 4914 770 4934
rect 731 4839 770 4914
rect 954 4932 1010 4937
rect 954 4912 961 4932
rect 981 4912 1010 4932
rect 954 4905 1010 4912
rect 954 4904 989 4905
rect 1494 4844 1533 4857
rect 1494 4839 1499 4844
rect 731 4822 1499 4839
rect 1523 4839 1533 4844
rect 1523 4822 1534 4839
rect 731 4814 1534 4822
rect 733 4813 1019 4814
rect 2055 4790 2082 6490
rect 2390 6244 2419 6929
rect 3350 6910 3636 6911
rect 2835 6902 3638 6910
rect 2835 6885 2846 6902
rect 2836 6880 2846 6885
rect 2870 6885 3638 6902
rect 2870 6880 2875 6885
rect 2836 6867 2875 6880
rect 3380 6819 3415 6820
rect 3359 6812 3415 6819
rect 3359 6792 3388 6812
rect 3408 6792 3415 6812
rect 3359 6787 3415 6792
rect 3599 6810 3638 6885
rect 5132 6888 5171 6963
rect 5355 6981 5411 6986
rect 5355 6961 5362 6981
rect 5382 6961 5411 6981
rect 5355 6954 5411 6961
rect 5355 6953 5390 6954
rect 5895 6893 5934 6906
rect 5895 6888 5900 6893
rect 5132 6871 5900 6888
rect 5924 6888 5934 6893
rect 5924 6871 5935 6888
rect 5132 6863 5935 6871
rect 5134 6862 5420 6863
rect 6351 6844 6380 7529
rect 6792 7462 6824 8271
rect 7100 8236 7126 8271
rect 6885 8230 6920 8231
rect 6864 8223 6920 8230
rect 6864 8203 6893 8223
rect 6913 8203 6920 8223
rect 6864 8198 6920 8203
rect 7096 8227 7132 8236
rect 7096 8210 7104 8227
rect 7123 8210 7132 8227
rect 7096 8201 7132 8210
rect 7761 8218 7795 8424
rect 9534 8421 9569 8428
rect 7829 8397 8414 8403
rect 7829 8377 7845 8397
rect 7865 8396 8414 8397
rect 7865 8377 8385 8396
rect 7829 8376 8385 8377
rect 8405 8376 8414 8396
rect 7829 8368 8414 8376
rect 9534 8401 9542 8421
rect 9562 8401 9569 8421
rect 9534 8328 9569 8401
rect 9748 8423 9804 8428
rect 9748 8403 9755 8423
rect 9775 8403 9804 8423
rect 9748 8396 9804 8403
rect 9839 8530 9869 8532
rect 10568 8530 10601 8531
rect 9839 8504 10602 8530
rect 9748 8395 9783 8396
rect 9839 8329 9869 8504
rect 10568 8483 10602 8504
rect 10567 8478 10602 8483
rect 10567 8458 10574 8478
rect 10594 8458 10602 8478
rect 10567 8450 10602 8458
rect 9834 8328 9869 8329
rect 9533 8301 9869 8328
rect 9839 8300 9869 8301
rect 9949 8292 10534 8300
rect 9949 8272 9958 8292
rect 9978 8291 10534 8292
rect 9978 8272 10498 8291
rect 9949 8271 10498 8272
rect 10518 8271 10534 8291
rect 9949 8265 10534 8271
rect 9773 8255 9805 8256
rect 9770 8250 9805 8255
rect 9770 8230 9777 8250
rect 9797 8230 9805 8250
rect 10568 8244 10602 8450
rect 11340 8414 11374 8620
rect 12137 8614 12145 8634
rect 12165 8614 12172 8634
rect 12137 8609 12172 8614
rect 12137 8608 12169 8609
rect 11408 8593 11993 8599
rect 11408 8573 11424 8593
rect 11444 8592 11993 8593
rect 11444 8573 11964 8592
rect 11408 8572 11964 8573
rect 11984 8572 11993 8592
rect 11408 8564 11993 8572
rect 12073 8563 12103 8564
rect 12073 8536 12409 8563
rect 12073 8535 12108 8536
rect 11340 8406 11375 8414
rect 11340 8386 11348 8406
rect 11368 8386 11375 8406
rect 11340 8381 11375 8386
rect 11340 8360 11374 8381
rect 12073 8360 12103 8535
rect 12159 8468 12194 8469
rect 11340 8334 12103 8360
rect 11341 8333 11374 8334
rect 12073 8332 12103 8334
rect 12138 8461 12194 8468
rect 12138 8441 12167 8461
rect 12187 8441 12194 8461
rect 12138 8436 12194 8441
rect 12373 8463 12408 8536
rect 12373 8443 12380 8463
rect 12400 8443 12408 8463
rect 13515 8489 14100 8497
rect 13515 8469 13524 8489
rect 13544 8488 14100 8489
rect 13544 8469 14064 8488
rect 13515 8468 14064 8469
rect 14084 8468 14100 8488
rect 13515 8462 14100 8468
rect 12373 8436 12408 8443
rect 14134 8441 14168 8647
rect 15704 8658 15760 8665
rect 15704 8638 15733 8658
rect 15753 8638 15760 8658
rect 15704 8633 15760 8638
rect 15937 8661 15971 8668
rect 15937 8643 15945 8661
rect 15964 8643 15971 8661
rect 15937 8635 15971 8643
rect 16501 8655 16535 8861
rect 16741 8860 16780 8864
rect 20767 8860 20823 8867
rect 20767 8840 20796 8860
rect 20816 8840 20823 8860
rect 16569 8834 17154 8840
rect 16569 8814 16585 8834
rect 16605 8833 17154 8834
rect 16605 8814 17125 8833
rect 16569 8813 17125 8814
rect 17145 8813 17154 8833
rect 16569 8805 17154 8813
rect 20767 8835 20823 8840
rect 21007 8858 21046 8933
rect 24608 8941 24618 8946
rect 24642 8946 25410 8963
rect 28984 8958 28995 8975
rect 24642 8941 24647 8946
rect 24608 8928 24647 8941
rect 25152 8880 25187 8881
rect 21007 8838 21018 8858
rect 21038 8838 21046 8858
rect 19851 8699 20233 8704
rect 19851 8680 19859 8699
rect 19880 8680 20233 8699
rect 19851 8672 20233 8680
rect 16501 8647 16536 8655
rect 18402 8654 18434 8655
rect 9770 8222 9805 8230
rect 7761 8210 7796 8218
rect 6864 7992 6898 8198
rect 7761 8190 7769 8210
rect 7789 8190 7796 8210
rect 7761 8185 7796 8190
rect 7761 8184 7793 8185
rect 6932 8171 7517 8177
rect 6932 8151 6948 8171
rect 6968 8170 7517 8171
rect 6968 8151 7488 8170
rect 6932 8150 7488 8151
rect 7508 8150 7517 8170
rect 6932 8142 7517 8150
rect 9152 8064 9737 8072
rect 9152 8044 9161 8064
rect 9181 8063 9737 8064
rect 9181 8044 9701 8063
rect 9152 8043 9701 8044
rect 9721 8043 9737 8063
rect 9152 8037 9737 8043
rect 9526 8013 9565 8017
rect 9771 8016 9805 8222
rect 10334 8237 10369 8243
rect 10334 8218 10339 8237
rect 10360 8218 10369 8237
rect 10334 8209 10369 8218
rect 10546 8239 10602 8244
rect 10546 8219 10553 8239
rect 10573 8219 10602 8239
rect 10546 8212 10602 8219
rect 11169 8283 11503 8311
rect 10546 8211 10581 8212
rect 10338 8141 10367 8209
rect 10338 8107 10684 8141
rect 9526 7993 9534 8013
rect 9554 7993 9565 8013
rect 6864 7984 6899 7992
rect 6864 7964 6872 7984
rect 6892 7976 6899 7984
rect 6892 7964 6903 7976
rect 6864 7727 6903 7964
rect 7734 7941 8020 7942
rect 7219 7933 8022 7941
rect 7219 7916 7230 7933
rect 7220 7911 7230 7916
rect 7254 7916 8022 7933
rect 7254 7911 7259 7916
rect 7220 7898 7259 7911
rect 7764 7850 7799 7851
rect 7743 7843 7799 7850
rect 7743 7823 7772 7843
rect 7792 7823 7799 7843
rect 7743 7818 7799 7823
rect 7983 7841 8022 7916
rect 9526 7918 9565 7993
rect 9749 8011 9805 8016
rect 9749 7991 9756 8011
rect 9776 7991 9805 8011
rect 9749 7984 9805 7991
rect 9749 7983 9784 7984
rect 10289 7923 10328 7936
rect 10289 7918 10294 7923
rect 9526 7901 10294 7918
rect 10318 7918 10328 7923
rect 10318 7901 10329 7918
rect 9526 7893 10329 7901
rect 9528 7892 9814 7893
rect 10645 7870 10684 8107
rect 10645 7858 10656 7870
rect 10649 7850 10656 7858
rect 10676 7850 10684 7870
rect 10649 7842 10684 7850
rect 7983 7821 7994 7841
rect 8014 7821 8022 7841
rect 6864 7693 7210 7727
rect 7181 7625 7210 7693
rect 6967 7622 7002 7623
rect 6792 7444 6795 7462
rect 6817 7444 6824 7462
rect 6792 7432 6824 7444
rect 6946 7615 7002 7622
rect 6946 7595 6975 7615
rect 6995 7595 7002 7615
rect 6946 7590 7002 7595
rect 7179 7616 7214 7625
rect 7179 7597 7188 7616
rect 7209 7597 7214 7616
rect 7179 7591 7214 7597
rect 7743 7612 7777 7818
rect 7983 7817 8022 7821
rect 7811 7791 8396 7797
rect 7811 7771 7827 7791
rect 7847 7790 8396 7791
rect 7847 7771 8367 7790
rect 7811 7770 8367 7771
rect 8387 7770 8396 7790
rect 7811 7762 8396 7770
rect 10031 7684 10616 7692
rect 10031 7664 10040 7684
rect 10060 7683 10616 7684
rect 10060 7664 10580 7683
rect 10031 7663 10580 7664
rect 10600 7663 10616 7683
rect 10031 7657 10616 7663
rect 9755 7649 9787 7650
rect 9752 7644 9787 7649
rect 9752 7624 9759 7644
rect 9779 7624 9787 7644
rect 10650 7636 10684 7842
rect 9752 7616 9787 7624
rect 7743 7604 7778 7612
rect 6946 7384 6980 7590
rect 7743 7584 7751 7604
rect 7771 7584 7778 7604
rect 7743 7579 7778 7584
rect 7743 7578 7775 7579
rect 7014 7563 7599 7569
rect 7014 7543 7030 7563
rect 7050 7562 7599 7563
rect 7050 7543 7570 7562
rect 7014 7542 7570 7543
rect 7590 7542 7599 7562
rect 7014 7534 7599 7542
rect 7679 7533 7709 7534
rect 7679 7506 8015 7533
rect 7679 7505 7714 7506
rect 6946 7376 6981 7384
rect 6946 7356 6954 7376
rect 6974 7356 6981 7376
rect 6946 7351 6981 7356
rect 6946 7330 6980 7351
rect 7679 7330 7709 7505
rect 7765 7438 7800 7439
rect 6946 7304 7709 7330
rect 6947 7303 6980 7304
rect 7679 7302 7709 7304
rect 7744 7431 7800 7438
rect 7744 7411 7773 7431
rect 7793 7411 7800 7431
rect 7744 7406 7800 7411
rect 7979 7433 8014 7506
rect 7979 7413 7986 7433
rect 8006 7413 8014 7433
rect 9134 7458 9719 7466
rect 9134 7438 9143 7458
rect 9163 7457 9719 7458
rect 9163 7438 9683 7457
rect 9134 7437 9683 7438
rect 9703 7437 9719 7457
rect 9134 7431 9719 7437
rect 7979 7406 8014 7413
rect 9753 7410 9787 7616
rect 10418 7630 10449 7636
rect 10418 7611 10423 7630
rect 10444 7611 10449 7630
rect 10418 7569 10449 7611
rect 10628 7631 10684 7636
rect 10628 7611 10635 7631
rect 10655 7611 10684 7631
rect 10628 7604 10684 7611
rect 10628 7603 10663 7604
rect 10418 7541 10757 7569
rect 6584 7270 7047 7278
rect 6584 7248 6596 7270
rect 6620 7248 7047 7270
rect 6584 7247 7047 7248
rect 6586 7235 6625 7247
rect 7020 7216 7047 7247
rect 6802 7214 6837 7215
rect 6781 7207 6837 7214
rect 6781 7187 6810 7207
rect 6830 7187 6837 7207
rect 6781 7182 6837 7187
rect 7016 7207 7049 7216
rect 7016 7185 7021 7207
rect 7044 7185 7049 7207
rect 6781 6976 6815 7182
rect 7016 7179 7049 7185
rect 7744 7200 7778 7406
rect 9517 7403 9552 7410
rect 7812 7379 8397 7385
rect 7812 7359 7828 7379
rect 7848 7378 8397 7379
rect 7848 7359 8368 7378
rect 7812 7358 8368 7359
rect 8388 7358 8397 7378
rect 7812 7350 8397 7358
rect 9517 7383 9525 7403
rect 9545 7383 9552 7403
rect 9517 7310 9552 7383
rect 9731 7405 9787 7410
rect 9731 7385 9738 7405
rect 9758 7385 9787 7405
rect 9731 7378 9787 7385
rect 9822 7512 9852 7514
rect 10551 7512 10584 7513
rect 9822 7486 10585 7512
rect 9731 7377 9766 7378
rect 9822 7311 9852 7486
rect 10551 7465 10585 7486
rect 10550 7460 10585 7465
rect 10550 7440 10557 7460
rect 10577 7440 10585 7460
rect 10550 7432 10585 7440
rect 9817 7310 9852 7311
rect 9516 7283 9852 7310
rect 9822 7282 9852 7283
rect 9932 7274 10517 7282
rect 9932 7254 9941 7274
rect 9961 7273 10517 7274
rect 9961 7254 10481 7273
rect 9932 7253 10481 7254
rect 10501 7253 10517 7273
rect 9932 7247 10517 7253
rect 9756 7237 9788 7238
rect 9753 7232 9788 7237
rect 9753 7212 9760 7232
rect 9780 7212 9788 7232
rect 10551 7226 10585 7432
rect 9753 7204 9788 7212
rect 7744 7192 7779 7200
rect 7744 7172 7752 7192
rect 7772 7172 7779 7192
rect 7744 7167 7779 7172
rect 7744 7166 7776 7167
rect 6849 7155 7434 7161
rect 6849 7135 6865 7155
rect 6885 7154 7434 7155
rect 6885 7135 7405 7154
rect 6849 7134 7405 7135
rect 7425 7134 7434 7154
rect 6849 7126 7434 7134
rect 9135 7046 9720 7054
rect 9135 7026 9144 7046
rect 9164 7045 9720 7046
rect 9164 7026 9684 7045
rect 9135 7025 9684 7026
rect 9704 7025 9720 7045
rect 9135 7019 9720 7025
rect 9509 6995 9548 6999
rect 9754 6998 9788 7204
rect 10318 7216 10352 7224
rect 10318 7198 10325 7216
rect 10344 7198 10352 7216
rect 10318 7191 10352 7198
rect 10529 7221 10585 7226
rect 10529 7201 10536 7221
rect 10556 7201 10585 7221
rect 10529 7194 10585 7201
rect 10529 7193 10564 7194
rect 10322 7161 10351 7191
rect 10322 7153 10704 7161
rect 10322 7134 10675 7153
rect 10696 7134 10704 7153
rect 10322 7129 10704 7134
rect 6781 6975 6816 6976
rect 6749 6968 6816 6975
rect 6749 6948 6789 6968
rect 6809 6948 6816 6968
rect 6749 6945 6816 6948
rect 9509 6975 9517 6995
rect 9537 6975 9548 6995
rect 6749 6942 6814 6945
rect 6320 6841 6385 6844
rect 6318 6838 6385 6841
rect 6318 6818 6325 6838
rect 6345 6818 6385 6838
rect 6318 6811 6385 6818
rect 6318 6810 6353 6811
rect 3599 6790 3610 6810
rect 3630 6790 3638 6810
rect 2443 6651 2825 6656
rect 2443 6632 2451 6651
rect 2472 6632 2825 6651
rect 2443 6624 2825 6632
rect 2796 6594 2825 6624
rect 2583 6591 2618 6592
rect 2562 6584 2618 6591
rect 2562 6564 2591 6584
rect 2611 6564 2618 6584
rect 2562 6559 2618 6564
rect 2795 6587 2829 6594
rect 2795 6569 2803 6587
rect 2822 6569 2829 6587
rect 2795 6561 2829 6569
rect 3359 6581 3393 6787
rect 3599 6786 3638 6790
rect 3427 6760 4012 6766
rect 3427 6740 3443 6760
rect 3463 6759 4012 6760
rect 3463 6740 3983 6759
rect 3427 6739 3983 6740
rect 4003 6739 4012 6759
rect 3427 6731 4012 6739
rect 5700 6652 6285 6660
rect 5700 6632 5709 6652
rect 5729 6651 6285 6652
rect 5729 6632 6249 6651
rect 5700 6631 6249 6632
rect 6269 6631 6285 6651
rect 5700 6625 6285 6631
rect 5358 6619 5390 6620
rect 5355 6614 5390 6619
rect 5355 6594 5362 6614
rect 5382 6594 5390 6614
rect 5355 6586 5390 6594
rect 3359 6573 3394 6581
rect 2562 6353 2596 6559
rect 3359 6553 3367 6573
rect 3387 6553 3394 6573
rect 3359 6548 3394 6553
rect 3359 6547 3391 6548
rect 2630 6532 3215 6538
rect 2630 6512 2646 6532
rect 2666 6531 3215 6532
rect 2666 6512 3186 6531
rect 2630 6511 3186 6512
rect 3206 6511 3215 6531
rect 2630 6503 3215 6511
rect 3295 6502 3325 6503
rect 3295 6475 3631 6502
rect 3295 6474 3330 6475
rect 2562 6345 2597 6353
rect 2562 6325 2570 6345
rect 2590 6325 2597 6345
rect 2562 6320 2597 6325
rect 2562 6299 2596 6320
rect 3295 6299 3325 6474
rect 3381 6407 3416 6408
rect 2562 6273 3325 6299
rect 2563 6272 2596 6273
rect 3295 6271 3325 6273
rect 3360 6400 3416 6407
rect 3360 6380 3389 6400
rect 3409 6380 3416 6400
rect 3360 6375 3416 6380
rect 3595 6402 3630 6475
rect 3595 6382 3602 6402
rect 3622 6382 3630 6402
rect 4737 6428 5322 6436
rect 4737 6408 4746 6428
rect 4766 6427 5322 6428
rect 4766 6408 5286 6427
rect 4737 6407 5286 6408
rect 5306 6407 5322 6427
rect 4737 6401 5322 6407
rect 3595 6375 3630 6382
rect 5356 6380 5390 6586
rect 6083 6596 6124 6607
rect 6319 6604 6353 6810
rect 6083 6578 6093 6596
rect 6111 6578 6124 6596
rect 6083 6570 6124 6578
rect 6297 6599 6353 6604
rect 6297 6579 6304 6599
rect 6324 6579 6353 6599
rect 6297 6572 6353 6579
rect 6297 6571 6332 6572
rect 6092 6540 6118 6570
rect 6092 6539 6430 6540
rect 6092 6503 6446 6539
rect 2390 6216 2729 6244
rect 2484 6181 2519 6182
rect 2463 6174 2519 6181
rect 2463 6154 2492 6174
rect 2512 6154 2519 6174
rect 2463 6149 2519 6154
rect 2698 6174 2729 6216
rect 2698 6155 2703 6174
rect 2724 6155 2729 6174
rect 2698 6149 2729 6155
rect 3360 6169 3394 6375
rect 5120 6373 5155 6380
rect 3428 6348 4013 6354
rect 3428 6328 3444 6348
rect 3464 6347 4013 6348
rect 3464 6328 3984 6347
rect 3428 6327 3984 6328
rect 4004 6327 4013 6347
rect 3428 6319 4013 6327
rect 5120 6353 5128 6373
rect 5148 6353 5155 6373
rect 5120 6280 5155 6353
rect 5334 6375 5390 6380
rect 5334 6355 5341 6375
rect 5361 6355 5390 6375
rect 5334 6348 5390 6355
rect 5425 6482 5455 6484
rect 6154 6482 6187 6483
rect 5425 6456 6188 6482
rect 5334 6347 5369 6348
rect 5425 6281 5455 6456
rect 6154 6435 6188 6456
rect 6153 6430 6188 6435
rect 6153 6410 6160 6430
rect 6180 6410 6188 6430
rect 6153 6402 6188 6410
rect 5420 6280 5455 6281
rect 5119 6253 5455 6280
rect 5425 6252 5455 6253
rect 5535 6244 6120 6252
rect 5535 6224 5544 6244
rect 5564 6243 6120 6244
rect 5564 6224 6084 6243
rect 5535 6223 6084 6224
rect 6104 6223 6120 6243
rect 5535 6217 6120 6223
rect 5359 6207 5391 6208
rect 5356 6202 5391 6207
rect 5356 6182 5363 6202
rect 5383 6182 5391 6202
rect 6154 6196 6188 6402
rect 5356 6174 5391 6182
rect 3360 6161 3395 6169
rect 2463 5943 2497 6149
rect 3360 6141 3368 6161
rect 3388 6141 3395 6161
rect 3360 6136 3395 6141
rect 3360 6135 3392 6136
rect 2531 6122 3116 6128
rect 2531 6102 2547 6122
rect 2567 6121 3116 6122
rect 2567 6102 3087 6121
rect 2531 6101 3087 6102
rect 3107 6101 3116 6121
rect 2531 6093 3116 6101
rect 4738 6016 5323 6024
rect 4738 5996 4747 6016
rect 4767 6015 5323 6016
rect 4767 5996 5287 6015
rect 4738 5995 5287 5996
rect 5307 5995 5323 6015
rect 4738 5989 5323 5995
rect 5112 5965 5151 5969
rect 5357 5968 5391 6174
rect 5920 6189 5955 6195
rect 5920 6170 5925 6189
rect 5946 6170 5955 6189
rect 5920 6161 5955 6170
rect 6132 6191 6188 6196
rect 6132 6171 6139 6191
rect 6159 6171 6188 6191
rect 6132 6164 6188 6171
rect 6132 6163 6167 6164
rect 5924 6093 5953 6161
rect 5924 6059 6270 6093
rect 5112 5945 5120 5965
rect 5140 5945 5151 5965
rect 2463 5935 2498 5943
rect 2463 5915 2471 5935
rect 2491 5927 2498 5935
rect 2491 5915 2502 5927
rect 2463 5678 2502 5915
rect 3333 5892 3619 5893
rect 2818 5884 3621 5892
rect 2818 5867 2829 5884
rect 2819 5862 2829 5867
rect 2853 5867 3621 5884
rect 2853 5862 2858 5867
rect 2819 5849 2858 5862
rect 3363 5801 3398 5802
rect 3342 5794 3398 5801
rect 3342 5774 3371 5794
rect 3391 5774 3398 5794
rect 3342 5769 3398 5774
rect 3582 5792 3621 5867
rect 5112 5870 5151 5945
rect 5335 5963 5391 5968
rect 5335 5943 5342 5963
rect 5362 5943 5391 5963
rect 5335 5936 5391 5943
rect 5335 5935 5370 5936
rect 5875 5875 5914 5888
rect 5875 5870 5880 5875
rect 5112 5853 5880 5870
rect 5904 5870 5914 5875
rect 5904 5853 5915 5870
rect 5112 5845 5915 5853
rect 5114 5844 5400 5845
rect 6231 5822 6270 6059
rect 6231 5810 6242 5822
rect 6235 5802 6242 5810
rect 6262 5802 6270 5822
rect 6235 5794 6270 5802
rect 3582 5772 3593 5792
rect 3613 5772 3621 5792
rect 2463 5644 2809 5678
rect 2780 5576 2809 5644
rect 2566 5573 2601 5574
rect 2545 5566 2601 5573
rect 2545 5546 2574 5566
rect 2594 5546 2601 5566
rect 2545 5541 2601 5546
rect 2778 5567 2813 5576
rect 2778 5548 2787 5567
rect 2808 5548 2813 5567
rect 2778 5542 2813 5548
rect 3342 5563 3376 5769
rect 3582 5768 3621 5772
rect 3410 5742 3995 5748
rect 3410 5722 3426 5742
rect 3446 5741 3995 5742
rect 3446 5722 3966 5741
rect 3410 5721 3966 5722
rect 3986 5721 3995 5741
rect 3410 5713 3995 5721
rect 5617 5636 6202 5644
rect 5617 5616 5626 5636
rect 5646 5635 6202 5636
rect 5646 5616 6166 5635
rect 5617 5615 6166 5616
rect 6186 5615 6202 5635
rect 5617 5609 6202 5615
rect 5341 5601 5373 5602
rect 5338 5596 5373 5601
rect 5338 5576 5345 5596
rect 5365 5576 5373 5596
rect 6236 5588 6270 5794
rect 5338 5568 5373 5576
rect 3342 5555 3377 5563
rect 2545 5335 2579 5541
rect 3342 5535 3350 5555
rect 3370 5535 3377 5555
rect 3342 5530 3377 5535
rect 3342 5529 3374 5530
rect 2613 5514 3198 5520
rect 2613 5494 2629 5514
rect 2649 5513 3198 5514
rect 2649 5494 3169 5513
rect 2613 5493 3169 5494
rect 3189 5493 3198 5513
rect 2613 5485 3198 5493
rect 3278 5484 3308 5485
rect 3278 5457 3614 5484
rect 3278 5456 3313 5457
rect 2545 5327 2580 5335
rect 2545 5307 2553 5327
rect 2573 5307 2580 5327
rect 2545 5302 2580 5307
rect 2545 5281 2579 5302
rect 3278 5281 3308 5456
rect 3364 5389 3399 5390
rect 2545 5255 3308 5281
rect 2546 5254 2579 5255
rect 3278 5253 3308 5255
rect 3343 5382 3399 5389
rect 3343 5362 3372 5382
rect 3392 5362 3399 5382
rect 3343 5357 3399 5362
rect 3578 5384 3613 5457
rect 3578 5364 3585 5384
rect 3605 5364 3613 5384
rect 4720 5410 5305 5418
rect 4720 5390 4729 5410
rect 4749 5409 5305 5410
rect 4749 5390 5269 5409
rect 4720 5389 5269 5390
rect 5289 5389 5305 5409
rect 4720 5383 5305 5389
rect 3578 5357 3613 5364
rect 5339 5362 5373 5568
rect 6002 5576 6038 5585
rect 6002 5559 6011 5576
rect 6030 5559 6038 5576
rect 6002 5550 6038 5559
rect 6214 5583 6270 5588
rect 6214 5563 6221 5583
rect 6241 5563 6270 5583
rect 6214 5556 6270 5563
rect 6214 5555 6249 5556
rect 6008 5515 6034 5550
rect 6316 5515 6348 5516
rect 6008 5510 6348 5515
rect 6008 5492 6323 5510
rect 6345 5492 6348 5510
rect 6008 5487 6348 5492
rect 6316 5486 6348 5487
rect 2197 5234 2514 5237
rect 2197 5207 2200 5234
rect 2227 5207 2514 5234
rect 2197 5201 2514 5207
rect 2197 5198 2233 5201
rect 2478 5171 2514 5201
rect 2262 5167 2297 5168
rect 2241 5160 2297 5167
rect 2241 5140 2270 5160
rect 2290 5140 2297 5160
rect 2241 5135 2297 5140
rect 2476 5165 2514 5171
rect 2476 5139 2482 5165
rect 2508 5139 2514 5165
rect 2241 4936 2275 5135
rect 2476 5131 2514 5139
rect 3343 5151 3377 5357
rect 5103 5355 5138 5362
rect 3411 5330 3996 5336
rect 3411 5310 3427 5330
rect 3447 5329 3996 5330
rect 3447 5310 3967 5329
rect 3411 5309 3967 5310
rect 3987 5309 3996 5329
rect 3411 5301 3996 5309
rect 5103 5335 5111 5355
rect 5131 5335 5138 5355
rect 5103 5262 5138 5335
rect 5317 5357 5373 5362
rect 5317 5337 5324 5357
rect 5344 5337 5373 5357
rect 5317 5330 5373 5337
rect 5408 5464 5438 5466
rect 6137 5464 6170 5465
rect 5408 5438 6171 5464
rect 5317 5329 5352 5330
rect 5408 5263 5438 5438
rect 6137 5417 6171 5438
rect 6136 5412 6171 5417
rect 6136 5392 6143 5412
rect 6163 5392 6171 5412
rect 6136 5384 6171 5392
rect 5403 5262 5438 5263
rect 5102 5235 5438 5262
rect 5408 5234 5438 5235
rect 5518 5226 6103 5234
rect 5518 5206 5527 5226
rect 5547 5225 6103 5226
rect 5547 5206 6067 5225
rect 5518 5205 6067 5206
rect 6087 5205 6103 5225
rect 5518 5199 6103 5205
rect 5342 5189 5374 5190
rect 5339 5184 5374 5189
rect 5339 5164 5346 5184
rect 5366 5164 5374 5184
rect 6137 5178 6171 5384
rect 5339 5156 5374 5164
rect 3343 5143 3378 5151
rect 3343 5123 3351 5143
rect 3371 5123 3378 5143
rect 3343 5118 3378 5123
rect 3343 5117 3375 5118
rect 2309 5108 2894 5114
rect 2309 5088 2325 5108
rect 2345 5107 2894 5108
rect 2345 5088 2865 5107
rect 2309 5087 2865 5088
rect 2885 5087 2894 5107
rect 2309 5079 2894 5087
rect 4721 4998 5306 5006
rect 4721 4978 4730 4998
rect 4750 4997 5306 4998
rect 4750 4978 5270 4997
rect 4721 4977 5270 4978
rect 5290 4977 5306 4997
rect 4721 4971 5306 4977
rect 5095 4947 5134 4951
rect 5340 4950 5374 5156
rect 5904 5168 5938 5176
rect 5904 5150 5911 5168
rect 5930 5150 5938 5168
rect 5904 5143 5938 5150
rect 6115 5173 6171 5178
rect 6115 5153 6122 5173
rect 6142 5153 6171 5173
rect 6115 5146 6171 5153
rect 6115 5145 6150 5146
rect 5908 5113 5937 5143
rect 5908 5105 6290 5113
rect 5908 5086 6261 5105
rect 6282 5086 6290 5105
rect 5908 5081 6290 5086
rect 2241 4921 2278 4936
rect 2241 4901 2249 4921
rect 2269 4901 2278 4921
rect 2241 4898 2278 4901
rect 2055 4787 2092 4790
rect 2055 4767 2064 4787
rect 2084 4767 2092 4787
rect 2055 4752 2092 4767
rect 1439 4601 2024 4609
rect 1439 4581 1448 4601
rect 1468 4600 2024 4601
rect 1468 4581 1988 4600
rect 1439 4580 1988 4581
rect 2008 4580 2024 4600
rect 1439 4574 2024 4580
rect 958 4570 990 4571
rect 955 4565 990 4570
rect 955 4545 962 4565
rect 982 4545 990 4565
rect 2058 4553 2092 4752
rect 2036 4548 2092 4553
rect 955 4537 990 4545
rect 337 4379 922 4387
rect 337 4359 346 4379
rect 366 4378 922 4379
rect 366 4359 886 4378
rect 337 4358 886 4359
rect 906 4358 922 4378
rect 337 4352 922 4358
rect 956 4331 990 4537
rect 1818 4546 1853 4548
rect 1818 4540 1856 4546
rect 1818 4517 1826 4540
rect 1849 4517 1856 4540
rect 2036 4528 2043 4548
rect 2063 4528 2092 4548
rect 2036 4521 2092 4528
rect 2036 4520 2071 4521
rect 1818 4511 1856 4517
rect 1818 4498 1853 4511
rect 1816 4440 1853 4498
rect 720 4324 755 4331
rect 720 4304 728 4324
rect 748 4304 755 4324
rect 720 4231 755 4304
rect 934 4326 990 4331
rect 934 4306 941 4326
rect 961 4306 990 4326
rect 934 4299 990 4306
rect 1025 4433 1055 4435
rect 1754 4433 1787 4434
rect 1025 4407 1788 4433
rect 934 4298 969 4299
rect 1025 4232 1055 4407
rect 1754 4386 1788 4407
rect 1816 4423 1851 4440
rect 1816 4422 2110 4423
rect 1816 4421 2153 4422
rect 1816 4414 2158 4421
rect 1816 4388 2118 4414
rect 2149 4388 2158 4414
rect 1753 4381 1788 4386
rect 2109 4385 2158 4388
rect 1753 4361 1760 4381
rect 1780 4361 1788 4381
rect 2115 4380 2158 4385
rect 1753 4353 1788 4361
rect 1020 4231 1055 4232
rect 719 4204 1055 4231
rect 1025 4203 1055 4204
rect 1135 4195 1720 4203
rect 1135 4175 1144 4195
rect 1164 4194 1720 4195
rect 1164 4175 1684 4194
rect 1135 4174 1684 4175
rect 1704 4174 1720 4194
rect 1135 4168 1720 4174
rect 959 4158 991 4159
rect 956 4153 991 4158
rect 956 4133 963 4153
rect 983 4133 991 4153
rect 1754 4147 1788 4353
rect 956 4125 991 4133
rect 338 3967 923 3975
rect 338 3947 347 3967
rect 367 3966 923 3967
rect 367 3947 887 3966
rect 338 3946 887 3947
rect 907 3946 923 3966
rect 338 3940 923 3946
rect 712 3916 751 3920
rect 957 3919 991 4125
rect 1520 4140 1555 4146
rect 1520 4121 1525 4140
rect 1546 4121 1555 4140
rect 1520 4112 1555 4121
rect 1732 4142 1788 4147
rect 1732 4122 1739 4142
rect 1759 4122 1788 4142
rect 1732 4115 1788 4122
rect 1732 4114 1767 4115
rect 1524 4044 1553 4112
rect 1524 4010 1870 4044
rect 712 3896 720 3916
rect 740 3896 751 3916
rect 712 3821 751 3896
rect 935 3914 991 3919
rect 935 3894 942 3914
rect 962 3894 991 3914
rect 935 3887 991 3894
rect 935 3886 970 3887
rect 1475 3826 1514 3839
rect 1475 3821 1480 3826
rect 712 3804 1480 3821
rect 1504 3821 1514 3826
rect 1504 3804 1515 3821
rect 712 3796 1515 3804
rect 714 3795 1000 3796
rect 1831 3773 1870 4010
rect 1831 3761 1842 3773
rect 1835 3753 1842 3761
rect 1862 3753 1870 3773
rect 1835 3745 1870 3753
rect 1217 3587 1802 3595
rect 1217 3567 1226 3587
rect 1246 3586 1802 3587
rect 1246 3567 1766 3586
rect 1217 3566 1766 3567
rect 1786 3566 1802 3586
rect 1217 3560 1802 3566
rect 941 3552 973 3553
rect 938 3547 973 3552
rect 938 3527 945 3547
rect 965 3527 973 3547
rect 1836 3539 1870 3745
rect 938 3519 973 3527
rect 320 3361 905 3369
rect 320 3341 329 3361
rect 349 3360 905 3361
rect 349 3341 869 3360
rect 320 3340 869 3341
rect 889 3340 905 3360
rect 320 3334 905 3340
rect 939 3313 973 3519
rect 1604 3533 1635 3539
rect 1604 3514 1609 3533
rect 1630 3514 1635 3533
rect 1604 3472 1635 3514
rect 1814 3534 1870 3539
rect 1814 3514 1821 3534
rect 1841 3514 1870 3534
rect 1814 3507 1870 3514
rect 1814 3506 1849 3507
rect 1604 3444 1943 3472
rect 703 3306 738 3313
rect 703 3286 711 3306
rect 731 3286 738 3306
rect 703 3213 738 3286
rect 917 3308 973 3313
rect 917 3288 924 3308
rect 944 3288 973 3308
rect 917 3281 973 3288
rect 1008 3415 1038 3417
rect 1737 3415 1770 3416
rect 1008 3389 1771 3415
rect 917 3280 952 3281
rect 1008 3214 1038 3389
rect 1737 3368 1771 3389
rect 1736 3363 1771 3368
rect 1736 3343 1743 3363
rect 1763 3343 1771 3363
rect 1736 3335 1771 3343
rect 1003 3213 1038 3214
rect 702 3186 1038 3213
rect 1008 3185 1038 3186
rect 1118 3177 1703 3185
rect 1118 3157 1127 3177
rect 1147 3176 1703 3177
rect 1147 3157 1667 3176
rect 1118 3156 1667 3157
rect 1687 3156 1703 3176
rect 1118 3150 1703 3156
rect 942 3140 974 3141
rect 939 3135 974 3140
rect 939 3115 946 3135
rect 966 3115 974 3135
rect 1737 3129 1771 3335
rect 939 3107 974 3115
rect 321 2949 906 2957
rect 321 2929 330 2949
rect 350 2948 906 2949
rect 350 2929 870 2948
rect 321 2928 870 2929
rect 890 2928 906 2948
rect 321 2922 906 2928
rect 695 2898 734 2902
rect 940 2901 974 3107
rect 1504 3119 1538 3127
rect 1504 3101 1511 3119
rect 1530 3101 1538 3119
rect 1504 3094 1538 3101
rect 1715 3124 1771 3129
rect 1715 3104 1722 3124
rect 1742 3104 1771 3124
rect 1715 3097 1771 3104
rect 1715 3096 1750 3097
rect 1508 3064 1537 3094
rect 1508 3056 1890 3064
rect 1508 3037 1861 3056
rect 1882 3037 1890 3056
rect 1508 3032 1890 3037
rect 695 2878 703 2898
rect 723 2878 734 2898
rect 695 2803 734 2878
rect 918 2896 974 2901
rect 918 2876 925 2896
rect 945 2876 974 2896
rect 918 2869 974 2876
rect 918 2868 953 2869
rect 1458 2808 1497 2821
rect 1458 2803 1463 2808
rect 695 2786 1463 2803
rect 1487 2803 1497 2808
rect 1487 2786 1498 2803
rect 695 2778 1498 2786
rect 697 2777 983 2778
rect 1914 2759 1943 3444
rect 2251 3198 2278 4898
rect 5095 4927 5103 4947
rect 5123 4927 5134 4947
rect 3314 4874 3600 4875
rect 2799 4866 3602 4874
rect 2799 4849 2810 4866
rect 2800 4844 2810 4849
rect 2834 4849 3602 4866
rect 2834 4844 2839 4849
rect 2800 4831 2839 4844
rect 3344 4783 3379 4784
rect 3323 4776 3379 4783
rect 3323 4756 3352 4776
rect 3372 4756 3379 4776
rect 3323 4751 3379 4756
rect 3563 4774 3602 4849
rect 5095 4852 5134 4927
rect 5318 4945 5374 4950
rect 5318 4925 5325 4945
rect 5345 4925 5374 4945
rect 5318 4918 5374 4925
rect 5318 4917 5353 4918
rect 5858 4857 5897 4870
rect 5858 4852 5863 4857
rect 5095 4835 5863 4852
rect 5887 4852 5897 4857
rect 5887 4835 5898 4852
rect 5095 4827 5898 4835
rect 5097 4826 5383 4827
rect 3563 4754 3574 4774
rect 3594 4754 3602 4774
rect 6419 4803 6446 6503
rect 6754 6257 6783 6942
rect 7714 6923 8000 6924
rect 7199 6915 8002 6923
rect 7199 6898 7210 6915
rect 7200 6893 7210 6898
rect 7234 6898 8002 6915
rect 7234 6893 7239 6898
rect 7200 6880 7239 6893
rect 7744 6832 7779 6833
rect 7723 6825 7779 6832
rect 7723 6805 7752 6825
rect 7772 6805 7779 6825
rect 7723 6800 7779 6805
rect 7963 6823 8002 6898
rect 9509 6900 9548 6975
rect 9732 6993 9788 6998
rect 9732 6973 9739 6993
rect 9759 6973 9788 6993
rect 9732 6966 9788 6973
rect 9732 6965 9767 6966
rect 10272 6905 10311 6918
rect 10272 6900 10277 6905
rect 9509 6883 10277 6900
rect 10301 6900 10311 6905
rect 10301 6883 10312 6900
rect 9509 6875 10312 6883
rect 9511 6874 9797 6875
rect 10728 6856 10757 7541
rect 11169 7474 11201 8283
rect 11477 8248 11503 8283
rect 11262 8242 11297 8243
rect 11241 8235 11297 8242
rect 11241 8215 11270 8235
rect 11290 8215 11297 8235
rect 11241 8210 11297 8215
rect 11473 8239 11509 8248
rect 11473 8222 11481 8239
rect 11500 8222 11509 8239
rect 11473 8213 11509 8222
rect 12138 8230 12172 8436
rect 13898 8434 13933 8441
rect 12206 8409 12791 8415
rect 12206 8389 12222 8409
rect 12242 8408 12791 8409
rect 12242 8389 12762 8408
rect 12206 8388 12762 8389
rect 12782 8388 12791 8408
rect 12206 8380 12791 8388
rect 13898 8414 13906 8434
rect 13926 8414 13933 8434
rect 13898 8341 13933 8414
rect 14112 8436 14168 8441
rect 14112 8416 14119 8436
rect 14139 8416 14168 8436
rect 14112 8409 14168 8416
rect 14203 8543 14233 8545
rect 14932 8543 14965 8544
rect 14203 8517 14966 8543
rect 14112 8408 14147 8409
rect 14203 8342 14233 8517
rect 14932 8496 14966 8517
rect 14931 8491 14966 8496
rect 14931 8471 14938 8491
rect 14958 8471 14966 8491
rect 14931 8463 14966 8471
rect 14198 8341 14233 8342
rect 13897 8314 14233 8341
rect 14203 8313 14233 8314
rect 14313 8305 14898 8313
rect 14313 8285 14322 8305
rect 14342 8304 14898 8305
rect 14342 8285 14862 8304
rect 14313 8284 14862 8285
rect 14882 8284 14898 8304
rect 14313 8278 14898 8284
rect 14137 8268 14169 8269
rect 14134 8263 14169 8268
rect 14134 8243 14141 8263
rect 14161 8243 14169 8263
rect 14932 8257 14966 8463
rect 15704 8427 15738 8633
rect 16501 8627 16509 8647
rect 16529 8627 16536 8647
rect 16501 8622 16536 8627
rect 18399 8649 18434 8654
rect 18399 8629 18406 8649
rect 18426 8629 18434 8649
rect 20204 8642 20233 8672
rect 19991 8639 20026 8640
rect 16501 8621 16533 8622
rect 18399 8621 18434 8629
rect 15772 8606 16357 8612
rect 15772 8586 15788 8606
rect 15808 8605 16357 8606
rect 15808 8586 16328 8605
rect 15772 8585 16328 8586
rect 16348 8585 16357 8605
rect 15772 8577 16357 8585
rect 16437 8576 16467 8577
rect 16437 8549 16773 8576
rect 16437 8548 16472 8549
rect 15704 8419 15739 8427
rect 15704 8399 15712 8419
rect 15732 8399 15739 8419
rect 15704 8394 15739 8399
rect 15704 8373 15738 8394
rect 16437 8373 16467 8548
rect 16523 8481 16558 8482
rect 15704 8347 16467 8373
rect 15705 8346 15738 8347
rect 16437 8345 16467 8347
rect 16502 8474 16558 8481
rect 16502 8454 16531 8474
rect 16551 8454 16558 8474
rect 16502 8449 16558 8454
rect 16737 8476 16772 8549
rect 16737 8456 16744 8476
rect 16764 8456 16772 8476
rect 16737 8449 16772 8456
rect 17781 8463 18366 8471
rect 14134 8235 14169 8243
rect 12138 8222 12173 8230
rect 11241 8004 11275 8210
rect 12138 8202 12146 8222
rect 12166 8202 12173 8222
rect 12138 8197 12173 8202
rect 12138 8196 12170 8197
rect 11309 8183 11894 8189
rect 11309 8163 11325 8183
rect 11345 8182 11894 8183
rect 11345 8163 11865 8182
rect 11309 8162 11865 8163
rect 11885 8162 11894 8182
rect 11309 8154 11894 8162
rect 13516 8077 14101 8085
rect 13516 8057 13525 8077
rect 13545 8076 14101 8077
rect 13545 8057 14065 8076
rect 13516 8056 14065 8057
rect 14085 8056 14101 8076
rect 13516 8050 14101 8056
rect 13890 8026 13929 8030
rect 14135 8029 14169 8235
rect 14698 8250 14733 8256
rect 14698 8231 14703 8250
rect 14724 8231 14733 8250
rect 14698 8222 14733 8231
rect 14910 8252 14966 8257
rect 14910 8232 14917 8252
rect 14937 8232 14966 8252
rect 14910 8225 14966 8232
rect 15533 8296 15867 8324
rect 14910 8224 14945 8225
rect 14702 8154 14731 8222
rect 14702 8120 15048 8154
rect 13890 8006 13898 8026
rect 13918 8006 13929 8026
rect 11241 7996 11276 8004
rect 11241 7976 11249 7996
rect 11269 7988 11276 7996
rect 11269 7976 11280 7988
rect 11241 7739 11280 7976
rect 12111 7953 12397 7954
rect 11596 7945 12399 7953
rect 11596 7928 11607 7945
rect 11597 7923 11607 7928
rect 11631 7928 12399 7945
rect 11631 7923 11636 7928
rect 11597 7910 11636 7923
rect 12141 7862 12176 7863
rect 12120 7855 12176 7862
rect 12120 7835 12149 7855
rect 12169 7835 12176 7855
rect 12120 7830 12176 7835
rect 12360 7853 12399 7928
rect 13890 7931 13929 8006
rect 14113 8024 14169 8029
rect 14113 8004 14120 8024
rect 14140 8004 14169 8024
rect 14113 7997 14169 8004
rect 14113 7996 14148 7997
rect 14653 7936 14692 7949
rect 14653 7931 14658 7936
rect 13890 7914 14658 7931
rect 14682 7931 14692 7936
rect 14682 7914 14693 7931
rect 13890 7906 14693 7914
rect 13892 7905 14178 7906
rect 15009 7883 15048 8120
rect 15009 7871 15020 7883
rect 15013 7863 15020 7871
rect 15040 7863 15048 7883
rect 15013 7855 15048 7863
rect 12360 7833 12371 7853
rect 12391 7833 12399 7853
rect 11241 7705 11587 7739
rect 11558 7637 11587 7705
rect 11344 7634 11379 7635
rect 11169 7456 11172 7474
rect 11194 7456 11201 7474
rect 11169 7444 11201 7456
rect 11323 7627 11379 7634
rect 11323 7607 11352 7627
rect 11372 7607 11379 7627
rect 11323 7602 11379 7607
rect 11556 7628 11591 7637
rect 11556 7609 11565 7628
rect 11586 7609 11591 7628
rect 11556 7603 11591 7609
rect 12120 7624 12154 7830
rect 12360 7829 12399 7833
rect 12188 7803 12773 7809
rect 12188 7783 12204 7803
rect 12224 7802 12773 7803
rect 12224 7783 12744 7802
rect 12188 7782 12744 7783
rect 12764 7782 12773 7802
rect 12188 7774 12773 7782
rect 14395 7697 14980 7705
rect 14395 7677 14404 7697
rect 14424 7696 14980 7697
rect 14424 7677 14944 7696
rect 14395 7676 14944 7677
rect 14964 7676 14980 7696
rect 14395 7670 14980 7676
rect 14119 7662 14151 7663
rect 14116 7657 14151 7662
rect 14116 7637 14123 7657
rect 14143 7637 14151 7657
rect 15014 7649 15048 7855
rect 14116 7629 14151 7637
rect 12120 7616 12155 7624
rect 11323 7396 11357 7602
rect 12120 7596 12128 7616
rect 12148 7596 12155 7616
rect 12120 7591 12155 7596
rect 12120 7590 12152 7591
rect 11391 7575 11976 7581
rect 11391 7555 11407 7575
rect 11427 7574 11976 7575
rect 11427 7555 11947 7574
rect 11391 7554 11947 7555
rect 11967 7554 11976 7574
rect 11391 7546 11976 7554
rect 12056 7545 12086 7546
rect 12056 7518 12392 7545
rect 12056 7517 12091 7518
rect 11323 7388 11358 7396
rect 11323 7368 11331 7388
rect 11351 7368 11358 7388
rect 11323 7363 11358 7368
rect 11323 7342 11357 7363
rect 12056 7342 12086 7517
rect 12142 7450 12177 7451
rect 11323 7316 12086 7342
rect 11324 7315 11357 7316
rect 12056 7314 12086 7316
rect 12121 7443 12177 7450
rect 12121 7423 12150 7443
rect 12170 7423 12177 7443
rect 12121 7418 12177 7423
rect 12356 7445 12391 7518
rect 12356 7425 12363 7445
rect 12383 7425 12391 7445
rect 13498 7471 14083 7479
rect 13498 7451 13507 7471
rect 13527 7470 14083 7471
rect 13527 7451 14047 7470
rect 13498 7450 14047 7451
rect 14067 7450 14083 7470
rect 13498 7444 14083 7450
rect 12356 7418 12391 7425
rect 14117 7423 14151 7629
rect 14782 7643 14813 7649
rect 14782 7624 14787 7643
rect 14808 7624 14813 7643
rect 14782 7582 14813 7624
rect 14992 7644 15048 7649
rect 14992 7624 14999 7644
rect 15019 7624 15048 7644
rect 14992 7617 15048 7624
rect 14992 7616 15027 7617
rect 14782 7554 15121 7582
rect 10961 7282 11424 7290
rect 10961 7260 10973 7282
rect 10997 7260 11424 7282
rect 10961 7259 11424 7260
rect 10963 7247 11002 7259
rect 11397 7228 11424 7259
rect 11179 7226 11214 7227
rect 11158 7219 11214 7226
rect 11158 7199 11187 7219
rect 11207 7199 11214 7219
rect 11158 7194 11214 7199
rect 11393 7219 11426 7228
rect 11393 7197 11398 7219
rect 11421 7197 11426 7219
rect 11158 6988 11192 7194
rect 11393 7191 11426 7197
rect 12121 7212 12155 7418
rect 13881 7416 13916 7423
rect 12189 7391 12774 7397
rect 12189 7371 12205 7391
rect 12225 7390 12774 7391
rect 12225 7371 12745 7390
rect 12189 7370 12745 7371
rect 12765 7370 12774 7390
rect 12189 7362 12774 7370
rect 13881 7396 13889 7416
rect 13909 7396 13916 7416
rect 13881 7323 13916 7396
rect 14095 7418 14151 7423
rect 14095 7398 14102 7418
rect 14122 7398 14151 7418
rect 14095 7391 14151 7398
rect 14186 7525 14216 7527
rect 14915 7525 14948 7526
rect 14186 7499 14949 7525
rect 14095 7390 14130 7391
rect 14186 7324 14216 7499
rect 14915 7478 14949 7499
rect 14914 7473 14949 7478
rect 14914 7453 14921 7473
rect 14941 7453 14949 7473
rect 14914 7445 14949 7453
rect 14181 7323 14216 7324
rect 13880 7296 14216 7323
rect 14186 7295 14216 7296
rect 14296 7287 14881 7295
rect 14296 7267 14305 7287
rect 14325 7286 14881 7287
rect 14325 7267 14845 7286
rect 14296 7266 14845 7267
rect 14865 7266 14881 7286
rect 14296 7260 14881 7266
rect 14120 7250 14152 7251
rect 14117 7245 14152 7250
rect 14117 7225 14124 7245
rect 14144 7225 14152 7245
rect 14915 7239 14949 7445
rect 14117 7217 14152 7225
rect 12121 7204 12156 7212
rect 12121 7184 12129 7204
rect 12149 7184 12156 7204
rect 12121 7179 12156 7184
rect 12121 7178 12153 7179
rect 11226 7167 11811 7173
rect 11226 7147 11242 7167
rect 11262 7166 11811 7167
rect 11262 7147 11782 7166
rect 11226 7146 11782 7147
rect 11802 7146 11811 7166
rect 11226 7138 11811 7146
rect 13499 7059 14084 7067
rect 13499 7039 13508 7059
rect 13528 7058 14084 7059
rect 13528 7039 14048 7058
rect 13499 7038 14048 7039
rect 14068 7038 14084 7058
rect 13499 7032 14084 7038
rect 13873 7008 13912 7012
rect 14118 7011 14152 7217
rect 14682 7229 14716 7237
rect 14682 7211 14689 7229
rect 14708 7211 14716 7229
rect 14682 7204 14716 7211
rect 14893 7234 14949 7239
rect 14893 7214 14900 7234
rect 14920 7214 14949 7234
rect 14893 7207 14949 7214
rect 14893 7206 14928 7207
rect 14686 7174 14715 7204
rect 14686 7166 15068 7174
rect 14686 7147 15039 7166
rect 15060 7147 15068 7166
rect 14686 7142 15068 7147
rect 13873 6988 13881 7008
rect 13901 6988 13912 7008
rect 11158 6987 11193 6988
rect 11126 6980 11193 6987
rect 11126 6960 11166 6980
rect 11186 6960 11193 6980
rect 11126 6957 11193 6960
rect 11126 6954 11191 6957
rect 10697 6853 10762 6856
rect 7963 6803 7974 6823
rect 7994 6803 8002 6823
rect 10695 6850 10762 6853
rect 10695 6830 10702 6850
rect 10722 6830 10762 6850
rect 10695 6823 10762 6830
rect 10695 6822 10730 6823
rect 6807 6664 7189 6669
rect 6807 6645 6815 6664
rect 6836 6645 7189 6664
rect 6807 6637 7189 6645
rect 7160 6607 7189 6637
rect 6947 6604 6982 6605
rect 6926 6597 6982 6604
rect 6926 6577 6955 6597
rect 6975 6577 6982 6597
rect 6926 6572 6982 6577
rect 7159 6600 7193 6607
rect 7159 6582 7167 6600
rect 7186 6582 7193 6600
rect 7159 6574 7193 6582
rect 7723 6594 7757 6800
rect 7963 6799 8002 6803
rect 7791 6773 8376 6779
rect 7791 6753 7807 6773
rect 7827 6772 8376 6773
rect 7827 6753 8347 6772
rect 7791 6752 8347 6753
rect 8367 6752 8376 6772
rect 7791 6744 8376 6752
rect 10077 6664 10662 6672
rect 10077 6644 10086 6664
rect 10106 6663 10662 6664
rect 10106 6644 10626 6663
rect 10077 6643 10626 6644
rect 10646 6643 10662 6663
rect 10077 6637 10662 6643
rect 9735 6631 9767 6632
rect 9732 6626 9767 6631
rect 9732 6606 9739 6626
rect 9759 6606 9767 6626
rect 9732 6598 9767 6606
rect 7723 6586 7758 6594
rect 6926 6366 6960 6572
rect 7723 6566 7731 6586
rect 7751 6566 7758 6586
rect 7723 6561 7758 6566
rect 7723 6560 7755 6561
rect 6994 6545 7579 6551
rect 6994 6525 7010 6545
rect 7030 6544 7579 6545
rect 7030 6525 7550 6544
rect 6994 6524 7550 6525
rect 7570 6524 7579 6544
rect 6994 6516 7579 6524
rect 7659 6515 7689 6516
rect 7659 6488 7995 6515
rect 7659 6487 7694 6488
rect 6926 6358 6961 6366
rect 6926 6338 6934 6358
rect 6954 6338 6961 6358
rect 6926 6333 6961 6338
rect 6926 6312 6960 6333
rect 7659 6312 7689 6487
rect 7745 6420 7780 6421
rect 6926 6286 7689 6312
rect 6927 6285 6960 6286
rect 7659 6284 7689 6286
rect 7724 6413 7780 6420
rect 7724 6393 7753 6413
rect 7773 6393 7780 6413
rect 7724 6388 7780 6393
rect 7959 6415 7994 6488
rect 7959 6395 7966 6415
rect 7986 6395 7994 6415
rect 9114 6440 9699 6448
rect 9114 6420 9123 6440
rect 9143 6439 9699 6440
rect 9143 6420 9663 6439
rect 9114 6419 9663 6420
rect 9683 6419 9699 6439
rect 9114 6413 9699 6419
rect 7959 6388 7994 6395
rect 9733 6392 9767 6598
rect 10460 6608 10501 6619
rect 10696 6616 10730 6822
rect 10460 6590 10470 6608
rect 10488 6590 10501 6608
rect 10460 6582 10501 6590
rect 10674 6611 10730 6616
rect 10674 6591 10681 6611
rect 10701 6591 10730 6611
rect 10674 6584 10730 6591
rect 10674 6583 10709 6584
rect 10469 6552 10495 6582
rect 10469 6551 10807 6552
rect 10469 6515 10823 6551
rect 6754 6229 7093 6257
rect 6848 6194 6883 6195
rect 6827 6187 6883 6194
rect 6827 6167 6856 6187
rect 6876 6167 6883 6187
rect 6827 6162 6883 6167
rect 7062 6187 7093 6229
rect 7062 6168 7067 6187
rect 7088 6168 7093 6187
rect 7062 6162 7093 6168
rect 7724 6182 7758 6388
rect 9497 6385 9532 6392
rect 7792 6361 8377 6367
rect 7792 6341 7808 6361
rect 7828 6360 8377 6361
rect 7828 6341 8348 6360
rect 7792 6340 8348 6341
rect 8368 6340 8377 6360
rect 7792 6332 8377 6340
rect 9497 6365 9505 6385
rect 9525 6365 9532 6385
rect 9497 6292 9532 6365
rect 9711 6387 9767 6392
rect 9711 6367 9718 6387
rect 9738 6367 9767 6387
rect 9711 6360 9767 6367
rect 9802 6494 9832 6496
rect 10531 6494 10564 6495
rect 9802 6468 10565 6494
rect 9711 6359 9746 6360
rect 9802 6293 9832 6468
rect 10531 6447 10565 6468
rect 10530 6442 10565 6447
rect 10530 6422 10537 6442
rect 10557 6422 10565 6442
rect 10530 6414 10565 6422
rect 9797 6292 9832 6293
rect 9496 6265 9832 6292
rect 9802 6264 9832 6265
rect 9912 6256 10497 6264
rect 9912 6236 9921 6256
rect 9941 6255 10497 6256
rect 9941 6236 10461 6255
rect 9912 6235 10461 6236
rect 10481 6235 10497 6255
rect 9912 6229 10497 6235
rect 9736 6219 9768 6220
rect 9733 6214 9768 6219
rect 9733 6194 9740 6214
rect 9760 6194 9768 6214
rect 10531 6208 10565 6414
rect 9733 6186 9768 6194
rect 7724 6174 7759 6182
rect 6827 5956 6861 6162
rect 7724 6154 7732 6174
rect 7752 6154 7759 6174
rect 7724 6149 7759 6154
rect 7724 6148 7756 6149
rect 6895 6135 7480 6141
rect 6895 6115 6911 6135
rect 6931 6134 7480 6135
rect 6931 6115 7451 6134
rect 6895 6114 7451 6115
rect 7471 6114 7480 6134
rect 6895 6106 7480 6114
rect 9115 6028 9700 6036
rect 9115 6008 9124 6028
rect 9144 6027 9700 6028
rect 9144 6008 9664 6027
rect 9115 6007 9664 6008
rect 9684 6007 9700 6027
rect 9115 6001 9700 6007
rect 9489 5977 9528 5981
rect 9734 5980 9768 6186
rect 10297 6201 10332 6207
rect 10297 6182 10302 6201
rect 10323 6182 10332 6201
rect 10297 6173 10332 6182
rect 10509 6203 10565 6208
rect 10509 6183 10516 6203
rect 10536 6183 10565 6203
rect 10509 6176 10565 6183
rect 10509 6175 10544 6176
rect 10301 6105 10330 6173
rect 10301 6071 10647 6105
rect 9489 5957 9497 5977
rect 9517 5957 9528 5977
rect 6827 5948 6862 5956
rect 6827 5928 6835 5948
rect 6855 5940 6862 5948
rect 6855 5928 6866 5940
rect 6827 5691 6866 5928
rect 7697 5905 7983 5906
rect 7182 5897 7985 5905
rect 7182 5880 7193 5897
rect 7183 5875 7193 5880
rect 7217 5880 7985 5897
rect 7217 5875 7222 5880
rect 7183 5862 7222 5875
rect 7727 5814 7762 5815
rect 7706 5807 7762 5814
rect 7706 5787 7735 5807
rect 7755 5787 7762 5807
rect 7706 5782 7762 5787
rect 7946 5805 7985 5880
rect 9489 5882 9528 5957
rect 9712 5975 9768 5980
rect 9712 5955 9719 5975
rect 9739 5955 9768 5975
rect 9712 5948 9768 5955
rect 9712 5947 9747 5948
rect 10252 5887 10291 5900
rect 10252 5882 10257 5887
rect 9489 5865 10257 5882
rect 10281 5882 10291 5887
rect 10281 5865 10292 5882
rect 9489 5857 10292 5865
rect 9491 5856 9777 5857
rect 10608 5834 10647 6071
rect 10608 5822 10619 5834
rect 10612 5814 10619 5822
rect 10639 5814 10647 5834
rect 10612 5806 10647 5814
rect 7946 5785 7957 5805
rect 7977 5785 7985 5805
rect 6827 5657 7173 5691
rect 7144 5589 7173 5657
rect 6930 5586 6965 5587
rect 6909 5579 6965 5586
rect 6909 5559 6938 5579
rect 6958 5559 6965 5579
rect 6909 5554 6965 5559
rect 7142 5580 7177 5589
rect 7142 5561 7151 5580
rect 7172 5561 7177 5580
rect 7142 5555 7177 5561
rect 7706 5576 7740 5782
rect 7946 5781 7985 5785
rect 7774 5755 8359 5761
rect 7774 5735 7790 5755
rect 7810 5754 8359 5755
rect 7810 5735 8330 5754
rect 7774 5734 8330 5735
rect 8350 5734 8359 5754
rect 7774 5726 8359 5734
rect 9994 5648 10579 5656
rect 9994 5628 10003 5648
rect 10023 5647 10579 5648
rect 10023 5628 10543 5647
rect 9994 5627 10543 5628
rect 10563 5627 10579 5647
rect 9994 5621 10579 5627
rect 9718 5613 9750 5614
rect 9715 5608 9750 5613
rect 9715 5588 9722 5608
rect 9742 5588 9750 5608
rect 10613 5600 10647 5806
rect 9715 5580 9750 5588
rect 7706 5568 7741 5576
rect 6909 5348 6943 5554
rect 7706 5548 7714 5568
rect 7734 5548 7741 5568
rect 7706 5543 7741 5548
rect 7706 5542 7738 5543
rect 6977 5527 7562 5533
rect 6977 5507 6993 5527
rect 7013 5526 7562 5527
rect 7013 5507 7533 5526
rect 6977 5506 7533 5507
rect 7553 5506 7562 5526
rect 6977 5498 7562 5506
rect 7642 5497 7672 5498
rect 7642 5470 7978 5497
rect 7642 5469 7677 5470
rect 6909 5340 6944 5348
rect 6909 5320 6917 5340
rect 6937 5320 6944 5340
rect 6909 5315 6944 5320
rect 6909 5294 6943 5315
rect 7642 5294 7672 5469
rect 7728 5402 7763 5403
rect 6909 5268 7672 5294
rect 6910 5267 6943 5268
rect 7642 5266 7672 5268
rect 7707 5395 7763 5402
rect 7707 5375 7736 5395
rect 7756 5375 7763 5395
rect 7707 5370 7763 5375
rect 7942 5397 7977 5470
rect 7942 5377 7949 5397
rect 7969 5377 7977 5397
rect 9097 5422 9682 5430
rect 9097 5402 9106 5422
rect 9126 5421 9682 5422
rect 9126 5402 9646 5421
rect 9097 5401 9646 5402
rect 9666 5401 9682 5421
rect 9097 5395 9682 5401
rect 7942 5370 7977 5377
rect 9716 5374 9750 5580
rect 10379 5588 10415 5597
rect 10379 5571 10388 5588
rect 10407 5571 10415 5588
rect 10379 5562 10415 5571
rect 10591 5595 10647 5600
rect 10591 5575 10598 5595
rect 10618 5575 10647 5595
rect 10591 5568 10647 5575
rect 10591 5567 10626 5568
rect 10385 5527 10411 5562
rect 10693 5527 10725 5528
rect 10385 5522 10725 5527
rect 10385 5504 10700 5522
rect 10722 5504 10725 5522
rect 10385 5499 10725 5504
rect 10693 5498 10725 5499
rect 6561 5247 6878 5250
rect 6561 5220 6564 5247
rect 6591 5220 6878 5247
rect 6561 5214 6878 5220
rect 6561 5211 6597 5214
rect 6842 5184 6878 5214
rect 6626 5180 6661 5181
rect 6605 5173 6661 5180
rect 6605 5153 6634 5173
rect 6654 5153 6661 5173
rect 6605 5148 6661 5153
rect 6840 5178 6878 5184
rect 6840 5152 6846 5178
rect 6872 5152 6878 5178
rect 6605 4949 6639 5148
rect 6840 5144 6878 5152
rect 7707 5164 7741 5370
rect 9480 5367 9515 5374
rect 7775 5343 8360 5349
rect 7775 5323 7791 5343
rect 7811 5342 8360 5343
rect 7811 5323 8331 5342
rect 7775 5322 8331 5323
rect 8351 5322 8360 5342
rect 7775 5314 8360 5322
rect 9480 5347 9488 5367
rect 9508 5347 9515 5367
rect 9480 5274 9515 5347
rect 9694 5369 9750 5374
rect 9694 5349 9701 5369
rect 9721 5349 9750 5369
rect 9694 5342 9750 5349
rect 9785 5476 9815 5478
rect 10514 5476 10547 5477
rect 9785 5450 10548 5476
rect 9694 5341 9729 5342
rect 9785 5275 9815 5450
rect 10514 5429 10548 5450
rect 10513 5424 10548 5429
rect 10513 5404 10520 5424
rect 10540 5404 10548 5424
rect 10513 5396 10548 5404
rect 9780 5274 9815 5275
rect 9479 5247 9815 5274
rect 9785 5246 9815 5247
rect 9895 5238 10480 5246
rect 9895 5218 9904 5238
rect 9924 5237 10480 5238
rect 9924 5218 10444 5237
rect 9895 5217 10444 5218
rect 10464 5217 10480 5237
rect 9895 5211 10480 5217
rect 9719 5201 9751 5202
rect 9716 5196 9751 5201
rect 9716 5176 9723 5196
rect 9743 5176 9751 5196
rect 10514 5190 10548 5396
rect 9716 5168 9751 5176
rect 7707 5156 7742 5164
rect 7707 5136 7715 5156
rect 7735 5136 7742 5156
rect 7707 5131 7742 5136
rect 7707 5130 7739 5131
rect 6673 5121 7258 5127
rect 6673 5101 6689 5121
rect 6709 5120 7258 5121
rect 6709 5101 7229 5120
rect 6673 5100 7229 5101
rect 7249 5100 7258 5120
rect 6673 5092 7258 5100
rect 9098 5010 9683 5018
rect 9098 4990 9107 5010
rect 9127 5009 9683 5010
rect 9127 4990 9647 5009
rect 9098 4989 9647 4990
rect 9667 4989 9683 5009
rect 9098 4983 9683 4989
rect 9472 4959 9511 4963
rect 9717 4962 9751 5168
rect 10281 5180 10315 5188
rect 10281 5162 10288 5180
rect 10307 5162 10315 5180
rect 10281 5155 10315 5162
rect 10492 5185 10548 5190
rect 10492 5165 10499 5185
rect 10519 5165 10548 5185
rect 10492 5158 10548 5165
rect 10492 5157 10527 5158
rect 10285 5125 10314 5155
rect 10285 5117 10667 5125
rect 10285 5098 10638 5117
rect 10659 5098 10667 5117
rect 10285 5093 10667 5098
rect 6605 4934 6642 4949
rect 6605 4914 6613 4934
rect 6633 4914 6642 4934
rect 6605 4911 6642 4914
rect 6419 4800 6456 4803
rect 6419 4780 6428 4800
rect 6448 4780 6456 4800
rect 6419 4765 6456 4780
rect 2407 4615 2789 4620
rect 2407 4596 2415 4615
rect 2436 4596 2789 4615
rect 2407 4588 2789 4596
rect 2760 4558 2789 4588
rect 2547 4555 2582 4556
rect 2526 4548 2582 4555
rect 2526 4528 2555 4548
rect 2575 4528 2582 4548
rect 2526 4523 2582 4528
rect 2759 4551 2793 4558
rect 2759 4533 2767 4551
rect 2786 4533 2793 4551
rect 2759 4525 2793 4533
rect 3323 4545 3357 4751
rect 3563 4750 3602 4754
rect 3391 4724 3976 4730
rect 3391 4704 3407 4724
rect 3427 4723 3976 4724
rect 3427 4704 3947 4723
rect 3391 4703 3947 4704
rect 3967 4703 3976 4723
rect 3391 4695 3976 4703
rect 5803 4614 6388 4622
rect 5803 4594 5812 4614
rect 5832 4613 6388 4614
rect 5832 4594 6352 4613
rect 5803 4593 6352 4594
rect 6372 4593 6388 4613
rect 5803 4587 6388 4593
rect 5322 4583 5354 4584
rect 5319 4578 5354 4583
rect 5319 4558 5326 4578
rect 5346 4558 5354 4578
rect 6422 4566 6456 4765
rect 6400 4561 6456 4566
rect 5319 4550 5354 4558
rect 3323 4537 3358 4545
rect 2526 4317 2560 4523
rect 3323 4517 3331 4537
rect 3351 4517 3358 4537
rect 3323 4512 3358 4517
rect 3323 4511 3355 4512
rect 2594 4496 3179 4502
rect 2594 4476 2610 4496
rect 2630 4495 3179 4496
rect 2630 4476 3150 4495
rect 2594 4475 3150 4476
rect 3170 4475 3179 4495
rect 2594 4467 3179 4475
rect 3259 4466 3289 4467
rect 3259 4439 3595 4466
rect 3259 4438 3294 4439
rect 2526 4309 2561 4317
rect 2526 4289 2534 4309
rect 2554 4289 2561 4309
rect 2526 4284 2561 4289
rect 2526 4263 2560 4284
rect 3259 4263 3289 4438
rect 3345 4371 3380 4372
rect 2526 4237 3289 4263
rect 2527 4236 2560 4237
rect 3259 4235 3289 4237
rect 3324 4364 3380 4371
rect 3324 4344 3353 4364
rect 3373 4344 3380 4364
rect 3324 4339 3380 4344
rect 3559 4366 3594 4439
rect 3559 4346 3566 4366
rect 3586 4346 3594 4366
rect 4701 4392 5286 4400
rect 4701 4372 4710 4392
rect 4730 4391 5286 4392
rect 4730 4372 5250 4391
rect 4701 4371 5250 4372
rect 5270 4371 5286 4391
rect 4701 4365 5286 4371
rect 3559 4339 3594 4346
rect 5320 4344 5354 4550
rect 6182 4559 6217 4561
rect 6182 4553 6220 4559
rect 6182 4530 6190 4553
rect 6213 4530 6220 4553
rect 6400 4541 6407 4561
rect 6427 4541 6456 4561
rect 6400 4534 6456 4541
rect 6400 4533 6435 4534
rect 6182 4524 6220 4530
rect 6182 4511 6217 4524
rect 6180 4453 6217 4511
rect 2349 4214 2381 4215
rect 2349 4209 2689 4214
rect 2349 4191 2352 4209
rect 2374 4191 2689 4209
rect 2349 4186 2689 4191
rect 2349 4185 2381 4186
rect 2663 4151 2689 4186
rect 2448 4145 2483 4146
rect 2427 4138 2483 4145
rect 2427 4118 2456 4138
rect 2476 4118 2483 4138
rect 2427 4113 2483 4118
rect 2659 4142 2695 4151
rect 2659 4125 2667 4142
rect 2686 4125 2695 4142
rect 2659 4116 2695 4125
rect 3324 4133 3358 4339
rect 5084 4337 5119 4344
rect 3392 4312 3977 4318
rect 3392 4292 3408 4312
rect 3428 4311 3977 4312
rect 3428 4292 3948 4311
rect 3392 4291 3948 4292
rect 3968 4291 3977 4311
rect 3392 4283 3977 4291
rect 5084 4317 5092 4337
rect 5112 4317 5119 4337
rect 5084 4244 5119 4317
rect 5298 4339 5354 4344
rect 5298 4319 5305 4339
rect 5325 4319 5354 4339
rect 5298 4312 5354 4319
rect 5389 4446 5419 4448
rect 6118 4446 6151 4447
rect 5389 4420 6152 4446
rect 5298 4311 5333 4312
rect 5389 4245 5419 4420
rect 6118 4399 6152 4420
rect 6180 4436 6215 4453
rect 6180 4435 6474 4436
rect 6180 4434 6517 4435
rect 6180 4427 6522 4434
rect 6180 4401 6482 4427
rect 6513 4401 6522 4427
rect 6117 4394 6152 4399
rect 6473 4398 6522 4401
rect 6117 4374 6124 4394
rect 6144 4374 6152 4394
rect 6479 4393 6522 4398
rect 6117 4366 6152 4374
rect 5384 4244 5419 4245
rect 5083 4217 5419 4244
rect 5389 4216 5419 4217
rect 5499 4208 6084 4216
rect 5499 4188 5508 4208
rect 5528 4207 6084 4208
rect 5528 4188 6048 4207
rect 5499 4187 6048 4188
rect 6068 4187 6084 4207
rect 5499 4181 6084 4187
rect 5323 4171 5355 4172
rect 5320 4166 5355 4171
rect 5320 4146 5327 4166
rect 5347 4146 5355 4166
rect 6118 4160 6152 4366
rect 5320 4138 5355 4146
rect 3324 4125 3359 4133
rect 2427 3907 2461 4113
rect 3324 4105 3332 4125
rect 3352 4105 3359 4125
rect 3324 4100 3359 4105
rect 3324 4099 3356 4100
rect 2495 4086 3080 4092
rect 2495 4066 2511 4086
rect 2531 4085 3080 4086
rect 2531 4066 3051 4085
rect 2495 4065 3051 4066
rect 3071 4065 3080 4085
rect 2495 4057 3080 4065
rect 4702 3980 5287 3988
rect 4702 3960 4711 3980
rect 4731 3979 5287 3980
rect 4731 3960 5251 3979
rect 4702 3959 5251 3960
rect 5271 3959 5287 3979
rect 4702 3953 5287 3959
rect 5076 3929 5115 3933
rect 5321 3932 5355 4138
rect 5884 4153 5919 4159
rect 5884 4134 5889 4153
rect 5910 4134 5919 4153
rect 5884 4125 5919 4134
rect 6096 4155 6152 4160
rect 6096 4135 6103 4155
rect 6123 4135 6152 4155
rect 6096 4128 6152 4135
rect 6096 4127 6131 4128
rect 5888 4057 5917 4125
rect 5888 4023 6234 4057
rect 5076 3909 5084 3929
rect 5104 3909 5115 3929
rect 2427 3899 2462 3907
rect 2427 3879 2435 3899
rect 2455 3891 2462 3899
rect 2455 3879 2466 3891
rect 2427 3642 2466 3879
rect 3297 3856 3583 3857
rect 2782 3848 3585 3856
rect 2782 3831 2793 3848
rect 2783 3826 2793 3831
rect 2817 3831 3585 3848
rect 2817 3826 2822 3831
rect 2783 3813 2822 3826
rect 3327 3765 3362 3766
rect 3306 3758 3362 3765
rect 3306 3738 3335 3758
rect 3355 3738 3362 3758
rect 3306 3733 3362 3738
rect 3546 3756 3585 3831
rect 5076 3834 5115 3909
rect 5299 3927 5355 3932
rect 5299 3907 5306 3927
rect 5326 3907 5355 3927
rect 5299 3900 5355 3907
rect 5299 3899 5334 3900
rect 5839 3839 5878 3852
rect 5839 3834 5844 3839
rect 5076 3817 5844 3834
rect 5868 3834 5878 3839
rect 5868 3817 5879 3834
rect 5076 3809 5879 3817
rect 5078 3808 5364 3809
rect 6195 3786 6234 4023
rect 6195 3774 6206 3786
rect 6199 3766 6206 3774
rect 6226 3766 6234 3786
rect 6199 3758 6234 3766
rect 3546 3736 3557 3756
rect 3577 3736 3585 3756
rect 2427 3608 2773 3642
rect 2744 3540 2773 3608
rect 2530 3537 2565 3538
rect 2509 3530 2565 3537
rect 2509 3510 2538 3530
rect 2558 3510 2565 3530
rect 2509 3505 2565 3510
rect 2742 3531 2777 3540
rect 2742 3512 2751 3531
rect 2772 3512 2777 3531
rect 2742 3506 2777 3512
rect 3306 3527 3340 3733
rect 3546 3732 3585 3736
rect 3374 3706 3959 3712
rect 3374 3686 3390 3706
rect 3410 3705 3959 3706
rect 3410 3686 3930 3705
rect 3374 3685 3930 3686
rect 3950 3685 3959 3705
rect 3374 3677 3959 3685
rect 5581 3600 6166 3608
rect 5581 3580 5590 3600
rect 5610 3599 6166 3600
rect 5610 3580 6130 3599
rect 5581 3579 6130 3580
rect 6150 3579 6166 3599
rect 5581 3573 6166 3579
rect 5305 3565 5337 3566
rect 5302 3560 5337 3565
rect 5302 3540 5309 3560
rect 5329 3540 5337 3560
rect 6200 3552 6234 3758
rect 5302 3532 5337 3540
rect 3306 3519 3341 3527
rect 2509 3299 2543 3505
rect 3306 3499 3314 3519
rect 3334 3499 3341 3519
rect 3306 3494 3341 3499
rect 3306 3493 3338 3494
rect 2577 3478 3162 3484
rect 2577 3458 2593 3478
rect 2613 3477 3162 3478
rect 2613 3458 3133 3477
rect 2577 3457 3133 3458
rect 3153 3457 3162 3477
rect 2577 3449 3162 3457
rect 3242 3448 3272 3449
rect 3242 3421 3578 3448
rect 3242 3420 3277 3421
rect 2509 3291 2544 3299
rect 2509 3271 2517 3291
rect 2537 3271 2544 3291
rect 2509 3266 2544 3271
rect 2509 3245 2543 3266
rect 3242 3245 3272 3420
rect 3328 3353 3363 3354
rect 2509 3219 3272 3245
rect 2510 3218 2543 3219
rect 3242 3217 3272 3219
rect 3307 3346 3363 3353
rect 3307 3326 3336 3346
rect 3356 3326 3363 3346
rect 3307 3321 3363 3326
rect 3542 3348 3577 3421
rect 3542 3328 3549 3348
rect 3569 3328 3577 3348
rect 4684 3374 5269 3382
rect 4684 3354 4693 3374
rect 4713 3373 5269 3374
rect 4713 3354 5233 3373
rect 4684 3353 5233 3354
rect 5253 3353 5269 3373
rect 4684 3347 5269 3353
rect 3542 3321 3577 3328
rect 5303 3326 5337 3532
rect 5968 3546 5999 3552
rect 5968 3527 5973 3546
rect 5994 3527 5999 3546
rect 5968 3485 5999 3527
rect 6178 3547 6234 3552
rect 6178 3527 6185 3547
rect 6205 3527 6234 3547
rect 6178 3520 6234 3527
rect 6178 3519 6213 3520
rect 5968 3457 6307 3485
rect 2251 3162 2605 3198
rect 2267 3161 2605 3162
rect 2579 3131 2605 3161
rect 2365 3129 2400 3130
rect 2344 3122 2400 3129
rect 2344 3102 2373 3122
rect 2393 3102 2400 3122
rect 2344 3097 2400 3102
rect 2573 3123 2614 3131
rect 2573 3105 2586 3123
rect 2604 3105 2614 3123
rect 2344 2891 2378 3097
rect 2573 3094 2614 3105
rect 3307 3115 3341 3321
rect 5067 3319 5102 3326
rect 3375 3294 3960 3300
rect 3375 3274 3391 3294
rect 3411 3293 3960 3294
rect 3411 3274 3931 3293
rect 3375 3273 3931 3274
rect 3951 3273 3960 3293
rect 3375 3265 3960 3273
rect 5067 3299 5075 3319
rect 5095 3299 5102 3319
rect 5067 3226 5102 3299
rect 5281 3321 5337 3326
rect 5281 3301 5288 3321
rect 5308 3301 5337 3321
rect 5281 3294 5337 3301
rect 5372 3428 5402 3430
rect 6101 3428 6134 3429
rect 5372 3402 6135 3428
rect 5281 3293 5316 3294
rect 5372 3227 5402 3402
rect 6101 3381 6135 3402
rect 6100 3376 6135 3381
rect 6100 3356 6107 3376
rect 6127 3356 6135 3376
rect 6100 3348 6135 3356
rect 5367 3226 5402 3227
rect 5066 3199 5402 3226
rect 5372 3198 5402 3199
rect 5482 3190 6067 3198
rect 5482 3170 5491 3190
rect 5511 3189 6067 3190
rect 5511 3170 6031 3189
rect 5482 3169 6031 3170
rect 6051 3169 6067 3189
rect 5482 3163 6067 3169
rect 5306 3153 5338 3154
rect 5303 3148 5338 3153
rect 5303 3128 5310 3148
rect 5330 3128 5338 3148
rect 6101 3142 6135 3348
rect 5303 3120 5338 3128
rect 3307 3107 3342 3115
rect 3307 3087 3315 3107
rect 3335 3087 3342 3107
rect 3307 3082 3342 3087
rect 3307 3081 3339 3082
rect 2412 3070 2997 3076
rect 2412 3050 2428 3070
rect 2448 3069 2997 3070
rect 2448 3050 2968 3069
rect 2412 3049 2968 3050
rect 2988 3049 2997 3069
rect 2412 3041 2997 3049
rect 4685 2962 5270 2970
rect 4685 2942 4694 2962
rect 4714 2961 5270 2962
rect 4714 2942 5234 2961
rect 4685 2941 5234 2942
rect 5254 2941 5270 2961
rect 4685 2935 5270 2941
rect 5059 2911 5098 2915
rect 5304 2914 5338 3120
rect 5868 3132 5902 3140
rect 5868 3114 5875 3132
rect 5894 3114 5902 3132
rect 5868 3107 5902 3114
rect 6079 3137 6135 3142
rect 6079 3117 6086 3137
rect 6106 3117 6135 3137
rect 6079 3110 6135 3117
rect 6079 3109 6114 3110
rect 5872 3077 5901 3107
rect 5872 3069 6254 3077
rect 5872 3050 6225 3069
rect 6246 3050 6254 3069
rect 5872 3045 6254 3050
rect 5059 2891 5067 2911
rect 5087 2891 5098 2911
rect 2344 2890 2379 2891
rect 2312 2883 2379 2890
rect 2312 2863 2352 2883
rect 2372 2863 2379 2883
rect 2312 2860 2379 2863
rect 2312 2857 2377 2860
rect 1883 2756 1948 2759
rect 1881 2753 1948 2756
rect 1881 2733 1888 2753
rect 1908 2733 1948 2753
rect 1881 2726 1948 2733
rect 1881 2725 1916 2726
rect 1263 2567 1848 2575
rect 1263 2547 1272 2567
rect 1292 2566 1848 2567
rect 1292 2547 1812 2566
rect 1263 2546 1812 2547
rect 1832 2546 1848 2566
rect 1263 2540 1848 2546
rect 921 2534 953 2535
rect 918 2529 953 2534
rect 918 2509 925 2529
rect 945 2509 953 2529
rect 918 2501 953 2509
rect 300 2343 885 2351
rect 300 2323 309 2343
rect 329 2342 885 2343
rect 329 2323 849 2342
rect 300 2322 849 2323
rect 869 2322 885 2342
rect 300 2316 885 2322
rect 919 2295 953 2501
rect 1648 2516 1681 2522
rect 1882 2519 1916 2725
rect 1648 2494 1653 2516
rect 1676 2494 1681 2516
rect 1648 2485 1681 2494
rect 1860 2514 1916 2519
rect 1860 2494 1867 2514
rect 1887 2494 1916 2514
rect 1860 2487 1916 2494
rect 1860 2486 1895 2487
rect 1650 2454 1677 2485
rect 2072 2454 2111 2466
rect 1650 2453 2113 2454
rect 1650 2431 2077 2453
rect 2101 2431 2113 2453
rect 1650 2423 2113 2431
rect 683 2288 718 2295
rect 683 2268 691 2288
rect 711 2268 718 2288
rect 683 2195 718 2268
rect 897 2290 953 2295
rect 897 2270 904 2290
rect 924 2270 953 2290
rect 897 2263 953 2270
rect 988 2397 1018 2399
rect 1717 2397 1750 2398
rect 988 2371 1751 2397
rect 897 2262 932 2263
rect 988 2196 1018 2371
rect 1717 2350 1751 2371
rect 1716 2345 1751 2350
rect 1716 2325 1723 2345
rect 1743 2325 1751 2345
rect 1716 2317 1751 2325
rect 983 2195 1018 2196
rect 682 2168 1018 2195
rect 988 2167 1018 2168
rect 1098 2159 1683 2167
rect 1098 2139 1107 2159
rect 1127 2158 1683 2159
rect 1127 2139 1647 2158
rect 1098 2138 1647 2139
rect 1667 2138 1683 2158
rect 1098 2132 1683 2138
rect 922 2122 954 2123
rect 919 2117 954 2122
rect 919 2097 926 2117
rect 946 2097 954 2117
rect 1717 2111 1751 2317
rect 919 2089 954 2097
rect 301 1931 886 1939
rect 301 1911 310 1931
rect 330 1930 886 1931
rect 330 1911 850 1930
rect 301 1910 850 1911
rect 870 1910 886 1930
rect 301 1904 886 1910
rect 675 1880 714 1884
rect 920 1883 954 2089
rect 1483 2104 1518 2110
rect 1483 2085 1488 2104
rect 1509 2085 1518 2104
rect 1483 2076 1518 2085
rect 1695 2106 1751 2111
rect 1695 2086 1702 2106
rect 1722 2086 1751 2106
rect 1695 2079 1751 2086
rect 1873 2257 1905 2269
rect 1873 2239 1880 2257
rect 1902 2239 1905 2257
rect 1695 2078 1730 2079
rect 1487 2008 1516 2076
rect 1487 1974 1833 2008
rect 675 1860 683 1880
rect 703 1860 714 1880
rect 675 1785 714 1860
rect 898 1878 954 1883
rect 898 1858 905 1878
rect 925 1858 954 1878
rect 898 1851 954 1858
rect 898 1850 933 1851
rect 1438 1790 1477 1803
rect 1438 1785 1443 1790
rect 675 1768 1443 1785
rect 1467 1785 1477 1790
rect 1467 1768 1478 1785
rect 675 1760 1478 1768
rect 677 1759 963 1760
rect 1794 1737 1833 1974
rect 1794 1725 1805 1737
rect 1798 1717 1805 1725
rect 1825 1717 1833 1737
rect 1798 1709 1833 1717
rect 1180 1551 1765 1559
rect 1180 1531 1189 1551
rect 1209 1550 1765 1551
rect 1209 1531 1729 1550
rect 1180 1530 1729 1531
rect 1749 1530 1765 1550
rect 1180 1524 1765 1530
rect 904 1516 936 1517
rect 901 1511 936 1516
rect 901 1491 908 1511
rect 928 1491 936 1511
rect 1799 1503 1833 1709
rect 901 1483 936 1491
rect 283 1325 868 1333
rect 283 1305 292 1325
rect 312 1324 868 1325
rect 312 1305 832 1324
rect 283 1304 832 1305
rect 852 1304 868 1324
rect 283 1298 868 1304
rect 902 1277 936 1483
rect 1565 1491 1601 1500
rect 1565 1474 1574 1491
rect 1593 1474 1601 1491
rect 1565 1465 1601 1474
rect 1777 1498 1833 1503
rect 1777 1478 1784 1498
rect 1804 1478 1833 1498
rect 1777 1471 1833 1478
rect 1777 1470 1812 1471
rect 1571 1430 1597 1465
rect 1873 1430 1905 2239
rect 2317 2172 2346 2857
rect 3277 2838 3563 2839
rect 2762 2830 3565 2838
rect 2762 2813 2773 2830
rect 2763 2808 2773 2813
rect 2797 2813 3565 2830
rect 2797 2808 2802 2813
rect 2763 2795 2802 2808
rect 3307 2747 3342 2748
rect 3286 2740 3342 2747
rect 3286 2720 3315 2740
rect 3335 2720 3342 2740
rect 3286 2715 3342 2720
rect 3526 2738 3565 2813
rect 5059 2816 5098 2891
rect 5282 2909 5338 2914
rect 5282 2889 5289 2909
rect 5309 2889 5338 2909
rect 5282 2882 5338 2889
rect 5282 2881 5317 2882
rect 5822 2821 5861 2834
rect 5822 2816 5827 2821
rect 5059 2799 5827 2816
rect 5851 2816 5861 2821
rect 5851 2799 5862 2816
rect 5059 2791 5862 2799
rect 5061 2790 5347 2791
rect 6278 2772 6307 3457
rect 6615 3211 6642 4911
rect 9472 4939 9480 4959
rect 9500 4939 9511 4959
rect 7678 4887 7964 4888
rect 7163 4879 7966 4887
rect 7163 4862 7174 4879
rect 7164 4857 7174 4862
rect 7198 4862 7966 4879
rect 7198 4857 7203 4862
rect 7164 4844 7203 4857
rect 7708 4796 7743 4797
rect 7687 4789 7743 4796
rect 7687 4769 7716 4789
rect 7736 4769 7743 4789
rect 7687 4764 7743 4769
rect 7927 4787 7966 4862
rect 9472 4864 9511 4939
rect 9695 4957 9751 4962
rect 9695 4937 9702 4957
rect 9722 4937 9751 4957
rect 9695 4930 9751 4937
rect 9695 4929 9730 4930
rect 10235 4869 10274 4882
rect 10235 4864 10240 4869
rect 9472 4847 10240 4864
rect 10264 4864 10274 4869
rect 10264 4847 10275 4864
rect 9472 4839 10275 4847
rect 9474 4838 9760 4839
rect 7927 4767 7938 4787
rect 7958 4767 7966 4787
rect 10796 4815 10823 6515
rect 11131 6269 11160 6954
rect 12091 6935 12377 6936
rect 11576 6927 12379 6935
rect 11576 6910 11587 6927
rect 11577 6905 11587 6910
rect 11611 6910 12379 6927
rect 11611 6905 11616 6910
rect 11577 6892 11616 6905
rect 12121 6844 12156 6845
rect 12100 6837 12156 6844
rect 12100 6817 12129 6837
rect 12149 6817 12156 6837
rect 12100 6812 12156 6817
rect 12340 6835 12379 6910
rect 13873 6913 13912 6988
rect 14096 7006 14152 7011
rect 14096 6986 14103 7006
rect 14123 6986 14152 7006
rect 14096 6979 14152 6986
rect 14096 6978 14131 6979
rect 14636 6918 14675 6931
rect 14636 6913 14641 6918
rect 13873 6896 14641 6913
rect 14665 6913 14675 6918
rect 14665 6896 14676 6913
rect 13873 6888 14676 6896
rect 13875 6887 14161 6888
rect 15092 6869 15121 7554
rect 15533 7487 15565 8296
rect 15841 8261 15867 8296
rect 15626 8255 15661 8256
rect 15605 8248 15661 8255
rect 15605 8228 15634 8248
rect 15654 8228 15661 8248
rect 15605 8223 15661 8228
rect 15837 8252 15873 8261
rect 15837 8235 15845 8252
rect 15864 8235 15873 8252
rect 15837 8226 15873 8235
rect 16502 8243 16536 8449
rect 17781 8443 17790 8463
rect 17810 8462 18366 8463
rect 17810 8443 18330 8462
rect 17781 8442 18330 8443
rect 18350 8442 18366 8462
rect 17781 8436 18366 8442
rect 16570 8422 17155 8428
rect 16570 8402 16586 8422
rect 16606 8421 17155 8422
rect 16606 8402 17126 8421
rect 16570 8401 17126 8402
rect 17146 8401 17155 8421
rect 18400 8415 18434 8621
rect 19970 8632 20026 8639
rect 19970 8612 19999 8632
rect 20019 8612 20026 8632
rect 19970 8607 20026 8612
rect 20203 8635 20237 8642
rect 20203 8617 20211 8635
rect 20230 8617 20237 8635
rect 20203 8609 20237 8617
rect 20767 8629 20801 8835
rect 21007 8834 21046 8838
rect 25131 8873 25187 8880
rect 25131 8853 25160 8873
rect 25180 8853 25187 8873
rect 25131 8848 25187 8853
rect 25371 8871 25410 8946
rect 28985 8953 28995 8958
rect 29019 8958 29787 8975
rect 33348 8971 33359 8988
rect 29019 8953 29024 8958
rect 28985 8940 29024 8953
rect 29529 8892 29564 8893
rect 25371 8851 25382 8871
rect 25402 8851 25410 8871
rect 20835 8808 21420 8814
rect 20835 8788 20851 8808
rect 20871 8807 21420 8808
rect 20871 8788 21391 8807
rect 20835 8787 21391 8788
rect 21411 8787 21420 8807
rect 20835 8779 21420 8787
rect 24215 8712 24597 8717
rect 24215 8693 24223 8712
rect 24244 8693 24597 8712
rect 24215 8685 24597 8693
rect 22766 8667 22798 8668
rect 22763 8662 22798 8667
rect 22763 8642 22770 8662
rect 22790 8642 22798 8662
rect 24568 8655 24597 8685
rect 24355 8652 24390 8653
rect 22763 8634 22798 8642
rect 20767 8621 20802 8629
rect 16570 8393 17155 8401
rect 18164 8408 18199 8415
rect 18164 8388 18172 8408
rect 18192 8388 18199 8408
rect 18164 8315 18199 8388
rect 18378 8410 18434 8415
rect 18378 8390 18385 8410
rect 18405 8390 18434 8410
rect 18378 8383 18434 8390
rect 18469 8517 18499 8519
rect 19198 8517 19231 8518
rect 18469 8491 19232 8517
rect 18378 8382 18413 8383
rect 18469 8316 18499 8491
rect 19198 8470 19232 8491
rect 19197 8465 19232 8470
rect 19197 8445 19204 8465
rect 19224 8445 19232 8465
rect 19197 8437 19232 8445
rect 18464 8315 18499 8316
rect 18163 8288 18499 8315
rect 18469 8287 18499 8288
rect 18579 8279 19164 8287
rect 18579 8259 18588 8279
rect 18608 8278 19164 8279
rect 18608 8259 19128 8278
rect 18579 8258 19128 8259
rect 19148 8258 19164 8278
rect 18579 8252 19164 8258
rect 16502 8235 16537 8243
rect 18403 8242 18435 8243
rect 15605 8017 15639 8223
rect 16502 8215 16510 8235
rect 16530 8215 16537 8235
rect 16502 8210 16537 8215
rect 18400 8237 18435 8242
rect 18400 8217 18407 8237
rect 18427 8217 18435 8237
rect 19198 8231 19232 8437
rect 19970 8401 20004 8607
rect 20767 8601 20775 8621
rect 20795 8601 20802 8621
rect 20767 8596 20802 8601
rect 20767 8595 20799 8596
rect 20038 8580 20623 8586
rect 20038 8560 20054 8580
rect 20074 8579 20623 8580
rect 20074 8560 20594 8579
rect 20038 8559 20594 8560
rect 20614 8559 20623 8579
rect 20038 8551 20623 8559
rect 20703 8550 20733 8551
rect 20703 8523 21039 8550
rect 20703 8522 20738 8523
rect 19970 8393 20005 8401
rect 19970 8373 19978 8393
rect 19998 8373 20005 8393
rect 19970 8368 20005 8373
rect 19970 8347 20004 8368
rect 20703 8347 20733 8522
rect 20789 8455 20824 8456
rect 19970 8321 20733 8347
rect 19971 8320 20004 8321
rect 20703 8319 20733 8321
rect 20768 8448 20824 8455
rect 20768 8428 20797 8448
rect 20817 8428 20824 8448
rect 20768 8423 20824 8428
rect 21003 8450 21038 8523
rect 21003 8430 21010 8450
rect 21030 8430 21038 8450
rect 22145 8476 22730 8484
rect 22145 8456 22154 8476
rect 22174 8475 22730 8476
rect 22174 8456 22694 8475
rect 22145 8455 22694 8456
rect 22714 8455 22730 8475
rect 22145 8449 22730 8455
rect 21003 8423 21038 8430
rect 22764 8428 22798 8634
rect 24334 8645 24390 8652
rect 24334 8625 24363 8645
rect 24383 8625 24390 8645
rect 24334 8620 24390 8625
rect 24567 8648 24601 8655
rect 24567 8630 24575 8648
rect 24594 8630 24601 8648
rect 24567 8622 24601 8630
rect 25131 8642 25165 8848
rect 25371 8847 25410 8851
rect 29508 8885 29564 8892
rect 29508 8865 29537 8885
rect 29557 8865 29564 8885
rect 29508 8860 29564 8865
rect 29748 8883 29787 8958
rect 33349 8966 33359 8971
rect 33383 8971 34151 8988
rect 33383 8966 33388 8971
rect 33349 8953 33388 8966
rect 33893 8905 33928 8906
rect 29748 8863 29759 8883
rect 29779 8863 29787 8883
rect 25199 8821 25784 8827
rect 25199 8801 25215 8821
rect 25235 8820 25784 8821
rect 25235 8801 25755 8820
rect 25199 8800 25755 8801
rect 25775 8800 25784 8820
rect 25199 8792 25784 8800
rect 28592 8724 28974 8729
rect 28592 8705 28600 8724
rect 28621 8705 28974 8724
rect 28592 8697 28974 8705
rect 27143 8679 27175 8680
rect 27140 8674 27175 8679
rect 27140 8654 27147 8674
rect 27167 8654 27175 8674
rect 28945 8667 28974 8697
rect 28732 8664 28767 8665
rect 27140 8646 27175 8654
rect 25131 8634 25166 8642
rect 16502 8209 16534 8210
rect 18400 8209 18435 8217
rect 15673 8196 16258 8202
rect 15673 8176 15689 8196
rect 15709 8195 16258 8196
rect 15709 8176 16229 8195
rect 15673 8175 16229 8176
rect 16249 8175 16258 8195
rect 15673 8167 16258 8175
rect 17782 8051 18367 8059
rect 17782 8031 17791 8051
rect 17811 8050 18367 8051
rect 17811 8031 18331 8050
rect 17782 8030 18331 8031
rect 18351 8030 18367 8050
rect 17782 8024 18367 8030
rect 15605 8009 15640 8017
rect 15605 7989 15613 8009
rect 15633 8001 15640 8009
rect 15633 7989 15644 8001
rect 15605 7752 15644 7989
rect 18156 8000 18195 8004
rect 18401 8003 18435 8209
rect 18964 8224 18999 8230
rect 18964 8205 18969 8224
rect 18990 8205 18999 8224
rect 18964 8196 18999 8205
rect 19176 8226 19232 8231
rect 19176 8206 19183 8226
rect 19203 8206 19232 8226
rect 19176 8199 19232 8206
rect 19799 8270 20133 8298
rect 19176 8198 19211 8199
rect 18968 8128 18997 8196
rect 18968 8094 19314 8128
rect 18156 7980 18164 8000
rect 18184 7980 18195 8000
rect 16475 7966 16761 7967
rect 15960 7958 16763 7966
rect 15960 7941 15971 7958
rect 15961 7936 15971 7941
rect 15995 7941 16763 7958
rect 15995 7936 16000 7941
rect 15961 7923 16000 7936
rect 16505 7875 16540 7876
rect 16484 7868 16540 7875
rect 16484 7848 16513 7868
rect 16533 7848 16540 7868
rect 16484 7843 16540 7848
rect 16724 7866 16763 7941
rect 18156 7905 18195 7980
rect 18379 7998 18435 8003
rect 18379 7978 18386 7998
rect 18406 7978 18435 7998
rect 18379 7971 18435 7978
rect 18379 7970 18414 7971
rect 18919 7910 18958 7923
rect 18919 7905 18924 7910
rect 18156 7888 18924 7905
rect 18948 7905 18958 7910
rect 18948 7888 18959 7905
rect 18156 7880 18959 7888
rect 18158 7879 18444 7880
rect 16724 7846 16735 7866
rect 16755 7846 16763 7866
rect 15605 7718 15951 7752
rect 15922 7650 15951 7718
rect 15708 7647 15743 7648
rect 15533 7469 15536 7487
rect 15558 7469 15565 7487
rect 15533 7457 15565 7469
rect 15687 7640 15743 7647
rect 15687 7620 15716 7640
rect 15736 7620 15743 7640
rect 15687 7615 15743 7620
rect 15920 7641 15955 7650
rect 15920 7622 15929 7641
rect 15950 7622 15955 7641
rect 15920 7616 15955 7622
rect 16484 7637 16518 7843
rect 16724 7842 16763 7846
rect 19275 7857 19314 8094
rect 19275 7845 19286 7857
rect 19279 7837 19286 7845
rect 19306 7837 19314 7857
rect 19279 7829 19314 7837
rect 16552 7816 17137 7822
rect 16552 7796 16568 7816
rect 16588 7815 17137 7816
rect 16588 7796 17108 7815
rect 16552 7795 17108 7796
rect 17128 7795 17137 7815
rect 16552 7787 17137 7795
rect 18661 7671 19246 7679
rect 18661 7651 18670 7671
rect 18690 7670 19246 7671
rect 18690 7651 19210 7670
rect 18661 7650 19210 7651
rect 19230 7650 19246 7670
rect 18661 7644 19246 7650
rect 16484 7629 16519 7637
rect 18385 7636 18417 7637
rect 15687 7409 15721 7615
rect 16484 7609 16492 7629
rect 16512 7609 16519 7629
rect 16484 7604 16519 7609
rect 18382 7631 18417 7636
rect 18382 7611 18389 7631
rect 18409 7611 18417 7631
rect 19280 7623 19314 7829
rect 16484 7603 16516 7604
rect 18382 7603 18417 7611
rect 15755 7588 16340 7594
rect 15755 7568 15771 7588
rect 15791 7587 16340 7588
rect 15791 7568 16311 7587
rect 15755 7567 16311 7568
rect 16331 7567 16340 7587
rect 15755 7559 16340 7567
rect 16420 7558 16450 7559
rect 16420 7531 16756 7558
rect 16420 7530 16455 7531
rect 15687 7401 15722 7409
rect 15687 7381 15695 7401
rect 15715 7381 15722 7401
rect 15687 7376 15722 7381
rect 15687 7355 15721 7376
rect 16420 7355 16450 7530
rect 16506 7463 16541 7464
rect 15687 7329 16450 7355
rect 15688 7328 15721 7329
rect 16420 7327 16450 7329
rect 16485 7456 16541 7463
rect 16485 7436 16514 7456
rect 16534 7436 16541 7456
rect 16485 7431 16541 7436
rect 16720 7458 16755 7531
rect 16720 7438 16727 7458
rect 16747 7438 16755 7458
rect 16720 7431 16755 7438
rect 17764 7445 18349 7453
rect 15325 7295 15788 7303
rect 15325 7273 15337 7295
rect 15361 7273 15788 7295
rect 15325 7272 15788 7273
rect 15327 7260 15366 7272
rect 15761 7241 15788 7272
rect 15543 7239 15578 7240
rect 15522 7232 15578 7239
rect 15522 7212 15551 7232
rect 15571 7212 15578 7232
rect 15522 7207 15578 7212
rect 15757 7232 15790 7241
rect 15757 7210 15762 7232
rect 15785 7210 15790 7232
rect 15522 7001 15556 7207
rect 15757 7204 15790 7210
rect 16485 7225 16519 7431
rect 17764 7425 17773 7445
rect 17793 7444 18349 7445
rect 17793 7425 18313 7444
rect 17764 7424 18313 7425
rect 18333 7424 18349 7444
rect 17764 7418 18349 7424
rect 16553 7404 17138 7410
rect 16553 7384 16569 7404
rect 16589 7403 17138 7404
rect 16589 7384 17109 7403
rect 16553 7383 17109 7384
rect 17129 7383 17138 7403
rect 18383 7397 18417 7603
rect 19048 7617 19079 7623
rect 19048 7598 19053 7617
rect 19074 7598 19079 7617
rect 19048 7556 19079 7598
rect 19258 7618 19314 7623
rect 19258 7598 19265 7618
rect 19285 7598 19314 7618
rect 19258 7591 19314 7598
rect 19258 7590 19293 7591
rect 19048 7528 19387 7556
rect 16553 7375 17138 7383
rect 18147 7390 18182 7397
rect 18147 7370 18155 7390
rect 18175 7370 18182 7390
rect 18147 7297 18182 7370
rect 18361 7392 18417 7397
rect 18361 7372 18368 7392
rect 18388 7372 18417 7392
rect 18361 7365 18417 7372
rect 18452 7499 18482 7501
rect 19181 7499 19214 7500
rect 18452 7473 19215 7499
rect 18361 7364 18396 7365
rect 18452 7298 18482 7473
rect 19181 7452 19215 7473
rect 19180 7447 19215 7452
rect 19180 7427 19187 7447
rect 19207 7427 19215 7447
rect 19180 7419 19215 7427
rect 18447 7297 18482 7298
rect 18146 7270 18482 7297
rect 18452 7269 18482 7270
rect 18562 7261 19147 7269
rect 18562 7241 18571 7261
rect 18591 7260 19147 7261
rect 18591 7241 19111 7260
rect 18562 7240 19111 7241
rect 19131 7240 19147 7260
rect 18562 7234 19147 7240
rect 16485 7217 16520 7225
rect 18386 7224 18418 7225
rect 16485 7197 16493 7217
rect 16513 7197 16520 7217
rect 16485 7192 16520 7197
rect 18383 7219 18418 7224
rect 18383 7199 18390 7219
rect 18410 7199 18418 7219
rect 19181 7213 19215 7419
rect 16485 7191 16517 7192
rect 18383 7191 18418 7199
rect 15590 7180 16175 7186
rect 15590 7160 15606 7180
rect 15626 7179 16175 7180
rect 15626 7160 16146 7179
rect 15590 7159 16146 7160
rect 16166 7159 16175 7179
rect 15590 7151 16175 7159
rect 17765 7033 18350 7041
rect 17765 7013 17774 7033
rect 17794 7032 18350 7033
rect 17794 7013 18314 7032
rect 17765 7012 18314 7013
rect 18334 7012 18350 7032
rect 17765 7006 18350 7012
rect 15522 7000 15557 7001
rect 15490 6993 15557 7000
rect 15490 6973 15530 6993
rect 15550 6973 15557 6993
rect 15490 6970 15557 6973
rect 18139 6982 18178 6986
rect 18384 6985 18418 7191
rect 18948 7203 18982 7211
rect 18948 7185 18955 7203
rect 18974 7185 18982 7203
rect 18948 7178 18982 7185
rect 19159 7208 19215 7213
rect 19159 7188 19166 7208
rect 19186 7188 19215 7208
rect 19159 7181 19215 7188
rect 19159 7180 19194 7181
rect 18952 7148 18981 7178
rect 18952 7140 19334 7148
rect 18952 7121 19305 7140
rect 19326 7121 19334 7140
rect 18952 7116 19334 7121
rect 15490 6967 15555 6970
rect 15061 6866 15126 6869
rect 15059 6863 15126 6866
rect 15059 6843 15066 6863
rect 15086 6843 15126 6863
rect 15059 6836 15126 6843
rect 15059 6835 15094 6836
rect 12340 6815 12351 6835
rect 12371 6815 12379 6835
rect 11184 6676 11566 6681
rect 11184 6657 11192 6676
rect 11213 6657 11566 6676
rect 11184 6649 11566 6657
rect 11537 6619 11566 6649
rect 11324 6616 11359 6617
rect 11303 6609 11359 6616
rect 11303 6589 11332 6609
rect 11352 6589 11359 6609
rect 11303 6584 11359 6589
rect 11536 6612 11570 6619
rect 11536 6594 11544 6612
rect 11563 6594 11570 6612
rect 11536 6586 11570 6594
rect 12100 6606 12134 6812
rect 12340 6811 12379 6815
rect 12168 6785 12753 6791
rect 12168 6765 12184 6785
rect 12204 6784 12753 6785
rect 12204 6765 12724 6784
rect 12168 6764 12724 6765
rect 12744 6764 12753 6784
rect 12168 6756 12753 6764
rect 14441 6677 15026 6685
rect 14441 6657 14450 6677
rect 14470 6676 15026 6677
rect 14470 6657 14990 6676
rect 14441 6656 14990 6657
rect 15010 6656 15026 6676
rect 14441 6650 15026 6656
rect 14099 6644 14131 6645
rect 14096 6639 14131 6644
rect 14096 6619 14103 6639
rect 14123 6619 14131 6639
rect 14096 6611 14131 6619
rect 12100 6598 12135 6606
rect 11303 6378 11337 6584
rect 12100 6578 12108 6598
rect 12128 6578 12135 6598
rect 12100 6573 12135 6578
rect 12100 6572 12132 6573
rect 11371 6557 11956 6563
rect 11371 6537 11387 6557
rect 11407 6556 11956 6557
rect 11407 6537 11927 6556
rect 11371 6536 11927 6537
rect 11947 6536 11956 6556
rect 11371 6528 11956 6536
rect 12036 6527 12066 6528
rect 12036 6500 12372 6527
rect 12036 6499 12071 6500
rect 11303 6370 11338 6378
rect 11303 6350 11311 6370
rect 11331 6350 11338 6370
rect 11303 6345 11338 6350
rect 11303 6324 11337 6345
rect 12036 6324 12066 6499
rect 12122 6432 12157 6433
rect 11303 6298 12066 6324
rect 11304 6297 11337 6298
rect 12036 6296 12066 6298
rect 12101 6425 12157 6432
rect 12101 6405 12130 6425
rect 12150 6405 12157 6425
rect 12101 6400 12157 6405
rect 12336 6427 12371 6500
rect 12336 6407 12343 6427
rect 12363 6407 12371 6427
rect 13478 6453 14063 6461
rect 13478 6433 13487 6453
rect 13507 6452 14063 6453
rect 13507 6433 14027 6452
rect 13478 6432 14027 6433
rect 14047 6432 14063 6452
rect 13478 6426 14063 6432
rect 12336 6400 12371 6407
rect 14097 6405 14131 6611
rect 14824 6621 14865 6632
rect 15060 6629 15094 6835
rect 14824 6603 14834 6621
rect 14852 6603 14865 6621
rect 14824 6595 14865 6603
rect 15038 6624 15094 6629
rect 15038 6604 15045 6624
rect 15065 6604 15094 6624
rect 15038 6597 15094 6604
rect 15038 6596 15073 6597
rect 14833 6565 14859 6595
rect 14833 6564 15171 6565
rect 14833 6528 15187 6564
rect 11131 6241 11470 6269
rect 11225 6206 11260 6207
rect 11204 6199 11260 6206
rect 11204 6179 11233 6199
rect 11253 6179 11260 6199
rect 11204 6174 11260 6179
rect 11439 6199 11470 6241
rect 11439 6180 11444 6199
rect 11465 6180 11470 6199
rect 11439 6174 11470 6180
rect 12101 6194 12135 6400
rect 13861 6398 13896 6405
rect 12169 6373 12754 6379
rect 12169 6353 12185 6373
rect 12205 6372 12754 6373
rect 12205 6353 12725 6372
rect 12169 6352 12725 6353
rect 12745 6352 12754 6372
rect 12169 6344 12754 6352
rect 13861 6378 13869 6398
rect 13889 6378 13896 6398
rect 13861 6305 13896 6378
rect 14075 6400 14131 6405
rect 14075 6380 14082 6400
rect 14102 6380 14131 6400
rect 14075 6373 14131 6380
rect 14166 6507 14196 6509
rect 14895 6507 14928 6508
rect 14166 6481 14929 6507
rect 14075 6372 14110 6373
rect 14166 6306 14196 6481
rect 14895 6460 14929 6481
rect 14894 6455 14929 6460
rect 14894 6435 14901 6455
rect 14921 6435 14929 6455
rect 14894 6427 14929 6435
rect 14161 6305 14196 6306
rect 13860 6278 14196 6305
rect 14166 6277 14196 6278
rect 14276 6269 14861 6277
rect 14276 6249 14285 6269
rect 14305 6268 14861 6269
rect 14305 6249 14825 6268
rect 14276 6248 14825 6249
rect 14845 6248 14861 6268
rect 14276 6242 14861 6248
rect 14100 6232 14132 6233
rect 14097 6227 14132 6232
rect 14097 6207 14104 6227
rect 14124 6207 14132 6227
rect 14895 6221 14929 6427
rect 14097 6199 14132 6207
rect 12101 6186 12136 6194
rect 11204 5968 11238 6174
rect 12101 6166 12109 6186
rect 12129 6166 12136 6186
rect 12101 6161 12136 6166
rect 12101 6160 12133 6161
rect 11272 6147 11857 6153
rect 11272 6127 11288 6147
rect 11308 6146 11857 6147
rect 11308 6127 11828 6146
rect 11272 6126 11828 6127
rect 11848 6126 11857 6146
rect 11272 6118 11857 6126
rect 13479 6041 14064 6049
rect 13479 6021 13488 6041
rect 13508 6040 14064 6041
rect 13508 6021 14028 6040
rect 13479 6020 14028 6021
rect 14048 6020 14064 6040
rect 13479 6014 14064 6020
rect 13853 5990 13892 5994
rect 14098 5993 14132 6199
rect 14661 6214 14696 6220
rect 14661 6195 14666 6214
rect 14687 6195 14696 6214
rect 14661 6186 14696 6195
rect 14873 6216 14929 6221
rect 14873 6196 14880 6216
rect 14900 6196 14929 6216
rect 14873 6189 14929 6196
rect 14873 6188 14908 6189
rect 14665 6118 14694 6186
rect 14665 6084 15011 6118
rect 13853 5970 13861 5990
rect 13881 5970 13892 5990
rect 11204 5960 11239 5968
rect 11204 5940 11212 5960
rect 11232 5952 11239 5960
rect 11232 5940 11243 5952
rect 11204 5703 11243 5940
rect 12074 5917 12360 5918
rect 11559 5909 12362 5917
rect 11559 5892 11570 5909
rect 11560 5887 11570 5892
rect 11594 5892 12362 5909
rect 11594 5887 11599 5892
rect 11560 5874 11599 5887
rect 12104 5826 12139 5827
rect 12083 5819 12139 5826
rect 12083 5799 12112 5819
rect 12132 5799 12139 5819
rect 12083 5794 12139 5799
rect 12323 5817 12362 5892
rect 13853 5895 13892 5970
rect 14076 5988 14132 5993
rect 14076 5968 14083 5988
rect 14103 5968 14132 5988
rect 14076 5961 14132 5968
rect 14076 5960 14111 5961
rect 14616 5900 14655 5913
rect 14616 5895 14621 5900
rect 13853 5878 14621 5895
rect 14645 5895 14655 5900
rect 14645 5878 14656 5895
rect 13853 5870 14656 5878
rect 13855 5869 14141 5870
rect 14972 5847 15011 6084
rect 14972 5835 14983 5847
rect 14976 5827 14983 5835
rect 15003 5827 15011 5847
rect 14976 5819 15011 5827
rect 12323 5797 12334 5817
rect 12354 5797 12362 5817
rect 11204 5669 11550 5703
rect 11521 5601 11550 5669
rect 11307 5598 11342 5599
rect 11286 5591 11342 5598
rect 11286 5571 11315 5591
rect 11335 5571 11342 5591
rect 11286 5566 11342 5571
rect 11519 5592 11554 5601
rect 11519 5573 11528 5592
rect 11549 5573 11554 5592
rect 11519 5567 11554 5573
rect 12083 5588 12117 5794
rect 12323 5793 12362 5797
rect 12151 5767 12736 5773
rect 12151 5747 12167 5767
rect 12187 5766 12736 5767
rect 12187 5747 12707 5766
rect 12151 5746 12707 5747
rect 12727 5746 12736 5766
rect 12151 5738 12736 5746
rect 14358 5661 14943 5669
rect 14358 5641 14367 5661
rect 14387 5660 14943 5661
rect 14387 5641 14907 5660
rect 14358 5640 14907 5641
rect 14927 5640 14943 5660
rect 14358 5634 14943 5640
rect 14082 5626 14114 5627
rect 14079 5621 14114 5626
rect 14079 5601 14086 5621
rect 14106 5601 14114 5621
rect 14977 5613 15011 5819
rect 14079 5593 14114 5601
rect 12083 5580 12118 5588
rect 11286 5360 11320 5566
rect 12083 5560 12091 5580
rect 12111 5560 12118 5580
rect 12083 5555 12118 5560
rect 12083 5554 12115 5555
rect 11354 5539 11939 5545
rect 11354 5519 11370 5539
rect 11390 5538 11939 5539
rect 11390 5519 11910 5538
rect 11354 5518 11910 5519
rect 11930 5518 11939 5538
rect 11354 5510 11939 5518
rect 12019 5509 12049 5510
rect 12019 5482 12355 5509
rect 12019 5481 12054 5482
rect 11286 5352 11321 5360
rect 11286 5332 11294 5352
rect 11314 5332 11321 5352
rect 11286 5327 11321 5332
rect 11286 5306 11320 5327
rect 12019 5306 12049 5481
rect 12105 5414 12140 5415
rect 11286 5280 12049 5306
rect 11287 5279 11320 5280
rect 12019 5278 12049 5280
rect 12084 5407 12140 5414
rect 12084 5387 12113 5407
rect 12133 5387 12140 5407
rect 12084 5382 12140 5387
rect 12319 5409 12354 5482
rect 12319 5389 12326 5409
rect 12346 5389 12354 5409
rect 13461 5435 14046 5443
rect 13461 5415 13470 5435
rect 13490 5434 14046 5435
rect 13490 5415 14010 5434
rect 13461 5414 14010 5415
rect 14030 5414 14046 5434
rect 13461 5408 14046 5414
rect 12319 5382 12354 5389
rect 14080 5387 14114 5593
rect 14743 5601 14779 5610
rect 14743 5584 14752 5601
rect 14771 5584 14779 5601
rect 14743 5575 14779 5584
rect 14955 5608 15011 5613
rect 14955 5588 14962 5608
rect 14982 5588 15011 5608
rect 14955 5581 15011 5588
rect 14955 5580 14990 5581
rect 14749 5540 14775 5575
rect 15057 5540 15089 5541
rect 14749 5535 15089 5540
rect 14749 5517 15064 5535
rect 15086 5517 15089 5535
rect 14749 5512 15089 5517
rect 15057 5511 15089 5512
rect 10938 5259 11255 5262
rect 10938 5232 10941 5259
rect 10968 5232 11255 5259
rect 10938 5226 11255 5232
rect 10938 5223 10974 5226
rect 11219 5196 11255 5226
rect 11003 5192 11038 5193
rect 10982 5185 11038 5192
rect 10982 5165 11011 5185
rect 11031 5165 11038 5185
rect 10982 5160 11038 5165
rect 11217 5190 11255 5196
rect 11217 5164 11223 5190
rect 11249 5164 11255 5190
rect 10982 4961 11016 5160
rect 11217 5156 11255 5164
rect 12084 5176 12118 5382
rect 13844 5380 13879 5387
rect 12152 5355 12737 5361
rect 12152 5335 12168 5355
rect 12188 5354 12737 5355
rect 12188 5335 12708 5354
rect 12152 5334 12708 5335
rect 12728 5334 12737 5354
rect 12152 5326 12737 5334
rect 13844 5360 13852 5380
rect 13872 5360 13879 5380
rect 13844 5287 13879 5360
rect 14058 5382 14114 5387
rect 14058 5362 14065 5382
rect 14085 5362 14114 5382
rect 14058 5355 14114 5362
rect 14149 5489 14179 5491
rect 14878 5489 14911 5490
rect 14149 5463 14912 5489
rect 14058 5354 14093 5355
rect 14149 5288 14179 5463
rect 14878 5442 14912 5463
rect 14877 5437 14912 5442
rect 14877 5417 14884 5437
rect 14904 5417 14912 5437
rect 14877 5409 14912 5417
rect 14144 5287 14179 5288
rect 13843 5260 14179 5287
rect 14149 5259 14179 5260
rect 14259 5251 14844 5259
rect 14259 5231 14268 5251
rect 14288 5250 14844 5251
rect 14288 5231 14808 5250
rect 14259 5230 14808 5231
rect 14828 5230 14844 5250
rect 14259 5224 14844 5230
rect 14083 5214 14115 5215
rect 14080 5209 14115 5214
rect 14080 5189 14087 5209
rect 14107 5189 14115 5209
rect 14878 5203 14912 5409
rect 14080 5181 14115 5189
rect 12084 5168 12119 5176
rect 12084 5148 12092 5168
rect 12112 5148 12119 5168
rect 12084 5143 12119 5148
rect 12084 5142 12116 5143
rect 11050 5133 11635 5139
rect 11050 5113 11066 5133
rect 11086 5132 11635 5133
rect 11086 5113 11606 5132
rect 11050 5112 11606 5113
rect 11626 5112 11635 5132
rect 11050 5104 11635 5112
rect 13462 5023 14047 5031
rect 13462 5003 13471 5023
rect 13491 5022 14047 5023
rect 13491 5003 14011 5022
rect 13462 5002 14011 5003
rect 14031 5002 14047 5022
rect 13462 4996 14047 5002
rect 13836 4972 13875 4976
rect 14081 4975 14115 5181
rect 14645 5193 14679 5201
rect 14645 5175 14652 5193
rect 14671 5175 14679 5193
rect 14645 5168 14679 5175
rect 14856 5198 14912 5203
rect 14856 5178 14863 5198
rect 14883 5178 14912 5198
rect 14856 5171 14912 5178
rect 14856 5170 14891 5171
rect 14649 5138 14678 5168
rect 14649 5130 15031 5138
rect 14649 5111 15002 5130
rect 15023 5111 15031 5130
rect 14649 5106 15031 5111
rect 10982 4946 11019 4961
rect 10982 4926 10990 4946
rect 11010 4926 11019 4946
rect 10982 4923 11019 4926
rect 10796 4812 10833 4815
rect 10796 4792 10805 4812
rect 10825 4792 10833 4812
rect 10796 4777 10833 4792
rect 6771 4628 7153 4633
rect 6771 4609 6779 4628
rect 6800 4609 7153 4628
rect 6771 4601 7153 4609
rect 7124 4571 7153 4601
rect 6911 4568 6946 4569
rect 6890 4561 6946 4568
rect 6890 4541 6919 4561
rect 6939 4541 6946 4561
rect 6890 4536 6946 4541
rect 7123 4564 7157 4571
rect 7123 4546 7131 4564
rect 7150 4546 7157 4564
rect 7123 4538 7157 4546
rect 7687 4558 7721 4764
rect 7927 4763 7966 4767
rect 7755 4737 8340 4743
rect 7755 4717 7771 4737
rect 7791 4736 8340 4737
rect 7791 4717 8311 4736
rect 7755 4716 8311 4717
rect 8331 4716 8340 4736
rect 7755 4708 8340 4716
rect 10180 4626 10765 4634
rect 10180 4606 10189 4626
rect 10209 4625 10765 4626
rect 10209 4606 10729 4625
rect 10180 4605 10729 4606
rect 10749 4605 10765 4625
rect 10180 4599 10765 4605
rect 9699 4595 9731 4596
rect 9696 4590 9731 4595
rect 9696 4570 9703 4590
rect 9723 4570 9731 4590
rect 10799 4578 10833 4777
rect 10777 4573 10833 4578
rect 9696 4562 9731 4570
rect 7687 4550 7722 4558
rect 6890 4330 6924 4536
rect 7687 4530 7695 4550
rect 7715 4530 7722 4550
rect 7687 4525 7722 4530
rect 7687 4524 7719 4525
rect 6958 4509 7543 4515
rect 6958 4489 6974 4509
rect 6994 4508 7543 4509
rect 6994 4489 7514 4508
rect 6958 4488 7514 4489
rect 7534 4488 7543 4508
rect 6958 4480 7543 4488
rect 7623 4479 7653 4480
rect 7623 4452 7959 4479
rect 7623 4451 7658 4452
rect 6890 4322 6925 4330
rect 6890 4302 6898 4322
rect 6918 4302 6925 4322
rect 6890 4297 6925 4302
rect 6890 4276 6924 4297
rect 7623 4276 7653 4451
rect 7709 4384 7744 4385
rect 6890 4250 7653 4276
rect 6891 4249 6924 4250
rect 7623 4248 7653 4250
rect 7688 4377 7744 4384
rect 7688 4357 7717 4377
rect 7737 4357 7744 4377
rect 7688 4352 7744 4357
rect 7923 4379 7958 4452
rect 7923 4359 7930 4379
rect 7950 4359 7958 4379
rect 9078 4404 9663 4412
rect 9078 4384 9087 4404
rect 9107 4403 9663 4404
rect 9107 4384 9627 4403
rect 9078 4383 9627 4384
rect 9647 4383 9663 4403
rect 9078 4377 9663 4383
rect 7923 4352 7958 4359
rect 9697 4356 9731 4562
rect 10559 4571 10594 4573
rect 10559 4565 10597 4571
rect 10559 4542 10567 4565
rect 10590 4542 10597 4565
rect 10777 4553 10784 4573
rect 10804 4553 10833 4573
rect 10777 4546 10833 4553
rect 10777 4545 10812 4546
rect 10559 4536 10597 4542
rect 10559 4523 10594 4536
rect 10557 4465 10594 4523
rect 6713 4227 6745 4228
rect 6713 4222 7053 4227
rect 6713 4204 6716 4222
rect 6738 4204 7053 4222
rect 6713 4199 7053 4204
rect 6713 4198 6745 4199
rect 7027 4164 7053 4199
rect 6812 4158 6847 4159
rect 6791 4151 6847 4158
rect 6791 4131 6820 4151
rect 6840 4131 6847 4151
rect 6791 4126 6847 4131
rect 7023 4155 7059 4164
rect 7023 4138 7031 4155
rect 7050 4138 7059 4155
rect 7023 4129 7059 4138
rect 7688 4146 7722 4352
rect 9461 4349 9496 4356
rect 7756 4325 8341 4331
rect 7756 4305 7772 4325
rect 7792 4324 8341 4325
rect 7792 4305 8312 4324
rect 7756 4304 8312 4305
rect 8332 4304 8341 4324
rect 7756 4296 8341 4304
rect 9461 4329 9469 4349
rect 9489 4329 9496 4349
rect 9461 4256 9496 4329
rect 9675 4351 9731 4356
rect 9675 4331 9682 4351
rect 9702 4331 9731 4351
rect 9675 4324 9731 4331
rect 9766 4458 9796 4460
rect 10495 4458 10528 4459
rect 9766 4432 10529 4458
rect 9675 4323 9710 4324
rect 9766 4257 9796 4432
rect 10495 4411 10529 4432
rect 10557 4448 10592 4465
rect 10557 4447 10851 4448
rect 10557 4446 10894 4447
rect 10557 4439 10899 4446
rect 10557 4413 10859 4439
rect 10890 4413 10899 4439
rect 10494 4406 10529 4411
rect 10850 4410 10899 4413
rect 10494 4386 10501 4406
rect 10521 4386 10529 4406
rect 10856 4405 10899 4410
rect 10494 4378 10529 4386
rect 9761 4256 9796 4257
rect 9460 4229 9796 4256
rect 9766 4228 9796 4229
rect 9876 4220 10461 4228
rect 9876 4200 9885 4220
rect 9905 4219 10461 4220
rect 9905 4200 10425 4219
rect 9876 4199 10425 4200
rect 10445 4199 10461 4219
rect 9876 4193 10461 4199
rect 9700 4183 9732 4184
rect 9697 4178 9732 4183
rect 9697 4158 9704 4178
rect 9724 4158 9732 4178
rect 10495 4172 10529 4378
rect 9697 4150 9732 4158
rect 7688 4138 7723 4146
rect 6791 3920 6825 4126
rect 7688 4118 7696 4138
rect 7716 4118 7723 4138
rect 7688 4113 7723 4118
rect 7688 4112 7720 4113
rect 6859 4099 7444 4105
rect 6859 4079 6875 4099
rect 6895 4098 7444 4099
rect 6895 4079 7415 4098
rect 6859 4078 7415 4079
rect 7435 4078 7444 4098
rect 6859 4070 7444 4078
rect 9079 3992 9664 4000
rect 9079 3972 9088 3992
rect 9108 3991 9664 3992
rect 9108 3972 9628 3991
rect 9079 3971 9628 3972
rect 9648 3971 9664 3991
rect 9079 3965 9664 3971
rect 9453 3941 9492 3945
rect 9698 3944 9732 4150
rect 10261 4165 10296 4171
rect 10261 4146 10266 4165
rect 10287 4146 10296 4165
rect 10261 4137 10296 4146
rect 10473 4167 10529 4172
rect 10473 4147 10480 4167
rect 10500 4147 10529 4167
rect 10473 4140 10529 4147
rect 10473 4139 10508 4140
rect 10265 4069 10294 4137
rect 10265 4035 10611 4069
rect 9453 3921 9461 3941
rect 9481 3921 9492 3941
rect 6791 3912 6826 3920
rect 6791 3892 6799 3912
rect 6819 3904 6826 3912
rect 6819 3892 6830 3904
rect 6791 3655 6830 3892
rect 7661 3869 7947 3870
rect 7146 3861 7949 3869
rect 7146 3844 7157 3861
rect 7147 3839 7157 3844
rect 7181 3844 7949 3861
rect 7181 3839 7186 3844
rect 7147 3826 7186 3839
rect 7691 3778 7726 3779
rect 7670 3771 7726 3778
rect 7670 3751 7699 3771
rect 7719 3751 7726 3771
rect 7670 3746 7726 3751
rect 7910 3769 7949 3844
rect 9453 3846 9492 3921
rect 9676 3939 9732 3944
rect 9676 3919 9683 3939
rect 9703 3919 9732 3939
rect 9676 3912 9732 3919
rect 9676 3911 9711 3912
rect 10216 3851 10255 3864
rect 10216 3846 10221 3851
rect 9453 3829 10221 3846
rect 10245 3846 10255 3851
rect 10245 3829 10256 3846
rect 9453 3821 10256 3829
rect 9455 3820 9741 3821
rect 10572 3798 10611 4035
rect 10572 3786 10583 3798
rect 10576 3778 10583 3786
rect 10603 3778 10611 3798
rect 10576 3770 10611 3778
rect 7910 3749 7921 3769
rect 7941 3749 7949 3769
rect 6791 3621 7137 3655
rect 7108 3553 7137 3621
rect 6894 3550 6929 3551
rect 6873 3543 6929 3550
rect 6873 3523 6902 3543
rect 6922 3523 6929 3543
rect 6873 3518 6929 3523
rect 7106 3544 7141 3553
rect 7106 3525 7115 3544
rect 7136 3525 7141 3544
rect 7106 3519 7141 3525
rect 7670 3540 7704 3746
rect 7910 3745 7949 3749
rect 7738 3719 8323 3725
rect 7738 3699 7754 3719
rect 7774 3718 8323 3719
rect 7774 3699 8294 3718
rect 7738 3698 8294 3699
rect 8314 3698 8323 3718
rect 7738 3690 8323 3698
rect 9958 3612 10543 3620
rect 9958 3592 9967 3612
rect 9987 3611 10543 3612
rect 9987 3592 10507 3611
rect 9958 3591 10507 3592
rect 10527 3591 10543 3611
rect 9958 3585 10543 3591
rect 9682 3577 9714 3578
rect 9679 3572 9714 3577
rect 9679 3552 9686 3572
rect 9706 3552 9714 3572
rect 10577 3564 10611 3770
rect 9679 3544 9714 3552
rect 7670 3532 7705 3540
rect 6873 3312 6907 3518
rect 7670 3512 7678 3532
rect 7698 3512 7705 3532
rect 7670 3507 7705 3512
rect 7670 3506 7702 3507
rect 6941 3491 7526 3497
rect 6941 3471 6957 3491
rect 6977 3490 7526 3491
rect 6977 3471 7497 3490
rect 6941 3470 7497 3471
rect 7517 3470 7526 3490
rect 6941 3462 7526 3470
rect 7606 3461 7636 3462
rect 7606 3434 7942 3461
rect 7606 3433 7641 3434
rect 6873 3304 6908 3312
rect 6873 3284 6881 3304
rect 6901 3284 6908 3304
rect 6873 3279 6908 3284
rect 6873 3258 6907 3279
rect 7606 3258 7636 3433
rect 7692 3366 7727 3367
rect 6873 3232 7636 3258
rect 6874 3231 6907 3232
rect 7606 3230 7636 3232
rect 7671 3359 7727 3366
rect 7671 3339 7700 3359
rect 7720 3339 7727 3359
rect 7671 3334 7727 3339
rect 7906 3361 7941 3434
rect 7906 3341 7913 3361
rect 7933 3341 7941 3361
rect 9061 3386 9646 3394
rect 9061 3366 9070 3386
rect 9090 3385 9646 3386
rect 9090 3366 9610 3385
rect 9061 3365 9610 3366
rect 9630 3365 9646 3385
rect 9061 3359 9646 3365
rect 7906 3334 7941 3341
rect 9680 3338 9714 3544
rect 10345 3558 10376 3564
rect 10345 3539 10350 3558
rect 10371 3539 10376 3558
rect 10345 3497 10376 3539
rect 10555 3559 10611 3564
rect 10555 3539 10562 3559
rect 10582 3539 10611 3559
rect 10555 3532 10611 3539
rect 10555 3531 10590 3532
rect 10345 3469 10684 3497
rect 6615 3175 6969 3211
rect 6631 3174 6969 3175
rect 6943 3144 6969 3174
rect 6729 3142 6764 3143
rect 6708 3135 6764 3142
rect 6708 3115 6737 3135
rect 6757 3115 6764 3135
rect 6708 3110 6764 3115
rect 6937 3136 6978 3144
rect 6937 3118 6950 3136
rect 6968 3118 6978 3136
rect 6708 2904 6742 3110
rect 6937 3107 6978 3118
rect 7671 3128 7705 3334
rect 9444 3331 9479 3338
rect 7739 3307 8324 3313
rect 7739 3287 7755 3307
rect 7775 3306 8324 3307
rect 7775 3287 8295 3306
rect 7739 3286 8295 3287
rect 8315 3286 8324 3306
rect 7739 3278 8324 3286
rect 9444 3311 9452 3331
rect 9472 3311 9479 3331
rect 9444 3238 9479 3311
rect 9658 3333 9714 3338
rect 9658 3313 9665 3333
rect 9685 3313 9714 3333
rect 9658 3306 9714 3313
rect 9749 3440 9779 3442
rect 10478 3440 10511 3441
rect 9749 3414 10512 3440
rect 9658 3305 9693 3306
rect 9749 3239 9779 3414
rect 10478 3393 10512 3414
rect 10477 3388 10512 3393
rect 10477 3368 10484 3388
rect 10504 3368 10512 3388
rect 10477 3360 10512 3368
rect 9744 3238 9779 3239
rect 9443 3211 9779 3238
rect 9749 3210 9779 3211
rect 9859 3202 10444 3210
rect 9859 3182 9868 3202
rect 9888 3201 10444 3202
rect 9888 3182 10408 3201
rect 9859 3181 10408 3182
rect 10428 3181 10444 3201
rect 9859 3175 10444 3181
rect 9683 3165 9715 3166
rect 9680 3160 9715 3165
rect 9680 3140 9687 3160
rect 9707 3140 9715 3160
rect 10478 3154 10512 3360
rect 9680 3132 9715 3140
rect 7671 3120 7706 3128
rect 7671 3100 7679 3120
rect 7699 3100 7706 3120
rect 7671 3095 7706 3100
rect 7671 3094 7703 3095
rect 6776 3083 7361 3089
rect 6776 3063 6792 3083
rect 6812 3082 7361 3083
rect 6812 3063 7332 3082
rect 6776 3062 7332 3063
rect 7352 3062 7361 3082
rect 6776 3054 7361 3062
rect 9062 2974 9647 2982
rect 9062 2954 9071 2974
rect 9091 2973 9647 2974
rect 9091 2954 9611 2973
rect 9062 2953 9611 2954
rect 9631 2953 9647 2973
rect 9062 2947 9647 2953
rect 9436 2923 9475 2927
rect 9681 2926 9715 3132
rect 10245 3144 10279 3152
rect 10245 3126 10252 3144
rect 10271 3126 10279 3144
rect 10245 3119 10279 3126
rect 10456 3149 10512 3154
rect 10456 3129 10463 3149
rect 10483 3129 10512 3149
rect 10456 3122 10512 3129
rect 10456 3121 10491 3122
rect 10249 3089 10278 3119
rect 10249 3081 10631 3089
rect 10249 3062 10602 3081
rect 10623 3062 10631 3081
rect 10249 3057 10631 3062
rect 6708 2903 6743 2904
rect 6676 2896 6743 2903
rect 6676 2876 6716 2896
rect 6736 2876 6743 2896
rect 6676 2873 6743 2876
rect 9436 2903 9444 2923
rect 9464 2903 9475 2923
rect 6676 2870 6741 2873
rect 6247 2769 6312 2772
rect 6245 2766 6312 2769
rect 6245 2746 6252 2766
rect 6272 2746 6312 2766
rect 6245 2739 6312 2746
rect 6245 2738 6280 2739
rect 3526 2718 3537 2738
rect 3557 2718 3565 2738
rect 2370 2579 2752 2584
rect 2370 2560 2378 2579
rect 2399 2560 2752 2579
rect 2370 2552 2752 2560
rect 2723 2522 2752 2552
rect 2510 2519 2545 2520
rect 2489 2512 2545 2519
rect 2489 2492 2518 2512
rect 2538 2492 2545 2512
rect 2489 2487 2545 2492
rect 2722 2515 2756 2522
rect 2722 2497 2730 2515
rect 2749 2497 2756 2515
rect 2722 2489 2756 2497
rect 3286 2509 3320 2715
rect 3526 2714 3565 2718
rect 3354 2688 3939 2694
rect 3354 2668 3370 2688
rect 3390 2687 3939 2688
rect 3390 2668 3910 2687
rect 3354 2667 3910 2668
rect 3930 2667 3939 2687
rect 3354 2659 3939 2667
rect 5627 2580 6212 2588
rect 5627 2560 5636 2580
rect 5656 2579 6212 2580
rect 5656 2560 6176 2579
rect 5627 2559 6176 2560
rect 6196 2559 6212 2579
rect 5627 2553 6212 2559
rect 5285 2547 5317 2548
rect 5282 2542 5317 2547
rect 5282 2522 5289 2542
rect 5309 2522 5317 2542
rect 5282 2514 5317 2522
rect 3286 2501 3321 2509
rect 2489 2281 2523 2487
rect 3286 2481 3294 2501
rect 3314 2481 3321 2501
rect 3286 2476 3321 2481
rect 3286 2475 3318 2476
rect 2557 2460 3142 2466
rect 2557 2440 2573 2460
rect 2593 2459 3142 2460
rect 2593 2440 3113 2459
rect 2557 2439 3113 2440
rect 3133 2439 3142 2459
rect 2557 2431 3142 2439
rect 3222 2430 3252 2431
rect 3222 2403 3558 2430
rect 3222 2402 3257 2403
rect 2489 2273 2524 2281
rect 2489 2253 2497 2273
rect 2517 2253 2524 2273
rect 2489 2248 2524 2253
rect 2489 2227 2523 2248
rect 3222 2227 3252 2402
rect 3308 2335 3343 2336
rect 2489 2201 3252 2227
rect 2490 2200 2523 2201
rect 3222 2199 3252 2201
rect 3287 2328 3343 2335
rect 3287 2308 3316 2328
rect 3336 2308 3343 2328
rect 3287 2303 3343 2308
rect 3522 2330 3557 2403
rect 3522 2310 3529 2330
rect 3549 2310 3557 2330
rect 4664 2356 5249 2364
rect 4664 2336 4673 2356
rect 4693 2355 5249 2356
rect 4693 2336 5213 2355
rect 4664 2335 5213 2336
rect 5233 2335 5249 2355
rect 4664 2329 5249 2335
rect 3522 2303 3557 2310
rect 5283 2308 5317 2514
rect 6012 2529 6045 2535
rect 6246 2532 6280 2738
rect 6012 2507 6017 2529
rect 6040 2507 6045 2529
rect 6012 2498 6045 2507
rect 6224 2527 6280 2532
rect 6224 2507 6231 2527
rect 6251 2507 6280 2527
rect 6224 2500 6280 2507
rect 6224 2499 6259 2500
rect 6014 2467 6041 2498
rect 6436 2467 6475 2479
rect 6014 2466 6477 2467
rect 6014 2444 6441 2466
rect 6465 2444 6477 2466
rect 6014 2436 6477 2444
rect 2317 2144 2656 2172
rect 2411 2109 2446 2110
rect 2390 2102 2446 2109
rect 2390 2082 2419 2102
rect 2439 2082 2446 2102
rect 2390 2077 2446 2082
rect 2625 2102 2656 2144
rect 2625 2083 2630 2102
rect 2651 2083 2656 2102
rect 2625 2077 2656 2083
rect 3287 2097 3321 2303
rect 5047 2301 5082 2308
rect 3355 2276 3940 2282
rect 3355 2256 3371 2276
rect 3391 2275 3940 2276
rect 3391 2256 3911 2275
rect 3355 2255 3911 2256
rect 3931 2255 3940 2275
rect 3355 2247 3940 2255
rect 5047 2281 5055 2301
rect 5075 2281 5082 2301
rect 5047 2208 5082 2281
rect 5261 2303 5317 2308
rect 5261 2283 5268 2303
rect 5288 2283 5317 2303
rect 5261 2276 5317 2283
rect 5352 2410 5382 2412
rect 6081 2410 6114 2411
rect 5352 2384 6115 2410
rect 5261 2275 5296 2276
rect 5352 2209 5382 2384
rect 6081 2363 6115 2384
rect 6080 2358 6115 2363
rect 6080 2338 6087 2358
rect 6107 2338 6115 2358
rect 6080 2330 6115 2338
rect 5347 2208 5382 2209
rect 5046 2181 5382 2208
rect 5352 2180 5382 2181
rect 5462 2172 6047 2180
rect 5462 2152 5471 2172
rect 5491 2171 6047 2172
rect 5491 2152 6011 2171
rect 5462 2151 6011 2152
rect 6031 2151 6047 2171
rect 5462 2145 6047 2151
rect 5286 2135 5318 2136
rect 5283 2130 5318 2135
rect 5283 2110 5290 2130
rect 5310 2110 5318 2130
rect 6081 2124 6115 2330
rect 5283 2102 5318 2110
rect 3287 2089 3322 2097
rect 2390 1871 2424 2077
rect 3287 2069 3295 2089
rect 3315 2069 3322 2089
rect 3287 2064 3322 2069
rect 3287 2063 3319 2064
rect 2458 2050 3043 2056
rect 2458 2030 2474 2050
rect 2494 2049 3043 2050
rect 2494 2030 3014 2049
rect 2458 2029 3014 2030
rect 3034 2029 3043 2049
rect 2458 2021 3043 2029
rect 4665 1944 5250 1952
rect 4665 1924 4674 1944
rect 4694 1943 5250 1944
rect 4694 1924 5214 1943
rect 4665 1923 5214 1924
rect 5234 1923 5250 1943
rect 4665 1917 5250 1923
rect 5039 1893 5078 1897
rect 5284 1896 5318 2102
rect 5847 2117 5882 2123
rect 5847 2098 5852 2117
rect 5873 2098 5882 2117
rect 5847 2089 5882 2098
rect 6059 2119 6115 2124
rect 6059 2099 6066 2119
rect 6086 2099 6115 2119
rect 6059 2092 6115 2099
rect 6237 2270 6269 2282
rect 6237 2252 6244 2270
rect 6266 2252 6269 2270
rect 6059 2091 6094 2092
rect 5851 2021 5880 2089
rect 5851 1987 6197 2021
rect 5039 1873 5047 1893
rect 5067 1873 5078 1893
rect 2390 1863 2425 1871
rect 2390 1843 2398 1863
rect 2418 1855 2425 1863
rect 2418 1843 2429 1855
rect 2390 1606 2429 1843
rect 3260 1820 3546 1821
rect 2745 1812 3548 1820
rect 2745 1795 2756 1812
rect 2746 1790 2756 1795
rect 2780 1795 3548 1812
rect 2780 1790 2785 1795
rect 2746 1777 2785 1790
rect 3290 1729 3325 1730
rect 3269 1722 3325 1729
rect 3269 1702 3298 1722
rect 3318 1702 3325 1722
rect 3269 1697 3325 1702
rect 3509 1720 3548 1795
rect 5039 1798 5078 1873
rect 5262 1891 5318 1896
rect 5262 1871 5269 1891
rect 5289 1871 5318 1891
rect 5262 1864 5318 1871
rect 5262 1863 5297 1864
rect 5802 1803 5841 1816
rect 5802 1798 5807 1803
rect 5039 1781 5807 1798
rect 5831 1798 5841 1803
rect 5831 1781 5842 1798
rect 5039 1773 5842 1781
rect 5041 1772 5327 1773
rect 6158 1750 6197 1987
rect 6158 1738 6169 1750
rect 6162 1730 6169 1738
rect 6189 1730 6197 1750
rect 6162 1722 6197 1730
rect 3509 1700 3520 1720
rect 3540 1700 3548 1720
rect 2390 1572 2736 1606
rect 2707 1504 2736 1572
rect 2493 1501 2528 1502
rect 1571 1402 1905 1430
rect 2472 1494 2528 1501
rect 2472 1474 2501 1494
rect 2521 1474 2528 1494
rect 2472 1469 2528 1474
rect 2705 1495 2740 1504
rect 2705 1476 2714 1495
rect 2735 1476 2740 1495
rect 2705 1470 2740 1476
rect 3269 1491 3303 1697
rect 3509 1696 3548 1700
rect 3337 1670 3922 1676
rect 3337 1650 3353 1670
rect 3373 1669 3922 1670
rect 3373 1650 3893 1669
rect 3337 1649 3893 1650
rect 3913 1649 3922 1669
rect 3337 1641 3922 1649
rect 5544 1564 6129 1572
rect 5544 1544 5553 1564
rect 5573 1563 6129 1564
rect 5573 1544 6093 1563
rect 5544 1543 6093 1544
rect 6113 1543 6129 1563
rect 5544 1537 6129 1543
rect 5268 1529 5300 1530
rect 5265 1524 5300 1529
rect 5265 1504 5272 1524
rect 5292 1504 5300 1524
rect 6163 1516 6197 1722
rect 5265 1496 5300 1504
rect 3269 1483 3304 1491
rect 666 1270 701 1277
rect 666 1250 674 1270
rect 694 1250 701 1270
rect 666 1177 701 1250
rect 880 1272 936 1277
rect 880 1252 887 1272
rect 907 1252 936 1272
rect 880 1245 936 1252
rect 971 1379 1001 1381
rect 1700 1379 1733 1380
rect 971 1353 1734 1379
rect 880 1244 915 1245
rect 971 1178 1001 1353
rect 1700 1332 1734 1353
rect 1699 1327 1734 1332
rect 1699 1307 1706 1327
rect 1726 1307 1734 1327
rect 1699 1299 1734 1307
rect 966 1177 1001 1178
rect 665 1150 1001 1177
rect 971 1149 1001 1150
rect 1081 1141 1666 1149
rect 1081 1121 1090 1141
rect 1110 1140 1666 1141
rect 1110 1121 1630 1140
rect 1081 1120 1630 1121
rect 1650 1120 1666 1140
rect 1081 1114 1666 1120
rect 905 1104 937 1105
rect 902 1099 937 1104
rect 902 1079 909 1099
rect 929 1079 937 1099
rect 1700 1093 1734 1299
rect 2472 1263 2506 1469
rect 3269 1463 3277 1483
rect 3297 1463 3304 1483
rect 3269 1458 3304 1463
rect 3269 1457 3301 1458
rect 2540 1442 3125 1448
rect 2540 1422 2556 1442
rect 2576 1441 3125 1442
rect 2576 1422 3096 1441
rect 2540 1421 3096 1422
rect 3116 1421 3125 1441
rect 2540 1413 3125 1421
rect 3205 1412 3235 1413
rect 3205 1385 3541 1412
rect 3205 1384 3240 1385
rect 2472 1255 2507 1263
rect 2472 1235 2480 1255
rect 2500 1235 2507 1255
rect 2472 1230 2507 1235
rect 2472 1209 2506 1230
rect 3205 1209 3235 1384
rect 3291 1317 3326 1318
rect 2472 1183 3235 1209
rect 2473 1182 2506 1183
rect 3205 1181 3235 1183
rect 3270 1310 3326 1317
rect 3270 1290 3299 1310
rect 3319 1290 3326 1310
rect 3270 1285 3326 1290
rect 3505 1312 3540 1385
rect 3505 1292 3512 1312
rect 3532 1292 3540 1312
rect 4647 1338 5232 1346
rect 4647 1318 4656 1338
rect 4676 1337 5232 1338
rect 4676 1318 5196 1337
rect 4647 1317 5196 1318
rect 5216 1317 5232 1337
rect 4647 1311 5232 1317
rect 3505 1285 3540 1292
rect 5266 1290 5300 1496
rect 5929 1504 5965 1513
rect 5929 1487 5938 1504
rect 5957 1487 5965 1504
rect 5929 1478 5965 1487
rect 6141 1511 6197 1516
rect 6141 1491 6148 1511
rect 6168 1491 6197 1511
rect 6141 1484 6197 1491
rect 6141 1483 6176 1484
rect 5935 1443 5961 1478
rect 6237 1443 6269 2252
rect 6681 2185 6710 2870
rect 7641 2851 7927 2852
rect 7126 2843 7929 2851
rect 7126 2826 7137 2843
rect 7127 2821 7137 2826
rect 7161 2826 7929 2843
rect 7161 2821 7166 2826
rect 7127 2808 7166 2821
rect 7671 2760 7706 2761
rect 7650 2753 7706 2760
rect 7650 2733 7679 2753
rect 7699 2733 7706 2753
rect 7650 2728 7706 2733
rect 7890 2751 7929 2826
rect 9436 2828 9475 2903
rect 9659 2921 9715 2926
rect 9659 2901 9666 2921
rect 9686 2901 9715 2921
rect 9659 2894 9715 2901
rect 9659 2893 9694 2894
rect 10199 2833 10238 2846
rect 10199 2828 10204 2833
rect 9436 2811 10204 2828
rect 10228 2828 10238 2833
rect 10228 2811 10239 2828
rect 9436 2803 10239 2811
rect 9438 2802 9724 2803
rect 10655 2784 10684 3469
rect 10992 3223 11019 4923
rect 13836 4952 13844 4972
rect 13864 4952 13875 4972
rect 12055 4899 12341 4900
rect 11540 4891 12343 4899
rect 11540 4874 11551 4891
rect 11541 4869 11551 4874
rect 11575 4874 12343 4891
rect 11575 4869 11580 4874
rect 11541 4856 11580 4869
rect 12085 4808 12120 4809
rect 12064 4801 12120 4808
rect 12064 4781 12093 4801
rect 12113 4781 12120 4801
rect 12064 4776 12120 4781
rect 12304 4799 12343 4874
rect 13836 4877 13875 4952
rect 14059 4970 14115 4975
rect 14059 4950 14066 4970
rect 14086 4950 14115 4970
rect 14059 4943 14115 4950
rect 14059 4942 14094 4943
rect 14599 4882 14638 4895
rect 14599 4877 14604 4882
rect 13836 4860 14604 4877
rect 14628 4877 14638 4882
rect 14628 4860 14639 4877
rect 13836 4852 14639 4860
rect 13838 4851 14124 4852
rect 12304 4779 12315 4799
rect 12335 4779 12343 4799
rect 15160 4828 15187 6528
rect 15495 6282 15524 6967
rect 18139 6962 18147 6982
rect 18167 6962 18178 6982
rect 16455 6948 16741 6949
rect 15940 6940 16743 6948
rect 15940 6923 15951 6940
rect 15941 6918 15951 6923
rect 15975 6923 16743 6940
rect 15975 6918 15980 6923
rect 15941 6905 15980 6918
rect 16485 6857 16520 6858
rect 16464 6850 16520 6857
rect 16464 6830 16493 6850
rect 16513 6830 16520 6850
rect 16464 6825 16520 6830
rect 16704 6848 16743 6923
rect 18139 6887 18178 6962
rect 18362 6980 18418 6985
rect 18362 6960 18369 6980
rect 18389 6960 18418 6980
rect 18362 6953 18418 6960
rect 18362 6952 18397 6953
rect 18902 6892 18941 6905
rect 18902 6887 18907 6892
rect 18139 6870 18907 6887
rect 18931 6887 18941 6892
rect 18931 6870 18942 6887
rect 18139 6862 18942 6870
rect 18141 6861 18427 6862
rect 16704 6828 16715 6848
rect 16735 6828 16743 6848
rect 19358 6843 19387 7528
rect 19799 7461 19831 8270
rect 20107 8235 20133 8270
rect 19892 8229 19927 8230
rect 19871 8222 19927 8229
rect 19871 8202 19900 8222
rect 19920 8202 19927 8222
rect 19871 8197 19927 8202
rect 20103 8226 20139 8235
rect 20103 8209 20111 8226
rect 20130 8209 20139 8226
rect 20103 8200 20139 8209
rect 20768 8217 20802 8423
rect 22528 8421 22563 8428
rect 20836 8396 21421 8402
rect 20836 8376 20852 8396
rect 20872 8395 21421 8396
rect 20872 8376 21392 8395
rect 20836 8375 21392 8376
rect 21412 8375 21421 8395
rect 20836 8367 21421 8375
rect 22528 8401 22536 8421
rect 22556 8401 22563 8421
rect 22528 8328 22563 8401
rect 22742 8423 22798 8428
rect 22742 8403 22749 8423
rect 22769 8403 22798 8423
rect 22742 8396 22798 8403
rect 22833 8530 22863 8532
rect 23562 8530 23595 8531
rect 22833 8504 23596 8530
rect 22742 8395 22777 8396
rect 22833 8329 22863 8504
rect 23562 8483 23596 8504
rect 23561 8478 23596 8483
rect 23561 8458 23568 8478
rect 23588 8458 23596 8478
rect 23561 8450 23596 8458
rect 22828 8328 22863 8329
rect 22527 8301 22863 8328
rect 22833 8300 22863 8301
rect 22943 8292 23528 8300
rect 22943 8272 22952 8292
rect 22972 8291 23528 8292
rect 22972 8272 23492 8291
rect 22943 8271 23492 8272
rect 23512 8271 23528 8291
rect 22943 8265 23528 8271
rect 22767 8255 22799 8256
rect 22764 8250 22799 8255
rect 22764 8230 22771 8250
rect 22791 8230 22799 8250
rect 23562 8244 23596 8450
rect 24334 8414 24368 8620
rect 25131 8614 25139 8634
rect 25159 8614 25166 8634
rect 25131 8609 25166 8614
rect 25131 8608 25163 8609
rect 24402 8593 24987 8599
rect 24402 8573 24418 8593
rect 24438 8592 24987 8593
rect 24438 8573 24958 8592
rect 24402 8572 24958 8573
rect 24978 8572 24987 8592
rect 24402 8564 24987 8572
rect 25067 8563 25097 8564
rect 25067 8536 25403 8563
rect 25067 8535 25102 8536
rect 24334 8406 24369 8414
rect 24334 8386 24342 8406
rect 24362 8386 24369 8406
rect 24334 8381 24369 8386
rect 24334 8360 24368 8381
rect 25067 8360 25097 8535
rect 25153 8468 25188 8469
rect 24334 8334 25097 8360
rect 24335 8333 24368 8334
rect 25067 8332 25097 8334
rect 25132 8461 25188 8468
rect 25132 8441 25161 8461
rect 25181 8441 25188 8461
rect 25132 8436 25188 8441
rect 25367 8463 25402 8536
rect 25367 8443 25374 8463
rect 25394 8443 25402 8463
rect 26522 8488 27107 8496
rect 26522 8468 26531 8488
rect 26551 8487 27107 8488
rect 26551 8468 27071 8487
rect 26522 8467 27071 8468
rect 27091 8467 27107 8487
rect 26522 8461 27107 8467
rect 25367 8436 25402 8443
rect 27141 8440 27175 8646
rect 28711 8657 28767 8664
rect 28711 8637 28740 8657
rect 28760 8637 28767 8657
rect 28711 8632 28767 8637
rect 28944 8660 28978 8667
rect 28944 8642 28952 8660
rect 28971 8642 28978 8660
rect 28944 8634 28978 8642
rect 29508 8654 29542 8860
rect 29748 8859 29787 8863
rect 33872 8898 33928 8905
rect 33872 8878 33901 8898
rect 33921 8878 33928 8898
rect 33872 8873 33928 8878
rect 34112 8896 34151 8971
rect 34112 8876 34123 8896
rect 34143 8876 34151 8896
rect 29576 8833 30161 8839
rect 29576 8813 29592 8833
rect 29612 8832 30161 8833
rect 29612 8813 30132 8832
rect 29576 8812 30132 8813
rect 30152 8812 30161 8832
rect 29576 8804 30161 8812
rect 32956 8737 33338 8742
rect 32956 8718 32964 8737
rect 32985 8718 33338 8737
rect 32956 8710 33338 8718
rect 31507 8692 31539 8693
rect 31504 8687 31539 8692
rect 31504 8667 31511 8687
rect 31531 8667 31539 8687
rect 33309 8680 33338 8710
rect 33096 8677 33131 8678
rect 31504 8659 31539 8667
rect 29508 8646 29543 8654
rect 22764 8222 22799 8230
rect 20768 8209 20803 8217
rect 19871 7991 19905 8197
rect 20768 8189 20776 8209
rect 20796 8189 20803 8209
rect 20768 8184 20803 8189
rect 20768 8183 20800 8184
rect 19939 8170 20524 8176
rect 19939 8150 19955 8170
rect 19975 8169 20524 8170
rect 19975 8150 20495 8169
rect 19939 8149 20495 8150
rect 20515 8149 20524 8169
rect 19939 8141 20524 8149
rect 22146 8064 22731 8072
rect 22146 8044 22155 8064
rect 22175 8063 22731 8064
rect 22175 8044 22695 8063
rect 22146 8043 22695 8044
rect 22715 8043 22731 8063
rect 22146 8037 22731 8043
rect 22520 8013 22559 8017
rect 22765 8016 22799 8222
rect 23328 8237 23363 8243
rect 23328 8218 23333 8237
rect 23354 8218 23363 8237
rect 23328 8209 23363 8218
rect 23540 8239 23596 8244
rect 23540 8219 23547 8239
rect 23567 8219 23596 8239
rect 23540 8212 23596 8219
rect 24163 8283 24497 8311
rect 23540 8211 23575 8212
rect 23332 8141 23361 8209
rect 23332 8107 23678 8141
rect 22520 7993 22528 8013
rect 22548 7993 22559 8013
rect 19871 7983 19906 7991
rect 19871 7963 19879 7983
rect 19899 7975 19906 7983
rect 19899 7963 19910 7975
rect 19871 7726 19910 7963
rect 20741 7940 21027 7941
rect 20226 7932 21029 7940
rect 20226 7915 20237 7932
rect 20227 7910 20237 7915
rect 20261 7915 21029 7932
rect 20261 7910 20266 7915
rect 20227 7897 20266 7910
rect 20771 7849 20806 7850
rect 20750 7842 20806 7849
rect 20750 7822 20779 7842
rect 20799 7822 20806 7842
rect 20750 7817 20806 7822
rect 20990 7840 21029 7915
rect 22520 7918 22559 7993
rect 22743 8011 22799 8016
rect 22743 7991 22750 8011
rect 22770 7991 22799 8011
rect 22743 7984 22799 7991
rect 22743 7983 22778 7984
rect 23283 7923 23322 7936
rect 23283 7918 23288 7923
rect 22520 7901 23288 7918
rect 23312 7918 23322 7923
rect 23312 7901 23323 7918
rect 22520 7893 23323 7901
rect 22522 7892 22808 7893
rect 23639 7870 23678 8107
rect 23639 7858 23650 7870
rect 23643 7850 23650 7858
rect 23670 7850 23678 7870
rect 23643 7842 23678 7850
rect 20990 7820 21001 7840
rect 21021 7820 21029 7840
rect 19871 7692 20217 7726
rect 20188 7624 20217 7692
rect 19974 7621 20009 7622
rect 19799 7443 19802 7461
rect 19824 7443 19831 7461
rect 19799 7431 19831 7443
rect 19953 7614 20009 7621
rect 19953 7594 19982 7614
rect 20002 7594 20009 7614
rect 19953 7589 20009 7594
rect 20186 7615 20221 7624
rect 20186 7596 20195 7615
rect 20216 7596 20221 7615
rect 20186 7590 20221 7596
rect 20750 7611 20784 7817
rect 20990 7816 21029 7820
rect 20818 7790 21403 7796
rect 20818 7770 20834 7790
rect 20854 7789 21403 7790
rect 20854 7770 21374 7789
rect 20818 7769 21374 7770
rect 21394 7769 21403 7789
rect 20818 7761 21403 7769
rect 23025 7684 23610 7692
rect 23025 7664 23034 7684
rect 23054 7683 23610 7684
rect 23054 7664 23574 7683
rect 23025 7663 23574 7664
rect 23594 7663 23610 7683
rect 23025 7657 23610 7663
rect 22749 7649 22781 7650
rect 22746 7644 22781 7649
rect 22746 7624 22753 7644
rect 22773 7624 22781 7644
rect 23644 7636 23678 7842
rect 22746 7616 22781 7624
rect 20750 7603 20785 7611
rect 19953 7383 19987 7589
rect 20750 7583 20758 7603
rect 20778 7583 20785 7603
rect 20750 7578 20785 7583
rect 20750 7577 20782 7578
rect 20021 7562 20606 7568
rect 20021 7542 20037 7562
rect 20057 7561 20606 7562
rect 20057 7542 20577 7561
rect 20021 7541 20577 7542
rect 20597 7541 20606 7561
rect 20021 7533 20606 7541
rect 20686 7532 20716 7533
rect 20686 7505 21022 7532
rect 20686 7504 20721 7505
rect 19953 7375 19988 7383
rect 19953 7355 19961 7375
rect 19981 7355 19988 7375
rect 19953 7350 19988 7355
rect 19953 7329 19987 7350
rect 20686 7329 20716 7504
rect 20772 7437 20807 7438
rect 19953 7303 20716 7329
rect 19954 7302 19987 7303
rect 20686 7301 20716 7303
rect 20751 7430 20807 7437
rect 20751 7410 20780 7430
rect 20800 7410 20807 7430
rect 20751 7405 20807 7410
rect 20986 7432 21021 7505
rect 20986 7412 20993 7432
rect 21013 7412 21021 7432
rect 22128 7458 22713 7466
rect 22128 7438 22137 7458
rect 22157 7457 22713 7458
rect 22157 7438 22677 7457
rect 22128 7437 22677 7438
rect 22697 7437 22713 7457
rect 22128 7431 22713 7437
rect 20986 7405 21021 7412
rect 22747 7410 22781 7616
rect 23412 7630 23443 7636
rect 23412 7611 23417 7630
rect 23438 7611 23443 7630
rect 23412 7569 23443 7611
rect 23622 7631 23678 7636
rect 23622 7611 23629 7631
rect 23649 7611 23678 7631
rect 23622 7604 23678 7611
rect 23622 7603 23657 7604
rect 23412 7541 23751 7569
rect 19591 7269 20054 7277
rect 19591 7247 19603 7269
rect 19627 7247 20054 7269
rect 19591 7246 20054 7247
rect 19593 7234 19632 7246
rect 20027 7215 20054 7246
rect 19809 7213 19844 7214
rect 19788 7206 19844 7213
rect 19788 7186 19817 7206
rect 19837 7186 19844 7206
rect 19788 7181 19844 7186
rect 20023 7206 20056 7215
rect 20023 7184 20028 7206
rect 20051 7184 20056 7206
rect 19788 6975 19822 7181
rect 20023 7178 20056 7184
rect 20751 7199 20785 7405
rect 22511 7403 22546 7410
rect 20819 7378 21404 7384
rect 20819 7358 20835 7378
rect 20855 7377 21404 7378
rect 20855 7358 21375 7377
rect 20819 7357 21375 7358
rect 21395 7357 21404 7377
rect 20819 7349 21404 7357
rect 22511 7383 22519 7403
rect 22539 7383 22546 7403
rect 22511 7310 22546 7383
rect 22725 7405 22781 7410
rect 22725 7385 22732 7405
rect 22752 7385 22781 7405
rect 22725 7378 22781 7385
rect 22816 7512 22846 7514
rect 23545 7512 23578 7513
rect 22816 7486 23579 7512
rect 22725 7377 22760 7378
rect 22816 7311 22846 7486
rect 23545 7465 23579 7486
rect 23544 7460 23579 7465
rect 23544 7440 23551 7460
rect 23571 7440 23579 7460
rect 23544 7432 23579 7440
rect 22811 7310 22846 7311
rect 22510 7283 22846 7310
rect 22816 7282 22846 7283
rect 22926 7274 23511 7282
rect 22926 7254 22935 7274
rect 22955 7273 23511 7274
rect 22955 7254 23475 7273
rect 22926 7253 23475 7254
rect 23495 7253 23511 7273
rect 22926 7247 23511 7253
rect 22750 7237 22782 7238
rect 22747 7232 22782 7237
rect 22747 7212 22754 7232
rect 22774 7212 22782 7232
rect 23545 7226 23579 7432
rect 22747 7204 22782 7212
rect 20751 7191 20786 7199
rect 20751 7171 20759 7191
rect 20779 7171 20786 7191
rect 20751 7166 20786 7171
rect 20751 7165 20783 7166
rect 19856 7154 20441 7160
rect 19856 7134 19872 7154
rect 19892 7153 20441 7154
rect 19892 7134 20412 7153
rect 19856 7133 20412 7134
rect 20432 7133 20441 7153
rect 19856 7125 20441 7133
rect 22129 7046 22714 7054
rect 22129 7026 22138 7046
rect 22158 7045 22714 7046
rect 22158 7026 22678 7045
rect 22129 7025 22678 7026
rect 22698 7025 22714 7045
rect 22129 7019 22714 7025
rect 22503 6995 22542 6999
rect 22748 6998 22782 7204
rect 23312 7216 23346 7224
rect 23312 7198 23319 7216
rect 23338 7198 23346 7216
rect 23312 7191 23346 7198
rect 23523 7221 23579 7226
rect 23523 7201 23530 7221
rect 23550 7201 23579 7221
rect 23523 7194 23579 7201
rect 23523 7193 23558 7194
rect 23316 7161 23345 7191
rect 23316 7153 23698 7161
rect 23316 7134 23669 7153
rect 23690 7134 23698 7153
rect 23316 7129 23698 7134
rect 22503 6975 22511 6995
rect 22531 6975 22542 6995
rect 19788 6974 19823 6975
rect 19756 6967 19823 6974
rect 19756 6947 19796 6967
rect 19816 6947 19823 6967
rect 19756 6944 19823 6947
rect 19756 6941 19821 6944
rect 19327 6840 19392 6843
rect 15548 6689 15930 6694
rect 15548 6670 15556 6689
rect 15577 6670 15930 6689
rect 15548 6662 15930 6670
rect 15901 6632 15930 6662
rect 15688 6629 15723 6630
rect 15667 6622 15723 6629
rect 15667 6602 15696 6622
rect 15716 6602 15723 6622
rect 15667 6597 15723 6602
rect 15900 6625 15934 6632
rect 15900 6607 15908 6625
rect 15927 6607 15934 6625
rect 15900 6599 15934 6607
rect 16464 6619 16498 6825
rect 16704 6824 16743 6828
rect 19325 6837 19392 6840
rect 19325 6817 19332 6837
rect 19352 6817 19392 6837
rect 19325 6810 19392 6817
rect 19325 6809 19360 6810
rect 16532 6798 17117 6804
rect 16532 6778 16548 6798
rect 16568 6797 17117 6798
rect 16568 6778 17088 6797
rect 16532 6777 17088 6778
rect 17108 6777 17117 6797
rect 16532 6769 17117 6777
rect 18707 6651 19292 6659
rect 18707 6631 18716 6651
rect 18736 6650 19292 6651
rect 18736 6631 19256 6650
rect 18707 6630 19256 6631
rect 19276 6630 19292 6650
rect 18707 6624 19292 6630
rect 16464 6611 16499 6619
rect 18365 6618 18397 6619
rect 15667 6391 15701 6597
rect 16464 6591 16472 6611
rect 16492 6591 16499 6611
rect 16464 6586 16499 6591
rect 18362 6613 18397 6618
rect 18362 6593 18369 6613
rect 18389 6593 18397 6613
rect 16464 6585 16496 6586
rect 18362 6585 18397 6593
rect 15735 6570 16320 6576
rect 15735 6550 15751 6570
rect 15771 6569 16320 6570
rect 15771 6550 16291 6569
rect 15735 6549 16291 6550
rect 16311 6549 16320 6569
rect 15735 6541 16320 6549
rect 16400 6540 16430 6541
rect 16400 6513 16736 6540
rect 16400 6512 16435 6513
rect 15667 6383 15702 6391
rect 15667 6363 15675 6383
rect 15695 6363 15702 6383
rect 15667 6358 15702 6363
rect 15667 6337 15701 6358
rect 16400 6337 16430 6512
rect 16486 6445 16521 6446
rect 15667 6311 16430 6337
rect 15668 6310 15701 6311
rect 16400 6309 16430 6311
rect 16465 6438 16521 6445
rect 16465 6418 16494 6438
rect 16514 6418 16521 6438
rect 16465 6413 16521 6418
rect 16700 6440 16735 6513
rect 16700 6420 16707 6440
rect 16727 6420 16735 6440
rect 16700 6413 16735 6420
rect 17744 6427 18329 6435
rect 15495 6254 15834 6282
rect 15589 6219 15624 6220
rect 15568 6212 15624 6219
rect 15568 6192 15597 6212
rect 15617 6192 15624 6212
rect 15568 6187 15624 6192
rect 15803 6212 15834 6254
rect 15803 6193 15808 6212
rect 15829 6193 15834 6212
rect 15803 6187 15834 6193
rect 16465 6207 16499 6413
rect 17744 6407 17753 6427
rect 17773 6426 18329 6427
rect 17773 6407 18293 6426
rect 17744 6406 18293 6407
rect 18313 6406 18329 6426
rect 17744 6400 18329 6406
rect 16533 6386 17118 6392
rect 16533 6366 16549 6386
rect 16569 6385 17118 6386
rect 16569 6366 17089 6385
rect 16533 6365 17089 6366
rect 17109 6365 17118 6385
rect 18363 6379 18397 6585
rect 19090 6595 19131 6606
rect 19326 6603 19360 6809
rect 19090 6577 19100 6595
rect 19118 6577 19131 6595
rect 19090 6569 19131 6577
rect 19304 6598 19360 6603
rect 19304 6578 19311 6598
rect 19331 6578 19360 6598
rect 19304 6571 19360 6578
rect 19304 6570 19339 6571
rect 19099 6539 19125 6569
rect 19099 6538 19437 6539
rect 19099 6502 19453 6538
rect 16533 6357 17118 6365
rect 18127 6372 18162 6379
rect 18127 6352 18135 6372
rect 18155 6352 18162 6372
rect 18127 6279 18162 6352
rect 18341 6374 18397 6379
rect 18341 6354 18348 6374
rect 18368 6354 18397 6374
rect 18341 6347 18397 6354
rect 18432 6481 18462 6483
rect 19161 6481 19194 6482
rect 18432 6455 19195 6481
rect 18341 6346 18376 6347
rect 18432 6280 18462 6455
rect 19161 6434 19195 6455
rect 19160 6429 19195 6434
rect 19160 6409 19167 6429
rect 19187 6409 19195 6429
rect 19160 6401 19195 6409
rect 18427 6279 18462 6280
rect 18126 6252 18462 6279
rect 18432 6251 18462 6252
rect 18542 6243 19127 6251
rect 18542 6223 18551 6243
rect 18571 6242 19127 6243
rect 18571 6223 19091 6242
rect 18542 6222 19091 6223
rect 19111 6222 19127 6242
rect 18542 6216 19127 6222
rect 16465 6199 16500 6207
rect 18366 6206 18398 6207
rect 15568 5981 15602 6187
rect 16465 6179 16473 6199
rect 16493 6179 16500 6199
rect 16465 6174 16500 6179
rect 18363 6201 18398 6206
rect 18363 6181 18370 6201
rect 18390 6181 18398 6201
rect 19161 6195 19195 6401
rect 16465 6173 16497 6174
rect 18363 6173 18398 6181
rect 15636 6160 16221 6166
rect 15636 6140 15652 6160
rect 15672 6159 16221 6160
rect 15672 6140 16192 6159
rect 15636 6139 16192 6140
rect 16212 6139 16221 6159
rect 15636 6131 16221 6139
rect 17745 6015 18330 6023
rect 17745 5995 17754 6015
rect 17774 6014 18330 6015
rect 17774 5995 18294 6014
rect 17745 5994 18294 5995
rect 18314 5994 18330 6014
rect 17745 5988 18330 5994
rect 15568 5973 15603 5981
rect 15568 5953 15576 5973
rect 15596 5965 15603 5973
rect 15596 5953 15607 5965
rect 15568 5716 15607 5953
rect 18119 5964 18158 5968
rect 18364 5967 18398 6173
rect 18927 6188 18962 6194
rect 18927 6169 18932 6188
rect 18953 6169 18962 6188
rect 18927 6160 18962 6169
rect 19139 6190 19195 6195
rect 19139 6170 19146 6190
rect 19166 6170 19195 6190
rect 19139 6163 19195 6170
rect 19139 6162 19174 6163
rect 18931 6092 18960 6160
rect 18931 6058 19277 6092
rect 18119 5944 18127 5964
rect 18147 5944 18158 5964
rect 16438 5930 16724 5931
rect 15923 5922 16726 5930
rect 15923 5905 15934 5922
rect 15924 5900 15934 5905
rect 15958 5905 16726 5922
rect 15958 5900 15963 5905
rect 15924 5887 15963 5900
rect 16468 5839 16503 5840
rect 16447 5832 16503 5839
rect 16447 5812 16476 5832
rect 16496 5812 16503 5832
rect 16447 5807 16503 5812
rect 16687 5830 16726 5905
rect 18119 5869 18158 5944
rect 18342 5962 18398 5967
rect 18342 5942 18349 5962
rect 18369 5942 18398 5962
rect 18342 5935 18398 5942
rect 18342 5934 18377 5935
rect 18882 5874 18921 5887
rect 18882 5869 18887 5874
rect 18119 5852 18887 5869
rect 18911 5869 18921 5874
rect 18911 5852 18922 5869
rect 18119 5844 18922 5852
rect 18121 5843 18407 5844
rect 16687 5810 16698 5830
rect 16718 5810 16726 5830
rect 15568 5682 15914 5716
rect 15885 5614 15914 5682
rect 15671 5611 15706 5612
rect 15650 5604 15706 5611
rect 15650 5584 15679 5604
rect 15699 5584 15706 5604
rect 15650 5579 15706 5584
rect 15883 5605 15918 5614
rect 15883 5586 15892 5605
rect 15913 5586 15918 5605
rect 15883 5580 15918 5586
rect 16447 5601 16481 5807
rect 16687 5806 16726 5810
rect 19238 5821 19277 6058
rect 19238 5809 19249 5821
rect 19242 5801 19249 5809
rect 19269 5801 19277 5821
rect 19242 5793 19277 5801
rect 16515 5780 17100 5786
rect 16515 5760 16531 5780
rect 16551 5779 17100 5780
rect 16551 5760 17071 5779
rect 16515 5759 17071 5760
rect 17091 5759 17100 5779
rect 16515 5751 17100 5759
rect 18624 5635 19209 5643
rect 18624 5615 18633 5635
rect 18653 5634 19209 5635
rect 18653 5615 19173 5634
rect 18624 5614 19173 5615
rect 19193 5614 19209 5634
rect 18624 5608 19209 5614
rect 16447 5593 16482 5601
rect 18348 5600 18380 5601
rect 15650 5373 15684 5579
rect 16447 5573 16455 5593
rect 16475 5573 16482 5593
rect 16447 5568 16482 5573
rect 18345 5595 18380 5600
rect 18345 5575 18352 5595
rect 18372 5575 18380 5595
rect 19243 5587 19277 5793
rect 16447 5567 16479 5568
rect 18345 5567 18380 5575
rect 15718 5552 16303 5558
rect 15718 5532 15734 5552
rect 15754 5551 16303 5552
rect 15754 5532 16274 5551
rect 15718 5531 16274 5532
rect 16294 5531 16303 5551
rect 15718 5523 16303 5531
rect 16383 5522 16413 5523
rect 16383 5495 16719 5522
rect 16383 5494 16418 5495
rect 15650 5365 15685 5373
rect 15650 5345 15658 5365
rect 15678 5345 15685 5365
rect 15650 5340 15685 5345
rect 15650 5319 15684 5340
rect 16383 5319 16413 5494
rect 16469 5427 16504 5428
rect 15650 5293 16413 5319
rect 15651 5292 15684 5293
rect 16383 5291 16413 5293
rect 16448 5420 16504 5427
rect 16448 5400 16477 5420
rect 16497 5400 16504 5420
rect 16448 5395 16504 5400
rect 16683 5422 16718 5495
rect 16683 5402 16690 5422
rect 16710 5402 16718 5422
rect 16683 5395 16718 5402
rect 17727 5409 18312 5417
rect 15302 5272 15619 5275
rect 15302 5245 15305 5272
rect 15332 5245 15619 5272
rect 15302 5239 15619 5245
rect 15302 5236 15338 5239
rect 15583 5209 15619 5239
rect 15367 5205 15402 5206
rect 15346 5198 15402 5205
rect 15346 5178 15375 5198
rect 15395 5178 15402 5198
rect 15346 5173 15402 5178
rect 15581 5203 15619 5209
rect 15581 5177 15587 5203
rect 15613 5177 15619 5203
rect 15346 4974 15380 5173
rect 15581 5169 15619 5177
rect 16448 5189 16482 5395
rect 17727 5389 17736 5409
rect 17756 5408 18312 5409
rect 17756 5389 18276 5408
rect 17727 5388 18276 5389
rect 18296 5388 18312 5408
rect 17727 5382 18312 5388
rect 16516 5368 17101 5374
rect 16516 5348 16532 5368
rect 16552 5367 17101 5368
rect 16552 5348 17072 5367
rect 16516 5347 17072 5348
rect 17092 5347 17101 5367
rect 18346 5361 18380 5567
rect 19009 5575 19045 5584
rect 19009 5558 19018 5575
rect 19037 5558 19045 5575
rect 19009 5549 19045 5558
rect 19221 5582 19277 5587
rect 19221 5562 19228 5582
rect 19248 5562 19277 5582
rect 19221 5555 19277 5562
rect 19221 5554 19256 5555
rect 19015 5514 19041 5549
rect 19323 5514 19355 5515
rect 19015 5509 19355 5514
rect 19015 5491 19330 5509
rect 19352 5491 19355 5509
rect 19015 5486 19355 5491
rect 19323 5485 19355 5486
rect 16516 5339 17101 5347
rect 18110 5354 18145 5361
rect 18110 5334 18118 5354
rect 18138 5334 18145 5354
rect 18110 5261 18145 5334
rect 18324 5356 18380 5361
rect 18324 5336 18331 5356
rect 18351 5336 18380 5356
rect 18324 5329 18380 5336
rect 18415 5463 18445 5465
rect 19144 5463 19177 5464
rect 18415 5437 19178 5463
rect 18324 5328 18359 5329
rect 18415 5262 18445 5437
rect 19144 5416 19178 5437
rect 19143 5411 19178 5416
rect 19143 5391 19150 5411
rect 19170 5391 19178 5411
rect 19143 5383 19178 5391
rect 18410 5261 18445 5262
rect 18109 5234 18445 5261
rect 18415 5233 18445 5234
rect 18525 5225 19110 5233
rect 18525 5205 18534 5225
rect 18554 5224 19110 5225
rect 18554 5205 19074 5224
rect 18525 5204 19074 5205
rect 19094 5204 19110 5224
rect 18525 5198 19110 5204
rect 16448 5181 16483 5189
rect 18349 5188 18381 5189
rect 16448 5161 16456 5181
rect 16476 5161 16483 5181
rect 16448 5156 16483 5161
rect 18346 5183 18381 5188
rect 18346 5163 18353 5183
rect 18373 5163 18381 5183
rect 19144 5177 19178 5383
rect 16448 5155 16480 5156
rect 18346 5155 18381 5163
rect 15414 5146 15999 5152
rect 15414 5126 15430 5146
rect 15450 5145 15999 5146
rect 15450 5126 15970 5145
rect 15414 5125 15970 5126
rect 15990 5125 15999 5145
rect 15414 5117 15999 5125
rect 17728 4997 18313 5005
rect 17728 4977 17737 4997
rect 17757 4996 18313 4997
rect 17757 4977 18277 4996
rect 17728 4976 18277 4977
rect 18297 4976 18313 4996
rect 15346 4959 15383 4974
rect 17728 4970 18313 4976
rect 15346 4939 15354 4959
rect 15374 4939 15383 4959
rect 15346 4936 15383 4939
rect 15160 4825 15197 4828
rect 15160 4805 15169 4825
rect 15189 4805 15197 4825
rect 15160 4790 15197 4805
rect 11148 4640 11530 4645
rect 11148 4621 11156 4640
rect 11177 4621 11530 4640
rect 11148 4613 11530 4621
rect 11501 4583 11530 4613
rect 11288 4580 11323 4581
rect 11267 4573 11323 4580
rect 11267 4553 11296 4573
rect 11316 4553 11323 4573
rect 11267 4548 11323 4553
rect 11500 4576 11534 4583
rect 11500 4558 11508 4576
rect 11527 4558 11534 4576
rect 11500 4550 11534 4558
rect 12064 4570 12098 4776
rect 12304 4775 12343 4779
rect 12132 4749 12717 4755
rect 12132 4729 12148 4749
rect 12168 4748 12717 4749
rect 12168 4729 12688 4748
rect 12132 4728 12688 4729
rect 12708 4728 12717 4748
rect 12132 4720 12717 4728
rect 14544 4639 15129 4647
rect 14544 4619 14553 4639
rect 14573 4638 15129 4639
rect 14573 4619 15093 4638
rect 14544 4618 15093 4619
rect 15113 4618 15129 4638
rect 14544 4612 15129 4618
rect 14063 4608 14095 4609
rect 14060 4603 14095 4608
rect 14060 4583 14067 4603
rect 14087 4583 14095 4603
rect 15163 4591 15197 4790
rect 15141 4586 15197 4591
rect 14060 4575 14095 4583
rect 12064 4562 12099 4570
rect 11267 4342 11301 4548
rect 12064 4542 12072 4562
rect 12092 4542 12099 4562
rect 12064 4537 12099 4542
rect 12064 4536 12096 4537
rect 11335 4521 11920 4527
rect 11335 4501 11351 4521
rect 11371 4520 11920 4521
rect 11371 4501 11891 4520
rect 11335 4500 11891 4501
rect 11911 4500 11920 4520
rect 11335 4492 11920 4500
rect 12000 4491 12030 4492
rect 12000 4464 12336 4491
rect 12000 4463 12035 4464
rect 11267 4334 11302 4342
rect 11267 4314 11275 4334
rect 11295 4314 11302 4334
rect 11267 4309 11302 4314
rect 11267 4288 11301 4309
rect 12000 4288 12030 4463
rect 12086 4396 12121 4397
rect 11267 4262 12030 4288
rect 11268 4261 11301 4262
rect 12000 4260 12030 4262
rect 12065 4389 12121 4396
rect 12065 4369 12094 4389
rect 12114 4369 12121 4389
rect 12065 4364 12121 4369
rect 12300 4391 12335 4464
rect 12300 4371 12307 4391
rect 12327 4371 12335 4391
rect 13442 4417 14027 4425
rect 13442 4397 13451 4417
rect 13471 4416 14027 4417
rect 13471 4397 13991 4416
rect 13442 4396 13991 4397
rect 14011 4396 14027 4416
rect 13442 4390 14027 4396
rect 12300 4364 12335 4371
rect 14061 4369 14095 4575
rect 14923 4584 14958 4586
rect 14923 4578 14961 4584
rect 14923 4555 14931 4578
rect 14954 4555 14961 4578
rect 15141 4566 15148 4586
rect 15168 4566 15197 4586
rect 15141 4559 15197 4566
rect 15141 4558 15176 4559
rect 14923 4549 14961 4555
rect 14923 4536 14958 4549
rect 14921 4478 14958 4536
rect 11090 4239 11122 4240
rect 11090 4234 11430 4239
rect 11090 4216 11093 4234
rect 11115 4216 11430 4234
rect 11090 4211 11430 4216
rect 11090 4210 11122 4211
rect 11404 4176 11430 4211
rect 11189 4170 11224 4171
rect 11168 4163 11224 4170
rect 11168 4143 11197 4163
rect 11217 4143 11224 4163
rect 11168 4138 11224 4143
rect 11400 4167 11436 4176
rect 11400 4150 11408 4167
rect 11427 4150 11436 4167
rect 11400 4141 11436 4150
rect 12065 4158 12099 4364
rect 13825 4362 13860 4369
rect 12133 4337 12718 4343
rect 12133 4317 12149 4337
rect 12169 4336 12718 4337
rect 12169 4317 12689 4336
rect 12133 4316 12689 4317
rect 12709 4316 12718 4336
rect 12133 4308 12718 4316
rect 13825 4342 13833 4362
rect 13853 4342 13860 4362
rect 13825 4269 13860 4342
rect 14039 4364 14095 4369
rect 14039 4344 14046 4364
rect 14066 4344 14095 4364
rect 14039 4337 14095 4344
rect 14130 4471 14160 4473
rect 14859 4471 14892 4472
rect 14130 4445 14893 4471
rect 14039 4336 14074 4337
rect 14130 4270 14160 4445
rect 14859 4424 14893 4445
rect 14921 4461 14956 4478
rect 14921 4460 15215 4461
rect 14921 4459 15258 4460
rect 14921 4452 15263 4459
rect 14921 4426 15223 4452
rect 15254 4426 15263 4452
rect 14858 4419 14893 4424
rect 15214 4423 15263 4426
rect 14858 4399 14865 4419
rect 14885 4399 14893 4419
rect 15220 4418 15263 4423
rect 14858 4391 14893 4399
rect 14125 4269 14160 4270
rect 13824 4242 14160 4269
rect 14130 4241 14160 4242
rect 14240 4233 14825 4241
rect 14240 4213 14249 4233
rect 14269 4232 14825 4233
rect 14269 4213 14789 4232
rect 14240 4212 14789 4213
rect 14809 4212 14825 4232
rect 14240 4206 14825 4212
rect 14064 4196 14096 4197
rect 14061 4191 14096 4196
rect 14061 4171 14068 4191
rect 14088 4171 14096 4191
rect 14859 4185 14893 4391
rect 14061 4163 14096 4171
rect 12065 4150 12100 4158
rect 11168 3932 11202 4138
rect 12065 4130 12073 4150
rect 12093 4130 12100 4150
rect 12065 4125 12100 4130
rect 12065 4124 12097 4125
rect 11236 4111 11821 4117
rect 11236 4091 11252 4111
rect 11272 4110 11821 4111
rect 11272 4091 11792 4110
rect 11236 4090 11792 4091
rect 11812 4090 11821 4110
rect 11236 4082 11821 4090
rect 13443 4005 14028 4013
rect 13443 3985 13452 4005
rect 13472 4004 14028 4005
rect 13472 3985 13992 4004
rect 13443 3984 13992 3985
rect 14012 3984 14028 4004
rect 13443 3978 14028 3984
rect 13817 3954 13856 3958
rect 14062 3957 14096 4163
rect 14625 4178 14660 4184
rect 14625 4159 14630 4178
rect 14651 4159 14660 4178
rect 14625 4150 14660 4159
rect 14837 4180 14893 4185
rect 14837 4160 14844 4180
rect 14864 4160 14893 4180
rect 14837 4153 14893 4160
rect 14837 4152 14872 4153
rect 14629 4082 14658 4150
rect 14629 4048 14975 4082
rect 13817 3934 13825 3954
rect 13845 3934 13856 3954
rect 11168 3924 11203 3932
rect 11168 3904 11176 3924
rect 11196 3916 11203 3924
rect 11196 3904 11207 3916
rect 11168 3667 11207 3904
rect 12038 3881 12324 3882
rect 11523 3873 12326 3881
rect 11523 3856 11534 3873
rect 11524 3851 11534 3856
rect 11558 3856 12326 3873
rect 11558 3851 11563 3856
rect 11524 3838 11563 3851
rect 12068 3790 12103 3791
rect 12047 3783 12103 3790
rect 12047 3763 12076 3783
rect 12096 3763 12103 3783
rect 12047 3758 12103 3763
rect 12287 3781 12326 3856
rect 13817 3859 13856 3934
rect 14040 3952 14096 3957
rect 14040 3932 14047 3952
rect 14067 3932 14096 3952
rect 14040 3925 14096 3932
rect 14040 3924 14075 3925
rect 14580 3864 14619 3877
rect 14580 3859 14585 3864
rect 13817 3842 14585 3859
rect 14609 3859 14619 3864
rect 14609 3842 14620 3859
rect 13817 3834 14620 3842
rect 13819 3833 14105 3834
rect 14936 3811 14975 4048
rect 14936 3799 14947 3811
rect 14940 3791 14947 3799
rect 14967 3791 14975 3811
rect 14940 3783 14975 3791
rect 12287 3761 12298 3781
rect 12318 3761 12326 3781
rect 11168 3633 11514 3667
rect 11485 3565 11514 3633
rect 11271 3562 11306 3563
rect 11250 3555 11306 3562
rect 11250 3535 11279 3555
rect 11299 3535 11306 3555
rect 11250 3530 11306 3535
rect 11483 3556 11518 3565
rect 11483 3537 11492 3556
rect 11513 3537 11518 3556
rect 11483 3531 11518 3537
rect 12047 3552 12081 3758
rect 12287 3757 12326 3761
rect 12115 3731 12700 3737
rect 12115 3711 12131 3731
rect 12151 3730 12700 3731
rect 12151 3711 12671 3730
rect 12115 3710 12671 3711
rect 12691 3710 12700 3730
rect 12115 3702 12700 3710
rect 14322 3625 14907 3633
rect 14322 3605 14331 3625
rect 14351 3624 14907 3625
rect 14351 3605 14871 3624
rect 14322 3604 14871 3605
rect 14891 3604 14907 3624
rect 14322 3598 14907 3604
rect 14046 3590 14078 3591
rect 14043 3585 14078 3590
rect 14043 3565 14050 3585
rect 14070 3565 14078 3585
rect 14941 3577 14975 3783
rect 14043 3557 14078 3565
rect 12047 3544 12082 3552
rect 11250 3324 11284 3530
rect 12047 3524 12055 3544
rect 12075 3524 12082 3544
rect 12047 3519 12082 3524
rect 12047 3518 12079 3519
rect 11318 3503 11903 3509
rect 11318 3483 11334 3503
rect 11354 3502 11903 3503
rect 11354 3483 11874 3502
rect 11318 3482 11874 3483
rect 11894 3482 11903 3502
rect 11318 3474 11903 3482
rect 11983 3473 12013 3474
rect 11983 3446 12319 3473
rect 11983 3445 12018 3446
rect 11250 3316 11285 3324
rect 11250 3296 11258 3316
rect 11278 3296 11285 3316
rect 11250 3291 11285 3296
rect 11250 3270 11284 3291
rect 11983 3270 12013 3445
rect 12069 3378 12104 3379
rect 11250 3244 12013 3270
rect 11251 3243 11284 3244
rect 11983 3242 12013 3244
rect 12048 3371 12104 3378
rect 12048 3351 12077 3371
rect 12097 3351 12104 3371
rect 12048 3346 12104 3351
rect 12283 3373 12318 3446
rect 12283 3353 12290 3373
rect 12310 3353 12318 3373
rect 13425 3399 14010 3407
rect 13425 3379 13434 3399
rect 13454 3398 14010 3399
rect 13454 3379 13974 3398
rect 13425 3378 13974 3379
rect 13994 3378 14010 3398
rect 13425 3372 14010 3378
rect 12283 3346 12318 3353
rect 14044 3351 14078 3557
rect 14709 3571 14740 3577
rect 14709 3552 14714 3571
rect 14735 3552 14740 3571
rect 14709 3510 14740 3552
rect 14919 3572 14975 3577
rect 14919 3552 14926 3572
rect 14946 3552 14975 3572
rect 14919 3545 14975 3552
rect 14919 3544 14954 3545
rect 14709 3482 15048 3510
rect 10992 3187 11346 3223
rect 11008 3186 11346 3187
rect 11320 3156 11346 3186
rect 11106 3154 11141 3155
rect 11085 3147 11141 3154
rect 11085 3127 11114 3147
rect 11134 3127 11141 3147
rect 11085 3122 11141 3127
rect 11314 3148 11355 3156
rect 11314 3130 11327 3148
rect 11345 3130 11355 3148
rect 11085 2916 11119 3122
rect 11314 3119 11355 3130
rect 12048 3140 12082 3346
rect 13808 3344 13843 3351
rect 12116 3319 12701 3325
rect 12116 3299 12132 3319
rect 12152 3318 12701 3319
rect 12152 3299 12672 3318
rect 12116 3298 12672 3299
rect 12692 3298 12701 3318
rect 12116 3290 12701 3298
rect 13808 3324 13816 3344
rect 13836 3324 13843 3344
rect 13808 3251 13843 3324
rect 14022 3346 14078 3351
rect 14022 3326 14029 3346
rect 14049 3326 14078 3346
rect 14022 3319 14078 3326
rect 14113 3453 14143 3455
rect 14842 3453 14875 3454
rect 14113 3427 14876 3453
rect 14022 3318 14057 3319
rect 14113 3252 14143 3427
rect 14842 3406 14876 3427
rect 14841 3401 14876 3406
rect 14841 3381 14848 3401
rect 14868 3381 14876 3401
rect 14841 3373 14876 3381
rect 14108 3251 14143 3252
rect 13807 3224 14143 3251
rect 14113 3223 14143 3224
rect 14223 3215 14808 3223
rect 14223 3195 14232 3215
rect 14252 3214 14808 3215
rect 14252 3195 14772 3214
rect 14223 3194 14772 3195
rect 14792 3194 14808 3214
rect 14223 3188 14808 3194
rect 14047 3178 14079 3179
rect 14044 3173 14079 3178
rect 14044 3153 14051 3173
rect 14071 3153 14079 3173
rect 14842 3167 14876 3373
rect 14044 3145 14079 3153
rect 12048 3132 12083 3140
rect 12048 3112 12056 3132
rect 12076 3112 12083 3132
rect 12048 3107 12083 3112
rect 12048 3106 12080 3107
rect 11153 3095 11738 3101
rect 11153 3075 11169 3095
rect 11189 3094 11738 3095
rect 11189 3075 11709 3094
rect 11153 3074 11709 3075
rect 11729 3074 11738 3094
rect 11153 3066 11738 3074
rect 13426 2987 14011 2995
rect 13426 2967 13435 2987
rect 13455 2986 14011 2987
rect 13455 2967 13975 2986
rect 13426 2966 13975 2967
rect 13995 2966 14011 2986
rect 13426 2960 14011 2966
rect 13800 2936 13839 2940
rect 14045 2939 14079 3145
rect 14609 3157 14643 3165
rect 14609 3139 14616 3157
rect 14635 3139 14643 3157
rect 14609 3132 14643 3139
rect 14820 3162 14876 3167
rect 14820 3142 14827 3162
rect 14847 3142 14876 3162
rect 14820 3135 14876 3142
rect 14820 3134 14855 3135
rect 14613 3102 14642 3132
rect 14613 3094 14995 3102
rect 14613 3075 14966 3094
rect 14987 3075 14995 3094
rect 14613 3070 14995 3075
rect 13800 2916 13808 2936
rect 13828 2916 13839 2936
rect 11085 2915 11120 2916
rect 11053 2908 11120 2915
rect 11053 2888 11093 2908
rect 11113 2888 11120 2908
rect 11053 2885 11120 2888
rect 11053 2882 11118 2885
rect 10624 2781 10689 2784
rect 7890 2731 7901 2751
rect 7921 2731 7929 2751
rect 10622 2778 10689 2781
rect 10622 2758 10629 2778
rect 10649 2758 10689 2778
rect 10622 2751 10689 2758
rect 10622 2750 10657 2751
rect 6734 2592 7116 2597
rect 6734 2573 6742 2592
rect 6763 2573 7116 2592
rect 6734 2565 7116 2573
rect 7087 2535 7116 2565
rect 6874 2532 6909 2533
rect 6853 2525 6909 2532
rect 6853 2505 6882 2525
rect 6902 2505 6909 2525
rect 6853 2500 6909 2505
rect 7086 2528 7120 2535
rect 7086 2510 7094 2528
rect 7113 2510 7120 2528
rect 7086 2502 7120 2510
rect 7650 2522 7684 2728
rect 7890 2727 7929 2731
rect 7718 2701 8303 2707
rect 7718 2681 7734 2701
rect 7754 2700 8303 2701
rect 7754 2681 8274 2700
rect 7718 2680 8274 2681
rect 8294 2680 8303 2700
rect 7718 2672 8303 2680
rect 10004 2592 10589 2600
rect 10004 2572 10013 2592
rect 10033 2591 10589 2592
rect 10033 2572 10553 2591
rect 10004 2571 10553 2572
rect 10573 2571 10589 2591
rect 10004 2565 10589 2571
rect 9662 2559 9694 2560
rect 9659 2554 9694 2559
rect 9659 2534 9666 2554
rect 9686 2534 9694 2554
rect 9659 2526 9694 2534
rect 7650 2514 7685 2522
rect 6853 2294 6887 2500
rect 7650 2494 7658 2514
rect 7678 2494 7685 2514
rect 7650 2489 7685 2494
rect 7650 2488 7682 2489
rect 6921 2473 7506 2479
rect 6921 2453 6937 2473
rect 6957 2472 7506 2473
rect 6957 2453 7477 2472
rect 6921 2452 7477 2453
rect 7497 2452 7506 2472
rect 6921 2444 7506 2452
rect 7586 2443 7616 2444
rect 7586 2416 7922 2443
rect 7586 2415 7621 2416
rect 6853 2286 6888 2294
rect 6853 2266 6861 2286
rect 6881 2266 6888 2286
rect 6853 2261 6888 2266
rect 6853 2240 6887 2261
rect 7586 2240 7616 2415
rect 7672 2348 7707 2349
rect 6853 2214 7616 2240
rect 6854 2213 6887 2214
rect 7586 2212 7616 2214
rect 7651 2341 7707 2348
rect 7651 2321 7680 2341
rect 7700 2321 7707 2341
rect 7651 2316 7707 2321
rect 7886 2343 7921 2416
rect 7886 2323 7893 2343
rect 7913 2323 7921 2343
rect 9041 2368 9626 2376
rect 9041 2348 9050 2368
rect 9070 2367 9626 2368
rect 9070 2348 9590 2367
rect 9041 2347 9590 2348
rect 9610 2347 9626 2367
rect 9041 2341 9626 2347
rect 7886 2316 7921 2323
rect 9660 2320 9694 2526
rect 10389 2541 10422 2547
rect 10623 2544 10657 2750
rect 10389 2519 10394 2541
rect 10417 2519 10422 2541
rect 10389 2510 10422 2519
rect 10601 2539 10657 2544
rect 10601 2519 10608 2539
rect 10628 2519 10657 2539
rect 10601 2512 10657 2519
rect 10601 2511 10636 2512
rect 10391 2479 10418 2510
rect 10813 2479 10852 2491
rect 10391 2478 10854 2479
rect 10391 2456 10818 2478
rect 10842 2456 10854 2478
rect 10391 2448 10854 2456
rect 6681 2157 7020 2185
rect 6775 2122 6810 2123
rect 6754 2115 6810 2122
rect 6754 2095 6783 2115
rect 6803 2095 6810 2115
rect 6754 2090 6810 2095
rect 6989 2115 7020 2157
rect 6989 2096 6994 2115
rect 7015 2096 7020 2115
rect 6989 2090 7020 2096
rect 7651 2110 7685 2316
rect 9424 2313 9459 2320
rect 7719 2289 8304 2295
rect 7719 2269 7735 2289
rect 7755 2288 8304 2289
rect 7755 2269 8275 2288
rect 7719 2268 8275 2269
rect 8295 2268 8304 2288
rect 7719 2260 8304 2268
rect 9424 2293 9432 2313
rect 9452 2293 9459 2313
rect 9424 2220 9459 2293
rect 9638 2315 9694 2320
rect 9638 2295 9645 2315
rect 9665 2295 9694 2315
rect 9638 2288 9694 2295
rect 9729 2422 9759 2424
rect 10458 2422 10491 2423
rect 9729 2396 10492 2422
rect 9638 2287 9673 2288
rect 9729 2221 9759 2396
rect 10458 2375 10492 2396
rect 10457 2370 10492 2375
rect 10457 2350 10464 2370
rect 10484 2350 10492 2370
rect 10457 2342 10492 2350
rect 9724 2220 9759 2221
rect 9423 2193 9759 2220
rect 9729 2192 9759 2193
rect 9839 2184 10424 2192
rect 9839 2164 9848 2184
rect 9868 2183 10424 2184
rect 9868 2164 10388 2183
rect 9839 2163 10388 2164
rect 10408 2163 10424 2183
rect 9839 2157 10424 2163
rect 9663 2147 9695 2148
rect 9660 2142 9695 2147
rect 9660 2122 9667 2142
rect 9687 2122 9695 2142
rect 10458 2136 10492 2342
rect 9660 2114 9695 2122
rect 7651 2102 7686 2110
rect 6754 1884 6788 2090
rect 7651 2082 7659 2102
rect 7679 2082 7686 2102
rect 7651 2077 7686 2082
rect 7651 2076 7683 2077
rect 6822 2063 7407 2069
rect 6822 2043 6838 2063
rect 6858 2062 7407 2063
rect 6858 2043 7378 2062
rect 6822 2042 7378 2043
rect 7398 2042 7407 2062
rect 6822 2034 7407 2042
rect 9042 1956 9627 1964
rect 9042 1936 9051 1956
rect 9071 1955 9627 1956
rect 9071 1936 9591 1955
rect 9042 1935 9591 1936
rect 9611 1935 9627 1955
rect 9042 1929 9627 1935
rect 9416 1905 9455 1909
rect 9661 1908 9695 2114
rect 10224 2129 10259 2135
rect 10224 2110 10229 2129
rect 10250 2110 10259 2129
rect 10224 2101 10259 2110
rect 10436 2131 10492 2136
rect 10436 2111 10443 2131
rect 10463 2111 10492 2131
rect 10436 2104 10492 2111
rect 10614 2282 10646 2294
rect 10614 2264 10621 2282
rect 10643 2264 10646 2282
rect 10436 2103 10471 2104
rect 10228 2033 10257 2101
rect 10228 1999 10574 2033
rect 9416 1885 9424 1905
rect 9444 1885 9455 1905
rect 6754 1876 6789 1884
rect 6754 1856 6762 1876
rect 6782 1868 6789 1876
rect 6782 1856 6793 1868
rect 6754 1619 6793 1856
rect 7624 1833 7910 1834
rect 7109 1825 7912 1833
rect 7109 1808 7120 1825
rect 7110 1803 7120 1808
rect 7144 1808 7912 1825
rect 7144 1803 7149 1808
rect 7110 1790 7149 1803
rect 7654 1742 7689 1743
rect 7633 1735 7689 1742
rect 7633 1715 7662 1735
rect 7682 1715 7689 1735
rect 7633 1710 7689 1715
rect 7873 1733 7912 1808
rect 9416 1810 9455 1885
rect 9639 1903 9695 1908
rect 9639 1883 9646 1903
rect 9666 1883 9695 1903
rect 9639 1876 9695 1883
rect 9639 1875 9674 1876
rect 10179 1815 10218 1828
rect 10179 1810 10184 1815
rect 9416 1793 10184 1810
rect 10208 1810 10218 1815
rect 10208 1793 10219 1810
rect 9416 1785 10219 1793
rect 9418 1784 9704 1785
rect 10535 1762 10574 1999
rect 10535 1750 10546 1762
rect 10539 1742 10546 1750
rect 10566 1742 10574 1762
rect 10539 1734 10574 1742
rect 7873 1713 7884 1733
rect 7904 1713 7912 1733
rect 6754 1585 7100 1619
rect 7071 1517 7100 1585
rect 6857 1514 6892 1515
rect 5935 1415 6269 1443
rect 6836 1507 6892 1514
rect 6836 1487 6865 1507
rect 6885 1487 6892 1507
rect 6836 1482 6892 1487
rect 7069 1508 7104 1517
rect 7069 1489 7078 1508
rect 7099 1489 7104 1508
rect 7069 1483 7104 1489
rect 7633 1504 7667 1710
rect 7873 1709 7912 1713
rect 7701 1683 8286 1689
rect 7701 1663 7717 1683
rect 7737 1682 8286 1683
rect 7737 1663 8257 1682
rect 7701 1662 8257 1663
rect 8277 1662 8286 1682
rect 7701 1654 8286 1662
rect 9921 1576 10506 1584
rect 9921 1556 9930 1576
rect 9950 1575 10506 1576
rect 9950 1556 10470 1575
rect 9921 1555 10470 1556
rect 10490 1555 10506 1575
rect 9921 1549 10506 1555
rect 9645 1541 9677 1542
rect 9642 1536 9677 1541
rect 9642 1516 9649 1536
rect 9669 1516 9677 1536
rect 10540 1528 10574 1734
rect 9642 1508 9677 1516
rect 7633 1496 7668 1504
rect 902 1071 937 1079
rect 284 913 869 921
rect 284 893 293 913
rect 313 912 869 913
rect 313 893 833 912
rect 284 892 833 893
rect 853 892 869 912
rect 284 886 869 892
rect 658 862 697 866
rect 903 865 937 1071
rect 1467 1083 1501 1091
rect 1467 1065 1474 1083
rect 1493 1065 1501 1083
rect 1467 1058 1501 1065
rect 1678 1088 1734 1093
rect 1678 1068 1685 1088
rect 1705 1068 1734 1088
rect 1678 1061 1734 1068
rect 3270 1079 3304 1285
rect 5030 1283 5065 1290
rect 3338 1258 3923 1264
rect 3338 1238 3354 1258
rect 3374 1257 3923 1258
rect 3374 1238 3894 1257
rect 3338 1237 3894 1238
rect 3914 1237 3923 1257
rect 3338 1229 3923 1237
rect 5030 1263 5038 1283
rect 5058 1263 5065 1283
rect 5030 1190 5065 1263
rect 5244 1285 5300 1290
rect 5244 1265 5251 1285
rect 5271 1265 5300 1285
rect 5244 1258 5300 1265
rect 5335 1392 5365 1394
rect 6064 1392 6097 1393
rect 5335 1366 6098 1392
rect 5244 1257 5279 1258
rect 5335 1191 5365 1366
rect 6064 1345 6098 1366
rect 6063 1340 6098 1345
rect 6063 1320 6070 1340
rect 6090 1320 6098 1340
rect 6063 1312 6098 1320
rect 5330 1190 5365 1191
rect 5029 1163 5365 1190
rect 5335 1162 5365 1163
rect 5445 1154 6030 1162
rect 5445 1134 5454 1154
rect 5474 1153 6030 1154
rect 5474 1134 5994 1153
rect 5445 1133 5994 1134
rect 6014 1133 6030 1153
rect 5445 1127 6030 1133
rect 5269 1117 5301 1118
rect 5266 1112 5301 1117
rect 5266 1092 5273 1112
rect 5293 1092 5301 1112
rect 6064 1106 6098 1312
rect 6836 1276 6870 1482
rect 7633 1476 7641 1496
rect 7661 1476 7668 1496
rect 7633 1471 7668 1476
rect 7633 1470 7665 1471
rect 6904 1455 7489 1461
rect 6904 1435 6920 1455
rect 6940 1454 7489 1455
rect 6940 1435 7460 1454
rect 6904 1434 7460 1435
rect 7480 1434 7489 1454
rect 6904 1426 7489 1434
rect 7569 1425 7599 1426
rect 7569 1398 7905 1425
rect 7569 1397 7604 1398
rect 6836 1268 6871 1276
rect 6836 1248 6844 1268
rect 6864 1248 6871 1268
rect 6836 1243 6871 1248
rect 6836 1222 6870 1243
rect 7569 1222 7599 1397
rect 7655 1330 7690 1331
rect 6836 1196 7599 1222
rect 6837 1195 6870 1196
rect 7569 1194 7599 1196
rect 7634 1323 7690 1330
rect 7634 1303 7663 1323
rect 7683 1303 7690 1323
rect 7634 1298 7690 1303
rect 7869 1325 7904 1398
rect 7869 1305 7876 1325
rect 7896 1305 7904 1325
rect 9024 1350 9609 1358
rect 9024 1330 9033 1350
rect 9053 1349 9609 1350
rect 9053 1330 9573 1349
rect 9024 1329 9573 1330
rect 9593 1329 9609 1349
rect 9024 1323 9609 1329
rect 7869 1298 7904 1305
rect 9643 1302 9677 1508
rect 10306 1516 10342 1525
rect 10306 1499 10315 1516
rect 10334 1499 10342 1516
rect 10306 1490 10342 1499
rect 10518 1523 10574 1528
rect 10518 1503 10525 1523
rect 10545 1503 10574 1523
rect 10518 1496 10574 1503
rect 10518 1495 10553 1496
rect 10312 1455 10338 1490
rect 10614 1455 10646 2264
rect 11058 2197 11087 2882
rect 12018 2863 12304 2864
rect 11503 2855 12306 2863
rect 11503 2838 11514 2855
rect 11504 2833 11514 2838
rect 11538 2838 12306 2855
rect 11538 2833 11543 2838
rect 11504 2820 11543 2833
rect 12048 2772 12083 2773
rect 12027 2765 12083 2772
rect 12027 2745 12056 2765
rect 12076 2745 12083 2765
rect 12027 2740 12083 2745
rect 12267 2763 12306 2838
rect 13800 2841 13839 2916
rect 14023 2934 14079 2939
rect 14023 2914 14030 2934
rect 14050 2914 14079 2934
rect 14023 2907 14079 2914
rect 14023 2906 14058 2907
rect 14563 2846 14602 2859
rect 14563 2841 14568 2846
rect 13800 2824 14568 2841
rect 14592 2841 14602 2846
rect 14592 2824 14603 2841
rect 13800 2816 14603 2824
rect 13802 2815 14088 2816
rect 15019 2797 15048 3482
rect 15356 3236 15383 4936
rect 18102 4946 18141 4950
rect 18347 4949 18381 5155
rect 18911 5167 18945 5175
rect 18911 5149 18918 5167
rect 18937 5149 18945 5167
rect 18911 5142 18945 5149
rect 19122 5172 19178 5177
rect 19122 5152 19129 5172
rect 19149 5152 19178 5172
rect 19122 5145 19178 5152
rect 19122 5144 19157 5145
rect 18915 5112 18944 5142
rect 18915 5104 19297 5112
rect 18915 5085 19268 5104
rect 19289 5085 19297 5104
rect 18915 5080 19297 5085
rect 18102 4926 18110 4946
rect 18130 4926 18141 4946
rect 16419 4912 16705 4913
rect 15904 4904 16707 4912
rect 15904 4887 15915 4904
rect 15905 4882 15915 4887
rect 15939 4887 16707 4904
rect 15939 4882 15944 4887
rect 15905 4869 15944 4882
rect 16449 4821 16484 4822
rect 16428 4814 16484 4821
rect 16428 4794 16457 4814
rect 16477 4794 16484 4814
rect 16428 4789 16484 4794
rect 16668 4812 16707 4887
rect 18102 4851 18141 4926
rect 18325 4944 18381 4949
rect 18325 4924 18332 4944
rect 18352 4924 18381 4944
rect 18325 4917 18381 4924
rect 18325 4916 18360 4917
rect 18865 4856 18904 4869
rect 18865 4851 18870 4856
rect 18102 4834 18870 4851
rect 18894 4851 18904 4856
rect 18894 4834 18905 4851
rect 18102 4826 18905 4834
rect 18104 4825 18390 4826
rect 16668 4792 16679 4812
rect 16699 4792 16707 4812
rect 15512 4653 15894 4658
rect 15512 4634 15520 4653
rect 15541 4634 15894 4653
rect 15512 4626 15894 4634
rect 15865 4596 15894 4626
rect 15652 4593 15687 4594
rect 15631 4586 15687 4593
rect 15631 4566 15660 4586
rect 15680 4566 15687 4586
rect 15631 4561 15687 4566
rect 15864 4589 15898 4596
rect 15864 4571 15872 4589
rect 15891 4571 15898 4589
rect 15864 4563 15898 4571
rect 16428 4583 16462 4789
rect 16668 4788 16707 4792
rect 19426 4802 19453 6502
rect 19761 6256 19790 6941
rect 20721 6922 21007 6923
rect 20206 6914 21009 6922
rect 20206 6897 20217 6914
rect 20207 6892 20217 6897
rect 20241 6897 21009 6914
rect 20241 6892 20246 6897
rect 20207 6879 20246 6892
rect 20751 6831 20786 6832
rect 20730 6824 20786 6831
rect 20730 6804 20759 6824
rect 20779 6804 20786 6824
rect 20730 6799 20786 6804
rect 20970 6822 21009 6897
rect 22503 6900 22542 6975
rect 22726 6993 22782 6998
rect 22726 6973 22733 6993
rect 22753 6973 22782 6993
rect 22726 6966 22782 6973
rect 22726 6965 22761 6966
rect 23266 6905 23305 6918
rect 23266 6900 23271 6905
rect 22503 6883 23271 6900
rect 23295 6900 23305 6905
rect 23295 6883 23306 6900
rect 22503 6875 23306 6883
rect 22505 6874 22791 6875
rect 23722 6856 23751 7541
rect 24163 7474 24195 8283
rect 24471 8248 24497 8283
rect 24256 8242 24291 8243
rect 24235 8235 24291 8242
rect 24235 8215 24264 8235
rect 24284 8215 24291 8235
rect 24235 8210 24291 8215
rect 24467 8239 24503 8248
rect 24467 8222 24475 8239
rect 24494 8222 24503 8239
rect 24467 8213 24503 8222
rect 25132 8230 25166 8436
rect 26905 8433 26940 8440
rect 25200 8409 25785 8415
rect 25200 8389 25216 8409
rect 25236 8408 25785 8409
rect 25236 8389 25756 8408
rect 25200 8388 25756 8389
rect 25776 8388 25785 8408
rect 25200 8380 25785 8388
rect 26905 8413 26913 8433
rect 26933 8413 26940 8433
rect 26905 8340 26940 8413
rect 27119 8435 27175 8440
rect 27119 8415 27126 8435
rect 27146 8415 27175 8435
rect 27119 8408 27175 8415
rect 27210 8542 27240 8544
rect 27939 8542 27972 8543
rect 27210 8516 27973 8542
rect 27119 8407 27154 8408
rect 27210 8341 27240 8516
rect 27939 8495 27973 8516
rect 27938 8490 27973 8495
rect 27938 8470 27945 8490
rect 27965 8470 27973 8490
rect 27938 8462 27973 8470
rect 27205 8340 27240 8341
rect 26904 8313 27240 8340
rect 27210 8312 27240 8313
rect 27320 8304 27905 8312
rect 27320 8284 27329 8304
rect 27349 8303 27905 8304
rect 27349 8284 27869 8303
rect 27320 8283 27869 8284
rect 27889 8283 27905 8303
rect 27320 8277 27905 8283
rect 27144 8267 27176 8268
rect 27141 8262 27176 8267
rect 27141 8242 27148 8262
rect 27168 8242 27176 8262
rect 27939 8256 27973 8462
rect 28711 8426 28745 8632
rect 29508 8626 29516 8646
rect 29536 8626 29543 8646
rect 29508 8621 29543 8626
rect 29508 8620 29540 8621
rect 28779 8605 29364 8611
rect 28779 8585 28795 8605
rect 28815 8604 29364 8605
rect 28815 8585 29335 8604
rect 28779 8584 29335 8585
rect 29355 8584 29364 8604
rect 28779 8576 29364 8584
rect 29444 8575 29474 8576
rect 29444 8548 29780 8575
rect 29444 8547 29479 8548
rect 28711 8418 28746 8426
rect 28711 8398 28719 8418
rect 28739 8398 28746 8418
rect 28711 8393 28746 8398
rect 28711 8372 28745 8393
rect 29444 8372 29474 8547
rect 29530 8480 29565 8481
rect 28711 8346 29474 8372
rect 28712 8345 28745 8346
rect 29444 8344 29474 8346
rect 29509 8473 29565 8480
rect 29509 8453 29538 8473
rect 29558 8453 29565 8473
rect 29509 8448 29565 8453
rect 29744 8475 29779 8548
rect 29744 8455 29751 8475
rect 29771 8455 29779 8475
rect 30886 8501 31471 8509
rect 30886 8481 30895 8501
rect 30915 8500 31471 8501
rect 30915 8481 31435 8500
rect 30886 8480 31435 8481
rect 31455 8480 31471 8500
rect 30886 8474 31471 8480
rect 29744 8448 29779 8455
rect 31505 8453 31539 8659
rect 33075 8670 33131 8677
rect 33075 8650 33104 8670
rect 33124 8650 33131 8670
rect 33075 8645 33131 8650
rect 33308 8673 33342 8680
rect 33308 8655 33316 8673
rect 33335 8655 33342 8673
rect 33308 8647 33342 8655
rect 33872 8667 33906 8873
rect 34112 8872 34151 8876
rect 33940 8846 34525 8852
rect 33940 8826 33956 8846
rect 33976 8845 34525 8846
rect 33976 8826 34496 8845
rect 33940 8825 34496 8826
rect 34516 8825 34525 8845
rect 33940 8817 34525 8825
rect 33872 8659 33907 8667
rect 27141 8234 27176 8242
rect 25132 8222 25167 8230
rect 24235 8004 24269 8210
rect 25132 8202 25140 8222
rect 25160 8202 25167 8222
rect 25132 8197 25167 8202
rect 25132 8196 25164 8197
rect 24303 8183 24888 8189
rect 24303 8163 24319 8183
rect 24339 8182 24888 8183
rect 24339 8163 24859 8182
rect 24303 8162 24859 8163
rect 24879 8162 24888 8182
rect 24303 8154 24888 8162
rect 26523 8076 27108 8084
rect 26523 8056 26532 8076
rect 26552 8075 27108 8076
rect 26552 8056 27072 8075
rect 26523 8055 27072 8056
rect 27092 8055 27108 8075
rect 26523 8049 27108 8055
rect 26897 8025 26936 8029
rect 27142 8028 27176 8234
rect 27705 8249 27740 8255
rect 27705 8230 27710 8249
rect 27731 8230 27740 8249
rect 27705 8221 27740 8230
rect 27917 8251 27973 8256
rect 27917 8231 27924 8251
rect 27944 8231 27973 8251
rect 27917 8224 27973 8231
rect 28540 8295 28874 8323
rect 27917 8223 27952 8224
rect 27709 8153 27738 8221
rect 27709 8119 28055 8153
rect 26897 8005 26905 8025
rect 26925 8005 26936 8025
rect 24235 7996 24270 8004
rect 24235 7976 24243 7996
rect 24263 7988 24270 7996
rect 24263 7976 24274 7988
rect 24235 7739 24274 7976
rect 25105 7953 25391 7954
rect 24590 7945 25393 7953
rect 24590 7928 24601 7945
rect 24591 7923 24601 7928
rect 24625 7928 25393 7945
rect 24625 7923 24630 7928
rect 24591 7910 24630 7923
rect 25135 7862 25170 7863
rect 25114 7855 25170 7862
rect 25114 7835 25143 7855
rect 25163 7835 25170 7855
rect 25114 7830 25170 7835
rect 25354 7853 25393 7928
rect 26897 7930 26936 8005
rect 27120 8023 27176 8028
rect 27120 8003 27127 8023
rect 27147 8003 27176 8023
rect 27120 7996 27176 8003
rect 27120 7995 27155 7996
rect 27660 7935 27699 7948
rect 27660 7930 27665 7935
rect 26897 7913 27665 7930
rect 27689 7930 27699 7935
rect 27689 7913 27700 7930
rect 26897 7905 27700 7913
rect 26899 7904 27185 7905
rect 28016 7882 28055 8119
rect 28016 7870 28027 7882
rect 28020 7862 28027 7870
rect 28047 7862 28055 7882
rect 28020 7854 28055 7862
rect 25354 7833 25365 7853
rect 25385 7833 25393 7853
rect 24235 7705 24581 7739
rect 24552 7637 24581 7705
rect 24338 7634 24373 7635
rect 24163 7456 24166 7474
rect 24188 7456 24195 7474
rect 24163 7444 24195 7456
rect 24317 7627 24373 7634
rect 24317 7607 24346 7627
rect 24366 7607 24373 7627
rect 24317 7602 24373 7607
rect 24550 7628 24585 7637
rect 24550 7609 24559 7628
rect 24580 7609 24585 7628
rect 24550 7603 24585 7609
rect 25114 7624 25148 7830
rect 25354 7829 25393 7833
rect 25182 7803 25767 7809
rect 25182 7783 25198 7803
rect 25218 7802 25767 7803
rect 25218 7783 25738 7802
rect 25182 7782 25738 7783
rect 25758 7782 25767 7802
rect 25182 7774 25767 7782
rect 27402 7696 27987 7704
rect 27402 7676 27411 7696
rect 27431 7695 27987 7696
rect 27431 7676 27951 7695
rect 27402 7675 27951 7676
rect 27971 7675 27987 7695
rect 27402 7669 27987 7675
rect 27126 7661 27158 7662
rect 27123 7656 27158 7661
rect 27123 7636 27130 7656
rect 27150 7636 27158 7656
rect 28021 7648 28055 7854
rect 27123 7628 27158 7636
rect 25114 7616 25149 7624
rect 24317 7396 24351 7602
rect 25114 7596 25122 7616
rect 25142 7596 25149 7616
rect 25114 7591 25149 7596
rect 25114 7590 25146 7591
rect 24385 7575 24970 7581
rect 24385 7555 24401 7575
rect 24421 7574 24970 7575
rect 24421 7555 24941 7574
rect 24385 7554 24941 7555
rect 24961 7554 24970 7574
rect 24385 7546 24970 7554
rect 25050 7545 25080 7546
rect 25050 7518 25386 7545
rect 25050 7517 25085 7518
rect 24317 7388 24352 7396
rect 24317 7368 24325 7388
rect 24345 7368 24352 7388
rect 24317 7363 24352 7368
rect 24317 7342 24351 7363
rect 25050 7342 25080 7517
rect 25136 7450 25171 7451
rect 24317 7316 25080 7342
rect 24318 7315 24351 7316
rect 25050 7314 25080 7316
rect 25115 7443 25171 7450
rect 25115 7423 25144 7443
rect 25164 7423 25171 7443
rect 25115 7418 25171 7423
rect 25350 7445 25385 7518
rect 25350 7425 25357 7445
rect 25377 7425 25385 7445
rect 26505 7470 27090 7478
rect 26505 7450 26514 7470
rect 26534 7469 27090 7470
rect 26534 7450 27054 7469
rect 26505 7449 27054 7450
rect 27074 7449 27090 7469
rect 26505 7443 27090 7449
rect 25350 7418 25385 7425
rect 27124 7422 27158 7628
rect 27789 7642 27820 7648
rect 27789 7623 27794 7642
rect 27815 7623 27820 7642
rect 27789 7581 27820 7623
rect 27999 7643 28055 7648
rect 27999 7623 28006 7643
rect 28026 7623 28055 7643
rect 27999 7616 28055 7623
rect 27999 7615 28034 7616
rect 27789 7553 28128 7581
rect 23955 7282 24418 7290
rect 23955 7260 23967 7282
rect 23991 7260 24418 7282
rect 23955 7259 24418 7260
rect 23957 7247 23996 7259
rect 24391 7228 24418 7259
rect 24173 7226 24208 7227
rect 24152 7219 24208 7226
rect 24152 7199 24181 7219
rect 24201 7199 24208 7219
rect 24152 7194 24208 7199
rect 24387 7219 24420 7228
rect 24387 7197 24392 7219
rect 24415 7197 24420 7219
rect 24152 6988 24186 7194
rect 24387 7191 24420 7197
rect 25115 7212 25149 7418
rect 26888 7415 26923 7422
rect 25183 7391 25768 7397
rect 25183 7371 25199 7391
rect 25219 7390 25768 7391
rect 25219 7371 25739 7390
rect 25183 7370 25739 7371
rect 25759 7370 25768 7390
rect 25183 7362 25768 7370
rect 26888 7395 26896 7415
rect 26916 7395 26923 7415
rect 26888 7322 26923 7395
rect 27102 7417 27158 7422
rect 27102 7397 27109 7417
rect 27129 7397 27158 7417
rect 27102 7390 27158 7397
rect 27193 7524 27223 7526
rect 27922 7524 27955 7525
rect 27193 7498 27956 7524
rect 27102 7389 27137 7390
rect 27193 7323 27223 7498
rect 27922 7477 27956 7498
rect 27921 7472 27956 7477
rect 27921 7452 27928 7472
rect 27948 7452 27956 7472
rect 27921 7444 27956 7452
rect 27188 7322 27223 7323
rect 26887 7295 27223 7322
rect 27193 7294 27223 7295
rect 27303 7286 27888 7294
rect 27303 7266 27312 7286
rect 27332 7285 27888 7286
rect 27332 7266 27852 7285
rect 27303 7265 27852 7266
rect 27872 7265 27888 7285
rect 27303 7259 27888 7265
rect 27127 7249 27159 7250
rect 27124 7244 27159 7249
rect 27124 7224 27131 7244
rect 27151 7224 27159 7244
rect 27922 7238 27956 7444
rect 27124 7216 27159 7224
rect 25115 7204 25150 7212
rect 25115 7184 25123 7204
rect 25143 7184 25150 7204
rect 25115 7179 25150 7184
rect 25115 7178 25147 7179
rect 24220 7167 24805 7173
rect 24220 7147 24236 7167
rect 24256 7166 24805 7167
rect 24256 7147 24776 7166
rect 24220 7146 24776 7147
rect 24796 7146 24805 7166
rect 24220 7138 24805 7146
rect 26506 7058 27091 7066
rect 26506 7038 26515 7058
rect 26535 7057 27091 7058
rect 26535 7038 27055 7057
rect 26506 7037 27055 7038
rect 27075 7037 27091 7057
rect 26506 7031 27091 7037
rect 26880 7007 26919 7011
rect 27125 7010 27159 7216
rect 27689 7228 27723 7236
rect 27689 7210 27696 7228
rect 27715 7210 27723 7228
rect 27689 7203 27723 7210
rect 27900 7233 27956 7238
rect 27900 7213 27907 7233
rect 27927 7213 27956 7233
rect 27900 7206 27956 7213
rect 27900 7205 27935 7206
rect 27693 7173 27722 7203
rect 27693 7165 28075 7173
rect 27693 7146 28046 7165
rect 28067 7146 28075 7165
rect 27693 7141 28075 7146
rect 24152 6987 24187 6988
rect 24120 6980 24187 6987
rect 24120 6960 24160 6980
rect 24180 6960 24187 6980
rect 24120 6957 24187 6960
rect 26880 6987 26888 7007
rect 26908 6987 26919 7007
rect 24120 6954 24185 6957
rect 23691 6853 23756 6856
rect 23689 6850 23756 6853
rect 23689 6830 23696 6850
rect 23716 6830 23756 6850
rect 23689 6823 23756 6830
rect 23689 6822 23724 6823
rect 20970 6802 20981 6822
rect 21001 6802 21009 6822
rect 19814 6663 20196 6668
rect 19814 6644 19822 6663
rect 19843 6644 20196 6663
rect 19814 6636 20196 6644
rect 20167 6606 20196 6636
rect 19954 6603 19989 6604
rect 19933 6596 19989 6603
rect 19933 6576 19962 6596
rect 19982 6576 19989 6596
rect 19933 6571 19989 6576
rect 20166 6599 20200 6606
rect 20166 6581 20174 6599
rect 20193 6581 20200 6599
rect 20166 6573 20200 6581
rect 20730 6593 20764 6799
rect 20970 6798 21009 6802
rect 20798 6772 21383 6778
rect 20798 6752 20814 6772
rect 20834 6771 21383 6772
rect 20834 6752 21354 6771
rect 20798 6751 21354 6752
rect 21374 6751 21383 6771
rect 20798 6743 21383 6751
rect 23071 6664 23656 6672
rect 23071 6644 23080 6664
rect 23100 6663 23656 6664
rect 23100 6644 23620 6663
rect 23071 6643 23620 6644
rect 23640 6643 23656 6663
rect 23071 6637 23656 6643
rect 22729 6631 22761 6632
rect 22726 6626 22761 6631
rect 22726 6606 22733 6626
rect 22753 6606 22761 6626
rect 22726 6598 22761 6606
rect 20730 6585 20765 6593
rect 19933 6365 19967 6571
rect 20730 6565 20738 6585
rect 20758 6565 20765 6585
rect 20730 6560 20765 6565
rect 20730 6559 20762 6560
rect 20001 6544 20586 6550
rect 20001 6524 20017 6544
rect 20037 6543 20586 6544
rect 20037 6524 20557 6543
rect 20001 6523 20557 6524
rect 20577 6523 20586 6543
rect 20001 6515 20586 6523
rect 20666 6514 20696 6515
rect 20666 6487 21002 6514
rect 20666 6486 20701 6487
rect 19933 6357 19968 6365
rect 19933 6337 19941 6357
rect 19961 6337 19968 6357
rect 19933 6332 19968 6337
rect 19933 6311 19967 6332
rect 20666 6311 20696 6486
rect 20752 6419 20787 6420
rect 19933 6285 20696 6311
rect 19934 6284 19967 6285
rect 20666 6283 20696 6285
rect 20731 6412 20787 6419
rect 20731 6392 20760 6412
rect 20780 6392 20787 6412
rect 20731 6387 20787 6392
rect 20966 6414 21001 6487
rect 20966 6394 20973 6414
rect 20993 6394 21001 6414
rect 22108 6440 22693 6448
rect 22108 6420 22117 6440
rect 22137 6439 22693 6440
rect 22137 6420 22657 6439
rect 22108 6419 22657 6420
rect 22677 6419 22693 6439
rect 22108 6413 22693 6419
rect 20966 6387 21001 6394
rect 22727 6392 22761 6598
rect 23454 6608 23495 6619
rect 23690 6616 23724 6822
rect 23454 6590 23464 6608
rect 23482 6590 23495 6608
rect 23454 6582 23495 6590
rect 23668 6611 23724 6616
rect 23668 6591 23675 6611
rect 23695 6591 23724 6611
rect 23668 6584 23724 6591
rect 23668 6583 23703 6584
rect 23463 6552 23489 6582
rect 23463 6551 23801 6552
rect 23463 6515 23817 6551
rect 19761 6228 20100 6256
rect 19855 6193 19890 6194
rect 19834 6186 19890 6193
rect 19834 6166 19863 6186
rect 19883 6166 19890 6186
rect 19834 6161 19890 6166
rect 20069 6186 20100 6228
rect 20069 6167 20074 6186
rect 20095 6167 20100 6186
rect 20069 6161 20100 6167
rect 20731 6181 20765 6387
rect 22491 6385 22526 6392
rect 20799 6360 21384 6366
rect 20799 6340 20815 6360
rect 20835 6359 21384 6360
rect 20835 6340 21355 6359
rect 20799 6339 21355 6340
rect 21375 6339 21384 6359
rect 20799 6331 21384 6339
rect 22491 6365 22499 6385
rect 22519 6365 22526 6385
rect 22491 6292 22526 6365
rect 22705 6387 22761 6392
rect 22705 6367 22712 6387
rect 22732 6367 22761 6387
rect 22705 6360 22761 6367
rect 22796 6494 22826 6496
rect 23525 6494 23558 6495
rect 22796 6468 23559 6494
rect 22705 6359 22740 6360
rect 22796 6293 22826 6468
rect 23525 6447 23559 6468
rect 23524 6442 23559 6447
rect 23524 6422 23531 6442
rect 23551 6422 23559 6442
rect 23524 6414 23559 6422
rect 22791 6292 22826 6293
rect 22490 6265 22826 6292
rect 22796 6264 22826 6265
rect 22906 6256 23491 6264
rect 22906 6236 22915 6256
rect 22935 6255 23491 6256
rect 22935 6236 23455 6255
rect 22906 6235 23455 6236
rect 23475 6235 23491 6255
rect 22906 6229 23491 6235
rect 22730 6219 22762 6220
rect 22727 6214 22762 6219
rect 22727 6194 22734 6214
rect 22754 6194 22762 6214
rect 23525 6208 23559 6414
rect 22727 6186 22762 6194
rect 20731 6173 20766 6181
rect 19834 5955 19868 6161
rect 20731 6153 20739 6173
rect 20759 6153 20766 6173
rect 20731 6148 20766 6153
rect 20731 6147 20763 6148
rect 19902 6134 20487 6140
rect 19902 6114 19918 6134
rect 19938 6133 20487 6134
rect 19938 6114 20458 6133
rect 19902 6113 20458 6114
rect 20478 6113 20487 6133
rect 19902 6105 20487 6113
rect 22109 6028 22694 6036
rect 22109 6008 22118 6028
rect 22138 6027 22694 6028
rect 22138 6008 22658 6027
rect 22109 6007 22658 6008
rect 22678 6007 22694 6027
rect 22109 6001 22694 6007
rect 22483 5977 22522 5981
rect 22728 5980 22762 6186
rect 23291 6201 23326 6207
rect 23291 6182 23296 6201
rect 23317 6182 23326 6201
rect 23291 6173 23326 6182
rect 23503 6203 23559 6208
rect 23503 6183 23510 6203
rect 23530 6183 23559 6203
rect 23503 6176 23559 6183
rect 23503 6175 23538 6176
rect 23295 6105 23324 6173
rect 23295 6071 23641 6105
rect 22483 5957 22491 5977
rect 22511 5957 22522 5977
rect 19834 5947 19869 5955
rect 19834 5927 19842 5947
rect 19862 5939 19869 5947
rect 19862 5927 19873 5939
rect 19834 5690 19873 5927
rect 20704 5904 20990 5905
rect 20189 5896 20992 5904
rect 20189 5879 20200 5896
rect 20190 5874 20200 5879
rect 20224 5879 20992 5896
rect 20224 5874 20229 5879
rect 20190 5861 20229 5874
rect 20734 5813 20769 5814
rect 20713 5806 20769 5813
rect 20713 5786 20742 5806
rect 20762 5786 20769 5806
rect 20713 5781 20769 5786
rect 20953 5804 20992 5879
rect 22483 5882 22522 5957
rect 22706 5975 22762 5980
rect 22706 5955 22713 5975
rect 22733 5955 22762 5975
rect 22706 5948 22762 5955
rect 22706 5947 22741 5948
rect 23246 5887 23285 5900
rect 23246 5882 23251 5887
rect 22483 5865 23251 5882
rect 23275 5882 23285 5887
rect 23275 5865 23286 5882
rect 22483 5857 23286 5865
rect 22485 5856 22771 5857
rect 23602 5834 23641 6071
rect 23602 5822 23613 5834
rect 23606 5814 23613 5822
rect 23633 5814 23641 5834
rect 23606 5806 23641 5814
rect 20953 5784 20964 5804
rect 20984 5784 20992 5804
rect 19834 5656 20180 5690
rect 20151 5588 20180 5656
rect 19937 5585 19972 5586
rect 19916 5578 19972 5585
rect 19916 5558 19945 5578
rect 19965 5558 19972 5578
rect 19916 5553 19972 5558
rect 20149 5579 20184 5588
rect 20149 5560 20158 5579
rect 20179 5560 20184 5579
rect 20149 5554 20184 5560
rect 20713 5575 20747 5781
rect 20953 5780 20992 5784
rect 20781 5754 21366 5760
rect 20781 5734 20797 5754
rect 20817 5753 21366 5754
rect 20817 5734 21337 5753
rect 20781 5733 21337 5734
rect 21357 5733 21366 5753
rect 20781 5725 21366 5733
rect 22988 5648 23573 5656
rect 22988 5628 22997 5648
rect 23017 5647 23573 5648
rect 23017 5628 23537 5647
rect 22988 5627 23537 5628
rect 23557 5627 23573 5647
rect 22988 5621 23573 5627
rect 22712 5613 22744 5614
rect 22709 5608 22744 5613
rect 22709 5588 22716 5608
rect 22736 5588 22744 5608
rect 23607 5600 23641 5806
rect 22709 5580 22744 5588
rect 20713 5567 20748 5575
rect 19916 5347 19950 5553
rect 20713 5547 20721 5567
rect 20741 5547 20748 5567
rect 20713 5542 20748 5547
rect 20713 5541 20745 5542
rect 19984 5526 20569 5532
rect 19984 5506 20000 5526
rect 20020 5525 20569 5526
rect 20020 5506 20540 5525
rect 19984 5505 20540 5506
rect 20560 5505 20569 5525
rect 19984 5497 20569 5505
rect 20649 5496 20679 5497
rect 20649 5469 20985 5496
rect 20649 5468 20684 5469
rect 19916 5339 19951 5347
rect 19916 5319 19924 5339
rect 19944 5319 19951 5339
rect 19916 5314 19951 5319
rect 19916 5293 19950 5314
rect 20649 5293 20679 5468
rect 20735 5401 20770 5402
rect 19916 5267 20679 5293
rect 19917 5266 19950 5267
rect 20649 5265 20679 5267
rect 20714 5394 20770 5401
rect 20714 5374 20743 5394
rect 20763 5374 20770 5394
rect 20714 5369 20770 5374
rect 20949 5396 20984 5469
rect 20949 5376 20956 5396
rect 20976 5376 20984 5396
rect 22091 5422 22676 5430
rect 22091 5402 22100 5422
rect 22120 5421 22676 5422
rect 22120 5402 22640 5421
rect 22091 5401 22640 5402
rect 22660 5401 22676 5421
rect 22091 5395 22676 5401
rect 20949 5369 20984 5376
rect 22710 5374 22744 5580
rect 23373 5588 23409 5597
rect 23373 5571 23382 5588
rect 23401 5571 23409 5588
rect 23373 5562 23409 5571
rect 23585 5595 23641 5600
rect 23585 5575 23592 5595
rect 23612 5575 23641 5595
rect 23585 5568 23641 5575
rect 23585 5567 23620 5568
rect 23379 5527 23405 5562
rect 23687 5527 23719 5528
rect 23379 5522 23719 5527
rect 23379 5504 23694 5522
rect 23716 5504 23719 5522
rect 23379 5499 23719 5504
rect 23687 5498 23719 5499
rect 19568 5246 19885 5249
rect 19568 5219 19571 5246
rect 19598 5219 19885 5246
rect 19568 5213 19885 5219
rect 19568 5210 19604 5213
rect 19849 5183 19885 5213
rect 19633 5179 19668 5180
rect 19612 5172 19668 5179
rect 19612 5152 19641 5172
rect 19661 5152 19668 5172
rect 19612 5147 19668 5152
rect 19847 5177 19885 5183
rect 19847 5151 19853 5177
rect 19879 5151 19885 5177
rect 19612 4948 19646 5147
rect 19847 5143 19885 5151
rect 20714 5163 20748 5369
rect 22474 5367 22509 5374
rect 20782 5342 21367 5348
rect 20782 5322 20798 5342
rect 20818 5341 21367 5342
rect 20818 5322 21338 5341
rect 20782 5321 21338 5322
rect 21358 5321 21367 5341
rect 20782 5313 21367 5321
rect 22474 5347 22482 5367
rect 22502 5347 22509 5367
rect 22474 5274 22509 5347
rect 22688 5369 22744 5374
rect 22688 5349 22695 5369
rect 22715 5349 22744 5369
rect 22688 5342 22744 5349
rect 22779 5476 22809 5478
rect 23508 5476 23541 5477
rect 22779 5450 23542 5476
rect 22688 5341 22723 5342
rect 22779 5275 22809 5450
rect 23508 5429 23542 5450
rect 23507 5424 23542 5429
rect 23507 5404 23514 5424
rect 23534 5404 23542 5424
rect 23507 5396 23542 5404
rect 22774 5274 22809 5275
rect 22473 5247 22809 5274
rect 22779 5246 22809 5247
rect 22889 5238 23474 5246
rect 22889 5218 22898 5238
rect 22918 5237 23474 5238
rect 22918 5218 23438 5237
rect 22889 5217 23438 5218
rect 23458 5217 23474 5237
rect 22889 5211 23474 5217
rect 22713 5201 22745 5202
rect 22710 5196 22745 5201
rect 22710 5176 22717 5196
rect 22737 5176 22745 5196
rect 23508 5190 23542 5396
rect 22710 5168 22745 5176
rect 20714 5155 20749 5163
rect 20714 5135 20722 5155
rect 20742 5135 20749 5155
rect 20714 5130 20749 5135
rect 20714 5129 20746 5130
rect 19680 5120 20265 5126
rect 19680 5100 19696 5120
rect 19716 5119 20265 5120
rect 19716 5100 20236 5119
rect 19680 5099 20236 5100
rect 20256 5099 20265 5119
rect 19680 5091 20265 5099
rect 22092 5010 22677 5018
rect 22092 4990 22101 5010
rect 22121 5009 22677 5010
rect 22121 4990 22641 5009
rect 22092 4989 22641 4990
rect 22661 4989 22677 5009
rect 22092 4983 22677 4989
rect 22466 4959 22505 4963
rect 22711 4962 22745 5168
rect 23275 5180 23309 5188
rect 23275 5162 23282 5180
rect 23301 5162 23309 5180
rect 23275 5155 23309 5162
rect 23486 5185 23542 5190
rect 23486 5165 23493 5185
rect 23513 5165 23542 5185
rect 23486 5158 23542 5165
rect 23486 5157 23521 5158
rect 23279 5125 23308 5155
rect 23279 5117 23661 5125
rect 23279 5098 23632 5117
rect 23653 5098 23661 5117
rect 23279 5093 23661 5098
rect 19612 4933 19649 4948
rect 19612 4913 19620 4933
rect 19640 4913 19649 4933
rect 19612 4910 19649 4913
rect 19426 4799 19463 4802
rect 19426 4779 19435 4799
rect 19455 4779 19463 4799
rect 16496 4762 17081 4768
rect 19426 4764 19463 4779
rect 16496 4742 16512 4762
rect 16532 4761 17081 4762
rect 16532 4742 17052 4761
rect 16496 4741 17052 4742
rect 17072 4741 17081 4761
rect 16496 4733 17081 4741
rect 18810 4613 19395 4621
rect 18810 4593 18819 4613
rect 18839 4612 19395 4613
rect 18839 4593 19359 4612
rect 18810 4592 19359 4593
rect 19379 4592 19395 4612
rect 18810 4586 19395 4592
rect 16428 4575 16463 4583
rect 18329 4582 18361 4583
rect 15631 4355 15665 4561
rect 16428 4555 16436 4575
rect 16456 4555 16463 4575
rect 16428 4550 16463 4555
rect 18326 4577 18361 4582
rect 18326 4557 18333 4577
rect 18353 4557 18361 4577
rect 19429 4565 19463 4764
rect 19407 4560 19463 4565
rect 16428 4549 16460 4550
rect 18326 4549 18361 4557
rect 15699 4534 16284 4540
rect 15699 4514 15715 4534
rect 15735 4533 16284 4534
rect 15735 4514 16255 4533
rect 15699 4513 16255 4514
rect 16275 4513 16284 4533
rect 15699 4505 16284 4513
rect 16364 4504 16394 4505
rect 16364 4477 16700 4504
rect 16364 4476 16399 4477
rect 15631 4347 15666 4355
rect 15631 4327 15639 4347
rect 15659 4327 15666 4347
rect 15631 4322 15666 4327
rect 15631 4301 15665 4322
rect 16364 4301 16394 4476
rect 16450 4409 16485 4410
rect 15631 4275 16394 4301
rect 15632 4274 15665 4275
rect 16364 4273 16394 4275
rect 16429 4402 16485 4409
rect 16429 4382 16458 4402
rect 16478 4382 16485 4402
rect 16429 4377 16485 4382
rect 16664 4404 16699 4477
rect 16664 4384 16671 4404
rect 16691 4384 16699 4404
rect 16664 4377 16699 4384
rect 17708 4391 18293 4399
rect 15454 4252 15486 4253
rect 15454 4247 15794 4252
rect 15454 4229 15457 4247
rect 15479 4229 15794 4247
rect 15454 4224 15794 4229
rect 15454 4223 15486 4224
rect 15768 4189 15794 4224
rect 15553 4183 15588 4184
rect 15532 4176 15588 4183
rect 15532 4156 15561 4176
rect 15581 4156 15588 4176
rect 15532 4151 15588 4156
rect 15764 4180 15800 4189
rect 15764 4163 15772 4180
rect 15791 4163 15800 4180
rect 15764 4154 15800 4163
rect 16429 4171 16463 4377
rect 17708 4371 17717 4391
rect 17737 4390 18293 4391
rect 17737 4371 18257 4390
rect 17708 4370 18257 4371
rect 18277 4370 18293 4390
rect 17708 4364 18293 4370
rect 16497 4350 17082 4356
rect 16497 4330 16513 4350
rect 16533 4349 17082 4350
rect 16533 4330 17053 4349
rect 16497 4329 17053 4330
rect 17073 4329 17082 4349
rect 18327 4343 18361 4549
rect 19189 4558 19224 4560
rect 19189 4552 19227 4558
rect 19189 4529 19197 4552
rect 19220 4529 19227 4552
rect 19407 4540 19414 4560
rect 19434 4540 19463 4560
rect 19407 4533 19463 4540
rect 19407 4532 19442 4533
rect 19189 4523 19227 4529
rect 19189 4510 19224 4523
rect 19187 4452 19224 4510
rect 16497 4321 17082 4329
rect 18091 4336 18126 4343
rect 18091 4316 18099 4336
rect 18119 4316 18126 4336
rect 18091 4243 18126 4316
rect 18305 4338 18361 4343
rect 18305 4318 18312 4338
rect 18332 4318 18361 4338
rect 18305 4311 18361 4318
rect 18396 4445 18426 4447
rect 19125 4445 19158 4446
rect 18396 4419 19159 4445
rect 18305 4310 18340 4311
rect 18396 4244 18426 4419
rect 19125 4398 19159 4419
rect 19187 4435 19222 4452
rect 19187 4434 19481 4435
rect 19187 4433 19524 4434
rect 19187 4426 19529 4433
rect 19187 4400 19489 4426
rect 19520 4400 19529 4426
rect 19124 4393 19159 4398
rect 19480 4397 19529 4400
rect 19124 4373 19131 4393
rect 19151 4373 19159 4393
rect 19486 4392 19529 4397
rect 19124 4365 19159 4373
rect 18391 4243 18426 4244
rect 18090 4216 18426 4243
rect 18396 4215 18426 4216
rect 18506 4207 19091 4215
rect 18506 4187 18515 4207
rect 18535 4206 19091 4207
rect 18535 4187 19055 4206
rect 18506 4186 19055 4187
rect 19075 4186 19091 4206
rect 18506 4180 19091 4186
rect 16429 4163 16464 4171
rect 18330 4170 18362 4171
rect 15532 3945 15566 4151
rect 16429 4143 16437 4163
rect 16457 4143 16464 4163
rect 16429 4138 16464 4143
rect 18327 4165 18362 4170
rect 18327 4145 18334 4165
rect 18354 4145 18362 4165
rect 19125 4159 19159 4365
rect 16429 4137 16461 4138
rect 18327 4137 18362 4145
rect 15600 4124 16185 4130
rect 15600 4104 15616 4124
rect 15636 4123 16185 4124
rect 15636 4104 16156 4123
rect 15600 4103 16156 4104
rect 16176 4103 16185 4123
rect 15600 4095 16185 4103
rect 17709 3979 18294 3987
rect 17709 3959 17718 3979
rect 17738 3978 18294 3979
rect 17738 3959 18258 3978
rect 17709 3958 18258 3959
rect 18278 3958 18294 3978
rect 17709 3952 18294 3958
rect 15532 3937 15567 3945
rect 15532 3917 15540 3937
rect 15560 3929 15567 3937
rect 15560 3917 15571 3929
rect 15532 3680 15571 3917
rect 18083 3928 18122 3932
rect 18328 3931 18362 4137
rect 18891 4152 18926 4158
rect 18891 4133 18896 4152
rect 18917 4133 18926 4152
rect 18891 4124 18926 4133
rect 19103 4154 19159 4159
rect 19103 4134 19110 4154
rect 19130 4134 19159 4154
rect 19103 4127 19159 4134
rect 19103 4126 19138 4127
rect 18895 4056 18924 4124
rect 18895 4022 19241 4056
rect 18083 3908 18091 3928
rect 18111 3908 18122 3928
rect 16402 3894 16688 3895
rect 15887 3886 16690 3894
rect 15887 3869 15898 3886
rect 15888 3864 15898 3869
rect 15922 3869 16690 3886
rect 15922 3864 15927 3869
rect 15888 3851 15927 3864
rect 16432 3803 16467 3804
rect 16411 3796 16467 3803
rect 16411 3776 16440 3796
rect 16460 3776 16467 3796
rect 16411 3771 16467 3776
rect 16651 3794 16690 3869
rect 18083 3833 18122 3908
rect 18306 3926 18362 3931
rect 18306 3906 18313 3926
rect 18333 3906 18362 3926
rect 18306 3899 18362 3906
rect 18306 3898 18341 3899
rect 18846 3838 18885 3851
rect 18846 3833 18851 3838
rect 18083 3816 18851 3833
rect 18875 3833 18885 3838
rect 18875 3816 18886 3833
rect 18083 3808 18886 3816
rect 18085 3807 18371 3808
rect 16651 3774 16662 3794
rect 16682 3774 16690 3794
rect 15532 3646 15878 3680
rect 15849 3578 15878 3646
rect 15635 3575 15670 3576
rect 15614 3568 15670 3575
rect 15614 3548 15643 3568
rect 15663 3548 15670 3568
rect 15614 3543 15670 3548
rect 15847 3569 15882 3578
rect 15847 3550 15856 3569
rect 15877 3550 15882 3569
rect 15847 3544 15882 3550
rect 16411 3565 16445 3771
rect 16651 3770 16690 3774
rect 19202 3785 19241 4022
rect 19202 3773 19213 3785
rect 19206 3765 19213 3773
rect 19233 3765 19241 3785
rect 19206 3757 19241 3765
rect 16479 3744 17064 3750
rect 16479 3724 16495 3744
rect 16515 3743 17064 3744
rect 16515 3724 17035 3743
rect 16479 3723 17035 3724
rect 17055 3723 17064 3743
rect 16479 3715 17064 3723
rect 18588 3599 19173 3607
rect 18588 3579 18597 3599
rect 18617 3598 19173 3599
rect 18617 3579 19137 3598
rect 18588 3578 19137 3579
rect 19157 3578 19173 3598
rect 18588 3572 19173 3578
rect 16411 3557 16446 3565
rect 18312 3564 18344 3565
rect 15614 3337 15648 3543
rect 16411 3537 16419 3557
rect 16439 3537 16446 3557
rect 16411 3532 16446 3537
rect 18309 3559 18344 3564
rect 18309 3539 18316 3559
rect 18336 3539 18344 3559
rect 19207 3551 19241 3757
rect 16411 3531 16443 3532
rect 18309 3531 18344 3539
rect 15682 3516 16267 3522
rect 15682 3496 15698 3516
rect 15718 3515 16267 3516
rect 15718 3496 16238 3515
rect 15682 3495 16238 3496
rect 16258 3495 16267 3515
rect 15682 3487 16267 3495
rect 16347 3486 16377 3487
rect 16347 3459 16683 3486
rect 16347 3458 16382 3459
rect 15614 3329 15649 3337
rect 15614 3309 15622 3329
rect 15642 3309 15649 3329
rect 15614 3304 15649 3309
rect 15614 3283 15648 3304
rect 16347 3283 16377 3458
rect 16433 3391 16468 3392
rect 15614 3257 16377 3283
rect 15615 3256 15648 3257
rect 16347 3255 16377 3257
rect 16412 3384 16468 3391
rect 16412 3364 16441 3384
rect 16461 3364 16468 3384
rect 16412 3359 16468 3364
rect 16647 3386 16682 3459
rect 16647 3366 16654 3386
rect 16674 3366 16682 3386
rect 16647 3359 16682 3366
rect 17691 3373 18276 3381
rect 15356 3200 15710 3236
rect 15372 3199 15710 3200
rect 15684 3169 15710 3199
rect 15470 3167 15505 3168
rect 15449 3160 15505 3167
rect 15449 3140 15478 3160
rect 15498 3140 15505 3160
rect 15449 3135 15505 3140
rect 15678 3161 15719 3169
rect 15678 3143 15691 3161
rect 15709 3143 15719 3161
rect 15449 2929 15483 3135
rect 15678 3132 15719 3143
rect 16412 3153 16446 3359
rect 17691 3353 17700 3373
rect 17720 3372 18276 3373
rect 17720 3353 18240 3372
rect 17691 3352 18240 3353
rect 18260 3352 18276 3372
rect 17691 3346 18276 3352
rect 16480 3332 17065 3338
rect 16480 3312 16496 3332
rect 16516 3331 17065 3332
rect 16516 3312 17036 3331
rect 16480 3311 17036 3312
rect 17056 3311 17065 3331
rect 18310 3325 18344 3531
rect 18975 3545 19006 3551
rect 18975 3526 18980 3545
rect 19001 3526 19006 3545
rect 18975 3484 19006 3526
rect 19185 3546 19241 3551
rect 19185 3526 19192 3546
rect 19212 3526 19241 3546
rect 19185 3519 19241 3526
rect 19185 3518 19220 3519
rect 18975 3456 19314 3484
rect 16480 3303 17065 3311
rect 18074 3318 18109 3325
rect 18074 3298 18082 3318
rect 18102 3298 18109 3318
rect 18074 3225 18109 3298
rect 18288 3320 18344 3325
rect 18288 3300 18295 3320
rect 18315 3300 18344 3320
rect 18288 3293 18344 3300
rect 18379 3427 18409 3429
rect 19108 3427 19141 3428
rect 18379 3401 19142 3427
rect 18288 3292 18323 3293
rect 18379 3226 18409 3401
rect 19108 3380 19142 3401
rect 19107 3375 19142 3380
rect 19107 3355 19114 3375
rect 19134 3355 19142 3375
rect 19107 3347 19142 3355
rect 18374 3225 18409 3226
rect 18073 3198 18409 3225
rect 18379 3197 18409 3198
rect 18489 3189 19074 3197
rect 18489 3169 18498 3189
rect 18518 3188 19074 3189
rect 18518 3169 19038 3188
rect 18489 3168 19038 3169
rect 19058 3168 19074 3188
rect 18489 3162 19074 3168
rect 16412 3145 16447 3153
rect 18313 3152 18345 3153
rect 16412 3125 16420 3145
rect 16440 3125 16447 3145
rect 16412 3120 16447 3125
rect 18310 3147 18345 3152
rect 18310 3127 18317 3147
rect 18337 3127 18345 3147
rect 19108 3141 19142 3347
rect 16412 3119 16444 3120
rect 18310 3119 18345 3127
rect 15517 3108 16102 3114
rect 15517 3088 15533 3108
rect 15553 3107 16102 3108
rect 15553 3088 16073 3107
rect 15517 3087 16073 3088
rect 16093 3087 16102 3107
rect 15517 3079 16102 3087
rect 17692 2961 18277 2969
rect 17692 2941 17701 2961
rect 17721 2960 18277 2961
rect 17721 2941 18241 2960
rect 17692 2940 18241 2941
rect 18261 2940 18277 2960
rect 17692 2934 18277 2940
rect 15449 2928 15484 2929
rect 15417 2921 15484 2928
rect 15417 2901 15457 2921
rect 15477 2901 15484 2921
rect 15417 2898 15484 2901
rect 18066 2910 18105 2914
rect 18311 2913 18345 3119
rect 18875 3131 18909 3139
rect 18875 3113 18882 3131
rect 18901 3113 18909 3131
rect 18875 3106 18909 3113
rect 19086 3136 19142 3141
rect 19086 3116 19093 3136
rect 19113 3116 19142 3136
rect 19086 3109 19142 3116
rect 19086 3108 19121 3109
rect 18879 3076 18908 3106
rect 18879 3068 19261 3076
rect 18879 3049 19232 3068
rect 19253 3049 19261 3068
rect 18879 3044 19261 3049
rect 15417 2895 15482 2898
rect 14988 2794 15053 2797
rect 14986 2791 15053 2794
rect 14986 2771 14993 2791
rect 15013 2771 15053 2791
rect 14986 2764 15053 2771
rect 14986 2763 15021 2764
rect 12267 2743 12278 2763
rect 12298 2743 12306 2763
rect 11111 2604 11493 2609
rect 11111 2585 11119 2604
rect 11140 2585 11493 2604
rect 11111 2577 11493 2585
rect 11464 2547 11493 2577
rect 11251 2544 11286 2545
rect 11230 2537 11286 2544
rect 11230 2517 11259 2537
rect 11279 2517 11286 2537
rect 11230 2512 11286 2517
rect 11463 2540 11497 2547
rect 11463 2522 11471 2540
rect 11490 2522 11497 2540
rect 11463 2514 11497 2522
rect 12027 2534 12061 2740
rect 12267 2739 12306 2743
rect 12095 2713 12680 2719
rect 12095 2693 12111 2713
rect 12131 2712 12680 2713
rect 12131 2693 12651 2712
rect 12095 2692 12651 2693
rect 12671 2692 12680 2712
rect 12095 2684 12680 2692
rect 14368 2605 14953 2613
rect 14368 2585 14377 2605
rect 14397 2604 14953 2605
rect 14397 2585 14917 2604
rect 14368 2584 14917 2585
rect 14937 2584 14953 2604
rect 14368 2578 14953 2584
rect 14026 2572 14058 2573
rect 14023 2567 14058 2572
rect 14023 2547 14030 2567
rect 14050 2547 14058 2567
rect 14023 2539 14058 2547
rect 12027 2526 12062 2534
rect 11230 2306 11264 2512
rect 12027 2506 12035 2526
rect 12055 2506 12062 2526
rect 12027 2501 12062 2506
rect 12027 2500 12059 2501
rect 11298 2485 11883 2491
rect 11298 2465 11314 2485
rect 11334 2484 11883 2485
rect 11334 2465 11854 2484
rect 11298 2464 11854 2465
rect 11874 2464 11883 2484
rect 11298 2456 11883 2464
rect 11963 2455 11993 2456
rect 11963 2428 12299 2455
rect 11963 2427 11998 2428
rect 11230 2298 11265 2306
rect 11230 2278 11238 2298
rect 11258 2278 11265 2298
rect 11230 2273 11265 2278
rect 11230 2252 11264 2273
rect 11963 2252 11993 2427
rect 12049 2360 12084 2361
rect 11230 2226 11993 2252
rect 11231 2225 11264 2226
rect 11963 2224 11993 2226
rect 12028 2353 12084 2360
rect 12028 2333 12057 2353
rect 12077 2333 12084 2353
rect 12028 2328 12084 2333
rect 12263 2355 12298 2428
rect 12263 2335 12270 2355
rect 12290 2335 12298 2355
rect 13405 2381 13990 2389
rect 13405 2361 13414 2381
rect 13434 2380 13990 2381
rect 13434 2361 13954 2380
rect 13405 2360 13954 2361
rect 13974 2360 13990 2380
rect 13405 2354 13990 2360
rect 12263 2328 12298 2335
rect 14024 2333 14058 2539
rect 14753 2554 14786 2560
rect 14987 2557 15021 2763
rect 14753 2532 14758 2554
rect 14781 2532 14786 2554
rect 14753 2523 14786 2532
rect 14965 2552 15021 2557
rect 14965 2532 14972 2552
rect 14992 2532 15021 2552
rect 14965 2525 15021 2532
rect 14965 2524 15000 2525
rect 14755 2492 14782 2523
rect 15177 2492 15216 2504
rect 14755 2491 15218 2492
rect 14755 2469 15182 2491
rect 15206 2469 15218 2491
rect 14755 2461 15218 2469
rect 11058 2169 11397 2197
rect 11152 2134 11187 2135
rect 11131 2127 11187 2134
rect 11131 2107 11160 2127
rect 11180 2107 11187 2127
rect 11131 2102 11187 2107
rect 11366 2127 11397 2169
rect 11366 2108 11371 2127
rect 11392 2108 11397 2127
rect 11366 2102 11397 2108
rect 12028 2122 12062 2328
rect 13788 2326 13823 2333
rect 12096 2301 12681 2307
rect 12096 2281 12112 2301
rect 12132 2300 12681 2301
rect 12132 2281 12652 2300
rect 12096 2280 12652 2281
rect 12672 2280 12681 2300
rect 12096 2272 12681 2280
rect 13788 2306 13796 2326
rect 13816 2306 13823 2326
rect 13788 2233 13823 2306
rect 14002 2328 14058 2333
rect 14002 2308 14009 2328
rect 14029 2308 14058 2328
rect 14002 2301 14058 2308
rect 14093 2435 14123 2437
rect 14822 2435 14855 2436
rect 14093 2409 14856 2435
rect 14002 2300 14037 2301
rect 14093 2234 14123 2409
rect 14822 2388 14856 2409
rect 14821 2383 14856 2388
rect 14821 2363 14828 2383
rect 14848 2363 14856 2383
rect 14821 2355 14856 2363
rect 14088 2233 14123 2234
rect 13787 2206 14123 2233
rect 14093 2205 14123 2206
rect 14203 2197 14788 2205
rect 14203 2177 14212 2197
rect 14232 2196 14788 2197
rect 14232 2177 14752 2196
rect 14203 2176 14752 2177
rect 14772 2176 14788 2196
rect 14203 2170 14788 2176
rect 14027 2160 14059 2161
rect 14024 2155 14059 2160
rect 14024 2135 14031 2155
rect 14051 2135 14059 2155
rect 14822 2149 14856 2355
rect 14024 2127 14059 2135
rect 12028 2114 12063 2122
rect 11131 1896 11165 2102
rect 12028 2094 12036 2114
rect 12056 2094 12063 2114
rect 12028 2089 12063 2094
rect 12028 2088 12060 2089
rect 11199 2075 11784 2081
rect 11199 2055 11215 2075
rect 11235 2074 11784 2075
rect 11235 2055 11755 2074
rect 11199 2054 11755 2055
rect 11775 2054 11784 2074
rect 11199 2046 11784 2054
rect 13406 1969 13991 1977
rect 13406 1949 13415 1969
rect 13435 1968 13991 1969
rect 13435 1949 13955 1968
rect 13406 1948 13955 1949
rect 13975 1948 13991 1968
rect 13406 1942 13991 1948
rect 13780 1918 13819 1922
rect 14025 1921 14059 2127
rect 14588 2142 14623 2148
rect 14588 2123 14593 2142
rect 14614 2123 14623 2142
rect 14588 2114 14623 2123
rect 14800 2144 14856 2149
rect 14800 2124 14807 2144
rect 14827 2124 14856 2144
rect 14800 2117 14856 2124
rect 14978 2295 15010 2307
rect 14978 2277 14985 2295
rect 15007 2277 15010 2295
rect 14800 2116 14835 2117
rect 14592 2046 14621 2114
rect 14592 2012 14938 2046
rect 13780 1898 13788 1918
rect 13808 1898 13819 1918
rect 11131 1888 11166 1896
rect 11131 1868 11139 1888
rect 11159 1880 11166 1888
rect 11159 1868 11170 1880
rect 11131 1631 11170 1868
rect 12001 1845 12287 1846
rect 11486 1837 12289 1845
rect 11486 1820 11497 1837
rect 11487 1815 11497 1820
rect 11521 1820 12289 1837
rect 11521 1815 11526 1820
rect 11487 1802 11526 1815
rect 12031 1754 12066 1755
rect 12010 1747 12066 1754
rect 12010 1727 12039 1747
rect 12059 1727 12066 1747
rect 12010 1722 12066 1727
rect 12250 1745 12289 1820
rect 13780 1823 13819 1898
rect 14003 1916 14059 1921
rect 14003 1896 14010 1916
rect 14030 1896 14059 1916
rect 14003 1889 14059 1896
rect 14003 1888 14038 1889
rect 14543 1828 14582 1841
rect 14543 1823 14548 1828
rect 13780 1806 14548 1823
rect 14572 1823 14582 1828
rect 14572 1806 14583 1823
rect 13780 1798 14583 1806
rect 13782 1797 14068 1798
rect 14899 1775 14938 2012
rect 14899 1763 14910 1775
rect 14903 1755 14910 1763
rect 14930 1755 14938 1775
rect 14903 1747 14938 1755
rect 12250 1725 12261 1745
rect 12281 1725 12289 1745
rect 11131 1597 11477 1631
rect 11448 1529 11477 1597
rect 11234 1526 11269 1527
rect 10312 1427 10646 1455
rect 11213 1519 11269 1526
rect 11213 1499 11242 1519
rect 11262 1499 11269 1519
rect 11213 1494 11269 1499
rect 11446 1520 11481 1529
rect 11446 1501 11455 1520
rect 11476 1501 11481 1520
rect 11446 1495 11481 1501
rect 12010 1516 12044 1722
rect 12250 1721 12289 1725
rect 12078 1695 12663 1701
rect 12078 1675 12094 1695
rect 12114 1694 12663 1695
rect 12114 1675 12634 1694
rect 12078 1674 12634 1675
rect 12654 1674 12663 1694
rect 12078 1666 12663 1674
rect 14285 1589 14870 1597
rect 14285 1569 14294 1589
rect 14314 1588 14870 1589
rect 14314 1569 14834 1588
rect 14285 1568 14834 1569
rect 14854 1568 14870 1588
rect 14285 1562 14870 1568
rect 14009 1554 14041 1555
rect 14006 1549 14041 1554
rect 14006 1529 14013 1549
rect 14033 1529 14041 1549
rect 14904 1541 14938 1747
rect 14006 1521 14041 1529
rect 12010 1508 12045 1516
rect 5266 1084 5301 1092
rect 3270 1071 3305 1079
rect 1678 1060 1713 1061
rect 1471 1028 1500 1058
rect 3270 1051 3278 1071
rect 3298 1051 3305 1071
rect 3270 1046 3305 1051
rect 3270 1045 3302 1046
rect 1471 1020 1853 1028
rect 1471 1001 1824 1020
rect 1845 1001 1853 1020
rect 1471 996 1853 1001
rect 4648 926 5233 934
rect 4648 906 4657 926
rect 4677 925 5233 926
rect 4677 906 5197 925
rect 4648 905 5197 906
rect 5217 905 5233 925
rect 4648 899 5233 905
rect 658 842 666 862
rect 686 842 697 862
rect 658 767 697 842
rect 881 860 937 865
rect 881 840 888 860
rect 908 840 937 860
rect 881 833 937 840
rect 5022 875 5061 879
rect 5267 878 5301 1084
rect 5831 1096 5865 1104
rect 5831 1078 5838 1096
rect 5857 1078 5865 1096
rect 5831 1071 5865 1078
rect 6042 1101 6098 1106
rect 6042 1081 6049 1101
rect 6069 1081 6098 1101
rect 6042 1074 6098 1081
rect 7634 1092 7668 1298
rect 9407 1295 9442 1302
rect 7702 1271 8287 1277
rect 7702 1251 7718 1271
rect 7738 1270 8287 1271
rect 7738 1251 8258 1270
rect 7702 1250 8258 1251
rect 8278 1250 8287 1270
rect 7702 1242 8287 1250
rect 9407 1275 9415 1295
rect 9435 1275 9442 1295
rect 9407 1202 9442 1275
rect 9621 1297 9677 1302
rect 9621 1277 9628 1297
rect 9648 1277 9677 1297
rect 9621 1270 9677 1277
rect 9712 1404 9742 1406
rect 10441 1404 10474 1405
rect 9712 1378 10475 1404
rect 9621 1269 9656 1270
rect 9712 1203 9742 1378
rect 10441 1357 10475 1378
rect 10440 1352 10475 1357
rect 10440 1332 10447 1352
rect 10467 1332 10475 1352
rect 10440 1324 10475 1332
rect 9707 1202 9742 1203
rect 9406 1175 9742 1202
rect 9712 1174 9742 1175
rect 9822 1166 10407 1174
rect 9822 1146 9831 1166
rect 9851 1165 10407 1166
rect 9851 1146 10371 1165
rect 9822 1145 10371 1146
rect 10391 1145 10407 1165
rect 9822 1139 10407 1145
rect 9646 1129 9678 1130
rect 9643 1124 9678 1129
rect 9643 1104 9650 1124
rect 9670 1104 9678 1124
rect 10441 1118 10475 1324
rect 11213 1288 11247 1494
rect 12010 1488 12018 1508
rect 12038 1488 12045 1508
rect 12010 1483 12045 1488
rect 12010 1482 12042 1483
rect 11281 1467 11866 1473
rect 11281 1447 11297 1467
rect 11317 1466 11866 1467
rect 11317 1447 11837 1466
rect 11281 1446 11837 1447
rect 11857 1446 11866 1466
rect 11281 1438 11866 1446
rect 11946 1437 11976 1438
rect 11946 1410 12282 1437
rect 11946 1409 11981 1410
rect 11213 1280 11248 1288
rect 11213 1260 11221 1280
rect 11241 1260 11248 1280
rect 11213 1255 11248 1260
rect 11213 1234 11247 1255
rect 11946 1234 11976 1409
rect 12032 1342 12067 1343
rect 11213 1208 11976 1234
rect 11214 1207 11247 1208
rect 11946 1206 11976 1208
rect 12011 1335 12067 1342
rect 12011 1315 12040 1335
rect 12060 1315 12067 1335
rect 12011 1310 12067 1315
rect 12246 1337 12281 1410
rect 12246 1317 12253 1337
rect 12273 1317 12281 1337
rect 13388 1363 13973 1371
rect 13388 1343 13397 1363
rect 13417 1362 13973 1363
rect 13417 1343 13937 1362
rect 13388 1342 13937 1343
rect 13957 1342 13973 1362
rect 13388 1336 13973 1342
rect 12246 1310 12281 1317
rect 14007 1315 14041 1521
rect 14670 1529 14706 1538
rect 14670 1512 14679 1529
rect 14698 1512 14706 1529
rect 14670 1503 14706 1512
rect 14882 1536 14938 1541
rect 14882 1516 14889 1536
rect 14909 1516 14938 1536
rect 14882 1509 14938 1516
rect 14882 1508 14917 1509
rect 14676 1468 14702 1503
rect 14978 1468 15010 2277
rect 15422 2210 15451 2895
rect 18066 2890 18074 2910
rect 18094 2890 18105 2910
rect 16382 2876 16668 2877
rect 15867 2868 16670 2876
rect 15867 2851 15878 2868
rect 15868 2846 15878 2851
rect 15902 2851 16670 2868
rect 15902 2846 15907 2851
rect 15868 2833 15907 2846
rect 16412 2785 16447 2786
rect 16391 2778 16447 2785
rect 16391 2758 16420 2778
rect 16440 2758 16447 2778
rect 16391 2753 16447 2758
rect 16631 2776 16670 2851
rect 18066 2815 18105 2890
rect 18289 2908 18345 2913
rect 18289 2888 18296 2908
rect 18316 2888 18345 2908
rect 18289 2881 18345 2888
rect 18289 2880 18324 2881
rect 18829 2820 18868 2833
rect 18829 2815 18834 2820
rect 18066 2798 18834 2815
rect 18858 2815 18868 2820
rect 18858 2798 18869 2815
rect 18066 2790 18869 2798
rect 18068 2789 18354 2790
rect 16631 2756 16642 2776
rect 16662 2756 16670 2776
rect 19285 2771 19314 3456
rect 19622 3210 19649 4910
rect 22466 4939 22474 4959
rect 22494 4939 22505 4959
rect 20685 4886 20971 4887
rect 20170 4878 20973 4886
rect 20170 4861 20181 4878
rect 20171 4856 20181 4861
rect 20205 4861 20973 4878
rect 20205 4856 20210 4861
rect 20171 4843 20210 4856
rect 20715 4795 20750 4796
rect 20694 4788 20750 4795
rect 20694 4768 20723 4788
rect 20743 4768 20750 4788
rect 20694 4763 20750 4768
rect 20934 4786 20973 4861
rect 22466 4864 22505 4939
rect 22689 4957 22745 4962
rect 22689 4937 22696 4957
rect 22716 4937 22745 4957
rect 22689 4930 22745 4937
rect 22689 4929 22724 4930
rect 23229 4869 23268 4882
rect 23229 4864 23234 4869
rect 22466 4847 23234 4864
rect 23258 4864 23268 4869
rect 23258 4847 23269 4864
rect 22466 4839 23269 4847
rect 22468 4838 22754 4839
rect 20934 4766 20945 4786
rect 20965 4766 20973 4786
rect 23790 4815 23817 6515
rect 24125 6269 24154 6954
rect 25085 6935 25371 6936
rect 24570 6927 25373 6935
rect 24570 6910 24581 6927
rect 24571 6905 24581 6910
rect 24605 6910 25373 6927
rect 24605 6905 24610 6910
rect 24571 6892 24610 6905
rect 25115 6844 25150 6845
rect 25094 6837 25150 6844
rect 25094 6817 25123 6837
rect 25143 6817 25150 6837
rect 25094 6812 25150 6817
rect 25334 6835 25373 6910
rect 26880 6912 26919 6987
rect 27103 7005 27159 7010
rect 27103 6985 27110 7005
rect 27130 6985 27159 7005
rect 27103 6978 27159 6985
rect 27103 6977 27138 6978
rect 27643 6917 27682 6930
rect 27643 6912 27648 6917
rect 26880 6895 27648 6912
rect 27672 6912 27682 6917
rect 27672 6895 27683 6912
rect 26880 6887 27683 6895
rect 26882 6886 27168 6887
rect 28099 6868 28128 7553
rect 28540 7486 28572 8295
rect 28848 8260 28874 8295
rect 28633 8254 28668 8255
rect 28612 8247 28668 8254
rect 28612 8227 28641 8247
rect 28661 8227 28668 8247
rect 28612 8222 28668 8227
rect 28844 8251 28880 8260
rect 28844 8234 28852 8251
rect 28871 8234 28880 8251
rect 28844 8225 28880 8234
rect 29509 8242 29543 8448
rect 31269 8446 31304 8453
rect 29577 8421 30162 8427
rect 29577 8401 29593 8421
rect 29613 8420 30162 8421
rect 29613 8401 30133 8420
rect 29577 8400 30133 8401
rect 30153 8400 30162 8420
rect 29577 8392 30162 8400
rect 31269 8426 31277 8446
rect 31297 8426 31304 8446
rect 31269 8353 31304 8426
rect 31483 8448 31539 8453
rect 31483 8428 31490 8448
rect 31510 8428 31539 8448
rect 31483 8421 31539 8428
rect 31574 8555 31604 8557
rect 32303 8555 32336 8556
rect 31574 8529 32337 8555
rect 31483 8420 31518 8421
rect 31574 8354 31604 8529
rect 32303 8508 32337 8529
rect 32302 8503 32337 8508
rect 32302 8483 32309 8503
rect 32329 8483 32337 8503
rect 32302 8475 32337 8483
rect 31569 8353 31604 8354
rect 31268 8326 31604 8353
rect 31574 8325 31604 8326
rect 31684 8317 32269 8325
rect 31684 8297 31693 8317
rect 31713 8316 32269 8317
rect 31713 8297 32233 8316
rect 31684 8296 32233 8297
rect 32253 8296 32269 8316
rect 31684 8290 32269 8296
rect 31508 8280 31540 8281
rect 31505 8275 31540 8280
rect 31505 8255 31512 8275
rect 31532 8255 31540 8275
rect 32303 8269 32337 8475
rect 33075 8439 33109 8645
rect 33872 8639 33880 8659
rect 33900 8639 33907 8659
rect 33872 8634 33907 8639
rect 33872 8633 33904 8634
rect 33143 8618 33728 8624
rect 33143 8598 33159 8618
rect 33179 8617 33728 8618
rect 33179 8598 33699 8617
rect 33143 8597 33699 8598
rect 33719 8597 33728 8617
rect 33143 8589 33728 8597
rect 33808 8588 33838 8589
rect 33808 8561 34144 8588
rect 33808 8560 33843 8561
rect 33075 8431 33110 8439
rect 33075 8411 33083 8431
rect 33103 8411 33110 8431
rect 33075 8406 33110 8411
rect 33075 8385 33109 8406
rect 33808 8385 33838 8560
rect 33894 8493 33929 8494
rect 33075 8359 33838 8385
rect 33076 8358 33109 8359
rect 33808 8357 33838 8359
rect 33873 8486 33929 8493
rect 33873 8466 33902 8486
rect 33922 8466 33929 8486
rect 33873 8461 33929 8466
rect 34108 8488 34143 8561
rect 34108 8468 34115 8488
rect 34135 8468 34143 8488
rect 34108 8461 34143 8468
rect 31505 8247 31540 8255
rect 29509 8234 29544 8242
rect 28612 8016 28646 8222
rect 29509 8214 29517 8234
rect 29537 8214 29544 8234
rect 29509 8209 29544 8214
rect 29509 8208 29541 8209
rect 28680 8195 29265 8201
rect 28680 8175 28696 8195
rect 28716 8194 29265 8195
rect 28716 8175 29236 8194
rect 28680 8174 29236 8175
rect 29256 8174 29265 8194
rect 28680 8166 29265 8174
rect 30887 8089 31472 8097
rect 30887 8069 30896 8089
rect 30916 8088 31472 8089
rect 30916 8069 31436 8088
rect 30887 8068 31436 8069
rect 31456 8068 31472 8088
rect 30887 8062 31472 8068
rect 31261 8038 31300 8042
rect 31506 8041 31540 8247
rect 32069 8262 32104 8268
rect 32069 8243 32074 8262
rect 32095 8243 32104 8262
rect 32069 8234 32104 8243
rect 32281 8264 32337 8269
rect 32281 8244 32288 8264
rect 32308 8244 32337 8264
rect 32281 8237 32337 8244
rect 32904 8308 33238 8336
rect 32281 8236 32316 8237
rect 32073 8166 32102 8234
rect 32073 8132 32419 8166
rect 31261 8018 31269 8038
rect 31289 8018 31300 8038
rect 28612 8008 28647 8016
rect 28612 7988 28620 8008
rect 28640 8000 28647 8008
rect 28640 7988 28651 8000
rect 28612 7751 28651 7988
rect 29482 7965 29768 7966
rect 28967 7957 29770 7965
rect 28967 7940 28978 7957
rect 28968 7935 28978 7940
rect 29002 7940 29770 7957
rect 29002 7935 29007 7940
rect 28968 7922 29007 7935
rect 29512 7874 29547 7875
rect 29491 7867 29547 7874
rect 29491 7847 29520 7867
rect 29540 7847 29547 7867
rect 29491 7842 29547 7847
rect 29731 7865 29770 7940
rect 31261 7943 31300 8018
rect 31484 8036 31540 8041
rect 31484 8016 31491 8036
rect 31511 8016 31540 8036
rect 31484 8009 31540 8016
rect 31484 8008 31519 8009
rect 32024 7948 32063 7961
rect 32024 7943 32029 7948
rect 31261 7926 32029 7943
rect 32053 7943 32063 7948
rect 32053 7926 32064 7943
rect 31261 7918 32064 7926
rect 31263 7917 31549 7918
rect 32380 7895 32419 8132
rect 32380 7883 32391 7895
rect 32384 7875 32391 7883
rect 32411 7875 32419 7895
rect 32384 7867 32419 7875
rect 29731 7845 29742 7865
rect 29762 7845 29770 7865
rect 28612 7717 28958 7751
rect 28929 7649 28958 7717
rect 28715 7646 28750 7647
rect 28540 7468 28543 7486
rect 28565 7468 28572 7486
rect 28540 7456 28572 7468
rect 28694 7639 28750 7646
rect 28694 7619 28723 7639
rect 28743 7619 28750 7639
rect 28694 7614 28750 7619
rect 28927 7640 28962 7649
rect 28927 7621 28936 7640
rect 28957 7621 28962 7640
rect 28927 7615 28962 7621
rect 29491 7636 29525 7842
rect 29731 7841 29770 7845
rect 29559 7815 30144 7821
rect 29559 7795 29575 7815
rect 29595 7814 30144 7815
rect 29595 7795 30115 7814
rect 29559 7794 30115 7795
rect 30135 7794 30144 7814
rect 29559 7786 30144 7794
rect 31766 7709 32351 7717
rect 31766 7689 31775 7709
rect 31795 7708 32351 7709
rect 31795 7689 32315 7708
rect 31766 7688 32315 7689
rect 32335 7688 32351 7708
rect 31766 7682 32351 7688
rect 31490 7674 31522 7675
rect 31487 7669 31522 7674
rect 31487 7649 31494 7669
rect 31514 7649 31522 7669
rect 32385 7661 32419 7867
rect 31487 7641 31522 7649
rect 29491 7628 29526 7636
rect 28694 7408 28728 7614
rect 29491 7608 29499 7628
rect 29519 7608 29526 7628
rect 29491 7603 29526 7608
rect 29491 7602 29523 7603
rect 28762 7587 29347 7593
rect 28762 7567 28778 7587
rect 28798 7586 29347 7587
rect 28798 7567 29318 7586
rect 28762 7566 29318 7567
rect 29338 7566 29347 7586
rect 28762 7558 29347 7566
rect 29427 7557 29457 7558
rect 29427 7530 29763 7557
rect 29427 7529 29462 7530
rect 28694 7400 28729 7408
rect 28694 7380 28702 7400
rect 28722 7380 28729 7400
rect 28694 7375 28729 7380
rect 28694 7354 28728 7375
rect 29427 7354 29457 7529
rect 29513 7462 29548 7463
rect 28694 7328 29457 7354
rect 28695 7327 28728 7328
rect 29427 7326 29457 7328
rect 29492 7455 29548 7462
rect 29492 7435 29521 7455
rect 29541 7435 29548 7455
rect 29492 7430 29548 7435
rect 29727 7457 29762 7530
rect 29727 7437 29734 7457
rect 29754 7437 29762 7457
rect 30869 7483 31454 7491
rect 30869 7463 30878 7483
rect 30898 7482 31454 7483
rect 30898 7463 31418 7482
rect 30869 7462 31418 7463
rect 31438 7462 31454 7482
rect 30869 7456 31454 7462
rect 29727 7430 29762 7437
rect 31488 7435 31522 7641
rect 32153 7655 32184 7661
rect 32153 7636 32158 7655
rect 32179 7636 32184 7655
rect 32153 7594 32184 7636
rect 32363 7656 32419 7661
rect 32363 7636 32370 7656
rect 32390 7636 32419 7656
rect 32363 7629 32419 7636
rect 32363 7628 32398 7629
rect 32153 7566 32492 7594
rect 28332 7294 28795 7302
rect 28332 7272 28344 7294
rect 28368 7272 28795 7294
rect 28332 7271 28795 7272
rect 28334 7259 28373 7271
rect 28768 7240 28795 7271
rect 28550 7238 28585 7239
rect 28529 7231 28585 7238
rect 28529 7211 28558 7231
rect 28578 7211 28585 7231
rect 28529 7206 28585 7211
rect 28764 7231 28797 7240
rect 28764 7209 28769 7231
rect 28792 7209 28797 7231
rect 28529 7000 28563 7206
rect 28764 7203 28797 7209
rect 29492 7224 29526 7430
rect 31252 7428 31287 7435
rect 29560 7403 30145 7409
rect 29560 7383 29576 7403
rect 29596 7402 30145 7403
rect 29596 7383 30116 7402
rect 29560 7382 30116 7383
rect 30136 7382 30145 7402
rect 29560 7374 30145 7382
rect 31252 7408 31260 7428
rect 31280 7408 31287 7428
rect 31252 7335 31287 7408
rect 31466 7430 31522 7435
rect 31466 7410 31473 7430
rect 31493 7410 31522 7430
rect 31466 7403 31522 7410
rect 31557 7537 31587 7539
rect 32286 7537 32319 7538
rect 31557 7511 32320 7537
rect 31466 7402 31501 7403
rect 31557 7336 31587 7511
rect 32286 7490 32320 7511
rect 32285 7485 32320 7490
rect 32285 7465 32292 7485
rect 32312 7465 32320 7485
rect 32285 7457 32320 7465
rect 31552 7335 31587 7336
rect 31251 7308 31587 7335
rect 31557 7307 31587 7308
rect 31667 7299 32252 7307
rect 31667 7279 31676 7299
rect 31696 7298 32252 7299
rect 31696 7279 32216 7298
rect 31667 7278 32216 7279
rect 32236 7278 32252 7298
rect 31667 7272 32252 7278
rect 31491 7262 31523 7263
rect 31488 7257 31523 7262
rect 31488 7237 31495 7257
rect 31515 7237 31523 7257
rect 32286 7251 32320 7457
rect 31488 7229 31523 7237
rect 29492 7216 29527 7224
rect 29492 7196 29500 7216
rect 29520 7196 29527 7216
rect 29492 7191 29527 7196
rect 29492 7190 29524 7191
rect 28597 7179 29182 7185
rect 28597 7159 28613 7179
rect 28633 7178 29182 7179
rect 28633 7159 29153 7178
rect 28597 7158 29153 7159
rect 29173 7158 29182 7178
rect 28597 7150 29182 7158
rect 30870 7071 31455 7079
rect 30870 7051 30879 7071
rect 30899 7070 31455 7071
rect 30899 7051 31419 7070
rect 30870 7050 31419 7051
rect 31439 7050 31455 7070
rect 30870 7044 31455 7050
rect 31244 7020 31283 7024
rect 31489 7023 31523 7229
rect 32053 7241 32087 7249
rect 32053 7223 32060 7241
rect 32079 7223 32087 7241
rect 32053 7216 32087 7223
rect 32264 7246 32320 7251
rect 32264 7226 32271 7246
rect 32291 7226 32320 7246
rect 32264 7219 32320 7226
rect 32264 7218 32299 7219
rect 32057 7186 32086 7216
rect 32057 7178 32439 7186
rect 32057 7159 32410 7178
rect 32431 7159 32439 7178
rect 32057 7154 32439 7159
rect 31244 7000 31252 7020
rect 31272 7000 31283 7020
rect 28529 6999 28564 7000
rect 28497 6992 28564 6999
rect 28497 6972 28537 6992
rect 28557 6972 28564 6992
rect 28497 6969 28564 6972
rect 28497 6966 28562 6969
rect 28068 6865 28133 6868
rect 25334 6815 25345 6835
rect 25365 6815 25373 6835
rect 28066 6862 28133 6865
rect 28066 6842 28073 6862
rect 28093 6842 28133 6862
rect 28066 6835 28133 6842
rect 28066 6834 28101 6835
rect 24178 6676 24560 6681
rect 24178 6657 24186 6676
rect 24207 6657 24560 6676
rect 24178 6649 24560 6657
rect 24531 6619 24560 6649
rect 24318 6616 24353 6617
rect 24297 6609 24353 6616
rect 24297 6589 24326 6609
rect 24346 6589 24353 6609
rect 24297 6584 24353 6589
rect 24530 6612 24564 6619
rect 24530 6594 24538 6612
rect 24557 6594 24564 6612
rect 24530 6586 24564 6594
rect 25094 6606 25128 6812
rect 25334 6811 25373 6815
rect 25162 6785 25747 6791
rect 25162 6765 25178 6785
rect 25198 6784 25747 6785
rect 25198 6765 25718 6784
rect 25162 6764 25718 6765
rect 25738 6764 25747 6784
rect 25162 6756 25747 6764
rect 27448 6676 28033 6684
rect 27448 6656 27457 6676
rect 27477 6675 28033 6676
rect 27477 6656 27997 6675
rect 27448 6655 27997 6656
rect 28017 6655 28033 6675
rect 27448 6649 28033 6655
rect 27106 6643 27138 6644
rect 27103 6638 27138 6643
rect 27103 6618 27110 6638
rect 27130 6618 27138 6638
rect 27103 6610 27138 6618
rect 25094 6598 25129 6606
rect 24297 6378 24331 6584
rect 25094 6578 25102 6598
rect 25122 6578 25129 6598
rect 25094 6573 25129 6578
rect 25094 6572 25126 6573
rect 24365 6557 24950 6563
rect 24365 6537 24381 6557
rect 24401 6556 24950 6557
rect 24401 6537 24921 6556
rect 24365 6536 24921 6537
rect 24941 6536 24950 6556
rect 24365 6528 24950 6536
rect 25030 6527 25060 6528
rect 25030 6500 25366 6527
rect 25030 6499 25065 6500
rect 24297 6370 24332 6378
rect 24297 6350 24305 6370
rect 24325 6350 24332 6370
rect 24297 6345 24332 6350
rect 24297 6324 24331 6345
rect 25030 6324 25060 6499
rect 25116 6432 25151 6433
rect 24297 6298 25060 6324
rect 24298 6297 24331 6298
rect 25030 6296 25060 6298
rect 25095 6425 25151 6432
rect 25095 6405 25124 6425
rect 25144 6405 25151 6425
rect 25095 6400 25151 6405
rect 25330 6427 25365 6500
rect 25330 6407 25337 6427
rect 25357 6407 25365 6427
rect 26485 6452 27070 6460
rect 26485 6432 26494 6452
rect 26514 6451 27070 6452
rect 26514 6432 27034 6451
rect 26485 6431 27034 6432
rect 27054 6431 27070 6451
rect 26485 6425 27070 6431
rect 25330 6400 25365 6407
rect 27104 6404 27138 6610
rect 27831 6620 27872 6631
rect 28067 6628 28101 6834
rect 27831 6602 27841 6620
rect 27859 6602 27872 6620
rect 27831 6594 27872 6602
rect 28045 6623 28101 6628
rect 28045 6603 28052 6623
rect 28072 6603 28101 6623
rect 28045 6596 28101 6603
rect 28045 6595 28080 6596
rect 27840 6564 27866 6594
rect 27840 6563 28178 6564
rect 27840 6527 28194 6563
rect 24125 6241 24464 6269
rect 24219 6206 24254 6207
rect 24198 6199 24254 6206
rect 24198 6179 24227 6199
rect 24247 6179 24254 6199
rect 24198 6174 24254 6179
rect 24433 6199 24464 6241
rect 24433 6180 24438 6199
rect 24459 6180 24464 6199
rect 24433 6174 24464 6180
rect 25095 6194 25129 6400
rect 26868 6397 26903 6404
rect 25163 6373 25748 6379
rect 25163 6353 25179 6373
rect 25199 6372 25748 6373
rect 25199 6353 25719 6372
rect 25163 6352 25719 6353
rect 25739 6352 25748 6372
rect 25163 6344 25748 6352
rect 26868 6377 26876 6397
rect 26896 6377 26903 6397
rect 26868 6304 26903 6377
rect 27082 6399 27138 6404
rect 27082 6379 27089 6399
rect 27109 6379 27138 6399
rect 27082 6372 27138 6379
rect 27173 6506 27203 6508
rect 27902 6506 27935 6507
rect 27173 6480 27936 6506
rect 27082 6371 27117 6372
rect 27173 6305 27203 6480
rect 27902 6459 27936 6480
rect 27901 6454 27936 6459
rect 27901 6434 27908 6454
rect 27928 6434 27936 6454
rect 27901 6426 27936 6434
rect 27168 6304 27203 6305
rect 26867 6277 27203 6304
rect 27173 6276 27203 6277
rect 27283 6268 27868 6276
rect 27283 6248 27292 6268
rect 27312 6267 27868 6268
rect 27312 6248 27832 6267
rect 27283 6247 27832 6248
rect 27852 6247 27868 6267
rect 27283 6241 27868 6247
rect 27107 6231 27139 6232
rect 27104 6226 27139 6231
rect 27104 6206 27111 6226
rect 27131 6206 27139 6226
rect 27902 6220 27936 6426
rect 27104 6198 27139 6206
rect 25095 6186 25130 6194
rect 24198 5968 24232 6174
rect 25095 6166 25103 6186
rect 25123 6166 25130 6186
rect 25095 6161 25130 6166
rect 25095 6160 25127 6161
rect 24266 6147 24851 6153
rect 24266 6127 24282 6147
rect 24302 6146 24851 6147
rect 24302 6127 24822 6146
rect 24266 6126 24822 6127
rect 24842 6126 24851 6146
rect 24266 6118 24851 6126
rect 26486 6040 27071 6048
rect 26486 6020 26495 6040
rect 26515 6039 27071 6040
rect 26515 6020 27035 6039
rect 26486 6019 27035 6020
rect 27055 6019 27071 6039
rect 26486 6013 27071 6019
rect 26860 5989 26899 5993
rect 27105 5992 27139 6198
rect 27668 6213 27703 6219
rect 27668 6194 27673 6213
rect 27694 6194 27703 6213
rect 27668 6185 27703 6194
rect 27880 6215 27936 6220
rect 27880 6195 27887 6215
rect 27907 6195 27936 6215
rect 27880 6188 27936 6195
rect 27880 6187 27915 6188
rect 27672 6117 27701 6185
rect 27672 6083 28018 6117
rect 26860 5969 26868 5989
rect 26888 5969 26899 5989
rect 24198 5960 24233 5968
rect 24198 5940 24206 5960
rect 24226 5952 24233 5960
rect 24226 5940 24237 5952
rect 24198 5703 24237 5940
rect 25068 5917 25354 5918
rect 24553 5909 25356 5917
rect 24553 5892 24564 5909
rect 24554 5887 24564 5892
rect 24588 5892 25356 5909
rect 24588 5887 24593 5892
rect 24554 5874 24593 5887
rect 25098 5826 25133 5827
rect 25077 5819 25133 5826
rect 25077 5799 25106 5819
rect 25126 5799 25133 5819
rect 25077 5794 25133 5799
rect 25317 5817 25356 5892
rect 26860 5894 26899 5969
rect 27083 5987 27139 5992
rect 27083 5967 27090 5987
rect 27110 5967 27139 5987
rect 27083 5960 27139 5967
rect 27083 5959 27118 5960
rect 27623 5899 27662 5912
rect 27623 5894 27628 5899
rect 26860 5877 27628 5894
rect 27652 5894 27662 5899
rect 27652 5877 27663 5894
rect 26860 5869 27663 5877
rect 26862 5868 27148 5869
rect 27979 5846 28018 6083
rect 27979 5834 27990 5846
rect 27983 5826 27990 5834
rect 28010 5826 28018 5846
rect 27983 5818 28018 5826
rect 25317 5797 25328 5817
rect 25348 5797 25356 5817
rect 24198 5669 24544 5703
rect 24515 5601 24544 5669
rect 24301 5598 24336 5599
rect 24280 5591 24336 5598
rect 24280 5571 24309 5591
rect 24329 5571 24336 5591
rect 24280 5566 24336 5571
rect 24513 5592 24548 5601
rect 24513 5573 24522 5592
rect 24543 5573 24548 5592
rect 24513 5567 24548 5573
rect 25077 5588 25111 5794
rect 25317 5793 25356 5797
rect 25145 5767 25730 5773
rect 25145 5747 25161 5767
rect 25181 5766 25730 5767
rect 25181 5747 25701 5766
rect 25145 5746 25701 5747
rect 25721 5746 25730 5766
rect 25145 5738 25730 5746
rect 27365 5660 27950 5668
rect 27365 5640 27374 5660
rect 27394 5659 27950 5660
rect 27394 5640 27914 5659
rect 27365 5639 27914 5640
rect 27934 5639 27950 5659
rect 27365 5633 27950 5639
rect 27089 5625 27121 5626
rect 27086 5620 27121 5625
rect 27086 5600 27093 5620
rect 27113 5600 27121 5620
rect 27984 5612 28018 5818
rect 27086 5592 27121 5600
rect 25077 5580 25112 5588
rect 24280 5360 24314 5566
rect 25077 5560 25085 5580
rect 25105 5560 25112 5580
rect 25077 5555 25112 5560
rect 25077 5554 25109 5555
rect 24348 5539 24933 5545
rect 24348 5519 24364 5539
rect 24384 5538 24933 5539
rect 24384 5519 24904 5538
rect 24348 5518 24904 5519
rect 24924 5518 24933 5538
rect 24348 5510 24933 5518
rect 25013 5509 25043 5510
rect 25013 5482 25349 5509
rect 25013 5481 25048 5482
rect 24280 5352 24315 5360
rect 24280 5332 24288 5352
rect 24308 5332 24315 5352
rect 24280 5327 24315 5332
rect 24280 5306 24314 5327
rect 25013 5306 25043 5481
rect 25099 5414 25134 5415
rect 24280 5280 25043 5306
rect 24281 5279 24314 5280
rect 25013 5278 25043 5280
rect 25078 5407 25134 5414
rect 25078 5387 25107 5407
rect 25127 5387 25134 5407
rect 25078 5382 25134 5387
rect 25313 5409 25348 5482
rect 25313 5389 25320 5409
rect 25340 5389 25348 5409
rect 26468 5434 27053 5442
rect 26468 5414 26477 5434
rect 26497 5433 27053 5434
rect 26497 5414 27017 5433
rect 26468 5413 27017 5414
rect 27037 5413 27053 5433
rect 26468 5407 27053 5413
rect 25313 5382 25348 5389
rect 27087 5386 27121 5592
rect 27750 5600 27786 5609
rect 27750 5583 27759 5600
rect 27778 5583 27786 5600
rect 27750 5574 27786 5583
rect 27962 5607 28018 5612
rect 27962 5587 27969 5607
rect 27989 5587 28018 5607
rect 27962 5580 28018 5587
rect 27962 5579 27997 5580
rect 27756 5539 27782 5574
rect 28064 5539 28096 5540
rect 27756 5534 28096 5539
rect 27756 5516 28071 5534
rect 28093 5516 28096 5534
rect 27756 5511 28096 5516
rect 28064 5510 28096 5511
rect 23932 5259 24249 5262
rect 23932 5232 23935 5259
rect 23962 5232 24249 5259
rect 23932 5226 24249 5232
rect 23932 5223 23968 5226
rect 24213 5196 24249 5226
rect 23997 5192 24032 5193
rect 23976 5185 24032 5192
rect 23976 5165 24005 5185
rect 24025 5165 24032 5185
rect 23976 5160 24032 5165
rect 24211 5190 24249 5196
rect 24211 5164 24217 5190
rect 24243 5164 24249 5190
rect 23976 4961 24010 5160
rect 24211 5156 24249 5164
rect 25078 5176 25112 5382
rect 26851 5379 26886 5386
rect 25146 5355 25731 5361
rect 25146 5335 25162 5355
rect 25182 5354 25731 5355
rect 25182 5335 25702 5354
rect 25146 5334 25702 5335
rect 25722 5334 25731 5354
rect 25146 5326 25731 5334
rect 26851 5359 26859 5379
rect 26879 5359 26886 5379
rect 26851 5286 26886 5359
rect 27065 5381 27121 5386
rect 27065 5361 27072 5381
rect 27092 5361 27121 5381
rect 27065 5354 27121 5361
rect 27156 5488 27186 5490
rect 27885 5488 27918 5489
rect 27156 5462 27919 5488
rect 27065 5353 27100 5354
rect 27156 5287 27186 5462
rect 27885 5441 27919 5462
rect 27884 5436 27919 5441
rect 27884 5416 27891 5436
rect 27911 5416 27919 5436
rect 27884 5408 27919 5416
rect 27151 5286 27186 5287
rect 26850 5259 27186 5286
rect 27156 5258 27186 5259
rect 27266 5250 27851 5258
rect 27266 5230 27275 5250
rect 27295 5249 27851 5250
rect 27295 5230 27815 5249
rect 27266 5229 27815 5230
rect 27835 5229 27851 5249
rect 27266 5223 27851 5229
rect 27090 5213 27122 5214
rect 27087 5208 27122 5213
rect 27087 5188 27094 5208
rect 27114 5188 27122 5208
rect 27885 5202 27919 5408
rect 27087 5180 27122 5188
rect 25078 5168 25113 5176
rect 25078 5148 25086 5168
rect 25106 5148 25113 5168
rect 25078 5143 25113 5148
rect 25078 5142 25110 5143
rect 24044 5133 24629 5139
rect 24044 5113 24060 5133
rect 24080 5132 24629 5133
rect 24080 5113 24600 5132
rect 24044 5112 24600 5113
rect 24620 5112 24629 5132
rect 24044 5104 24629 5112
rect 26469 5022 27054 5030
rect 26469 5002 26478 5022
rect 26498 5021 27054 5022
rect 26498 5002 27018 5021
rect 26469 5001 27018 5002
rect 27038 5001 27054 5021
rect 26469 4995 27054 5001
rect 26843 4971 26882 4975
rect 27088 4974 27122 5180
rect 27652 5192 27686 5200
rect 27652 5174 27659 5192
rect 27678 5174 27686 5192
rect 27652 5167 27686 5174
rect 27863 5197 27919 5202
rect 27863 5177 27870 5197
rect 27890 5177 27919 5197
rect 27863 5170 27919 5177
rect 27863 5169 27898 5170
rect 27656 5137 27685 5167
rect 27656 5129 28038 5137
rect 27656 5110 28009 5129
rect 28030 5110 28038 5129
rect 27656 5105 28038 5110
rect 23976 4946 24013 4961
rect 23976 4926 23984 4946
rect 24004 4926 24013 4946
rect 23976 4923 24013 4926
rect 23790 4812 23827 4815
rect 23790 4792 23799 4812
rect 23819 4792 23827 4812
rect 23790 4777 23827 4792
rect 19778 4627 20160 4632
rect 19778 4608 19786 4627
rect 19807 4608 20160 4627
rect 19778 4600 20160 4608
rect 20131 4570 20160 4600
rect 19918 4567 19953 4568
rect 19897 4560 19953 4567
rect 19897 4540 19926 4560
rect 19946 4540 19953 4560
rect 19897 4535 19953 4540
rect 20130 4563 20164 4570
rect 20130 4545 20138 4563
rect 20157 4545 20164 4563
rect 20130 4537 20164 4545
rect 20694 4557 20728 4763
rect 20934 4762 20973 4766
rect 20762 4736 21347 4742
rect 20762 4716 20778 4736
rect 20798 4735 21347 4736
rect 20798 4716 21318 4735
rect 20762 4715 21318 4716
rect 21338 4715 21347 4735
rect 20762 4707 21347 4715
rect 23174 4626 23759 4634
rect 23174 4606 23183 4626
rect 23203 4625 23759 4626
rect 23203 4606 23723 4625
rect 23174 4605 23723 4606
rect 23743 4605 23759 4625
rect 23174 4599 23759 4605
rect 22693 4595 22725 4596
rect 22690 4590 22725 4595
rect 22690 4570 22697 4590
rect 22717 4570 22725 4590
rect 23793 4578 23827 4777
rect 23771 4573 23827 4578
rect 22690 4562 22725 4570
rect 20694 4549 20729 4557
rect 19897 4329 19931 4535
rect 20694 4529 20702 4549
rect 20722 4529 20729 4549
rect 20694 4524 20729 4529
rect 20694 4523 20726 4524
rect 19965 4508 20550 4514
rect 19965 4488 19981 4508
rect 20001 4507 20550 4508
rect 20001 4488 20521 4507
rect 19965 4487 20521 4488
rect 20541 4487 20550 4507
rect 19965 4479 20550 4487
rect 20630 4478 20660 4479
rect 20630 4451 20966 4478
rect 20630 4450 20665 4451
rect 19897 4321 19932 4329
rect 19897 4301 19905 4321
rect 19925 4301 19932 4321
rect 19897 4296 19932 4301
rect 19897 4275 19931 4296
rect 20630 4275 20660 4450
rect 20716 4383 20751 4384
rect 19897 4249 20660 4275
rect 19898 4248 19931 4249
rect 20630 4247 20660 4249
rect 20695 4376 20751 4383
rect 20695 4356 20724 4376
rect 20744 4356 20751 4376
rect 20695 4351 20751 4356
rect 20930 4378 20965 4451
rect 20930 4358 20937 4378
rect 20957 4358 20965 4378
rect 22072 4404 22657 4412
rect 22072 4384 22081 4404
rect 22101 4403 22657 4404
rect 22101 4384 22621 4403
rect 22072 4383 22621 4384
rect 22641 4383 22657 4403
rect 22072 4377 22657 4383
rect 20930 4351 20965 4358
rect 22691 4356 22725 4562
rect 23553 4571 23588 4573
rect 23553 4565 23591 4571
rect 23553 4542 23561 4565
rect 23584 4542 23591 4565
rect 23771 4553 23778 4573
rect 23798 4553 23827 4573
rect 23771 4546 23827 4553
rect 23771 4545 23806 4546
rect 23553 4536 23591 4542
rect 23553 4523 23588 4536
rect 23551 4465 23588 4523
rect 19720 4226 19752 4227
rect 19720 4221 20060 4226
rect 19720 4203 19723 4221
rect 19745 4203 20060 4221
rect 19720 4198 20060 4203
rect 19720 4197 19752 4198
rect 20034 4163 20060 4198
rect 19819 4157 19854 4158
rect 19798 4150 19854 4157
rect 19798 4130 19827 4150
rect 19847 4130 19854 4150
rect 19798 4125 19854 4130
rect 20030 4154 20066 4163
rect 20030 4137 20038 4154
rect 20057 4137 20066 4154
rect 20030 4128 20066 4137
rect 20695 4145 20729 4351
rect 22455 4349 22490 4356
rect 20763 4324 21348 4330
rect 20763 4304 20779 4324
rect 20799 4323 21348 4324
rect 20799 4304 21319 4323
rect 20763 4303 21319 4304
rect 21339 4303 21348 4323
rect 20763 4295 21348 4303
rect 22455 4329 22463 4349
rect 22483 4329 22490 4349
rect 22455 4256 22490 4329
rect 22669 4351 22725 4356
rect 22669 4331 22676 4351
rect 22696 4331 22725 4351
rect 22669 4324 22725 4331
rect 22760 4458 22790 4460
rect 23489 4458 23522 4459
rect 22760 4432 23523 4458
rect 22669 4323 22704 4324
rect 22760 4257 22790 4432
rect 23489 4411 23523 4432
rect 23551 4448 23586 4465
rect 23551 4447 23845 4448
rect 23551 4446 23888 4447
rect 23551 4439 23893 4446
rect 23551 4413 23853 4439
rect 23884 4413 23893 4439
rect 23488 4406 23523 4411
rect 23844 4410 23893 4413
rect 23488 4386 23495 4406
rect 23515 4386 23523 4406
rect 23850 4405 23893 4410
rect 23488 4378 23523 4386
rect 22755 4256 22790 4257
rect 22454 4229 22790 4256
rect 22760 4228 22790 4229
rect 22870 4220 23455 4228
rect 22870 4200 22879 4220
rect 22899 4219 23455 4220
rect 22899 4200 23419 4219
rect 22870 4199 23419 4200
rect 23439 4199 23455 4219
rect 22870 4193 23455 4199
rect 22694 4183 22726 4184
rect 22691 4178 22726 4183
rect 22691 4158 22698 4178
rect 22718 4158 22726 4178
rect 23489 4172 23523 4378
rect 22691 4150 22726 4158
rect 20695 4137 20730 4145
rect 19798 3919 19832 4125
rect 20695 4117 20703 4137
rect 20723 4117 20730 4137
rect 20695 4112 20730 4117
rect 20695 4111 20727 4112
rect 19866 4098 20451 4104
rect 19866 4078 19882 4098
rect 19902 4097 20451 4098
rect 19902 4078 20422 4097
rect 19866 4077 20422 4078
rect 20442 4077 20451 4097
rect 19866 4069 20451 4077
rect 22073 3992 22658 4000
rect 22073 3972 22082 3992
rect 22102 3991 22658 3992
rect 22102 3972 22622 3991
rect 22073 3971 22622 3972
rect 22642 3971 22658 3991
rect 22073 3965 22658 3971
rect 22447 3941 22486 3945
rect 22692 3944 22726 4150
rect 23255 4165 23290 4171
rect 23255 4146 23260 4165
rect 23281 4146 23290 4165
rect 23255 4137 23290 4146
rect 23467 4167 23523 4172
rect 23467 4147 23474 4167
rect 23494 4147 23523 4167
rect 23467 4140 23523 4147
rect 23467 4139 23502 4140
rect 23259 4069 23288 4137
rect 23259 4035 23605 4069
rect 22447 3921 22455 3941
rect 22475 3921 22486 3941
rect 19798 3911 19833 3919
rect 19798 3891 19806 3911
rect 19826 3903 19833 3911
rect 19826 3891 19837 3903
rect 19798 3654 19837 3891
rect 20668 3868 20954 3869
rect 20153 3860 20956 3868
rect 20153 3843 20164 3860
rect 20154 3838 20164 3843
rect 20188 3843 20956 3860
rect 20188 3838 20193 3843
rect 20154 3825 20193 3838
rect 20698 3777 20733 3778
rect 20677 3770 20733 3777
rect 20677 3750 20706 3770
rect 20726 3750 20733 3770
rect 20677 3745 20733 3750
rect 20917 3768 20956 3843
rect 22447 3846 22486 3921
rect 22670 3939 22726 3944
rect 22670 3919 22677 3939
rect 22697 3919 22726 3939
rect 22670 3912 22726 3919
rect 22670 3911 22705 3912
rect 23210 3851 23249 3864
rect 23210 3846 23215 3851
rect 22447 3829 23215 3846
rect 23239 3846 23249 3851
rect 23239 3829 23250 3846
rect 22447 3821 23250 3829
rect 22449 3820 22735 3821
rect 23566 3798 23605 4035
rect 23566 3786 23577 3798
rect 23570 3778 23577 3786
rect 23597 3778 23605 3798
rect 23570 3770 23605 3778
rect 20917 3748 20928 3768
rect 20948 3748 20956 3768
rect 19798 3620 20144 3654
rect 20115 3552 20144 3620
rect 19901 3549 19936 3550
rect 19880 3542 19936 3549
rect 19880 3522 19909 3542
rect 19929 3522 19936 3542
rect 19880 3517 19936 3522
rect 20113 3543 20148 3552
rect 20113 3524 20122 3543
rect 20143 3524 20148 3543
rect 20113 3518 20148 3524
rect 20677 3539 20711 3745
rect 20917 3744 20956 3748
rect 20745 3718 21330 3724
rect 20745 3698 20761 3718
rect 20781 3717 21330 3718
rect 20781 3698 21301 3717
rect 20745 3697 21301 3698
rect 21321 3697 21330 3717
rect 20745 3689 21330 3697
rect 22952 3612 23537 3620
rect 22952 3592 22961 3612
rect 22981 3611 23537 3612
rect 22981 3592 23501 3611
rect 22952 3591 23501 3592
rect 23521 3591 23537 3611
rect 22952 3585 23537 3591
rect 22676 3577 22708 3578
rect 22673 3572 22708 3577
rect 22673 3552 22680 3572
rect 22700 3552 22708 3572
rect 23571 3564 23605 3770
rect 22673 3544 22708 3552
rect 20677 3531 20712 3539
rect 19880 3311 19914 3517
rect 20677 3511 20685 3531
rect 20705 3511 20712 3531
rect 20677 3506 20712 3511
rect 20677 3505 20709 3506
rect 19948 3490 20533 3496
rect 19948 3470 19964 3490
rect 19984 3489 20533 3490
rect 19984 3470 20504 3489
rect 19948 3469 20504 3470
rect 20524 3469 20533 3489
rect 19948 3461 20533 3469
rect 20613 3460 20643 3461
rect 20613 3433 20949 3460
rect 20613 3432 20648 3433
rect 19880 3303 19915 3311
rect 19880 3283 19888 3303
rect 19908 3283 19915 3303
rect 19880 3278 19915 3283
rect 19880 3257 19914 3278
rect 20613 3257 20643 3432
rect 20699 3365 20734 3366
rect 19880 3231 20643 3257
rect 19881 3230 19914 3231
rect 20613 3229 20643 3231
rect 20678 3358 20734 3365
rect 20678 3338 20707 3358
rect 20727 3338 20734 3358
rect 20678 3333 20734 3338
rect 20913 3360 20948 3433
rect 20913 3340 20920 3360
rect 20940 3340 20948 3360
rect 22055 3386 22640 3394
rect 22055 3366 22064 3386
rect 22084 3385 22640 3386
rect 22084 3366 22604 3385
rect 22055 3365 22604 3366
rect 22624 3365 22640 3385
rect 22055 3359 22640 3365
rect 20913 3333 20948 3340
rect 22674 3338 22708 3544
rect 23339 3558 23370 3564
rect 23339 3539 23344 3558
rect 23365 3539 23370 3558
rect 23339 3497 23370 3539
rect 23549 3559 23605 3564
rect 23549 3539 23556 3559
rect 23576 3539 23605 3559
rect 23549 3532 23605 3539
rect 23549 3531 23584 3532
rect 23339 3469 23678 3497
rect 19622 3174 19976 3210
rect 19638 3173 19976 3174
rect 19950 3143 19976 3173
rect 19736 3141 19771 3142
rect 19715 3134 19771 3141
rect 19715 3114 19744 3134
rect 19764 3114 19771 3134
rect 19715 3109 19771 3114
rect 19944 3135 19985 3143
rect 19944 3117 19957 3135
rect 19975 3117 19985 3135
rect 19715 2903 19749 3109
rect 19944 3106 19985 3117
rect 20678 3127 20712 3333
rect 22438 3331 22473 3338
rect 20746 3306 21331 3312
rect 20746 3286 20762 3306
rect 20782 3305 21331 3306
rect 20782 3286 21302 3305
rect 20746 3285 21302 3286
rect 21322 3285 21331 3305
rect 20746 3277 21331 3285
rect 22438 3311 22446 3331
rect 22466 3311 22473 3331
rect 22438 3238 22473 3311
rect 22652 3333 22708 3338
rect 22652 3313 22659 3333
rect 22679 3313 22708 3333
rect 22652 3306 22708 3313
rect 22743 3440 22773 3442
rect 23472 3440 23505 3441
rect 22743 3414 23506 3440
rect 22652 3305 22687 3306
rect 22743 3239 22773 3414
rect 23472 3393 23506 3414
rect 23471 3388 23506 3393
rect 23471 3368 23478 3388
rect 23498 3368 23506 3388
rect 23471 3360 23506 3368
rect 22738 3238 22773 3239
rect 22437 3211 22773 3238
rect 22743 3210 22773 3211
rect 22853 3202 23438 3210
rect 22853 3182 22862 3202
rect 22882 3201 23438 3202
rect 22882 3182 23402 3201
rect 22853 3181 23402 3182
rect 23422 3181 23438 3201
rect 22853 3175 23438 3181
rect 22677 3165 22709 3166
rect 22674 3160 22709 3165
rect 22674 3140 22681 3160
rect 22701 3140 22709 3160
rect 23472 3154 23506 3360
rect 22674 3132 22709 3140
rect 20678 3119 20713 3127
rect 20678 3099 20686 3119
rect 20706 3099 20713 3119
rect 20678 3094 20713 3099
rect 20678 3093 20710 3094
rect 19783 3082 20368 3088
rect 19783 3062 19799 3082
rect 19819 3081 20368 3082
rect 19819 3062 20339 3081
rect 19783 3061 20339 3062
rect 20359 3061 20368 3081
rect 19783 3053 20368 3061
rect 22056 2974 22641 2982
rect 22056 2954 22065 2974
rect 22085 2973 22641 2974
rect 22085 2954 22605 2973
rect 22056 2953 22605 2954
rect 22625 2953 22641 2973
rect 22056 2947 22641 2953
rect 22430 2923 22469 2927
rect 22675 2926 22709 3132
rect 23239 3144 23273 3152
rect 23239 3126 23246 3144
rect 23265 3126 23273 3144
rect 23239 3119 23273 3126
rect 23450 3149 23506 3154
rect 23450 3129 23457 3149
rect 23477 3129 23506 3149
rect 23450 3122 23506 3129
rect 23450 3121 23485 3122
rect 23243 3089 23272 3119
rect 23243 3081 23625 3089
rect 23243 3062 23596 3081
rect 23617 3062 23625 3081
rect 23243 3057 23625 3062
rect 22430 2903 22438 2923
rect 22458 2903 22469 2923
rect 19715 2902 19750 2903
rect 19683 2895 19750 2902
rect 19683 2875 19723 2895
rect 19743 2875 19750 2895
rect 19683 2872 19750 2875
rect 19683 2869 19748 2872
rect 19254 2768 19319 2771
rect 15475 2617 15857 2622
rect 15475 2598 15483 2617
rect 15504 2598 15857 2617
rect 15475 2590 15857 2598
rect 15828 2560 15857 2590
rect 15615 2557 15650 2558
rect 15594 2550 15650 2557
rect 15594 2530 15623 2550
rect 15643 2530 15650 2550
rect 15594 2525 15650 2530
rect 15827 2553 15861 2560
rect 15827 2535 15835 2553
rect 15854 2535 15861 2553
rect 15827 2527 15861 2535
rect 16391 2547 16425 2753
rect 16631 2752 16670 2756
rect 19252 2765 19319 2768
rect 19252 2745 19259 2765
rect 19279 2745 19319 2765
rect 19252 2738 19319 2745
rect 19252 2737 19287 2738
rect 16459 2726 17044 2732
rect 16459 2706 16475 2726
rect 16495 2725 17044 2726
rect 16495 2706 17015 2725
rect 16459 2705 17015 2706
rect 17035 2705 17044 2725
rect 16459 2697 17044 2705
rect 18634 2579 19219 2587
rect 18634 2559 18643 2579
rect 18663 2578 19219 2579
rect 18663 2559 19183 2578
rect 18634 2558 19183 2559
rect 19203 2558 19219 2578
rect 18634 2552 19219 2558
rect 16391 2539 16426 2547
rect 18292 2546 18324 2547
rect 15594 2319 15628 2525
rect 16391 2519 16399 2539
rect 16419 2519 16426 2539
rect 16391 2514 16426 2519
rect 18289 2541 18324 2546
rect 18289 2521 18296 2541
rect 18316 2521 18324 2541
rect 16391 2513 16423 2514
rect 18289 2513 18324 2521
rect 15662 2498 16247 2504
rect 15662 2478 15678 2498
rect 15698 2497 16247 2498
rect 15698 2478 16218 2497
rect 15662 2477 16218 2478
rect 16238 2477 16247 2497
rect 15662 2469 16247 2477
rect 16327 2468 16357 2469
rect 16327 2441 16663 2468
rect 16327 2440 16362 2441
rect 15594 2311 15629 2319
rect 15594 2291 15602 2311
rect 15622 2291 15629 2311
rect 15594 2286 15629 2291
rect 15594 2265 15628 2286
rect 16327 2265 16357 2440
rect 16413 2373 16448 2374
rect 15594 2239 16357 2265
rect 15595 2238 15628 2239
rect 16327 2237 16357 2239
rect 16392 2366 16448 2373
rect 16392 2346 16421 2366
rect 16441 2346 16448 2366
rect 16392 2341 16448 2346
rect 16627 2368 16662 2441
rect 16627 2348 16634 2368
rect 16654 2348 16662 2368
rect 16627 2341 16662 2348
rect 17671 2355 18256 2363
rect 15422 2182 15761 2210
rect 15516 2147 15551 2148
rect 15495 2140 15551 2147
rect 15495 2120 15524 2140
rect 15544 2120 15551 2140
rect 15495 2115 15551 2120
rect 15730 2140 15761 2182
rect 15730 2121 15735 2140
rect 15756 2121 15761 2140
rect 15730 2115 15761 2121
rect 16392 2135 16426 2341
rect 17671 2335 17680 2355
rect 17700 2354 18256 2355
rect 17700 2335 18220 2354
rect 17671 2334 18220 2335
rect 18240 2334 18256 2354
rect 17671 2328 18256 2334
rect 16460 2314 17045 2320
rect 16460 2294 16476 2314
rect 16496 2313 17045 2314
rect 16496 2294 17016 2313
rect 16460 2293 17016 2294
rect 17036 2293 17045 2313
rect 18290 2307 18324 2513
rect 19019 2528 19052 2534
rect 19253 2531 19287 2737
rect 19019 2506 19024 2528
rect 19047 2506 19052 2528
rect 19019 2497 19052 2506
rect 19231 2526 19287 2531
rect 19231 2506 19238 2526
rect 19258 2506 19287 2526
rect 19231 2499 19287 2506
rect 19231 2498 19266 2499
rect 19021 2466 19048 2497
rect 19443 2466 19482 2478
rect 19021 2465 19484 2466
rect 19021 2443 19448 2465
rect 19472 2443 19484 2465
rect 19021 2435 19484 2443
rect 16460 2285 17045 2293
rect 18054 2300 18089 2307
rect 18054 2280 18062 2300
rect 18082 2280 18089 2300
rect 18054 2207 18089 2280
rect 18268 2302 18324 2307
rect 18268 2282 18275 2302
rect 18295 2282 18324 2302
rect 18268 2275 18324 2282
rect 18359 2409 18389 2411
rect 19088 2409 19121 2410
rect 18359 2383 19122 2409
rect 18268 2274 18303 2275
rect 18359 2208 18389 2383
rect 19088 2362 19122 2383
rect 19087 2357 19122 2362
rect 19087 2337 19094 2357
rect 19114 2337 19122 2357
rect 19087 2329 19122 2337
rect 18354 2207 18389 2208
rect 18053 2180 18389 2207
rect 18359 2179 18389 2180
rect 18469 2171 19054 2179
rect 18469 2151 18478 2171
rect 18498 2170 19054 2171
rect 18498 2151 19018 2170
rect 18469 2150 19018 2151
rect 19038 2150 19054 2170
rect 18469 2144 19054 2150
rect 16392 2127 16427 2135
rect 18293 2134 18325 2135
rect 15495 1909 15529 2115
rect 16392 2107 16400 2127
rect 16420 2107 16427 2127
rect 16392 2102 16427 2107
rect 18290 2129 18325 2134
rect 18290 2109 18297 2129
rect 18317 2109 18325 2129
rect 19088 2123 19122 2329
rect 16392 2101 16424 2102
rect 18290 2101 18325 2109
rect 15563 2088 16148 2094
rect 15563 2068 15579 2088
rect 15599 2087 16148 2088
rect 15599 2068 16119 2087
rect 15563 2067 16119 2068
rect 16139 2067 16148 2087
rect 15563 2059 16148 2067
rect 17672 1943 18257 1951
rect 17672 1923 17681 1943
rect 17701 1942 18257 1943
rect 17701 1923 18221 1942
rect 17672 1922 18221 1923
rect 18241 1922 18257 1942
rect 17672 1916 18257 1922
rect 15495 1901 15530 1909
rect 15495 1881 15503 1901
rect 15523 1893 15530 1901
rect 15523 1881 15534 1893
rect 15495 1644 15534 1881
rect 18046 1892 18085 1896
rect 18291 1895 18325 2101
rect 18854 2116 18889 2122
rect 18854 2097 18859 2116
rect 18880 2097 18889 2116
rect 18854 2088 18889 2097
rect 19066 2118 19122 2123
rect 19066 2098 19073 2118
rect 19093 2098 19122 2118
rect 19066 2091 19122 2098
rect 19244 2269 19276 2281
rect 19244 2251 19251 2269
rect 19273 2251 19276 2269
rect 19066 2090 19101 2091
rect 18858 2020 18887 2088
rect 18858 1986 19204 2020
rect 18046 1872 18054 1892
rect 18074 1872 18085 1892
rect 16365 1858 16651 1859
rect 15850 1850 16653 1858
rect 15850 1833 15861 1850
rect 15851 1828 15861 1833
rect 15885 1833 16653 1850
rect 15885 1828 15890 1833
rect 15851 1815 15890 1828
rect 16395 1767 16430 1768
rect 16374 1760 16430 1767
rect 16374 1740 16403 1760
rect 16423 1740 16430 1760
rect 16374 1735 16430 1740
rect 16614 1758 16653 1833
rect 18046 1797 18085 1872
rect 18269 1890 18325 1895
rect 18269 1870 18276 1890
rect 18296 1870 18325 1890
rect 18269 1863 18325 1870
rect 18269 1862 18304 1863
rect 18809 1802 18848 1815
rect 18809 1797 18814 1802
rect 18046 1780 18814 1797
rect 18838 1797 18848 1802
rect 18838 1780 18849 1797
rect 18046 1772 18849 1780
rect 18048 1771 18334 1772
rect 16614 1738 16625 1758
rect 16645 1738 16653 1758
rect 15495 1610 15841 1644
rect 15812 1542 15841 1610
rect 15598 1539 15633 1540
rect 14676 1440 15010 1468
rect 15577 1532 15633 1539
rect 15577 1512 15606 1532
rect 15626 1512 15633 1532
rect 15577 1507 15633 1512
rect 15810 1533 15845 1542
rect 15810 1514 15819 1533
rect 15840 1514 15845 1533
rect 15810 1508 15845 1514
rect 16374 1529 16408 1735
rect 16614 1734 16653 1738
rect 19165 1749 19204 1986
rect 19165 1737 19176 1749
rect 19169 1729 19176 1737
rect 19196 1729 19204 1749
rect 19169 1721 19204 1729
rect 16442 1708 17027 1714
rect 16442 1688 16458 1708
rect 16478 1707 17027 1708
rect 16478 1688 16998 1707
rect 16442 1687 16998 1688
rect 17018 1687 17027 1707
rect 16442 1679 17027 1687
rect 18551 1563 19136 1571
rect 18551 1543 18560 1563
rect 18580 1562 19136 1563
rect 18580 1543 19100 1562
rect 18551 1542 19100 1543
rect 19120 1542 19136 1562
rect 18551 1536 19136 1542
rect 16374 1521 16409 1529
rect 18275 1528 18307 1529
rect 9643 1096 9678 1104
rect 7634 1084 7669 1092
rect 6042 1073 6077 1074
rect 5835 1041 5864 1071
rect 7634 1064 7642 1084
rect 7662 1064 7669 1084
rect 7634 1059 7669 1064
rect 7634 1058 7666 1059
rect 5835 1033 6217 1041
rect 5835 1014 6188 1033
rect 6209 1014 6217 1033
rect 5835 1009 6217 1014
rect 9025 938 9610 946
rect 9025 918 9034 938
rect 9054 937 9610 938
rect 9054 918 9574 937
rect 9025 917 9574 918
rect 9594 917 9610 937
rect 9025 911 9610 917
rect 5022 855 5030 875
rect 5050 855 5061 875
rect 881 832 916 833
rect 2116 785 2167 816
rect 1421 772 1460 785
rect 1421 767 1426 772
rect 658 750 1426 767
rect 1450 767 1460 772
rect 1450 750 1461 767
rect 658 742 1461 750
rect 2116 759 2133 785
rect 2161 759 2167 785
rect 660 741 946 742
rect 2116 736 2167 759
rect 2196 791 2242 822
rect 4040 820 4083 828
rect 2196 760 2210 791
rect 2238 760 2242 791
rect 2196 753 2242 760
rect 4034 813 4089 820
rect 4034 788 4047 813
rect 4079 788 4089 813
rect 498 725 559 734
rect 498 698 506 725
rect 542 719 559 725
rect 600 719 675 723
rect 542 717 675 719
rect 542 698 606 717
rect 498 681 606 698
rect 651 681 675 717
rect 498 679 675 681
rect 600 649 675 679
rect 2129 544 2160 736
rect 2115 523 2161 544
rect 2115 502 2122 523
rect 2143 502 2161 523
rect 2115 498 2161 502
rect 2115 495 2150 498
rect 1497 337 2082 345
rect 1497 317 1506 337
rect 1526 336 2082 337
rect 1526 317 2046 336
rect 1497 316 2046 317
rect 2066 316 2082 336
rect 1497 310 2082 316
rect 2116 289 2150 495
rect 2198 429 2232 753
rect 4034 696 4089 788
rect 5022 780 5061 855
rect 5245 873 5301 878
rect 5245 853 5252 873
rect 5272 853 5301 873
rect 5245 846 5301 853
rect 9399 887 9438 891
rect 9644 890 9678 1096
rect 10208 1108 10242 1116
rect 10208 1090 10215 1108
rect 10234 1090 10242 1108
rect 10208 1083 10242 1090
rect 10419 1113 10475 1118
rect 10419 1093 10426 1113
rect 10446 1093 10475 1113
rect 10419 1086 10475 1093
rect 12011 1104 12045 1310
rect 13771 1308 13806 1315
rect 12079 1283 12664 1289
rect 12079 1263 12095 1283
rect 12115 1282 12664 1283
rect 12115 1263 12635 1282
rect 12079 1262 12635 1263
rect 12655 1262 12664 1282
rect 12079 1254 12664 1262
rect 13771 1288 13779 1308
rect 13799 1288 13806 1308
rect 13771 1215 13806 1288
rect 13985 1310 14041 1315
rect 13985 1290 13992 1310
rect 14012 1290 14041 1310
rect 13985 1283 14041 1290
rect 14076 1417 14106 1419
rect 14805 1417 14838 1418
rect 14076 1391 14839 1417
rect 13985 1282 14020 1283
rect 14076 1216 14106 1391
rect 14805 1370 14839 1391
rect 14804 1365 14839 1370
rect 14804 1345 14811 1365
rect 14831 1345 14839 1365
rect 14804 1337 14839 1345
rect 14071 1215 14106 1216
rect 13770 1188 14106 1215
rect 14076 1187 14106 1188
rect 14186 1179 14771 1187
rect 14186 1159 14195 1179
rect 14215 1178 14771 1179
rect 14215 1159 14735 1178
rect 14186 1158 14735 1159
rect 14755 1158 14771 1178
rect 14186 1152 14771 1158
rect 14010 1142 14042 1143
rect 14007 1137 14042 1142
rect 14007 1117 14014 1137
rect 14034 1117 14042 1137
rect 14805 1131 14839 1337
rect 15577 1301 15611 1507
rect 16374 1501 16382 1521
rect 16402 1501 16409 1521
rect 16374 1496 16409 1501
rect 18272 1523 18307 1528
rect 18272 1503 18279 1523
rect 18299 1503 18307 1523
rect 19170 1515 19204 1721
rect 16374 1495 16406 1496
rect 18272 1495 18307 1503
rect 15645 1480 16230 1486
rect 15645 1460 15661 1480
rect 15681 1479 16230 1480
rect 15681 1460 16201 1479
rect 15645 1459 16201 1460
rect 16221 1459 16230 1479
rect 15645 1451 16230 1459
rect 16310 1450 16340 1451
rect 16310 1423 16646 1450
rect 16310 1422 16345 1423
rect 15577 1293 15612 1301
rect 15577 1273 15585 1293
rect 15605 1273 15612 1293
rect 15577 1268 15612 1273
rect 15577 1247 15611 1268
rect 16310 1247 16340 1422
rect 16396 1355 16431 1356
rect 15577 1221 16340 1247
rect 15578 1220 15611 1221
rect 16310 1219 16340 1221
rect 16375 1348 16431 1355
rect 16375 1328 16404 1348
rect 16424 1328 16431 1348
rect 16375 1323 16431 1328
rect 16610 1350 16645 1423
rect 16610 1330 16617 1350
rect 16637 1330 16645 1350
rect 16610 1323 16645 1330
rect 17654 1337 18239 1345
rect 14007 1109 14042 1117
rect 12011 1096 12046 1104
rect 10419 1085 10454 1086
rect 10212 1053 10241 1083
rect 12011 1076 12019 1096
rect 12039 1076 12046 1096
rect 12011 1071 12046 1076
rect 12011 1070 12043 1071
rect 10212 1045 10594 1053
rect 10212 1026 10565 1045
rect 10586 1026 10594 1045
rect 10212 1021 10594 1026
rect 13389 951 13974 959
rect 13389 931 13398 951
rect 13418 950 13974 951
rect 13418 931 13938 950
rect 13389 930 13938 931
rect 13958 930 13974 950
rect 13389 924 13974 930
rect 9399 867 9407 887
rect 9427 867 9438 887
rect 5245 845 5280 846
rect 6480 798 6531 829
rect 5785 785 5824 798
rect 5785 780 5790 785
rect 5022 763 5790 780
rect 5814 780 5824 785
rect 5814 763 5825 780
rect 5022 755 5825 763
rect 6480 772 6497 798
rect 6525 772 6531 798
rect 5024 754 5310 755
rect 6480 749 6531 772
rect 6560 804 6606 835
rect 8404 833 8447 841
rect 6560 773 6574 804
rect 6602 773 6606 804
rect 6560 766 6606 773
rect 8398 826 8453 833
rect 8398 801 8411 826
rect 8443 801 8453 826
rect 4034 664 4045 696
rect 4085 664 4089 696
rect 4862 738 4923 747
rect 4862 711 4870 738
rect 4906 732 4923 738
rect 4964 732 5039 736
rect 4906 730 5039 732
rect 4906 711 4970 730
rect 4862 694 4970 711
rect 5015 694 5039 730
rect 4862 692 5039 694
rect 4034 651 4089 664
rect 4964 662 5039 692
rect 6493 557 6524 749
rect 6479 536 6525 557
rect 6479 515 6486 536
rect 6507 515 6525 536
rect 6479 511 6525 515
rect 6479 508 6514 511
rect 4618 471 4649 476
rect 2198 409 2204 429
rect 2224 409 2232 429
rect 2198 403 2232 409
rect 3820 451 4654 471
rect 1877 283 1920 287
rect 1877 259 1888 283
rect 1911 259 1920 283
rect 1877 255 1920 259
rect 2094 284 2150 289
rect 2094 264 2101 284
rect 2121 264 2150 284
rect 2094 257 2150 264
rect 2094 256 2129 257
rect 1884 191 1915 255
rect 3820 191 3846 451
rect 4604 449 4650 451
rect 4604 428 4611 449
rect 4632 428 4650 449
rect 4684 441 5777 474
rect 4604 424 4650 428
rect 4604 421 4639 424
rect 3986 263 4571 271
rect 3986 243 3995 263
rect 4015 262 4571 263
rect 4015 243 4535 262
rect 3986 242 4535 243
rect 4555 242 4571 262
rect 3986 236 4571 242
rect 4605 215 4639 421
rect 4686 355 4729 441
rect 4686 335 4693 355
rect 4713 335 4729 355
rect 4686 324 4729 335
rect 4583 210 4639 215
rect 4373 205 4405 210
rect 1884 168 3847 191
rect 1892 166 3847 168
rect 4373 184 4380 205
rect 4397 184 4405 205
rect 4373 177 4405 184
rect 4583 190 4590 210
rect 4610 190 4639 210
rect 4583 183 4639 190
rect 5746 198 5775 441
rect 5861 350 6446 358
rect 5861 330 5870 350
rect 5890 349 6446 350
rect 5890 330 6410 349
rect 5861 329 6410 330
rect 6430 329 6446 349
rect 5861 323 6446 329
rect 6243 303 6286 305
rect 6239 297 6290 303
rect 6480 302 6514 508
rect 6562 442 6596 766
rect 8398 709 8453 801
rect 9399 792 9438 867
rect 9622 885 9678 890
rect 9622 865 9629 885
rect 9649 865 9678 885
rect 9622 858 9678 865
rect 13763 900 13802 904
rect 14008 903 14042 1109
rect 14572 1121 14606 1129
rect 14572 1103 14579 1121
rect 14598 1103 14606 1121
rect 14572 1096 14606 1103
rect 14783 1126 14839 1131
rect 14783 1106 14790 1126
rect 14810 1106 14839 1126
rect 14783 1099 14839 1106
rect 16375 1117 16409 1323
rect 17654 1317 17663 1337
rect 17683 1336 18239 1337
rect 17683 1317 18203 1336
rect 17654 1316 18203 1317
rect 18223 1316 18239 1336
rect 17654 1310 18239 1316
rect 16443 1296 17028 1302
rect 16443 1276 16459 1296
rect 16479 1295 17028 1296
rect 16479 1276 16999 1295
rect 16443 1275 16999 1276
rect 17019 1275 17028 1295
rect 18273 1289 18307 1495
rect 18936 1503 18972 1512
rect 18936 1486 18945 1503
rect 18964 1486 18972 1503
rect 18936 1477 18972 1486
rect 19148 1510 19204 1515
rect 19148 1490 19155 1510
rect 19175 1490 19204 1510
rect 19148 1483 19204 1490
rect 19148 1482 19183 1483
rect 18942 1442 18968 1477
rect 19244 1442 19276 2251
rect 19688 2184 19717 2869
rect 20648 2850 20934 2851
rect 20133 2842 20936 2850
rect 20133 2825 20144 2842
rect 20134 2820 20144 2825
rect 20168 2825 20936 2842
rect 20168 2820 20173 2825
rect 20134 2807 20173 2820
rect 20678 2759 20713 2760
rect 20657 2752 20713 2759
rect 20657 2732 20686 2752
rect 20706 2732 20713 2752
rect 20657 2727 20713 2732
rect 20897 2750 20936 2825
rect 22430 2828 22469 2903
rect 22653 2921 22709 2926
rect 22653 2901 22660 2921
rect 22680 2901 22709 2921
rect 22653 2894 22709 2901
rect 22653 2893 22688 2894
rect 23193 2833 23232 2846
rect 23193 2828 23198 2833
rect 22430 2811 23198 2828
rect 23222 2828 23232 2833
rect 23222 2811 23233 2828
rect 22430 2803 23233 2811
rect 22432 2802 22718 2803
rect 23649 2784 23678 3469
rect 23986 3223 24013 4923
rect 26843 4951 26851 4971
rect 26871 4951 26882 4971
rect 25049 4899 25335 4900
rect 24534 4891 25337 4899
rect 24534 4874 24545 4891
rect 24535 4869 24545 4874
rect 24569 4874 25337 4891
rect 24569 4869 24574 4874
rect 24535 4856 24574 4869
rect 25079 4808 25114 4809
rect 25058 4801 25114 4808
rect 25058 4781 25087 4801
rect 25107 4781 25114 4801
rect 25058 4776 25114 4781
rect 25298 4799 25337 4874
rect 26843 4876 26882 4951
rect 27066 4969 27122 4974
rect 27066 4949 27073 4969
rect 27093 4949 27122 4969
rect 27066 4942 27122 4949
rect 27066 4941 27101 4942
rect 27606 4881 27645 4894
rect 27606 4876 27611 4881
rect 26843 4859 27611 4876
rect 27635 4876 27645 4881
rect 27635 4859 27646 4876
rect 26843 4851 27646 4859
rect 26845 4850 27131 4851
rect 25298 4779 25309 4799
rect 25329 4779 25337 4799
rect 28167 4827 28194 6527
rect 28502 6281 28531 6966
rect 29462 6947 29748 6948
rect 28947 6939 29750 6947
rect 28947 6922 28958 6939
rect 28948 6917 28958 6922
rect 28982 6922 29750 6939
rect 28982 6917 28987 6922
rect 28948 6904 28987 6917
rect 29492 6856 29527 6857
rect 29471 6849 29527 6856
rect 29471 6829 29500 6849
rect 29520 6829 29527 6849
rect 29471 6824 29527 6829
rect 29711 6847 29750 6922
rect 31244 6925 31283 7000
rect 31467 7018 31523 7023
rect 31467 6998 31474 7018
rect 31494 6998 31523 7018
rect 31467 6991 31523 6998
rect 31467 6990 31502 6991
rect 32007 6930 32046 6943
rect 32007 6925 32012 6930
rect 31244 6908 32012 6925
rect 32036 6925 32046 6930
rect 32036 6908 32047 6925
rect 31244 6900 32047 6908
rect 31246 6899 31532 6900
rect 32463 6881 32492 7566
rect 32904 7499 32936 8308
rect 33212 8273 33238 8308
rect 32997 8267 33032 8268
rect 32976 8260 33032 8267
rect 32976 8240 33005 8260
rect 33025 8240 33032 8260
rect 32976 8235 33032 8240
rect 33208 8264 33244 8273
rect 33208 8247 33216 8264
rect 33235 8247 33244 8264
rect 33208 8238 33244 8247
rect 33873 8255 33907 8461
rect 33941 8434 34526 8440
rect 33941 8414 33957 8434
rect 33977 8433 34526 8434
rect 33977 8414 34497 8433
rect 33941 8413 34497 8414
rect 34517 8413 34526 8433
rect 33941 8405 34526 8413
rect 33873 8247 33908 8255
rect 32976 8029 33010 8235
rect 33873 8227 33881 8247
rect 33901 8227 33908 8247
rect 33873 8222 33908 8227
rect 33873 8221 33905 8222
rect 33044 8208 33629 8214
rect 33044 8188 33060 8208
rect 33080 8207 33629 8208
rect 33080 8188 33600 8207
rect 33044 8187 33600 8188
rect 33620 8187 33629 8207
rect 33044 8179 33629 8187
rect 32976 8021 33011 8029
rect 32976 8001 32984 8021
rect 33004 8013 33011 8021
rect 33004 8001 33015 8013
rect 32976 7764 33015 8001
rect 33846 7978 34132 7979
rect 33331 7970 34134 7978
rect 33331 7953 33342 7970
rect 33332 7948 33342 7953
rect 33366 7953 34134 7970
rect 33366 7948 33371 7953
rect 33332 7935 33371 7948
rect 33876 7887 33911 7888
rect 33855 7880 33911 7887
rect 33855 7860 33884 7880
rect 33904 7860 33911 7880
rect 33855 7855 33911 7860
rect 34095 7878 34134 7953
rect 34095 7858 34106 7878
rect 34126 7858 34134 7878
rect 32976 7730 33322 7764
rect 33293 7662 33322 7730
rect 33079 7659 33114 7660
rect 32904 7481 32907 7499
rect 32929 7481 32936 7499
rect 32904 7469 32936 7481
rect 33058 7652 33114 7659
rect 33058 7632 33087 7652
rect 33107 7632 33114 7652
rect 33058 7627 33114 7632
rect 33291 7653 33326 7662
rect 33291 7634 33300 7653
rect 33321 7634 33326 7653
rect 33291 7628 33326 7634
rect 33855 7649 33889 7855
rect 34095 7854 34134 7858
rect 33923 7828 34508 7834
rect 33923 7808 33939 7828
rect 33959 7827 34508 7828
rect 33959 7808 34479 7827
rect 33923 7807 34479 7808
rect 34499 7807 34508 7827
rect 33923 7799 34508 7807
rect 33855 7641 33890 7649
rect 33058 7421 33092 7627
rect 33855 7621 33863 7641
rect 33883 7621 33890 7641
rect 33855 7616 33890 7621
rect 33855 7615 33887 7616
rect 33126 7600 33711 7606
rect 33126 7580 33142 7600
rect 33162 7599 33711 7600
rect 33162 7580 33682 7599
rect 33126 7579 33682 7580
rect 33702 7579 33711 7599
rect 33126 7571 33711 7579
rect 33791 7570 33821 7571
rect 33791 7543 34127 7570
rect 33791 7542 33826 7543
rect 33058 7413 33093 7421
rect 33058 7393 33066 7413
rect 33086 7393 33093 7413
rect 33058 7388 33093 7393
rect 33058 7367 33092 7388
rect 33791 7367 33821 7542
rect 33877 7475 33912 7476
rect 33058 7341 33821 7367
rect 33059 7340 33092 7341
rect 33791 7339 33821 7341
rect 33856 7468 33912 7475
rect 33856 7448 33885 7468
rect 33905 7448 33912 7468
rect 33856 7443 33912 7448
rect 34091 7470 34126 7543
rect 34091 7450 34098 7470
rect 34118 7450 34126 7470
rect 34091 7443 34126 7450
rect 32696 7307 33159 7315
rect 32696 7285 32708 7307
rect 32732 7285 33159 7307
rect 32696 7284 33159 7285
rect 32698 7272 32737 7284
rect 33132 7253 33159 7284
rect 32914 7251 32949 7252
rect 32893 7244 32949 7251
rect 32893 7224 32922 7244
rect 32942 7224 32949 7244
rect 32893 7219 32949 7224
rect 33128 7244 33161 7253
rect 33128 7222 33133 7244
rect 33156 7222 33161 7244
rect 32893 7013 32927 7219
rect 33128 7216 33161 7222
rect 33856 7237 33890 7443
rect 33924 7416 34509 7422
rect 33924 7396 33940 7416
rect 33960 7415 34509 7416
rect 33960 7396 34480 7415
rect 33924 7395 34480 7396
rect 34500 7395 34509 7415
rect 33924 7387 34509 7395
rect 33856 7229 33891 7237
rect 33856 7209 33864 7229
rect 33884 7209 33891 7229
rect 33856 7204 33891 7209
rect 33856 7203 33888 7204
rect 32961 7192 33546 7198
rect 32961 7172 32977 7192
rect 32997 7191 33546 7192
rect 32997 7172 33517 7191
rect 32961 7171 33517 7172
rect 33537 7171 33546 7191
rect 32961 7163 33546 7171
rect 32893 7012 32928 7013
rect 32861 7005 32928 7012
rect 32861 6985 32901 7005
rect 32921 6985 32928 7005
rect 32861 6982 32928 6985
rect 32861 6979 32926 6982
rect 32432 6878 32497 6881
rect 32430 6875 32497 6878
rect 32430 6855 32437 6875
rect 32457 6855 32497 6875
rect 32430 6848 32497 6855
rect 32430 6847 32465 6848
rect 29711 6827 29722 6847
rect 29742 6827 29750 6847
rect 28555 6688 28937 6693
rect 28555 6669 28563 6688
rect 28584 6669 28937 6688
rect 28555 6661 28937 6669
rect 28908 6631 28937 6661
rect 28695 6628 28730 6629
rect 28674 6621 28730 6628
rect 28674 6601 28703 6621
rect 28723 6601 28730 6621
rect 28674 6596 28730 6601
rect 28907 6624 28941 6631
rect 28907 6606 28915 6624
rect 28934 6606 28941 6624
rect 28907 6598 28941 6606
rect 29471 6618 29505 6824
rect 29711 6823 29750 6827
rect 29539 6797 30124 6803
rect 29539 6777 29555 6797
rect 29575 6796 30124 6797
rect 29575 6777 30095 6796
rect 29539 6776 30095 6777
rect 30115 6776 30124 6796
rect 29539 6768 30124 6776
rect 31812 6689 32397 6697
rect 31812 6669 31821 6689
rect 31841 6688 32397 6689
rect 31841 6669 32361 6688
rect 31812 6668 32361 6669
rect 32381 6668 32397 6688
rect 31812 6662 32397 6668
rect 31470 6656 31502 6657
rect 31467 6651 31502 6656
rect 31467 6631 31474 6651
rect 31494 6631 31502 6651
rect 31467 6623 31502 6631
rect 29471 6610 29506 6618
rect 28674 6390 28708 6596
rect 29471 6590 29479 6610
rect 29499 6590 29506 6610
rect 29471 6585 29506 6590
rect 29471 6584 29503 6585
rect 28742 6569 29327 6575
rect 28742 6549 28758 6569
rect 28778 6568 29327 6569
rect 28778 6549 29298 6568
rect 28742 6548 29298 6549
rect 29318 6548 29327 6568
rect 28742 6540 29327 6548
rect 29407 6539 29437 6540
rect 29407 6512 29743 6539
rect 29407 6511 29442 6512
rect 28674 6382 28709 6390
rect 28674 6362 28682 6382
rect 28702 6362 28709 6382
rect 28674 6357 28709 6362
rect 28674 6336 28708 6357
rect 29407 6336 29437 6511
rect 29493 6444 29528 6445
rect 28674 6310 29437 6336
rect 28675 6309 28708 6310
rect 29407 6308 29437 6310
rect 29472 6437 29528 6444
rect 29472 6417 29501 6437
rect 29521 6417 29528 6437
rect 29472 6412 29528 6417
rect 29707 6439 29742 6512
rect 29707 6419 29714 6439
rect 29734 6419 29742 6439
rect 30849 6465 31434 6473
rect 30849 6445 30858 6465
rect 30878 6464 31434 6465
rect 30878 6445 31398 6464
rect 30849 6444 31398 6445
rect 31418 6444 31434 6464
rect 30849 6438 31434 6444
rect 29707 6412 29742 6419
rect 31468 6417 31502 6623
rect 32195 6633 32236 6644
rect 32431 6641 32465 6847
rect 32195 6615 32205 6633
rect 32223 6615 32236 6633
rect 32195 6607 32236 6615
rect 32409 6636 32465 6641
rect 32409 6616 32416 6636
rect 32436 6616 32465 6636
rect 32409 6609 32465 6616
rect 32409 6608 32444 6609
rect 32204 6577 32230 6607
rect 32204 6576 32542 6577
rect 32204 6540 32558 6576
rect 28502 6253 28841 6281
rect 28596 6218 28631 6219
rect 28575 6211 28631 6218
rect 28575 6191 28604 6211
rect 28624 6191 28631 6211
rect 28575 6186 28631 6191
rect 28810 6211 28841 6253
rect 28810 6192 28815 6211
rect 28836 6192 28841 6211
rect 28810 6186 28841 6192
rect 29472 6206 29506 6412
rect 31232 6410 31267 6417
rect 29540 6385 30125 6391
rect 29540 6365 29556 6385
rect 29576 6384 30125 6385
rect 29576 6365 30096 6384
rect 29540 6364 30096 6365
rect 30116 6364 30125 6384
rect 29540 6356 30125 6364
rect 31232 6390 31240 6410
rect 31260 6390 31267 6410
rect 31232 6317 31267 6390
rect 31446 6412 31502 6417
rect 31446 6392 31453 6412
rect 31473 6392 31502 6412
rect 31446 6385 31502 6392
rect 31537 6519 31567 6521
rect 32266 6519 32299 6520
rect 31537 6493 32300 6519
rect 31446 6384 31481 6385
rect 31537 6318 31567 6493
rect 32266 6472 32300 6493
rect 32265 6467 32300 6472
rect 32265 6447 32272 6467
rect 32292 6447 32300 6467
rect 32265 6439 32300 6447
rect 31532 6317 31567 6318
rect 31231 6290 31567 6317
rect 31537 6289 31567 6290
rect 31647 6281 32232 6289
rect 31647 6261 31656 6281
rect 31676 6280 32232 6281
rect 31676 6261 32196 6280
rect 31647 6260 32196 6261
rect 32216 6260 32232 6280
rect 31647 6254 32232 6260
rect 31471 6244 31503 6245
rect 31468 6239 31503 6244
rect 31468 6219 31475 6239
rect 31495 6219 31503 6239
rect 32266 6233 32300 6439
rect 31468 6211 31503 6219
rect 29472 6198 29507 6206
rect 28575 5980 28609 6186
rect 29472 6178 29480 6198
rect 29500 6178 29507 6198
rect 29472 6173 29507 6178
rect 29472 6172 29504 6173
rect 28643 6159 29228 6165
rect 28643 6139 28659 6159
rect 28679 6158 29228 6159
rect 28679 6139 29199 6158
rect 28643 6138 29199 6139
rect 29219 6138 29228 6158
rect 28643 6130 29228 6138
rect 30850 6053 31435 6061
rect 30850 6033 30859 6053
rect 30879 6052 31435 6053
rect 30879 6033 31399 6052
rect 30850 6032 31399 6033
rect 31419 6032 31435 6052
rect 30850 6026 31435 6032
rect 31224 6002 31263 6006
rect 31469 6005 31503 6211
rect 32032 6226 32067 6232
rect 32032 6207 32037 6226
rect 32058 6207 32067 6226
rect 32032 6198 32067 6207
rect 32244 6228 32300 6233
rect 32244 6208 32251 6228
rect 32271 6208 32300 6228
rect 32244 6201 32300 6208
rect 32244 6200 32279 6201
rect 32036 6130 32065 6198
rect 32036 6096 32382 6130
rect 31224 5982 31232 6002
rect 31252 5982 31263 6002
rect 28575 5972 28610 5980
rect 28575 5952 28583 5972
rect 28603 5964 28610 5972
rect 28603 5952 28614 5964
rect 28575 5715 28614 5952
rect 29445 5929 29731 5930
rect 28930 5921 29733 5929
rect 28930 5904 28941 5921
rect 28931 5899 28941 5904
rect 28965 5904 29733 5921
rect 28965 5899 28970 5904
rect 28931 5886 28970 5899
rect 29475 5838 29510 5839
rect 29454 5831 29510 5838
rect 29454 5811 29483 5831
rect 29503 5811 29510 5831
rect 29454 5806 29510 5811
rect 29694 5829 29733 5904
rect 31224 5907 31263 5982
rect 31447 6000 31503 6005
rect 31447 5980 31454 6000
rect 31474 5980 31503 6000
rect 31447 5973 31503 5980
rect 31447 5972 31482 5973
rect 31987 5912 32026 5925
rect 31987 5907 31992 5912
rect 31224 5890 31992 5907
rect 32016 5907 32026 5912
rect 32016 5890 32027 5907
rect 31224 5882 32027 5890
rect 31226 5881 31512 5882
rect 32343 5859 32382 6096
rect 32343 5847 32354 5859
rect 32347 5839 32354 5847
rect 32374 5839 32382 5859
rect 32347 5831 32382 5839
rect 29694 5809 29705 5829
rect 29725 5809 29733 5829
rect 28575 5681 28921 5715
rect 28892 5613 28921 5681
rect 28678 5610 28713 5611
rect 28657 5603 28713 5610
rect 28657 5583 28686 5603
rect 28706 5583 28713 5603
rect 28657 5578 28713 5583
rect 28890 5604 28925 5613
rect 28890 5585 28899 5604
rect 28920 5585 28925 5604
rect 28890 5579 28925 5585
rect 29454 5600 29488 5806
rect 29694 5805 29733 5809
rect 29522 5779 30107 5785
rect 29522 5759 29538 5779
rect 29558 5778 30107 5779
rect 29558 5759 30078 5778
rect 29522 5758 30078 5759
rect 30098 5758 30107 5778
rect 29522 5750 30107 5758
rect 31729 5673 32314 5681
rect 31729 5653 31738 5673
rect 31758 5672 32314 5673
rect 31758 5653 32278 5672
rect 31729 5652 32278 5653
rect 32298 5652 32314 5672
rect 31729 5646 32314 5652
rect 31453 5638 31485 5639
rect 31450 5633 31485 5638
rect 31450 5613 31457 5633
rect 31477 5613 31485 5633
rect 32348 5625 32382 5831
rect 31450 5605 31485 5613
rect 29454 5592 29489 5600
rect 28657 5372 28691 5578
rect 29454 5572 29462 5592
rect 29482 5572 29489 5592
rect 29454 5567 29489 5572
rect 29454 5566 29486 5567
rect 28725 5551 29310 5557
rect 28725 5531 28741 5551
rect 28761 5550 29310 5551
rect 28761 5531 29281 5550
rect 28725 5530 29281 5531
rect 29301 5530 29310 5550
rect 28725 5522 29310 5530
rect 29390 5521 29420 5522
rect 29390 5494 29726 5521
rect 29390 5493 29425 5494
rect 28657 5364 28692 5372
rect 28657 5344 28665 5364
rect 28685 5344 28692 5364
rect 28657 5339 28692 5344
rect 28657 5318 28691 5339
rect 29390 5318 29420 5493
rect 29476 5426 29511 5427
rect 28657 5292 29420 5318
rect 28658 5291 28691 5292
rect 29390 5290 29420 5292
rect 29455 5419 29511 5426
rect 29455 5399 29484 5419
rect 29504 5399 29511 5419
rect 29455 5394 29511 5399
rect 29690 5421 29725 5494
rect 29690 5401 29697 5421
rect 29717 5401 29725 5421
rect 30832 5447 31417 5455
rect 30832 5427 30841 5447
rect 30861 5446 31417 5447
rect 30861 5427 31381 5446
rect 30832 5426 31381 5427
rect 31401 5426 31417 5446
rect 30832 5420 31417 5426
rect 29690 5394 29725 5401
rect 31451 5399 31485 5605
rect 32114 5613 32150 5622
rect 32114 5596 32123 5613
rect 32142 5596 32150 5613
rect 32114 5587 32150 5596
rect 32326 5620 32382 5625
rect 32326 5600 32333 5620
rect 32353 5600 32382 5620
rect 32326 5593 32382 5600
rect 32326 5592 32361 5593
rect 32120 5552 32146 5587
rect 32428 5552 32460 5553
rect 32120 5547 32460 5552
rect 32120 5529 32435 5547
rect 32457 5529 32460 5547
rect 32120 5524 32460 5529
rect 32428 5523 32460 5524
rect 28309 5271 28626 5274
rect 28309 5244 28312 5271
rect 28339 5244 28626 5271
rect 28309 5238 28626 5244
rect 28309 5235 28345 5238
rect 28590 5208 28626 5238
rect 28374 5204 28409 5205
rect 28353 5197 28409 5204
rect 28353 5177 28382 5197
rect 28402 5177 28409 5197
rect 28353 5172 28409 5177
rect 28588 5202 28626 5208
rect 28588 5176 28594 5202
rect 28620 5176 28626 5202
rect 28353 4973 28387 5172
rect 28588 5168 28626 5176
rect 29455 5188 29489 5394
rect 31215 5392 31250 5399
rect 29523 5367 30108 5373
rect 29523 5347 29539 5367
rect 29559 5366 30108 5367
rect 29559 5347 30079 5366
rect 29523 5346 30079 5347
rect 30099 5346 30108 5366
rect 29523 5338 30108 5346
rect 31215 5372 31223 5392
rect 31243 5372 31250 5392
rect 31215 5299 31250 5372
rect 31429 5394 31485 5399
rect 31429 5374 31436 5394
rect 31456 5374 31485 5394
rect 31429 5367 31485 5374
rect 31520 5501 31550 5503
rect 32249 5501 32282 5502
rect 31520 5475 32283 5501
rect 31429 5366 31464 5367
rect 31520 5300 31550 5475
rect 32249 5454 32283 5475
rect 32248 5449 32283 5454
rect 32248 5429 32255 5449
rect 32275 5429 32283 5449
rect 32248 5421 32283 5429
rect 31515 5299 31550 5300
rect 31214 5272 31550 5299
rect 31520 5271 31550 5272
rect 31630 5263 32215 5271
rect 31630 5243 31639 5263
rect 31659 5262 32215 5263
rect 31659 5243 32179 5262
rect 31630 5242 32179 5243
rect 32199 5242 32215 5262
rect 31630 5236 32215 5242
rect 31454 5226 31486 5227
rect 31451 5221 31486 5226
rect 31451 5201 31458 5221
rect 31478 5201 31486 5221
rect 32249 5215 32283 5421
rect 31451 5193 31486 5201
rect 29455 5180 29490 5188
rect 29455 5160 29463 5180
rect 29483 5160 29490 5180
rect 29455 5155 29490 5160
rect 29455 5154 29487 5155
rect 28421 5145 29006 5151
rect 28421 5125 28437 5145
rect 28457 5144 29006 5145
rect 28457 5125 28977 5144
rect 28421 5124 28977 5125
rect 28997 5124 29006 5144
rect 28421 5116 29006 5124
rect 30833 5035 31418 5043
rect 30833 5015 30842 5035
rect 30862 5034 31418 5035
rect 30862 5015 31382 5034
rect 30833 5014 31382 5015
rect 31402 5014 31418 5034
rect 30833 5008 31418 5014
rect 31207 4984 31246 4988
rect 31452 4987 31486 5193
rect 32016 5205 32050 5213
rect 32016 5187 32023 5205
rect 32042 5187 32050 5205
rect 32016 5180 32050 5187
rect 32227 5210 32283 5215
rect 32227 5190 32234 5210
rect 32254 5190 32283 5210
rect 32227 5183 32283 5190
rect 32227 5182 32262 5183
rect 32020 5150 32049 5180
rect 32020 5142 32402 5150
rect 32020 5123 32373 5142
rect 32394 5123 32402 5142
rect 32020 5118 32402 5123
rect 28353 4958 28390 4973
rect 28353 4938 28361 4958
rect 28381 4938 28390 4958
rect 28353 4935 28390 4938
rect 28167 4824 28204 4827
rect 28167 4804 28176 4824
rect 28196 4804 28204 4824
rect 28167 4789 28204 4804
rect 24142 4640 24524 4645
rect 24142 4621 24150 4640
rect 24171 4621 24524 4640
rect 24142 4613 24524 4621
rect 24495 4583 24524 4613
rect 24282 4580 24317 4581
rect 24261 4573 24317 4580
rect 24261 4553 24290 4573
rect 24310 4553 24317 4573
rect 24261 4548 24317 4553
rect 24494 4576 24528 4583
rect 24494 4558 24502 4576
rect 24521 4558 24528 4576
rect 24494 4550 24528 4558
rect 25058 4570 25092 4776
rect 25298 4775 25337 4779
rect 25126 4749 25711 4755
rect 25126 4729 25142 4749
rect 25162 4748 25711 4749
rect 25162 4729 25682 4748
rect 25126 4728 25682 4729
rect 25702 4728 25711 4748
rect 25126 4720 25711 4728
rect 27551 4638 28136 4646
rect 27551 4618 27560 4638
rect 27580 4637 28136 4638
rect 27580 4618 28100 4637
rect 27551 4617 28100 4618
rect 28120 4617 28136 4637
rect 27551 4611 28136 4617
rect 27070 4607 27102 4608
rect 27067 4602 27102 4607
rect 27067 4582 27074 4602
rect 27094 4582 27102 4602
rect 28170 4590 28204 4789
rect 28148 4585 28204 4590
rect 27067 4574 27102 4582
rect 25058 4562 25093 4570
rect 24261 4342 24295 4548
rect 25058 4542 25066 4562
rect 25086 4542 25093 4562
rect 25058 4537 25093 4542
rect 25058 4536 25090 4537
rect 24329 4521 24914 4527
rect 24329 4501 24345 4521
rect 24365 4520 24914 4521
rect 24365 4501 24885 4520
rect 24329 4500 24885 4501
rect 24905 4500 24914 4520
rect 24329 4492 24914 4500
rect 24994 4491 25024 4492
rect 24994 4464 25330 4491
rect 24994 4463 25029 4464
rect 24261 4334 24296 4342
rect 24261 4314 24269 4334
rect 24289 4314 24296 4334
rect 24261 4309 24296 4314
rect 24261 4288 24295 4309
rect 24994 4288 25024 4463
rect 25080 4396 25115 4397
rect 24261 4262 25024 4288
rect 24262 4261 24295 4262
rect 24994 4260 25024 4262
rect 25059 4389 25115 4396
rect 25059 4369 25088 4389
rect 25108 4369 25115 4389
rect 25059 4364 25115 4369
rect 25294 4391 25329 4464
rect 25294 4371 25301 4391
rect 25321 4371 25329 4391
rect 26449 4416 27034 4424
rect 26449 4396 26458 4416
rect 26478 4415 27034 4416
rect 26478 4396 26998 4415
rect 26449 4395 26998 4396
rect 27018 4395 27034 4415
rect 26449 4389 27034 4395
rect 25294 4364 25329 4371
rect 27068 4368 27102 4574
rect 27930 4583 27965 4585
rect 27930 4577 27968 4583
rect 27930 4554 27938 4577
rect 27961 4554 27968 4577
rect 28148 4565 28155 4585
rect 28175 4565 28204 4585
rect 28148 4558 28204 4565
rect 28148 4557 28183 4558
rect 27930 4548 27968 4554
rect 27930 4535 27965 4548
rect 27928 4477 27965 4535
rect 24084 4239 24116 4240
rect 24084 4234 24424 4239
rect 24084 4216 24087 4234
rect 24109 4216 24424 4234
rect 24084 4211 24424 4216
rect 24084 4210 24116 4211
rect 24398 4176 24424 4211
rect 24183 4170 24218 4171
rect 24162 4163 24218 4170
rect 24162 4143 24191 4163
rect 24211 4143 24218 4163
rect 24162 4138 24218 4143
rect 24394 4167 24430 4176
rect 24394 4150 24402 4167
rect 24421 4150 24430 4167
rect 24394 4141 24430 4150
rect 25059 4158 25093 4364
rect 26832 4361 26867 4368
rect 25127 4337 25712 4343
rect 25127 4317 25143 4337
rect 25163 4336 25712 4337
rect 25163 4317 25683 4336
rect 25127 4316 25683 4317
rect 25703 4316 25712 4336
rect 25127 4308 25712 4316
rect 26832 4341 26840 4361
rect 26860 4341 26867 4361
rect 26832 4268 26867 4341
rect 27046 4363 27102 4368
rect 27046 4343 27053 4363
rect 27073 4343 27102 4363
rect 27046 4336 27102 4343
rect 27137 4470 27167 4472
rect 27866 4470 27899 4471
rect 27137 4444 27900 4470
rect 27046 4335 27081 4336
rect 27137 4269 27167 4444
rect 27866 4423 27900 4444
rect 27928 4460 27963 4477
rect 27928 4459 28222 4460
rect 27928 4458 28265 4459
rect 27928 4451 28270 4458
rect 27928 4425 28230 4451
rect 28261 4425 28270 4451
rect 27865 4418 27900 4423
rect 28221 4422 28270 4425
rect 27865 4398 27872 4418
rect 27892 4398 27900 4418
rect 28227 4417 28270 4422
rect 27865 4390 27900 4398
rect 27132 4268 27167 4269
rect 26831 4241 27167 4268
rect 27137 4240 27167 4241
rect 27247 4232 27832 4240
rect 27247 4212 27256 4232
rect 27276 4231 27832 4232
rect 27276 4212 27796 4231
rect 27247 4211 27796 4212
rect 27816 4211 27832 4231
rect 27247 4205 27832 4211
rect 27071 4195 27103 4196
rect 27068 4190 27103 4195
rect 27068 4170 27075 4190
rect 27095 4170 27103 4190
rect 27866 4184 27900 4390
rect 27068 4162 27103 4170
rect 25059 4150 25094 4158
rect 24162 3932 24196 4138
rect 25059 4130 25067 4150
rect 25087 4130 25094 4150
rect 25059 4125 25094 4130
rect 25059 4124 25091 4125
rect 24230 4111 24815 4117
rect 24230 4091 24246 4111
rect 24266 4110 24815 4111
rect 24266 4091 24786 4110
rect 24230 4090 24786 4091
rect 24806 4090 24815 4110
rect 24230 4082 24815 4090
rect 26450 4004 27035 4012
rect 26450 3984 26459 4004
rect 26479 4003 27035 4004
rect 26479 3984 26999 4003
rect 26450 3983 26999 3984
rect 27019 3983 27035 4003
rect 26450 3977 27035 3983
rect 26824 3953 26863 3957
rect 27069 3956 27103 4162
rect 27632 4177 27667 4183
rect 27632 4158 27637 4177
rect 27658 4158 27667 4177
rect 27632 4149 27667 4158
rect 27844 4179 27900 4184
rect 27844 4159 27851 4179
rect 27871 4159 27900 4179
rect 27844 4152 27900 4159
rect 27844 4151 27879 4152
rect 27636 4081 27665 4149
rect 27636 4047 27982 4081
rect 26824 3933 26832 3953
rect 26852 3933 26863 3953
rect 24162 3924 24197 3932
rect 24162 3904 24170 3924
rect 24190 3916 24197 3924
rect 24190 3904 24201 3916
rect 24162 3667 24201 3904
rect 25032 3881 25318 3882
rect 24517 3873 25320 3881
rect 24517 3856 24528 3873
rect 24518 3851 24528 3856
rect 24552 3856 25320 3873
rect 24552 3851 24557 3856
rect 24518 3838 24557 3851
rect 25062 3790 25097 3791
rect 25041 3783 25097 3790
rect 25041 3763 25070 3783
rect 25090 3763 25097 3783
rect 25041 3758 25097 3763
rect 25281 3781 25320 3856
rect 26824 3858 26863 3933
rect 27047 3951 27103 3956
rect 27047 3931 27054 3951
rect 27074 3931 27103 3951
rect 27047 3924 27103 3931
rect 27047 3923 27082 3924
rect 27587 3863 27626 3876
rect 27587 3858 27592 3863
rect 26824 3841 27592 3858
rect 27616 3858 27626 3863
rect 27616 3841 27627 3858
rect 26824 3833 27627 3841
rect 26826 3832 27112 3833
rect 27943 3810 27982 4047
rect 27943 3798 27954 3810
rect 27947 3790 27954 3798
rect 27974 3790 27982 3810
rect 27947 3782 27982 3790
rect 25281 3761 25292 3781
rect 25312 3761 25320 3781
rect 24162 3633 24508 3667
rect 24479 3565 24508 3633
rect 24265 3562 24300 3563
rect 24244 3555 24300 3562
rect 24244 3535 24273 3555
rect 24293 3535 24300 3555
rect 24244 3530 24300 3535
rect 24477 3556 24512 3565
rect 24477 3537 24486 3556
rect 24507 3537 24512 3556
rect 24477 3531 24512 3537
rect 25041 3552 25075 3758
rect 25281 3757 25320 3761
rect 25109 3731 25694 3737
rect 25109 3711 25125 3731
rect 25145 3730 25694 3731
rect 25145 3711 25665 3730
rect 25109 3710 25665 3711
rect 25685 3710 25694 3730
rect 25109 3702 25694 3710
rect 27329 3624 27914 3632
rect 27329 3604 27338 3624
rect 27358 3623 27914 3624
rect 27358 3604 27878 3623
rect 27329 3603 27878 3604
rect 27898 3603 27914 3623
rect 27329 3597 27914 3603
rect 27053 3589 27085 3590
rect 27050 3584 27085 3589
rect 27050 3564 27057 3584
rect 27077 3564 27085 3584
rect 27948 3576 27982 3782
rect 27050 3556 27085 3564
rect 25041 3544 25076 3552
rect 24244 3324 24278 3530
rect 25041 3524 25049 3544
rect 25069 3524 25076 3544
rect 25041 3519 25076 3524
rect 25041 3518 25073 3519
rect 24312 3503 24897 3509
rect 24312 3483 24328 3503
rect 24348 3502 24897 3503
rect 24348 3483 24868 3502
rect 24312 3482 24868 3483
rect 24888 3482 24897 3502
rect 24312 3474 24897 3482
rect 24977 3473 25007 3474
rect 24977 3446 25313 3473
rect 24977 3445 25012 3446
rect 24244 3316 24279 3324
rect 24244 3296 24252 3316
rect 24272 3296 24279 3316
rect 24244 3291 24279 3296
rect 24244 3270 24278 3291
rect 24977 3270 25007 3445
rect 25063 3378 25098 3379
rect 24244 3244 25007 3270
rect 24245 3243 24278 3244
rect 24977 3242 25007 3244
rect 25042 3371 25098 3378
rect 25042 3351 25071 3371
rect 25091 3351 25098 3371
rect 25042 3346 25098 3351
rect 25277 3373 25312 3446
rect 25277 3353 25284 3373
rect 25304 3353 25312 3373
rect 26432 3398 27017 3406
rect 26432 3378 26441 3398
rect 26461 3397 27017 3398
rect 26461 3378 26981 3397
rect 26432 3377 26981 3378
rect 27001 3377 27017 3397
rect 26432 3371 27017 3377
rect 25277 3346 25312 3353
rect 27051 3350 27085 3556
rect 27716 3570 27747 3576
rect 27716 3551 27721 3570
rect 27742 3551 27747 3570
rect 27716 3509 27747 3551
rect 27926 3571 27982 3576
rect 27926 3551 27933 3571
rect 27953 3551 27982 3571
rect 27926 3544 27982 3551
rect 27926 3543 27961 3544
rect 27716 3481 28055 3509
rect 23986 3187 24340 3223
rect 24002 3186 24340 3187
rect 24314 3156 24340 3186
rect 24100 3154 24135 3155
rect 24079 3147 24135 3154
rect 24079 3127 24108 3147
rect 24128 3127 24135 3147
rect 24079 3122 24135 3127
rect 24308 3148 24349 3156
rect 24308 3130 24321 3148
rect 24339 3130 24349 3148
rect 24079 2916 24113 3122
rect 24308 3119 24349 3130
rect 25042 3140 25076 3346
rect 26815 3343 26850 3350
rect 25110 3319 25695 3325
rect 25110 3299 25126 3319
rect 25146 3318 25695 3319
rect 25146 3299 25666 3318
rect 25110 3298 25666 3299
rect 25686 3298 25695 3318
rect 25110 3290 25695 3298
rect 26815 3323 26823 3343
rect 26843 3323 26850 3343
rect 26815 3250 26850 3323
rect 27029 3345 27085 3350
rect 27029 3325 27036 3345
rect 27056 3325 27085 3345
rect 27029 3318 27085 3325
rect 27120 3452 27150 3454
rect 27849 3452 27882 3453
rect 27120 3426 27883 3452
rect 27029 3317 27064 3318
rect 27120 3251 27150 3426
rect 27849 3405 27883 3426
rect 27848 3400 27883 3405
rect 27848 3380 27855 3400
rect 27875 3380 27883 3400
rect 27848 3372 27883 3380
rect 27115 3250 27150 3251
rect 26814 3223 27150 3250
rect 27120 3222 27150 3223
rect 27230 3214 27815 3222
rect 27230 3194 27239 3214
rect 27259 3213 27815 3214
rect 27259 3194 27779 3213
rect 27230 3193 27779 3194
rect 27799 3193 27815 3213
rect 27230 3187 27815 3193
rect 27054 3177 27086 3178
rect 27051 3172 27086 3177
rect 27051 3152 27058 3172
rect 27078 3152 27086 3172
rect 27849 3166 27883 3372
rect 27051 3144 27086 3152
rect 25042 3132 25077 3140
rect 25042 3112 25050 3132
rect 25070 3112 25077 3132
rect 25042 3107 25077 3112
rect 25042 3106 25074 3107
rect 24147 3095 24732 3101
rect 24147 3075 24163 3095
rect 24183 3094 24732 3095
rect 24183 3075 24703 3094
rect 24147 3074 24703 3075
rect 24723 3074 24732 3094
rect 24147 3066 24732 3074
rect 26433 2986 27018 2994
rect 26433 2966 26442 2986
rect 26462 2985 27018 2986
rect 26462 2966 26982 2985
rect 26433 2965 26982 2966
rect 27002 2965 27018 2985
rect 26433 2959 27018 2965
rect 26807 2935 26846 2939
rect 27052 2938 27086 3144
rect 27616 3156 27650 3164
rect 27616 3138 27623 3156
rect 27642 3138 27650 3156
rect 27616 3131 27650 3138
rect 27827 3161 27883 3166
rect 27827 3141 27834 3161
rect 27854 3141 27883 3161
rect 27827 3134 27883 3141
rect 27827 3133 27862 3134
rect 27620 3101 27649 3131
rect 27620 3093 28002 3101
rect 27620 3074 27973 3093
rect 27994 3074 28002 3093
rect 27620 3069 28002 3074
rect 24079 2915 24114 2916
rect 24047 2908 24114 2915
rect 24047 2888 24087 2908
rect 24107 2888 24114 2908
rect 24047 2885 24114 2888
rect 26807 2915 26815 2935
rect 26835 2915 26846 2935
rect 24047 2882 24112 2885
rect 23618 2781 23683 2784
rect 23616 2778 23683 2781
rect 23616 2758 23623 2778
rect 23643 2758 23683 2778
rect 23616 2751 23683 2758
rect 23616 2750 23651 2751
rect 20897 2730 20908 2750
rect 20928 2730 20936 2750
rect 19741 2591 20123 2596
rect 19741 2572 19749 2591
rect 19770 2572 20123 2591
rect 19741 2564 20123 2572
rect 20094 2534 20123 2564
rect 19881 2531 19916 2532
rect 19860 2524 19916 2531
rect 19860 2504 19889 2524
rect 19909 2504 19916 2524
rect 19860 2499 19916 2504
rect 20093 2527 20127 2534
rect 20093 2509 20101 2527
rect 20120 2509 20127 2527
rect 20093 2501 20127 2509
rect 20657 2521 20691 2727
rect 20897 2726 20936 2730
rect 20725 2700 21310 2706
rect 20725 2680 20741 2700
rect 20761 2699 21310 2700
rect 20761 2680 21281 2699
rect 20725 2679 21281 2680
rect 21301 2679 21310 2699
rect 20725 2671 21310 2679
rect 22998 2592 23583 2600
rect 22998 2572 23007 2592
rect 23027 2591 23583 2592
rect 23027 2572 23547 2591
rect 22998 2571 23547 2572
rect 23567 2571 23583 2591
rect 22998 2565 23583 2571
rect 22656 2559 22688 2560
rect 22653 2554 22688 2559
rect 22653 2534 22660 2554
rect 22680 2534 22688 2554
rect 22653 2526 22688 2534
rect 20657 2513 20692 2521
rect 19860 2293 19894 2499
rect 20657 2493 20665 2513
rect 20685 2493 20692 2513
rect 20657 2488 20692 2493
rect 20657 2487 20689 2488
rect 19928 2472 20513 2478
rect 19928 2452 19944 2472
rect 19964 2471 20513 2472
rect 19964 2452 20484 2471
rect 19928 2451 20484 2452
rect 20504 2451 20513 2471
rect 19928 2443 20513 2451
rect 20593 2442 20623 2443
rect 20593 2415 20929 2442
rect 20593 2414 20628 2415
rect 19860 2285 19895 2293
rect 19860 2265 19868 2285
rect 19888 2265 19895 2285
rect 19860 2260 19895 2265
rect 19860 2239 19894 2260
rect 20593 2239 20623 2414
rect 20679 2347 20714 2348
rect 19860 2213 20623 2239
rect 19861 2212 19894 2213
rect 20593 2211 20623 2213
rect 20658 2340 20714 2347
rect 20658 2320 20687 2340
rect 20707 2320 20714 2340
rect 20658 2315 20714 2320
rect 20893 2342 20928 2415
rect 20893 2322 20900 2342
rect 20920 2322 20928 2342
rect 22035 2368 22620 2376
rect 22035 2348 22044 2368
rect 22064 2367 22620 2368
rect 22064 2348 22584 2367
rect 22035 2347 22584 2348
rect 22604 2347 22620 2367
rect 22035 2341 22620 2347
rect 20893 2315 20928 2322
rect 22654 2320 22688 2526
rect 23383 2541 23416 2547
rect 23617 2544 23651 2750
rect 23383 2519 23388 2541
rect 23411 2519 23416 2541
rect 23383 2510 23416 2519
rect 23595 2539 23651 2544
rect 23595 2519 23602 2539
rect 23622 2519 23651 2539
rect 23595 2512 23651 2519
rect 23595 2511 23630 2512
rect 23385 2479 23412 2510
rect 23807 2479 23846 2491
rect 23385 2478 23848 2479
rect 23385 2456 23812 2478
rect 23836 2456 23848 2478
rect 23385 2448 23848 2456
rect 19688 2156 20027 2184
rect 19782 2121 19817 2122
rect 19761 2114 19817 2121
rect 19761 2094 19790 2114
rect 19810 2094 19817 2114
rect 19761 2089 19817 2094
rect 19996 2114 20027 2156
rect 19996 2095 20001 2114
rect 20022 2095 20027 2114
rect 19996 2089 20027 2095
rect 20658 2109 20692 2315
rect 22418 2313 22453 2320
rect 20726 2288 21311 2294
rect 20726 2268 20742 2288
rect 20762 2287 21311 2288
rect 20762 2268 21282 2287
rect 20726 2267 21282 2268
rect 21302 2267 21311 2287
rect 20726 2259 21311 2267
rect 22418 2293 22426 2313
rect 22446 2293 22453 2313
rect 22418 2220 22453 2293
rect 22632 2315 22688 2320
rect 22632 2295 22639 2315
rect 22659 2295 22688 2315
rect 22632 2288 22688 2295
rect 22723 2422 22753 2424
rect 23452 2422 23485 2423
rect 22723 2396 23486 2422
rect 22632 2287 22667 2288
rect 22723 2221 22753 2396
rect 23452 2375 23486 2396
rect 23451 2370 23486 2375
rect 23451 2350 23458 2370
rect 23478 2350 23486 2370
rect 23451 2342 23486 2350
rect 22718 2220 22753 2221
rect 22417 2193 22753 2220
rect 22723 2192 22753 2193
rect 22833 2184 23418 2192
rect 22833 2164 22842 2184
rect 22862 2183 23418 2184
rect 22862 2164 23382 2183
rect 22833 2163 23382 2164
rect 23402 2163 23418 2183
rect 22833 2157 23418 2163
rect 22657 2147 22689 2148
rect 22654 2142 22689 2147
rect 22654 2122 22661 2142
rect 22681 2122 22689 2142
rect 23452 2136 23486 2342
rect 22654 2114 22689 2122
rect 20658 2101 20693 2109
rect 19761 1883 19795 2089
rect 20658 2081 20666 2101
rect 20686 2081 20693 2101
rect 20658 2076 20693 2081
rect 20658 2075 20690 2076
rect 19829 2062 20414 2068
rect 19829 2042 19845 2062
rect 19865 2061 20414 2062
rect 19865 2042 20385 2061
rect 19829 2041 20385 2042
rect 20405 2041 20414 2061
rect 19829 2033 20414 2041
rect 22036 1956 22621 1964
rect 22036 1936 22045 1956
rect 22065 1955 22621 1956
rect 22065 1936 22585 1955
rect 22036 1935 22585 1936
rect 22605 1935 22621 1955
rect 22036 1929 22621 1935
rect 22410 1905 22449 1909
rect 22655 1908 22689 2114
rect 23218 2129 23253 2135
rect 23218 2110 23223 2129
rect 23244 2110 23253 2129
rect 23218 2101 23253 2110
rect 23430 2131 23486 2136
rect 23430 2111 23437 2131
rect 23457 2111 23486 2131
rect 23430 2104 23486 2111
rect 23608 2282 23640 2294
rect 23608 2264 23615 2282
rect 23637 2264 23640 2282
rect 23430 2103 23465 2104
rect 23222 2033 23251 2101
rect 23222 1999 23568 2033
rect 22410 1885 22418 1905
rect 22438 1885 22449 1905
rect 19761 1875 19796 1883
rect 19761 1855 19769 1875
rect 19789 1867 19796 1875
rect 19789 1855 19800 1867
rect 19761 1618 19800 1855
rect 20631 1832 20917 1833
rect 20116 1824 20919 1832
rect 20116 1807 20127 1824
rect 20117 1802 20127 1807
rect 20151 1807 20919 1824
rect 20151 1802 20156 1807
rect 20117 1789 20156 1802
rect 20661 1741 20696 1742
rect 20640 1734 20696 1741
rect 20640 1714 20669 1734
rect 20689 1714 20696 1734
rect 20640 1709 20696 1714
rect 20880 1732 20919 1807
rect 22410 1810 22449 1885
rect 22633 1903 22689 1908
rect 22633 1883 22640 1903
rect 22660 1883 22689 1903
rect 22633 1876 22689 1883
rect 22633 1875 22668 1876
rect 23173 1815 23212 1828
rect 23173 1810 23178 1815
rect 22410 1793 23178 1810
rect 23202 1810 23212 1815
rect 23202 1793 23213 1810
rect 22410 1785 23213 1793
rect 22412 1784 22698 1785
rect 23529 1762 23568 1999
rect 23529 1750 23540 1762
rect 23533 1742 23540 1750
rect 23560 1742 23568 1762
rect 23533 1734 23568 1742
rect 20880 1712 20891 1732
rect 20911 1712 20919 1732
rect 19761 1584 20107 1618
rect 20078 1516 20107 1584
rect 19864 1513 19899 1514
rect 18942 1414 19276 1442
rect 19843 1506 19899 1513
rect 19843 1486 19872 1506
rect 19892 1486 19899 1506
rect 19843 1481 19899 1486
rect 20076 1507 20111 1516
rect 20076 1488 20085 1507
rect 20106 1488 20111 1507
rect 20076 1482 20111 1488
rect 20640 1503 20674 1709
rect 20880 1708 20919 1712
rect 20708 1682 21293 1688
rect 20708 1662 20724 1682
rect 20744 1681 21293 1682
rect 20744 1662 21264 1681
rect 20708 1661 21264 1662
rect 21284 1661 21293 1681
rect 20708 1653 21293 1661
rect 22915 1576 23500 1584
rect 22915 1556 22924 1576
rect 22944 1575 23500 1576
rect 22944 1556 23464 1575
rect 22915 1555 23464 1556
rect 23484 1555 23500 1575
rect 22915 1549 23500 1555
rect 22639 1541 22671 1542
rect 22636 1536 22671 1541
rect 22636 1516 22643 1536
rect 22663 1516 22671 1536
rect 23534 1528 23568 1734
rect 22636 1508 22671 1516
rect 20640 1495 20675 1503
rect 16443 1267 17028 1275
rect 18037 1282 18072 1289
rect 18037 1262 18045 1282
rect 18065 1262 18072 1282
rect 18037 1189 18072 1262
rect 18251 1284 18307 1289
rect 18251 1264 18258 1284
rect 18278 1264 18307 1284
rect 18251 1257 18307 1264
rect 18342 1391 18372 1393
rect 19071 1391 19104 1392
rect 18342 1365 19105 1391
rect 18251 1256 18286 1257
rect 18342 1190 18372 1365
rect 19071 1344 19105 1365
rect 19070 1339 19105 1344
rect 19070 1319 19077 1339
rect 19097 1319 19105 1339
rect 19070 1311 19105 1319
rect 18337 1189 18372 1190
rect 18036 1162 18372 1189
rect 18342 1161 18372 1162
rect 18452 1153 19037 1161
rect 18452 1133 18461 1153
rect 18481 1152 19037 1153
rect 18481 1133 19001 1152
rect 18452 1132 19001 1133
rect 19021 1132 19037 1152
rect 18452 1126 19037 1132
rect 16375 1109 16410 1117
rect 18276 1116 18308 1117
rect 14783 1098 14818 1099
rect 14576 1066 14605 1096
rect 16375 1089 16383 1109
rect 16403 1089 16410 1109
rect 16375 1084 16410 1089
rect 18273 1111 18308 1116
rect 18273 1091 18280 1111
rect 18300 1091 18308 1111
rect 19071 1105 19105 1311
rect 19843 1275 19877 1481
rect 20640 1475 20648 1495
rect 20668 1475 20675 1495
rect 20640 1470 20675 1475
rect 20640 1469 20672 1470
rect 19911 1454 20496 1460
rect 19911 1434 19927 1454
rect 19947 1453 20496 1454
rect 19947 1434 20467 1453
rect 19911 1433 20467 1434
rect 20487 1433 20496 1453
rect 19911 1425 20496 1433
rect 20576 1424 20606 1425
rect 20576 1397 20912 1424
rect 20576 1396 20611 1397
rect 19843 1267 19878 1275
rect 19843 1247 19851 1267
rect 19871 1247 19878 1267
rect 19843 1242 19878 1247
rect 19843 1221 19877 1242
rect 20576 1221 20606 1396
rect 20662 1329 20697 1330
rect 19843 1195 20606 1221
rect 19844 1194 19877 1195
rect 20576 1193 20606 1195
rect 20641 1322 20697 1329
rect 20641 1302 20670 1322
rect 20690 1302 20697 1322
rect 20641 1297 20697 1302
rect 20876 1324 20911 1397
rect 20876 1304 20883 1324
rect 20903 1304 20911 1324
rect 22018 1350 22603 1358
rect 22018 1330 22027 1350
rect 22047 1349 22603 1350
rect 22047 1330 22567 1349
rect 22018 1329 22567 1330
rect 22587 1329 22603 1349
rect 22018 1323 22603 1329
rect 20876 1297 20911 1304
rect 22637 1302 22671 1508
rect 23300 1516 23336 1525
rect 23300 1499 23309 1516
rect 23328 1499 23336 1516
rect 23300 1490 23336 1499
rect 23512 1523 23568 1528
rect 23512 1503 23519 1523
rect 23539 1503 23568 1523
rect 23512 1496 23568 1503
rect 23512 1495 23547 1496
rect 23306 1455 23332 1490
rect 23608 1455 23640 2264
rect 24052 2197 24081 2882
rect 25012 2863 25298 2864
rect 24497 2855 25300 2863
rect 24497 2838 24508 2855
rect 24498 2833 24508 2838
rect 24532 2838 25300 2855
rect 24532 2833 24537 2838
rect 24498 2820 24537 2833
rect 25042 2772 25077 2773
rect 25021 2765 25077 2772
rect 25021 2745 25050 2765
rect 25070 2745 25077 2765
rect 25021 2740 25077 2745
rect 25261 2763 25300 2838
rect 26807 2840 26846 2915
rect 27030 2933 27086 2938
rect 27030 2913 27037 2933
rect 27057 2913 27086 2933
rect 27030 2906 27086 2913
rect 27030 2905 27065 2906
rect 27570 2845 27609 2858
rect 27570 2840 27575 2845
rect 26807 2823 27575 2840
rect 27599 2840 27609 2845
rect 27599 2823 27610 2840
rect 26807 2815 27610 2823
rect 26809 2814 27095 2815
rect 28026 2796 28055 3481
rect 28363 3235 28390 4935
rect 31207 4964 31215 4984
rect 31235 4964 31246 4984
rect 29426 4911 29712 4912
rect 28911 4903 29714 4911
rect 28911 4886 28922 4903
rect 28912 4881 28922 4886
rect 28946 4886 29714 4903
rect 28946 4881 28951 4886
rect 28912 4868 28951 4881
rect 29456 4820 29491 4821
rect 29435 4813 29491 4820
rect 29435 4793 29464 4813
rect 29484 4793 29491 4813
rect 29435 4788 29491 4793
rect 29675 4811 29714 4886
rect 31207 4889 31246 4964
rect 31430 4982 31486 4987
rect 31430 4962 31437 4982
rect 31457 4962 31486 4982
rect 31430 4955 31486 4962
rect 31430 4954 31465 4955
rect 31970 4894 32009 4907
rect 31970 4889 31975 4894
rect 31207 4872 31975 4889
rect 31999 4889 32009 4894
rect 31999 4872 32010 4889
rect 31207 4864 32010 4872
rect 31209 4863 31495 4864
rect 29675 4791 29686 4811
rect 29706 4791 29714 4811
rect 32531 4840 32558 6540
rect 32866 6294 32895 6979
rect 33826 6960 34112 6961
rect 33311 6952 34114 6960
rect 33311 6935 33322 6952
rect 33312 6930 33322 6935
rect 33346 6935 34114 6952
rect 33346 6930 33351 6935
rect 33312 6917 33351 6930
rect 33856 6869 33891 6870
rect 33835 6862 33891 6869
rect 33835 6842 33864 6862
rect 33884 6842 33891 6862
rect 33835 6837 33891 6842
rect 34075 6860 34114 6935
rect 34075 6840 34086 6860
rect 34106 6840 34114 6860
rect 32919 6701 33301 6706
rect 32919 6682 32927 6701
rect 32948 6682 33301 6701
rect 32919 6674 33301 6682
rect 33272 6644 33301 6674
rect 33059 6641 33094 6642
rect 33038 6634 33094 6641
rect 33038 6614 33067 6634
rect 33087 6614 33094 6634
rect 33038 6609 33094 6614
rect 33271 6637 33305 6644
rect 33271 6619 33279 6637
rect 33298 6619 33305 6637
rect 33271 6611 33305 6619
rect 33835 6631 33869 6837
rect 34075 6836 34114 6840
rect 33903 6810 34488 6816
rect 33903 6790 33919 6810
rect 33939 6809 34488 6810
rect 33939 6790 34459 6809
rect 33903 6789 34459 6790
rect 34479 6789 34488 6809
rect 33903 6781 34488 6789
rect 33835 6623 33870 6631
rect 33038 6403 33072 6609
rect 33835 6603 33843 6623
rect 33863 6603 33870 6623
rect 33835 6598 33870 6603
rect 33835 6597 33867 6598
rect 33106 6582 33691 6588
rect 33106 6562 33122 6582
rect 33142 6581 33691 6582
rect 33142 6562 33662 6581
rect 33106 6561 33662 6562
rect 33682 6561 33691 6581
rect 33106 6553 33691 6561
rect 33771 6552 33801 6553
rect 33771 6525 34107 6552
rect 33771 6524 33806 6525
rect 33038 6395 33073 6403
rect 33038 6375 33046 6395
rect 33066 6375 33073 6395
rect 33038 6370 33073 6375
rect 33038 6349 33072 6370
rect 33771 6349 33801 6524
rect 33857 6457 33892 6458
rect 33038 6323 33801 6349
rect 33039 6322 33072 6323
rect 33771 6321 33801 6323
rect 33836 6450 33892 6457
rect 33836 6430 33865 6450
rect 33885 6430 33892 6450
rect 33836 6425 33892 6430
rect 34071 6452 34106 6525
rect 34071 6432 34078 6452
rect 34098 6432 34106 6452
rect 34071 6425 34106 6432
rect 32866 6266 33205 6294
rect 32960 6231 32995 6232
rect 32939 6224 32995 6231
rect 32939 6204 32968 6224
rect 32988 6204 32995 6224
rect 32939 6199 32995 6204
rect 33174 6224 33205 6266
rect 33174 6205 33179 6224
rect 33200 6205 33205 6224
rect 33174 6199 33205 6205
rect 33836 6219 33870 6425
rect 33904 6398 34489 6404
rect 33904 6378 33920 6398
rect 33940 6397 34489 6398
rect 33940 6378 34460 6397
rect 33904 6377 34460 6378
rect 34480 6377 34489 6397
rect 33904 6369 34489 6377
rect 33836 6211 33871 6219
rect 32939 5993 32973 6199
rect 33836 6191 33844 6211
rect 33864 6191 33871 6211
rect 33836 6186 33871 6191
rect 33836 6185 33868 6186
rect 33007 6172 33592 6178
rect 33007 6152 33023 6172
rect 33043 6171 33592 6172
rect 33043 6152 33563 6171
rect 33007 6151 33563 6152
rect 33583 6151 33592 6171
rect 33007 6143 33592 6151
rect 32939 5985 32974 5993
rect 32939 5965 32947 5985
rect 32967 5977 32974 5985
rect 32967 5965 32978 5977
rect 32939 5728 32978 5965
rect 33809 5942 34095 5943
rect 33294 5934 34097 5942
rect 33294 5917 33305 5934
rect 33295 5912 33305 5917
rect 33329 5917 34097 5934
rect 33329 5912 33334 5917
rect 33295 5899 33334 5912
rect 33839 5851 33874 5852
rect 33818 5844 33874 5851
rect 33818 5824 33847 5844
rect 33867 5824 33874 5844
rect 33818 5819 33874 5824
rect 34058 5842 34097 5917
rect 34058 5822 34069 5842
rect 34089 5822 34097 5842
rect 32939 5694 33285 5728
rect 33256 5626 33285 5694
rect 33042 5623 33077 5624
rect 33021 5616 33077 5623
rect 33021 5596 33050 5616
rect 33070 5596 33077 5616
rect 33021 5591 33077 5596
rect 33254 5617 33289 5626
rect 33254 5598 33263 5617
rect 33284 5598 33289 5617
rect 33254 5592 33289 5598
rect 33818 5613 33852 5819
rect 34058 5818 34097 5822
rect 33886 5792 34471 5798
rect 33886 5772 33902 5792
rect 33922 5791 34471 5792
rect 33922 5772 34442 5791
rect 33886 5771 34442 5772
rect 34462 5771 34471 5791
rect 33886 5763 34471 5771
rect 33818 5605 33853 5613
rect 33021 5385 33055 5591
rect 33818 5585 33826 5605
rect 33846 5585 33853 5605
rect 33818 5580 33853 5585
rect 33818 5579 33850 5580
rect 33089 5564 33674 5570
rect 33089 5544 33105 5564
rect 33125 5563 33674 5564
rect 33125 5544 33645 5563
rect 33089 5543 33645 5544
rect 33665 5543 33674 5563
rect 33089 5535 33674 5543
rect 33754 5534 33784 5535
rect 33754 5507 34090 5534
rect 33754 5506 33789 5507
rect 33021 5377 33056 5385
rect 33021 5357 33029 5377
rect 33049 5357 33056 5377
rect 33021 5352 33056 5357
rect 33021 5331 33055 5352
rect 33754 5331 33784 5506
rect 33840 5439 33875 5440
rect 33021 5305 33784 5331
rect 33022 5304 33055 5305
rect 33754 5303 33784 5305
rect 33819 5432 33875 5439
rect 33819 5412 33848 5432
rect 33868 5412 33875 5432
rect 33819 5407 33875 5412
rect 34054 5434 34089 5507
rect 34054 5414 34061 5434
rect 34081 5414 34089 5434
rect 34054 5407 34089 5414
rect 32673 5284 32990 5287
rect 32673 5257 32676 5284
rect 32703 5257 32990 5284
rect 32673 5251 32990 5257
rect 32673 5248 32709 5251
rect 32954 5221 32990 5251
rect 32738 5217 32773 5218
rect 32717 5210 32773 5217
rect 32717 5190 32746 5210
rect 32766 5190 32773 5210
rect 32717 5185 32773 5190
rect 32952 5215 32990 5221
rect 32952 5189 32958 5215
rect 32984 5189 32990 5215
rect 32717 4986 32751 5185
rect 32952 5181 32990 5189
rect 33819 5201 33853 5407
rect 33887 5380 34472 5386
rect 33887 5360 33903 5380
rect 33923 5379 34472 5380
rect 33923 5360 34443 5379
rect 33887 5359 34443 5360
rect 34463 5359 34472 5379
rect 33887 5351 34472 5359
rect 33819 5193 33854 5201
rect 33819 5173 33827 5193
rect 33847 5173 33854 5193
rect 33819 5168 33854 5173
rect 33819 5167 33851 5168
rect 32785 5158 33370 5164
rect 32785 5138 32801 5158
rect 32821 5157 33370 5158
rect 32821 5138 33341 5157
rect 32785 5137 33341 5138
rect 33361 5137 33370 5157
rect 32785 5129 33370 5137
rect 32717 4971 32754 4986
rect 32717 4951 32725 4971
rect 32745 4951 32754 4971
rect 32717 4948 32754 4951
rect 32531 4837 32568 4840
rect 32531 4817 32540 4837
rect 32560 4817 32568 4837
rect 32531 4802 32568 4817
rect 28519 4652 28901 4657
rect 28519 4633 28527 4652
rect 28548 4633 28901 4652
rect 28519 4625 28901 4633
rect 28872 4595 28901 4625
rect 28659 4592 28694 4593
rect 28638 4585 28694 4592
rect 28638 4565 28667 4585
rect 28687 4565 28694 4585
rect 28638 4560 28694 4565
rect 28871 4588 28905 4595
rect 28871 4570 28879 4588
rect 28898 4570 28905 4588
rect 28871 4562 28905 4570
rect 29435 4582 29469 4788
rect 29675 4787 29714 4791
rect 29503 4761 30088 4767
rect 29503 4741 29519 4761
rect 29539 4760 30088 4761
rect 29539 4741 30059 4760
rect 29503 4740 30059 4741
rect 30079 4740 30088 4760
rect 29503 4732 30088 4740
rect 31915 4651 32500 4659
rect 31915 4631 31924 4651
rect 31944 4650 32500 4651
rect 31944 4631 32464 4650
rect 31915 4630 32464 4631
rect 32484 4630 32500 4650
rect 31915 4624 32500 4630
rect 31434 4620 31466 4621
rect 31431 4615 31466 4620
rect 31431 4595 31438 4615
rect 31458 4595 31466 4615
rect 32534 4603 32568 4802
rect 32512 4598 32568 4603
rect 31431 4587 31466 4595
rect 29435 4574 29470 4582
rect 28638 4354 28672 4560
rect 29435 4554 29443 4574
rect 29463 4554 29470 4574
rect 29435 4549 29470 4554
rect 29435 4548 29467 4549
rect 28706 4533 29291 4539
rect 28706 4513 28722 4533
rect 28742 4532 29291 4533
rect 28742 4513 29262 4532
rect 28706 4512 29262 4513
rect 29282 4512 29291 4532
rect 28706 4504 29291 4512
rect 29371 4503 29401 4504
rect 29371 4476 29707 4503
rect 29371 4475 29406 4476
rect 28638 4346 28673 4354
rect 28638 4326 28646 4346
rect 28666 4326 28673 4346
rect 28638 4321 28673 4326
rect 28638 4300 28672 4321
rect 29371 4300 29401 4475
rect 29457 4408 29492 4409
rect 28638 4274 29401 4300
rect 28639 4273 28672 4274
rect 29371 4272 29401 4274
rect 29436 4401 29492 4408
rect 29436 4381 29465 4401
rect 29485 4381 29492 4401
rect 29436 4376 29492 4381
rect 29671 4403 29706 4476
rect 29671 4383 29678 4403
rect 29698 4383 29706 4403
rect 30813 4429 31398 4437
rect 30813 4409 30822 4429
rect 30842 4428 31398 4429
rect 30842 4409 31362 4428
rect 30813 4408 31362 4409
rect 31382 4408 31398 4428
rect 30813 4402 31398 4408
rect 29671 4376 29706 4383
rect 31432 4381 31466 4587
rect 32294 4596 32329 4598
rect 32294 4590 32332 4596
rect 32294 4567 32302 4590
rect 32325 4567 32332 4590
rect 32512 4578 32519 4598
rect 32539 4578 32568 4598
rect 32512 4571 32568 4578
rect 32512 4570 32547 4571
rect 32294 4561 32332 4567
rect 32294 4548 32329 4561
rect 32292 4490 32329 4548
rect 28461 4251 28493 4252
rect 28461 4246 28801 4251
rect 28461 4228 28464 4246
rect 28486 4228 28801 4246
rect 28461 4223 28801 4228
rect 28461 4222 28493 4223
rect 28775 4188 28801 4223
rect 28560 4182 28595 4183
rect 28539 4175 28595 4182
rect 28539 4155 28568 4175
rect 28588 4155 28595 4175
rect 28539 4150 28595 4155
rect 28771 4179 28807 4188
rect 28771 4162 28779 4179
rect 28798 4162 28807 4179
rect 28771 4153 28807 4162
rect 29436 4170 29470 4376
rect 31196 4374 31231 4381
rect 29504 4349 30089 4355
rect 29504 4329 29520 4349
rect 29540 4348 30089 4349
rect 29540 4329 30060 4348
rect 29504 4328 30060 4329
rect 30080 4328 30089 4348
rect 29504 4320 30089 4328
rect 31196 4354 31204 4374
rect 31224 4354 31231 4374
rect 31196 4281 31231 4354
rect 31410 4376 31466 4381
rect 31410 4356 31417 4376
rect 31437 4356 31466 4376
rect 31410 4349 31466 4356
rect 31501 4483 31531 4485
rect 32230 4483 32263 4484
rect 31501 4457 32264 4483
rect 31410 4348 31445 4349
rect 31501 4282 31531 4457
rect 32230 4436 32264 4457
rect 32292 4473 32327 4490
rect 32292 4472 32586 4473
rect 32292 4471 32629 4472
rect 32292 4464 32634 4471
rect 32292 4438 32594 4464
rect 32625 4438 32634 4464
rect 32229 4431 32264 4436
rect 32585 4435 32634 4438
rect 32229 4411 32236 4431
rect 32256 4411 32264 4431
rect 32591 4430 32634 4435
rect 32229 4403 32264 4411
rect 31496 4281 31531 4282
rect 31195 4254 31531 4281
rect 31501 4253 31531 4254
rect 31611 4245 32196 4253
rect 31611 4225 31620 4245
rect 31640 4244 32196 4245
rect 31640 4225 32160 4244
rect 31611 4224 32160 4225
rect 32180 4224 32196 4244
rect 31611 4218 32196 4224
rect 31435 4208 31467 4209
rect 31432 4203 31467 4208
rect 31432 4183 31439 4203
rect 31459 4183 31467 4203
rect 32230 4197 32264 4403
rect 31432 4175 31467 4183
rect 29436 4162 29471 4170
rect 28539 3944 28573 4150
rect 29436 4142 29444 4162
rect 29464 4142 29471 4162
rect 29436 4137 29471 4142
rect 29436 4136 29468 4137
rect 28607 4123 29192 4129
rect 28607 4103 28623 4123
rect 28643 4122 29192 4123
rect 28643 4103 29163 4122
rect 28607 4102 29163 4103
rect 29183 4102 29192 4122
rect 28607 4094 29192 4102
rect 30814 4017 31399 4025
rect 30814 3997 30823 4017
rect 30843 4016 31399 4017
rect 30843 3997 31363 4016
rect 30814 3996 31363 3997
rect 31383 3996 31399 4016
rect 30814 3990 31399 3996
rect 31188 3966 31227 3970
rect 31433 3969 31467 4175
rect 31996 4190 32031 4196
rect 31996 4171 32001 4190
rect 32022 4171 32031 4190
rect 31996 4162 32031 4171
rect 32208 4192 32264 4197
rect 32208 4172 32215 4192
rect 32235 4172 32264 4192
rect 32208 4165 32264 4172
rect 32208 4164 32243 4165
rect 32000 4094 32029 4162
rect 32000 4060 32346 4094
rect 31188 3946 31196 3966
rect 31216 3946 31227 3966
rect 28539 3936 28574 3944
rect 28539 3916 28547 3936
rect 28567 3928 28574 3936
rect 28567 3916 28578 3928
rect 28539 3679 28578 3916
rect 29409 3893 29695 3894
rect 28894 3885 29697 3893
rect 28894 3868 28905 3885
rect 28895 3863 28905 3868
rect 28929 3868 29697 3885
rect 28929 3863 28934 3868
rect 28895 3850 28934 3863
rect 29439 3802 29474 3803
rect 29418 3795 29474 3802
rect 29418 3775 29447 3795
rect 29467 3775 29474 3795
rect 29418 3770 29474 3775
rect 29658 3793 29697 3868
rect 31188 3871 31227 3946
rect 31411 3964 31467 3969
rect 31411 3944 31418 3964
rect 31438 3944 31467 3964
rect 31411 3937 31467 3944
rect 31411 3936 31446 3937
rect 31951 3876 31990 3889
rect 31951 3871 31956 3876
rect 31188 3854 31956 3871
rect 31980 3871 31990 3876
rect 31980 3854 31991 3871
rect 31188 3846 31991 3854
rect 31190 3845 31476 3846
rect 32307 3823 32346 4060
rect 32307 3811 32318 3823
rect 32311 3803 32318 3811
rect 32338 3803 32346 3823
rect 32311 3795 32346 3803
rect 29658 3773 29669 3793
rect 29689 3773 29697 3793
rect 28539 3645 28885 3679
rect 28856 3577 28885 3645
rect 28642 3574 28677 3575
rect 28621 3567 28677 3574
rect 28621 3547 28650 3567
rect 28670 3547 28677 3567
rect 28621 3542 28677 3547
rect 28854 3568 28889 3577
rect 28854 3549 28863 3568
rect 28884 3549 28889 3568
rect 28854 3543 28889 3549
rect 29418 3564 29452 3770
rect 29658 3769 29697 3773
rect 29486 3743 30071 3749
rect 29486 3723 29502 3743
rect 29522 3742 30071 3743
rect 29522 3723 30042 3742
rect 29486 3722 30042 3723
rect 30062 3722 30071 3742
rect 29486 3714 30071 3722
rect 31693 3637 32278 3645
rect 31693 3617 31702 3637
rect 31722 3636 32278 3637
rect 31722 3617 32242 3636
rect 31693 3616 32242 3617
rect 32262 3616 32278 3636
rect 31693 3610 32278 3616
rect 31417 3602 31449 3603
rect 31414 3597 31449 3602
rect 31414 3577 31421 3597
rect 31441 3577 31449 3597
rect 32312 3589 32346 3795
rect 31414 3569 31449 3577
rect 29418 3556 29453 3564
rect 28621 3336 28655 3542
rect 29418 3536 29426 3556
rect 29446 3536 29453 3556
rect 29418 3531 29453 3536
rect 29418 3530 29450 3531
rect 28689 3515 29274 3521
rect 28689 3495 28705 3515
rect 28725 3514 29274 3515
rect 28725 3495 29245 3514
rect 28689 3494 29245 3495
rect 29265 3494 29274 3514
rect 28689 3486 29274 3494
rect 29354 3485 29384 3486
rect 29354 3458 29690 3485
rect 29354 3457 29389 3458
rect 28621 3328 28656 3336
rect 28621 3308 28629 3328
rect 28649 3308 28656 3328
rect 28621 3303 28656 3308
rect 28621 3282 28655 3303
rect 29354 3282 29384 3457
rect 29440 3390 29475 3391
rect 28621 3256 29384 3282
rect 28622 3255 28655 3256
rect 29354 3254 29384 3256
rect 29419 3383 29475 3390
rect 29419 3363 29448 3383
rect 29468 3363 29475 3383
rect 29419 3358 29475 3363
rect 29654 3385 29689 3458
rect 29654 3365 29661 3385
rect 29681 3365 29689 3385
rect 30796 3411 31381 3419
rect 30796 3391 30805 3411
rect 30825 3410 31381 3411
rect 30825 3391 31345 3410
rect 30796 3390 31345 3391
rect 31365 3390 31381 3410
rect 30796 3384 31381 3390
rect 29654 3358 29689 3365
rect 31415 3363 31449 3569
rect 32080 3583 32111 3589
rect 32080 3564 32085 3583
rect 32106 3564 32111 3583
rect 32080 3522 32111 3564
rect 32290 3584 32346 3589
rect 32290 3564 32297 3584
rect 32317 3564 32346 3584
rect 32290 3557 32346 3564
rect 32290 3556 32325 3557
rect 32080 3494 32419 3522
rect 28363 3199 28717 3235
rect 28379 3198 28717 3199
rect 28691 3168 28717 3198
rect 28477 3166 28512 3167
rect 28456 3159 28512 3166
rect 28456 3139 28485 3159
rect 28505 3139 28512 3159
rect 28456 3134 28512 3139
rect 28685 3160 28726 3168
rect 28685 3142 28698 3160
rect 28716 3142 28726 3160
rect 28456 2928 28490 3134
rect 28685 3131 28726 3142
rect 29419 3152 29453 3358
rect 31179 3356 31214 3363
rect 29487 3331 30072 3337
rect 29487 3311 29503 3331
rect 29523 3330 30072 3331
rect 29523 3311 30043 3330
rect 29487 3310 30043 3311
rect 30063 3310 30072 3330
rect 29487 3302 30072 3310
rect 31179 3336 31187 3356
rect 31207 3336 31214 3356
rect 31179 3263 31214 3336
rect 31393 3358 31449 3363
rect 31393 3338 31400 3358
rect 31420 3338 31449 3358
rect 31393 3331 31449 3338
rect 31484 3465 31514 3467
rect 32213 3465 32246 3466
rect 31484 3439 32247 3465
rect 31393 3330 31428 3331
rect 31484 3264 31514 3439
rect 32213 3418 32247 3439
rect 32212 3413 32247 3418
rect 32212 3393 32219 3413
rect 32239 3393 32247 3413
rect 32212 3385 32247 3393
rect 31479 3263 31514 3264
rect 31178 3236 31514 3263
rect 31484 3235 31514 3236
rect 31594 3227 32179 3235
rect 31594 3207 31603 3227
rect 31623 3226 32179 3227
rect 31623 3207 32143 3226
rect 31594 3206 32143 3207
rect 32163 3206 32179 3226
rect 31594 3200 32179 3206
rect 31418 3190 31450 3191
rect 31415 3185 31450 3190
rect 31415 3165 31422 3185
rect 31442 3165 31450 3185
rect 32213 3179 32247 3385
rect 31415 3157 31450 3165
rect 29419 3144 29454 3152
rect 29419 3124 29427 3144
rect 29447 3124 29454 3144
rect 29419 3119 29454 3124
rect 29419 3118 29451 3119
rect 28524 3107 29109 3113
rect 28524 3087 28540 3107
rect 28560 3106 29109 3107
rect 28560 3087 29080 3106
rect 28524 3086 29080 3087
rect 29100 3086 29109 3106
rect 28524 3078 29109 3086
rect 30797 2999 31382 3007
rect 30797 2979 30806 2999
rect 30826 2998 31382 2999
rect 30826 2979 31346 2998
rect 30797 2978 31346 2979
rect 31366 2978 31382 2998
rect 30797 2972 31382 2978
rect 31171 2948 31210 2952
rect 31416 2951 31450 3157
rect 31980 3169 32014 3177
rect 31980 3151 31987 3169
rect 32006 3151 32014 3169
rect 31980 3144 32014 3151
rect 32191 3174 32247 3179
rect 32191 3154 32198 3174
rect 32218 3154 32247 3174
rect 32191 3147 32247 3154
rect 32191 3146 32226 3147
rect 31984 3114 32013 3144
rect 31984 3106 32366 3114
rect 31984 3087 32337 3106
rect 32358 3087 32366 3106
rect 31984 3082 32366 3087
rect 31171 2928 31179 2948
rect 31199 2928 31210 2948
rect 28456 2927 28491 2928
rect 28424 2920 28491 2927
rect 28424 2900 28464 2920
rect 28484 2900 28491 2920
rect 28424 2897 28491 2900
rect 28424 2894 28489 2897
rect 27995 2793 28060 2796
rect 25261 2743 25272 2763
rect 25292 2743 25300 2763
rect 27993 2790 28060 2793
rect 27993 2770 28000 2790
rect 28020 2770 28060 2790
rect 27993 2763 28060 2770
rect 27993 2762 28028 2763
rect 24105 2604 24487 2609
rect 24105 2585 24113 2604
rect 24134 2585 24487 2604
rect 24105 2577 24487 2585
rect 24458 2547 24487 2577
rect 24245 2544 24280 2545
rect 24224 2537 24280 2544
rect 24224 2517 24253 2537
rect 24273 2517 24280 2537
rect 24224 2512 24280 2517
rect 24457 2540 24491 2547
rect 24457 2522 24465 2540
rect 24484 2522 24491 2540
rect 24457 2514 24491 2522
rect 25021 2534 25055 2740
rect 25261 2739 25300 2743
rect 25089 2713 25674 2719
rect 25089 2693 25105 2713
rect 25125 2712 25674 2713
rect 25125 2693 25645 2712
rect 25089 2692 25645 2693
rect 25665 2692 25674 2712
rect 25089 2684 25674 2692
rect 27375 2604 27960 2612
rect 27375 2584 27384 2604
rect 27404 2603 27960 2604
rect 27404 2584 27924 2603
rect 27375 2583 27924 2584
rect 27944 2583 27960 2603
rect 27375 2577 27960 2583
rect 27033 2571 27065 2572
rect 27030 2566 27065 2571
rect 27030 2546 27037 2566
rect 27057 2546 27065 2566
rect 27030 2538 27065 2546
rect 25021 2526 25056 2534
rect 24224 2306 24258 2512
rect 25021 2506 25029 2526
rect 25049 2506 25056 2526
rect 25021 2501 25056 2506
rect 25021 2500 25053 2501
rect 24292 2485 24877 2491
rect 24292 2465 24308 2485
rect 24328 2484 24877 2485
rect 24328 2465 24848 2484
rect 24292 2464 24848 2465
rect 24868 2464 24877 2484
rect 24292 2456 24877 2464
rect 24957 2455 24987 2456
rect 24957 2428 25293 2455
rect 24957 2427 24992 2428
rect 24224 2298 24259 2306
rect 24224 2278 24232 2298
rect 24252 2278 24259 2298
rect 24224 2273 24259 2278
rect 24224 2252 24258 2273
rect 24957 2252 24987 2427
rect 25043 2360 25078 2361
rect 24224 2226 24987 2252
rect 24225 2225 24258 2226
rect 24957 2224 24987 2226
rect 25022 2353 25078 2360
rect 25022 2333 25051 2353
rect 25071 2333 25078 2353
rect 25022 2328 25078 2333
rect 25257 2355 25292 2428
rect 25257 2335 25264 2355
rect 25284 2335 25292 2355
rect 26412 2380 26997 2388
rect 26412 2360 26421 2380
rect 26441 2379 26997 2380
rect 26441 2360 26961 2379
rect 26412 2359 26961 2360
rect 26981 2359 26997 2379
rect 26412 2353 26997 2359
rect 25257 2328 25292 2335
rect 27031 2332 27065 2538
rect 27760 2553 27793 2559
rect 27994 2556 28028 2762
rect 27760 2531 27765 2553
rect 27788 2531 27793 2553
rect 27760 2522 27793 2531
rect 27972 2551 28028 2556
rect 27972 2531 27979 2551
rect 27999 2531 28028 2551
rect 27972 2524 28028 2531
rect 27972 2523 28007 2524
rect 27762 2491 27789 2522
rect 28184 2491 28223 2503
rect 27762 2490 28225 2491
rect 27762 2468 28189 2490
rect 28213 2468 28225 2490
rect 27762 2460 28225 2468
rect 24052 2169 24391 2197
rect 24146 2134 24181 2135
rect 24125 2127 24181 2134
rect 24125 2107 24154 2127
rect 24174 2107 24181 2127
rect 24125 2102 24181 2107
rect 24360 2127 24391 2169
rect 24360 2108 24365 2127
rect 24386 2108 24391 2127
rect 24360 2102 24391 2108
rect 25022 2122 25056 2328
rect 26795 2325 26830 2332
rect 25090 2301 25675 2307
rect 25090 2281 25106 2301
rect 25126 2300 25675 2301
rect 25126 2281 25646 2300
rect 25090 2280 25646 2281
rect 25666 2280 25675 2300
rect 25090 2272 25675 2280
rect 26795 2305 26803 2325
rect 26823 2305 26830 2325
rect 26795 2232 26830 2305
rect 27009 2327 27065 2332
rect 27009 2307 27016 2327
rect 27036 2307 27065 2327
rect 27009 2300 27065 2307
rect 27100 2434 27130 2436
rect 27829 2434 27862 2435
rect 27100 2408 27863 2434
rect 27009 2299 27044 2300
rect 27100 2233 27130 2408
rect 27829 2387 27863 2408
rect 27828 2382 27863 2387
rect 27828 2362 27835 2382
rect 27855 2362 27863 2382
rect 27828 2354 27863 2362
rect 27095 2232 27130 2233
rect 26794 2205 27130 2232
rect 27100 2204 27130 2205
rect 27210 2196 27795 2204
rect 27210 2176 27219 2196
rect 27239 2195 27795 2196
rect 27239 2176 27759 2195
rect 27210 2175 27759 2176
rect 27779 2175 27795 2195
rect 27210 2169 27795 2175
rect 27034 2159 27066 2160
rect 27031 2154 27066 2159
rect 27031 2134 27038 2154
rect 27058 2134 27066 2154
rect 27829 2148 27863 2354
rect 27031 2126 27066 2134
rect 25022 2114 25057 2122
rect 24125 1896 24159 2102
rect 25022 2094 25030 2114
rect 25050 2094 25057 2114
rect 25022 2089 25057 2094
rect 25022 2088 25054 2089
rect 24193 2075 24778 2081
rect 24193 2055 24209 2075
rect 24229 2074 24778 2075
rect 24229 2055 24749 2074
rect 24193 2054 24749 2055
rect 24769 2054 24778 2074
rect 24193 2046 24778 2054
rect 26413 1968 26998 1976
rect 26413 1948 26422 1968
rect 26442 1967 26998 1968
rect 26442 1948 26962 1967
rect 26413 1947 26962 1948
rect 26982 1947 26998 1967
rect 26413 1941 26998 1947
rect 26787 1917 26826 1921
rect 27032 1920 27066 2126
rect 27595 2141 27630 2147
rect 27595 2122 27600 2141
rect 27621 2122 27630 2141
rect 27595 2113 27630 2122
rect 27807 2143 27863 2148
rect 27807 2123 27814 2143
rect 27834 2123 27863 2143
rect 27807 2116 27863 2123
rect 27985 2294 28017 2306
rect 27985 2276 27992 2294
rect 28014 2276 28017 2294
rect 27807 2115 27842 2116
rect 27599 2045 27628 2113
rect 27599 2011 27945 2045
rect 26787 1897 26795 1917
rect 26815 1897 26826 1917
rect 24125 1888 24160 1896
rect 24125 1868 24133 1888
rect 24153 1880 24160 1888
rect 24153 1868 24164 1880
rect 24125 1631 24164 1868
rect 24995 1845 25281 1846
rect 24480 1837 25283 1845
rect 24480 1820 24491 1837
rect 24481 1815 24491 1820
rect 24515 1820 25283 1837
rect 24515 1815 24520 1820
rect 24481 1802 24520 1815
rect 25025 1754 25060 1755
rect 25004 1747 25060 1754
rect 25004 1727 25033 1747
rect 25053 1727 25060 1747
rect 25004 1722 25060 1727
rect 25244 1745 25283 1820
rect 26787 1822 26826 1897
rect 27010 1915 27066 1920
rect 27010 1895 27017 1915
rect 27037 1895 27066 1915
rect 27010 1888 27066 1895
rect 27010 1887 27045 1888
rect 27550 1827 27589 1840
rect 27550 1822 27555 1827
rect 26787 1805 27555 1822
rect 27579 1822 27589 1827
rect 27579 1805 27590 1822
rect 26787 1797 27590 1805
rect 26789 1796 27075 1797
rect 27906 1774 27945 2011
rect 27906 1762 27917 1774
rect 27910 1754 27917 1762
rect 27937 1754 27945 1774
rect 27910 1746 27945 1754
rect 25244 1725 25255 1745
rect 25275 1725 25283 1745
rect 24125 1597 24471 1631
rect 24442 1529 24471 1597
rect 24228 1526 24263 1527
rect 23306 1427 23640 1455
rect 24207 1519 24263 1526
rect 24207 1499 24236 1519
rect 24256 1499 24263 1519
rect 24207 1494 24263 1499
rect 24440 1520 24475 1529
rect 24440 1501 24449 1520
rect 24470 1501 24475 1520
rect 24440 1495 24475 1501
rect 25004 1516 25038 1722
rect 25244 1721 25283 1725
rect 25072 1695 25657 1701
rect 25072 1675 25088 1695
rect 25108 1694 25657 1695
rect 25108 1675 25628 1694
rect 25072 1674 25628 1675
rect 25648 1674 25657 1694
rect 25072 1666 25657 1674
rect 27292 1588 27877 1596
rect 27292 1568 27301 1588
rect 27321 1587 27877 1588
rect 27321 1568 27841 1587
rect 27292 1567 27841 1568
rect 27861 1567 27877 1587
rect 27292 1561 27877 1567
rect 27016 1553 27048 1554
rect 27013 1548 27048 1553
rect 27013 1528 27020 1548
rect 27040 1528 27048 1548
rect 27911 1540 27945 1746
rect 27013 1520 27048 1528
rect 25004 1508 25039 1516
rect 16375 1083 16407 1084
rect 18273 1083 18308 1091
rect 14576 1058 14958 1066
rect 14576 1039 14929 1058
rect 14950 1039 14958 1058
rect 14576 1034 14958 1039
rect 13763 880 13771 900
rect 13791 880 13802 900
rect 9622 857 9657 858
rect 10857 810 10908 841
rect 10162 797 10201 810
rect 10162 792 10167 797
rect 9399 775 10167 792
rect 10191 792 10201 797
rect 10191 775 10202 792
rect 9399 767 10202 775
rect 10857 784 10874 810
rect 10902 784 10908 810
rect 9401 766 9687 767
rect 10857 761 10908 784
rect 10937 816 10983 847
rect 12781 845 12824 853
rect 10937 785 10951 816
rect 10979 785 10983 816
rect 10937 778 10983 785
rect 12775 838 12830 845
rect 12775 813 12788 838
rect 12820 813 12830 838
rect 8398 677 8409 709
rect 8449 677 8453 709
rect 9239 750 9300 759
rect 9239 723 9247 750
rect 9283 744 9300 750
rect 9341 744 9416 748
rect 9283 742 9416 744
rect 9283 723 9347 742
rect 9239 706 9347 723
rect 9392 706 9416 742
rect 9239 704 9416 706
rect 8398 664 8453 677
rect 9341 674 9416 704
rect 10870 569 10901 761
rect 10856 548 10902 569
rect 10856 527 10863 548
rect 10884 527 10902 548
rect 10856 523 10902 527
rect 10856 520 10891 523
rect 9066 495 9097 500
rect 6562 422 6568 442
rect 6588 422 6596 442
rect 6562 416 6596 422
rect 8268 475 9102 495
rect 6239 273 6255 297
rect 6278 273 6290 297
rect 6239 264 6290 273
rect 6458 297 6514 302
rect 6458 277 6465 297
rect 6485 277 6514 297
rect 6458 270 6514 277
rect 6458 269 6493 270
rect 6243 198 6286 264
rect 4583 182 4618 183
rect 4373 117 4401 177
rect 5746 170 6286 198
rect 5749 168 6286 170
rect 6243 166 6286 168
rect 8268 117 8294 475
rect 9052 473 9098 475
rect 9052 452 9059 473
rect 9080 452 9098 473
rect 9132 465 10061 498
rect 9052 448 9098 452
rect 9052 445 9087 448
rect 8434 287 9019 295
rect 8434 267 8443 287
rect 8463 286 9019 287
rect 8463 267 8983 286
rect 8434 266 8983 267
rect 9003 266 9019 286
rect 8434 260 9019 266
rect 9053 239 9087 445
rect 9134 379 9177 465
rect 9261 459 10061 465
rect 9134 359 9141 379
rect 9161 359 9177 379
rect 9134 348 9177 359
rect 8810 227 8856 237
rect 8810 209 8819 227
rect 8840 209 8856 227
rect 8810 204 8856 209
rect 9031 234 9087 239
rect 9031 214 9038 234
rect 9058 214 9087 234
rect 9031 207 9087 214
rect 9031 206 9066 207
rect 8815 141 8849 204
rect 8815 139 8850 141
rect 8815 128 8868 139
rect 8815 117 8824 128
rect 4373 83 8299 117
rect 8816 97 8824 117
rect 8853 97 8868 128
rect 8816 85 8868 97
rect 10022 46 10061 459
rect 10238 362 10823 370
rect 10238 342 10247 362
rect 10267 361 10823 362
rect 10267 342 10787 361
rect 10238 341 10787 342
rect 10807 341 10823 361
rect 10238 335 10823 341
rect 10857 314 10891 520
rect 10939 454 10973 778
rect 12775 721 12830 813
rect 13763 805 13802 880
rect 13986 898 14042 903
rect 17655 925 18240 933
rect 17655 905 17664 925
rect 17684 924 18240 925
rect 17684 905 18204 924
rect 17655 904 18204 905
rect 18224 904 18240 924
rect 17655 898 18240 904
rect 13986 878 13993 898
rect 14013 878 14042 898
rect 13986 871 14042 878
rect 18029 874 18068 878
rect 18274 877 18308 1083
rect 18838 1095 18872 1103
rect 18838 1077 18845 1095
rect 18864 1077 18872 1095
rect 18838 1070 18872 1077
rect 19049 1100 19105 1105
rect 19049 1080 19056 1100
rect 19076 1080 19105 1100
rect 19049 1073 19105 1080
rect 20641 1091 20675 1297
rect 22401 1295 22436 1302
rect 20709 1270 21294 1276
rect 20709 1250 20725 1270
rect 20745 1269 21294 1270
rect 20745 1250 21265 1269
rect 20709 1249 21265 1250
rect 21285 1249 21294 1269
rect 20709 1241 21294 1249
rect 22401 1275 22409 1295
rect 22429 1275 22436 1295
rect 22401 1202 22436 1275
rect 22615 1297 22671 1302
rect 22615 1277 22622 1297
rect 22642 1277 22671 1297
rect 22615 1270 22671 1277
rect 22706 1404 22736 1406
rect 23435 1404 23468 1405
rect 22706 1378 23469 1404
rect 22615 1269 22650 1270
rect 22706 1203 22736 1378
rect 23435 1357 23469 1378
rect 23434 1352 23469 1357
rect 23434 1332 23441 1352
rect 23461 1332 23469 1352
rect 23434 1324 23469 1332
rect 22701 1202 22736 1203
rect 22400 1175 22736 1202
rect 22706 1174 22736 1175
rect 22816 1166 23401 1174
rect 22816 1146 22825 1166
rect 22845 1165 23401 1166
rect 22845 1146 23365 1165
rect 22816 1145 23365 1146
rect 23385 1145 23401 1165
rect 22816 1139 23401 1145
rect 22640 1129 22672 1130
rect 22637 1124 22672 1129
rect 22637 1104 22644 1124
rect 22664 1104 22672 1124
rect 23435 1118 23469 1324
rect 24207 1288 24241 1494
rect 25004 1488 25012 1508
rect 25032 1488 25039 1508
rect 25004 1483 25039 1488
rect 25004 1482 25036 1483
rect 24275 1467 24860 1473
rect 24275 1447 24291 1467
rect 24311 1466 24860 1467
rect 24311 1447 24831 1466
rect 24275 1446 24831 1447
rect 24851 1446 24860 1466
rect 24275 1438 24860 1446
rect 24940 1437 24970 1438
rect 24940 1410 25276 1437
rect 24940 1409 24975 1410
rect 24207 1280 24242 1288
rect 24207 1260 24215 1280
rect 24235 1260 24242 1280
rect 24207 1255 24242 1260
rect 24207 1234 24241 1255
rect 24940 1234 24970 1409
rect 25026 1342 25061 1343
rect 24207 1208 24970 1234
rect 24208 1207 24241 1208
rect 24940 1206 24970 1208
rect 25005 1335 25061 1342
rect 25005 1315 25034 1335
rect 25054 1315 25061 1335
rect 25005 1310 25061 1315
rect 25240 1337 25275 1410
rect 25240 1317 25247 1337
rect 25267 1317 25275 1337
rect 26395 1362 26980 1370
rect 26395 1342 26404 1362
rect 26424 1361 26980 1362
rect 26424 1342 26944 1361
rect 26395 1341 26944 1342
rect 26964 1341 26980 1361
rect 26395 1335 26980 1341
rect 25240 1310 25275 1317
rect 27014 1314 27048 1520
rect 27677 1528 27713 1537
rect 27677 1511 27686 1528
rect 27705 1511 27713 1528
rect 27677 1502 27713 1511
rect 27889 1535 27945 1540
rect 27889 1515 27896 1535
rect 27916 1515 27945 1535
rect 27889 1508 27945 1515
rect 27889 1507 27924 1508
rect 27683 1467 27709 1502
rect 27985 1467 28017 2276
rect 28429 2209 28458 2894
rect 29389 2875 29675 2876
rect 28874 2867 29677 2875
rect 28874 2850 28885 2867
rect 28875 2845 28885 2850
rect 28909 2850 29677 2867
rect 28909 2845 28914 2850
rect 28875 2832 28914 2845
rect 29419 2784 29454 2785
rect 29398 2777 29454 2784
rect 29398 2757 29427 2777
rect 29447 2757 29454 2777
rect 29398 2752 29454 2757
rect 29638 2775 29677 2850
rect 31171 2853 31210 2928
rect 31394 2946 31450 2951
rect 31394 2926 31401 2946
rect 31421 2926 31450 2946
rect 31394 2919 31450 2926
rect 31394 2918 31429 2919
rect 31934 2858 31973 2871
rect 31934 2853 31939 2858
rect 31171 2836 31939 2853
rect 31963 2853 31973 2858
rect 31963 2836 31974 2853
rect 31171 2828 31974 2836
rect 31173 2827 31459 2828
rect 32390 2809 32419 3494
rect 32727 3248 32754 4948
rect 33790 4924 34076 4925
rect 33275 4916 34078 4924
rect 33275 4899 33286 4916
rect 33276 4894 33286 4899
rect 33310 4899 34078 4916
rect 33310 4894 33315 4899
rect 33276 4881 33315 4894
rect 33820 4833 33855 4834
rect 33799 4826 33855 4833
rect 33799 4806 33828 4826
rect 33848 4806 33855 4826
rect 33799 4801 33855 4806
rect 34039 4824 34078 4899
rect 34039 4804 34050 4824
rect 34070 4804 34078 4824
rect 32883 4665 33265 4670
rect 32883 4646 32891 4665
rect 32912 4646 33265 4665
rect 32883 4638 33265 4646
rect 33236 4608 33265 4638
rect 33023 4605 33058 4606
rect 33002 4598 33058 4605
rect 33002 4578 33031 4598
rect 33051 4578 33058 4598
rect 33002 4573 33058 4578
rect 33235 4601 33269 4608
rect 33235 4583 33243 4601
rect 33262 4583 33269 4601
rect 33235 4575 33269 4583
rect 33799 4595 33833 4801
rect 34039 4800 34078 4804
rect 33867 4774 34452 4780
rect 33867 4754 33883 4774
rect 33903 4773 34452 4774
rect 33903 4754 34423 4773
rect 33867 4753 34423 4754
rect 34443 4753 34452 4773
rect 33867 4745 34452 4753
rect 33799 4587 33834 4595
rect 33002 4367 33036 4573
rect 33799 4567 33807 4587
rect 33827 4567 33834 4587
rect 33799 4562 33834 4567
rect 33799 4561 33831 4562
rect 33070 4546 33655 4552
rect 33070 4526 33086 4546
rect 33106 4545 33655 4546
rect 33106 4526 33626 4545
rect 33070 4525 33626 4526
rect 33646 4525 33655 4545
rect 33070 4517 33655 4525
rect 33735 4516 33765 4517
rect 33735 4489 34071 4516
rect 33735 4488 33770 4489
rect 33002 4359 33037 4367
rect 33002 4339 33010 4359
rect 33030 4339 33037 4359
rect 33002 4334 33037 4339
rect 33002 4313 33036 4334
rect 33735 4313 33765 4488
rect 33821 4421 33856 4422
rect 33002 4287 33765 4313
rect 33003 4286 33036 4287
rect 33735 4285 33765 4287
rect 33800 4414 33856 4421
rect 33800 4394 33829 4414
rect 33849 4394 33856 4414
rect 33800 4389 33856 4394
rect 34035 4416 34070 4489
rect 34035 4396 34042 4416
rect 34062 4396 34070 4416
rect 34035 4389 34070 4396
rect 32825 4264 32857 4265
rect 32825 4259 33165 4264
rect 32825 4241 32828 4259
rect 32850 4241 33165 4259
rect 32825 4236 33165 4241
rect 32825 4235 32857 4236
rect 33139 4201 33165 4236
rect 32924 4195 32959 4196
rect 32903 4188 32959 4195
rect 32903 4168 32932 4188
rect 32952 4168 32959 4188
rect 32903 4163 32959 4168
rect 33135 4192 33171 4201
rect 33135 4175 33143 4192
rect 33162 4175 33171 4192
rect 33135 4166 33171 4175
rect 33800 4183 33834 4389
rect 33868 4362 34453 4368
rect 33868 4342 33884 4362
rect 33904 4361 34453 4362
rect 33904 4342 34424 4361
rect 33868 4341 34424 4342
rect 34444 4341 34453 4361
rect 33868 4333 34453 4341
rect 33800 4175 33835 4183
rect 32903 3957 32937 4163
rect 33800 4155 33808 4175
rect 33828 4155 33835 4175
rect 33800 4150 33835 4155
rect 33800 4149 33832 4150
rect 32971 4136 33556 4142
rect 32971 4116 32987 4136
rect 33007 4135 33556 4136
rect 33007 4116 33527 4135
rect 32971 4115 33527 4116
rect 33547 4115 33556 4135
rect 32971 4107 33556 4115
rect 32903 3949 32938 3957
rect 32903 3929 32911 3949
rect 32931 3941 32938 3949
rect 32931 3929 32942 3941
rect 32903 3692 32942 3929
rect 33773 3906 34059 3907
rect 33258 3898 34061 3906
rect 33258 3881 33269 3898
rect 33259 3876 33269 3881
rect 33293 3881 34061 3898
rect 33293 3876 33298 3881
rect 33259 3863 33298 3876
rect 33803 3815 33838 3816
rect 33782 3808 33838 3815
rect 33782 3788 33811 3808
rect 33831 3788 33838 3808
rect 33782 3783 33838 3788
rect 34022 3806 34061 3881
rect 34022 3786 34033 3806
rect 34053 3786 34061 3806
rect 32903 3658 33249 3692
rect 33220 3590 33249 3658
rect 33006 3587 33041 3588
rect 32985 3580 33041 3587
rect 32985 3560 33014 3580
rect 33034 3560 33041 3580
rect 32985 3555 33041 3560
rect 33218 3581 33253 3590
rect 33218 3562 33227 3581
rect 33248 3562 33253 3581
rect 33218 3556 33253 3562
rect 33782 3577 33816 3783
rect 34022 3782 34061 3786
rect 33850 3756 34435 3762
rect 33850 3736 33866 3756
rect 33886 3755 34435 3756
rect 33886 3736 34406 3755
rect 33850 3735 34406 3736
rect 34426 3735 34435 3755
rect 33850 3727 34435 3735
rect 33782 3569 33817 3577
rect 32985 3349 33019 3555
rect 33782 3549 33790 3569
rect 33810 3549 33817 3569
rect 33782 3544 33817 3549
rect 33782 3543 33814 3544
rect 33053 3528 33638 3534
rect 33053 3508 33069 3528
rect 33089 3527 33638 3528
rect 33089 3508 33609 3527
rect 33053 3507 33609 3508
rect 33629 3507 33638 3527
rect 33053 3499 33638 3507
rect 33718 3498 33748 3499
rect 33718 3471 34054 3498
rect 33718 3470 33753 3471
rect 32985 3341 33020 3349
rect 32985 3321 32993 3341
rect 33013 3321 33020 3341
rect 32985 3316 33020 3321
rect 32985 3295 33019 3316
rect 33718 3295 33748 3470
rect 33804 3403 33839 3404
rect 32985 3269 33748 3295
rect 32986 3268 33019 3269
rect 33718 3267 33748 3269
rect 33783 3396 33839 3403
rect 33783 3376 33812 3396
rect 33832 3376 33839 3396
rect 33783 3371 33839 3376
rect 34018 3398 34053 3471
rect 34018 3378 34025 3398
rect 34045 3378 34053 3398
rect 34018 3371 34053 3378
rect 32727 3212 33081 3248
rect 32743 3211 33081 3212
rect 33055 3181 33081 3211
rect 32841 3179 32876 3180
rect 32820 3172 32876 3179
rect 32820 3152 32849 3172
rect 32869 3152 32876 3172
rect 32820 3147 32876 3152
rect 33049 3173 33090 3181
rect 33049 3155 33062 3173
rect 33080 3155 33090 3173
rect 32820 2941 32854 3147
rect 33049 3144 33090 3155
rect 33783 3165 33817 3371
rect 33851 3344 34436 3350
rect 33851 3324 33867 3344
rect 33887 3343 34436 3344
rect 33887 3324 34407 3343
rect 33851 3323 34407 3324
rect 34427 3323 34436 3343
rect 33851 3315 34436 3323
rect 33783 3157 33818 3165
rect 33783 3137 33791 3157
rect 33811 3137 33818 3157
rect 33783 3132 33818 3137
rect 33783 3131 33815 3132
rect 32888 3120 33473 3126
rect 32888 3100 32904 3120
rect 32924 3119 33473 3120
rect 32924 3100 33444 3119
rect 32888 3099 33444 3100
rect 33464 3099 33473 3119
rect 32888 3091 33473 3099
rect 32820 2940 32855 2941
rect 32788 2933 32855 2940
rect 32788 2913 32828 2933
rect 32848 2913 32855 2933
rect 32788 2910 32855 2913
rect 32788 2907 32853 2910
rect 32359 2806 32424 2809
rect 32357 2803 32424 2806
rect 32357 2783 32364 2803
rect 32384 2783 32424 2803
rect 32357 2776 32424 2783
rect 32357 2775 32392 2776
rect 29638 2755 29649 2775
rect 29669 2755 29677 2775
rect 28482 2616 28864 2621
rect 28482 2597 28490 2616
rect 28511 2597 28864 2616
rect 28482 2589 28864 2597
rect 28835 2559 28864 2589
rect 28622 2556 28657 2557
rect 28601 2549 28657 2556
rect 28601 2529 28630 2549
rect 28650 2529 28657 2549
rect 28601 2524 28657 2529
rect 28834 2552 28868 2559
rect 28834 2534 28842 2552
rect 28861 2534 28868 2552
rect 28834 2526 28868 2534
rect 29398 2546 29432 2752
rect 29638 2751 29677 2755
rect 29466 2725 30051 2731
rect 29466 2705 29482 2725
rect 29502 2724 30051 2725
rect 29502 2705 30022 2724
rect 29466 2704 30022 2705
rect 30042 2704 30051 2724
rect 29466 2696 30051 2704
rect 31739 2617 32324 2625
rect 31739 2597 31748 2617
rect 31768 2616 32324 2617
rect 31768 2597 32288 2616
rect 31739 2596 32288 2597
rect 32308 2596 32324 2616
rect 31739 2590 32324 2596
rect 31397 2584 31429 2585
rect 31394 2579 31429 2584
rect 31394 2559 31401 2579
rect 31421 2559 31429 2579
rect 31394 2551 31429 2559
rect 29398 2538 29433 2546
rect 28601 2318 28635 2524
rect 29398 2518 29406 2538
rect 29426 2518 29433 2538
rect 29398 2513 29433 2518
rect 29398 2512 29430 2513
rect 28669 2497 29254 2503
rect 28669 2477 28685 2497
rect 28705 2496 29254 2497
rect 28705 2477 29225 2496
rect 28669 2476 29225 2477
rect 29245 2476 29254 2496
rect 28669 2468 29254 2476
rect 29334 2467 29364 2468
rect 29334 2440 29670 2467
rect 29334 2439 29369 2440
rect 28601 2310 28636 2318
rect 28601 2290 28609 2310
rect 28629 2290 28636 2310
rect 28601 2285 28636 2290
rect 28601 2264 28635 2285
rect 29334 2264 29364 2439
rect 29420 2372 29455 2373
rect 28601 2238 29364 2264
rect 28602 2237 28635 2238
rect 29334 2236 29364 2238
rect 29399 2365 29455 2372
rect 29399 2345 29428 2365
rect 29448 2345 29455 2365
rect 29399 2340 29455 2345
rect 29634 2367 29669 2440
rect 29634 2347 29641 2367
rect 29661 2347 29669 2367
rect 30776 2393 31361 2401
rect 30776 2373 30785 2393
rect 30805 2392 31361 2393
rect 30805 2373 31325 2392
rect 30776 2372 31325 2373
rect 31345 2372 31361 2392
rect 30776 2366 31361 2372
rect 29634 2340 29669 2347
rect 31395 2345 31429 2551
rect 32124 2566 32157 2572
rect 32358 2569 32392 2775
rect 32124 2544 32129 2566
rect 32152 2544 32157 2566
rect 32124 2535 32157 2544
rect 32336 2564 32392 2569
rect 32336 2544 32343 2564
rect 32363 2544 32392 2564
rect 32336 2537 32392 2544
rect 32336 2536 32371 2537
rect 32126 2504 32153 2535
rect 32548 2504 32587 2516
rect 32126 2503 32589 2504
rect 32126 2481 32553 2503
rect 32577 2481 32589 2503
rect 32126 2473 32589 2481
rect 28429 2181 28768 2209
rect 28523 2146 28558 2147
rect 28502 2139 28558 2146
rect 28502 2119 28531 2139
rect 28551 2119 28558 2139
rect 28502 2114 28558 2119
rect 28737 2139 28768 2181
rect 28737 2120 28742 2139
rect 28763 2120 28768 2139
rect 28737 2114 28768 2120
rect 29399 2134 29433 2340
rect 31159 2338 31194 2345
rect 29467 2313 30052 2319
rect 29467 2293 29483 2313
rect 29503 2312 30052 2313
rect 29503 2293 30023 2312
rect 29467 2292 30023 2293
rect 30043 2292 30052 2312
rect 29467 2284 30052 2292
rect 31159 2318 31167 2338
rect 31187 2318 31194 2338
rect 31159 2245 31194 2318
rect 31373 2340 31429 2345
rect 31373 2320 31380 2340
rect 31400 2320 31429 2340
rect 31373 2313 31429 2320
rect 31464 2447 31494 2449
rect 32193 2447 32226 2448
rect 31464 2421 32227 2447
rect 31373 2312 31408 2313
rect 31464 2246 31494 2421
rect 32193 2400 32227 2421
rect 32192 2395 32227 2400
rect 32192 2375 32199 2395
rect 32219 2375 32227 2395
rect 32192 2367 32227 2375
rect 31459 2245 31494 2246
rect 31158 2218 31494 2245
rect 31464 2217 31494 2218
rect 31574 2209 32159 2217
rect 31574 2189 31583 2209
rect 31603 2208 32159 2209
rect 31603 2189 32123 2208
rect 31574 2188 32123 2189
rect 32143 2188 32159 2208
rect 31574 2182 32159 2188
rect 31398 2172 31430 2173
rect 31395 2167 31430 2172
rect 31395 2147 31402 2167
rect 31422 2147 31430 2167
rect 32193 2161 32227 2367
rect 31395 2139 31430 2147
rect 29399 2126 29434 2134
rect 28502 1908 28536 2114
rect 29399 2106 29407 2126
rect 29427 2106 29434 2126
rect 29399 2101 29434 2106
rect 29399 2100 29431 2101
rect 28570 2087 29155 2093
rect 28570 2067 28586 2087
rect 28606 2086 29155 2087
rect 28606 2067 29126 2086
rect 28570 2066 29126 2067
rect 29146 2066 29155 2086
rect 28570 2058 29155 2066
rect 30777 1981 31362 1989
rect 30777 1961 30786 1981
rect 30806 1980 31362 1981
rect 30806 1961 31326 1980
rect 30777 1960 31326 1961
rect 31346 1960 31362 1980
rect 30777 1954 31362 1960
rect 31151 1930 31190 1934
rect 31396 1933 31430 2139
rect 31959 2154 31994 2160
rect 31959 2135 31964 2154
rect 31985 2135 31994 2154
rect 31959 2126 31994 2135
rect 32171 2156 32227 2161
rect 32171 2136 32178 2156
rect 32198 2136 32227 2156
rect 32171 2129 32227 2136
rect 32349 2307 32381 2319
rect 32349 2289 32356 2307
rect 32378 2289 32381 2307
rect 32171 2128 32206 2129
rect 31963 2058 31992 2126
rect 31963 2024 32309 2058
rect 31151 1910 31159 1930
rect 31179 1910 31190 1930
rect 28502 1900 28537 1908
rect 28502 1880 28510 1900
rect 28530 1892 28537 1900
rect 28530 1880 28541 1892
rect 28502 1643 28541 1880
rect 29372 1857 29658 1858
rect 28857 1849 29660 1857
rect 28857 1832 28868 1849
rect 28858 1827 28868 1832
rect 28892 1832 29660 1849
rect 28892 1827 28897 1832
rect 28858 1814 28897 1827
rect 29402 1766 29437 1767
rect 29381 1759 29437 1766
rect 29381 1739 29410 1759
rect 29430 1739 29437 1759
rect 29381 1734 29437 1739
rect 29621 1757 29660 1832
rect 31151 1835 31190 1910
rect 31374 1928 31430 1933
rect 31374 1908 31381 1928
rect 31401 1908 31430 1928
rect 31374 1901 31430 1908
rect 31374 1900 31409 1901
rect 31914 1840 31953 1853
rect 31914 1835 31919 1840
rect 31151 1818 31919 1835
rect 31943 1835 31953 1840
rect 31943 1818 31954 1835
rect 31151 1810 31954 1818
rect 31153 1809 31439 1810
rect 32270 1787 32309 2024
rect 32270 1775 32281 1787
rect 32274 1767 32281 1775
rect 32301 1767 32309 1787
rect 32274 1759 32309 1767
rect 29621 1737 29632 1757
rect 29652 1737 29660 1757
rect 28502 1609 28848 1643
rect 28819 1541 28848 1609
rect 28605 1538 28640 1539
rect 27683 1439 28017 1467
rect 28584 1531 28640 1538
rect 28584 1511 28613 1531
rect 28633 1511 28640 1531
rect 28584 1506 28640 1511
rect 28817 1532 28852 1541
rect 28817 1513 28826 1532
rect 28847 1513 28852 1532
rect 28817 1507 28852 1513
rect 29381 1528 29415 1734
rect 29621 1733 29660 1737
rect 29449 1707 30034 1713
rect 29449 1687 29465 1707
rect 29485 1706 30034 1707
rect 29485 1687 30005 1706
rect 29449 1686 30005 1687
rect 30025 1686 30034 1706
rect 29449 1678 30034 1686
rect 31656 1601 32241 1609
rect 31656 1581 31665 1601
rect 31685 1600 32241 1601
rect 31685 1581 32205 1600
rect 31656 1580 32205 1581
rect 32225 1580 32241 1600
rect 31656 1574 32241 1580
rect 31380 1566 31412 1567
rect 31377 1561 31412 1566
rect 31377 1541 31384 1561
rect 31404 1541 31412 1561
rect 32275 1553 32309 1759
rect 31377 1533 31412 1541
rect 29381 1520 29416 1528
rect 22637 1096 22672 1104
rect 20641 1083 20676 1091
rect 19049 1072 19084 1073
rect 18842 1040 18871 1070
rect 20641 1063 20649 1083
rect 20669 1063 20676 1083
rect 20641 1058 20676 1063
rect 20641 1057 20673 1058
rect 18842 1032 19224 1040
rect 18842 1013 19195 1032
rect 19216 1013 19224 1032
rect 18842 1008 19224 1013
rect 22019 938 22604 946
rect 22019 918 22028 938
rect 22048 937 22604 938
rect 22048 918 22568 937
rect 22019 917 22568 918
rect 22588 917 22604 937
rect 22019 911 22604 917
rect 13986 870 14021 871
rect 15221 823 15272 854
rect 14526 810 14565 823
rect 14526 805 14531 810
rect 13763 788 14531 805
rect 14555 805 14565 810
rect 14555 788 14566 805
rect 13763 780 14566 788
rect 15221 797 15238 823
rect 15266 797 15272 823
rect 13765 779 14051 780
rect 15221 774 15272 797
rect 15301 829 15347 860
rect 17145 858 17188 866
rect 15301 798 15315 829
rect 15343 798 15347 829
rect 15301 791 15347 798
rect 17139 851 17194 858
rect 17139 826 17152 851
rect 17184 826 17194 851
rect 12775 689 12786 721
rect 12826 689 12830 721
rect 13603 763 13664 772
rect 13603 736 13611 763
rect 13647 757 13664 763
rect 13705 757 13780 761
rect 13647 755 13780 757
rect 13647 736 13711 755
rect 13603 719 13711 736
rect 13756 719 13780 755
rect 13603 717 13780 719
rect 12775 676 12830 689
rect 13705 687 13780 717
rect 15234 582 15265 774
rect 15220 561 15266 582
rect 15220 540 15227 561
rect 15248 540 15266 561
rect 15220 536 15266 540
rect 15220 533 15255 536
rect 13359 496 13390 501
rect 10939 434 10945 454
rect 10965 434 10973 454
rect 10939 428 10973 434
rect 12561 476 13395 496
rect 10618 308 10661 312
rect 10618 284 10629 308
rect 10652 284 10661 308
rect 10618 280 10661 284
rect 10835 309 10891 314
rect 10835 289 10842 309
rect 10862 289 10891 309
rect 10835 282 10891 289
rect 10835 281 10870 282
rect 10625 216 10656 280
rect 12561 216 12587 476
rect 13345 474 13391 476
rect 13345 453 13352 474
rect 13373 453 13391 474
rect 13425 466 14518 499
rect 13345 449 13391 453
rect 13345 446 13380 449
rect 12727 288 13312 296
rect 12727 268 12736 288
rect 12756 287 13312 288
rect 12756 268 13276 287
rect 12727 267 13276 268
rect 13296 267 13312 287
rect 12727 261 13312 267
rect 13346 240 13380 446
rect 13427 380 13470 466
rect 13427 360 13434 380
rect 13454 360 13470 380
rect 13427 349 13470 360
rect 13105 233 13157 239
rect 10625 193 12588 216
rect 10633 191 12588 193
rect 13105 211 13117 233
rect 13138 211 13157 233
rect 13105 46 13157 211
rect 13324 235 13380 240
rect 13324 215 13331 235
rect 13351 215 13380 235
rect 13324 208 13380 215
rect 14487 223 14516 466
rect 14602 375 15187 383
rect 14602 355 14611 375
rect 14631 374 15187 375
rect 14631 355 15151 374
rect 14602 354 15151 355
rect 15171 354 15187 374
rect 14602 348 15187 354
rect 14984 328 15027 330
rect 14980 322 15031 328
rect 15221 327 15255 533
rect 15303 467 15337 791
rect 17139 734 17194 826
rect 18029 854 18037 874
rect 18057 854 18068 874
rect 18029 779 18068 854
rect 18252 872 18308 877
rect 18252 852 18259 872
rect 18279 852 18308 872
rect 18252 845 18308 852
rect 22393 887 22432 891
rect 22638 890 22672 1096
rect 23202 1108 23236 1116
rect 23202 1090 23209 1108
rect 23228 1090 23236 1108
rect 23202 1083 23236 1090
rect 23413 1113 23469 1118
rect 23413 1093 23420 1113
rect 23440 1093 23469 1113
rect 23413 1086 23469 1093
rect 25005 1104 25039 1310
rect 26778 1307 26813 1314
rect 25073 1283 25658 1289
rect 25073 1263 25089 1283
rect 25109 1282 25658 1283
rect 25109 1263 25629 1282
rect 25073 1262 25629 1263
rect 25649 1262 25658 1282
rect 25073 1254 25658 1262
rect 26778 1287 26786 1307
rect 26806 1287 26813 1307
rect 26778 1214 26813 1287
rect 26992 1309 27048 1314
rect 26992 1289 26999 1309
rect 27019 1289 27048 1309
rect 26992 1282 27048 1289
rect 27083 1416 27113 1418
rect 27812 1416 27845 1417
rect 27083 1390 27846 1416
rect 26992 1281 27027 1282
rect 27083 1215 27113 1390
rect 27812 1369 27846 1390
rect 27811 1364 27846 1369
rect 27811 1344 27818 1364
rect 27838 1344 27846 1364
rect 27811 1336 27846 1344
rect 27078 1214 27113 1215
rect 26777 1187 27113 1214
rect 27083 1186 27113 1187
rect 27193 1178 27778 1186
rect 27193 1158 27202 1178
rect 27222 1177 27778 1178
rect 27222 1158 27742 1177
rect 27193 1157 27742 1158
rect 27762 1157 27778 1177
rect 27193 1151 27778 1157
rect 27017 1141 27049 1142
rect 27014 1136 27049 1141
rect 27014 1116 27021 1136
rect 27041 1116 27049 1136
rect 27812 1130 27846 1336
rect 28584 1300 28618 1506
rect 29381 1500 29389 1520
rect 29409 1500 29416 1520
rect 29381 1495 29416 1500
rect 29381 1494 29413 1495
rect 28652 1479 29237 1485
rect 28652 1459 28668 1479
rect 28688 1478 29237 1479
rect 28688 1459 29208 1478
rect 28652 1458 29208 1459
rect 29228 1458 29237 1478
rect 28652 1450 29237 1458
rect 29317 1449 29347 1450
rect 29317 1422 29653 1449
rect 29317 1421 29352 1422
rect 28584 1292 28619 1300
rect 28584 1272 28592 1292
rect 28612 1272 28619 1292
rect 28584 1267 28619 1272
rect 28584 1246 28618 1267
rect 29317 1246 29347 1421
rect 29403 1354 29438 1355
rect 28584 1220 29347 1246
rect 28585 1219 28618 1220
rect 29317 1218 29347 1220
rect 29382 1347 29438 1354
rect 29382 1327 29411 1347
rect 29431 1327 29438 1347
rect 29382 1322 29438 1327
rect 29617 1349 29652 1422
rect 29617 1329 29624 1349
rect 29644 1329 29652 1349
rect 30759 1375 31344 1383
rect 30759 1355 30768 1375
rect 30788 1374 31344 1375
rect 30788 1355 31308 1374
rect 30759 1354 31308 1355
rect 31328 1354 31344 1374
rect 30759 1348 31344 1354
rect 29617 1322 29652 1329
rect 31378 1327 31412 1533
rect 32041 1541 32077 1550
rect 32041 1524 32050 1541
rect 32069 1524 32077 1541
rect 32041 1515 32077 1524
rect 32253 1548 32309 1553
rect 32253 1528 32260 1548
rect 32280 1528 32309 1548
rect 32253 1521 32309 1528
rect 32253 1520 32288 1521
rect 32047 1480 32073 1515
rect 32349 1480 32381 2289
rect 32793 2222 32822 2907
rect 33753 2888 34039 2889
rect 33238 2880 34041 2888
rect 33238 2863 33249 2880
rect 33239 2858 33249 2863
rect 33273 2863 34041 2880
rect 33273 2858 33278 2863
rect 33239 2845 33278 2858
rect 33783 2797 33818 2798
rect 33762 2790 33818 2797
rect 33762 2770 33791 2790
rect 33811 2770 33818 2790
rect 33762 2765 33818 2770
rect 34002 2788 34041 2863
rect 34002 2768 34013 2788
rect 34033 2768 34041 2788
rect 32846 2629 33228 2634
rect 32846 2610 32854 2629
rect 32875 2610 33228 2629
rect 32846 2602 33228 2610
rect 33199 2572 33228 2602
rect 32986 2569 33021 2570
rect 32965 2562 33021 2569
rect 32965 2542 32994 2562
rect 33014 2542 33021 2562
rect 32965 2537 33021 2542
rect 33198 2565 33232 2572
rect 33198 2547 33206 2565
rect 33225 2547 33232 2565
rect 33198 2539 33232 2547
rect 33762 2559 33796 2765
rect 34002 2764 34041 2768
rect 33830 2738 34415 2744
rect 33830 2718 33846 2738
rect 33866 2737 34415 2738
rect 33866 2718 34386 2737
rect 33830 2717 34386 2718
rect 34406 2717 34415 2737
rect 33830 2709 34415 2717
rect 33762 2551 33797 2559
rect 32965 2331 32999 2537
rect 33762 2531 33770 2551
rect 33790 2531 33797 2551
rect 33762 2526 33797 2531
rect 33762 2525 33794 2526
rect 33033 2510 33618 2516
rect 33033 2490 33049 2510
rect 33069 2509 33618 2510
rect 33069 2490 33589 2509
rect 33033 2489 33589 2490
rect 33609 2489 33618 2509
rect 33033 2481 33618 2489
rect 33698 2480 33728 2481
rect 33698 2453 34034 2480
rect 33698 2452 33733 2453
rect 32965 2323 33000 2331
rect 32965 2303 32973 2323
rect 32993 2303 33000 2323
rect 32965 2298 33000 2303
rect 32965 2277 32999 2298
rect 33698 2277 33728 2452
rect 33784 2385 33819 2386
rect 32965 2251 33728 2277
rect 32966 2250 32999 2251
rect 33698 2249 33728 2251
rect 33763 2378 33819 2385
rect 33763 2358 33792 2378
rect 33812 2358 33819 2378
rect 33763 2353 33819 2358
rect 33998 2380 34033 2453
rect 33998 2360 34005 2380
rect 34025 2360 34033 2380
rect 33998 2353 34033 2360
rect 32793 2194 33132 2222
rect 32887 2159 32922 2160
rect 32866 2152 32922 2159
rect 32866 2132 32895 2152
rect 32915 2132 32922 2152
rect 32866 2127 32922 2132
rect 33101 2152 33132 2194
rect 33101 2133 33106 2152
rect 33127 2133 33132 2152
rect 33101 2127 33132 2133
rect 33763 2147 33797 2353
rect 33831 2326 34416 2332
rect 33831 2306 33847 2326
rect 33867 2325 34416 2326
rect 33867 2306 34387 2325
rect 33831 2305 34387 2306
rect 34407 2305 34416 2325
rect 33831 2297 34416 2305
rect 33763 2139 33798 2147
rect 32866 1921 32900 2127
rect 33763 2119 33771 2139
rect 33791 2119 33798 2139
rect 33763 2114 33798 2119
rect 33763 2113 33795 2114
rect 32934 2100 33519 2106
rect 32934 2080 32950 2100
rect 32970 2099 33519 2100
rect 32970 2080 33490 2099
rect 32934 2079 33490 2080
rect 33510 2079 33519 2099
rect 32934 2071 33519 2079
rect 32866 1913 32901 1921
rect 32866 1893 32874 1913
rect 32894 1905 32901 1913
rect 32894 1893 32905 1905
rect 32866 1656 32905 1893
rect 33736 1870 34022 1871
rect 33221 1862 34024 1870
rect 33221 1845 33232 1862
rect 33222 1840 33232 1845
rect 33256 1845 34024 1862
rect 33256 1840 33261 1845
rect 33222 1827 33261 1840
rect 33766 1779 33801 1780
rect 33745 1772 33801 1779
rect 33745 1752 33774 1772
rect 33794 1752 33801 1772
rect 33745 1747 33801 1752
rect 33985 1770 34024 1845
rect 33985 1750 33996 1770
rect 34016 1750 34024 1770
rect 32866 1622 33212 1656
rect 33183 1554 33212 1622
rect 32969 1551 33004 1552
rect 32047 1452 32381 1480
rect 32948 1544 33004 1551
rect 32948 1524 32977 1544
rect 32997 1524 33004 1544
rect 32948 1519 33004 1524
rect 33181 1545 33216 1554
rect 33181 1526 33190 1545
rect 33211 1526 33216 1545
rect 33181 1520 33216 1526
rect 33745 1541 33779 1747
rect 33985 1746 34024 1750
rect 33813 1720 34398 1726
rect 33813 1700 33829 1720
rect 33849 1719 34398 1720
rect 33849 1700 34369 1719
rect 33813 1699 34369 1700
rect 34389 1699 34398 1719
rect 33813 1691 34398 1699
rect 33745 1533 33780 1541
rect 27014 1108 27049 1116
rect 25005 1096 25040 1104
rect 23413 1085 23448 1086
rect 23206 1053 23235 1083
rect 25005 1076 25013 1096
rect 25033 1076 25040 1096
rect 25005 1071 25040 1076
rect 25005 1070 25037 1071
rect 23206 1045 23588 1053
rect 23206 1026 23559 1045
rect 23580 1026 23588 1045
rect 23206 1021 23588 1026
rect 26396 950 26981 958
rect 26396 930 26405 950
rect 26425 949 26981 950
rect 26425 930 26945 949
rect 26396 929 26945 930
rect 26965 929 26981 949
rect 26396 923 26981 929
rect 22393 867 22401 887
rect 22421 867 22432 887
rect 18252 844 18287 845
rect 19487 797 19538 828
rect 18792 784 18831 797
rect 18792 779 18797 784
rect 18029 762 18797 779
rect 18821 779 18831 784
rect 18821 762 18832 779
rect 18029 754 18832 762
rect 19487 771 19504 797
rect 19532 771 19538 797
rect 18031 753 18317 754
rect 19487 748 19538 771
rect 19567 803 19613 834
rect 21411 832 21454 840
rect 19567 772 19581 803
rect 19609 772 19613 803
rect 19567 765 19613 772
rect 21405 825 21460 832
rect 21405 800 21418 825
rect 21450 800 21460 825
rect 17139 702 17150 734
rect 17190 702 17194 734
rect 17139 689 17194 702
rect 17869 737 17930 746
rect 17869 710 17877 737
rect 17913 731 17930 737
rect 17971 731 18046 735
rect 17913 729 18046 731
rect 17913 710 17977 729
rect 17869 693 17977 710
rect 18022 693 18046 729
rect 17869 691 18046 693
rect 17971 661 18046 691
rect 19500 556 19531 748
rect 19486 535 19532 556
rect 19486 514 19493 535
rect 19514 514 19532 535
rect 19486 510 19532 514
rect 19486 507 19521 510
rect 15303 447 15309 467
rect 15329 447 15337 467
rect 15303 441 15337 447
rect 17556 432 17587 437
rect 17893 435 17958 437
rect 14980 298 14996 322
rect 15019 298 15031 322
rect 14980 289 15031 298
rect 15199 322 15255 327
rect 15199 302 15206 322
rect 15226 302 15255 322
rect 15199 295 15255 302
rect 16758 412 17592 432
rect 17622 427 17958 435
rect 15199 294 15234 295
rect 14984 223 15027 289
rect 13324 207 13359 208
rect 14487 195 15027 223
rect 14490 193 15027 195
rect 14984 191 15027 193
rect 16758 130 16784 412
rect 17542 410 17588 412
rect 17542 389 17549 410
rect 17570 389 17588 410
rect 17622 402 17903 427
rect 17542 385 17588 389
rect 17542 382 17577 385
rect 16924 224 17509 232
rect 16924 204 16933 224
rect 16953 223 17509 224
rect 16953 204 17473 223
rect 16924 203 17473 204
rect 17493 203 17509 223
rect 16924 197 17509 203
rect 17543 176 17577 382
rect 17624 316 17667 402
rect 17751 396 17903 402
rect 17893 386 17903 396
rect 17943 386 17958 427
rect 17893 372 17958 386
rect 18868 349 19453 357
rect 18868 329 18877 349
rect 18897 348 19453 349
rect 18897 329 19417 348
rect 18868 328 19417 329
rect 19437 328 19453 348
rect 18868 322 19453 328
rect 17624 296 17631 316
rect 17651 296 17667 316
rect 19487 301 19521 507
rect 19569 441 19603 765
rect 21405 708 21460 800
rect 22393 792 22432 867
rect 22616 885 22672 890
rect 22616 865 22623 885
rect 22643 865 22672 885
rect 22616 858 22672 865
rect 26770 899 26809 903
rect 27015 902 27049 1108
rect 27579 1120 27613 1128
rect 27579 1102 27586 1120
rect 27605 1102 27613 1120
rect 27579 1095 27613 1102
rect 27790 1125 27846 1130
rect 27790 1105 27797 1125
rect 27817 1105 27846 1125
rect 27790 1098 27846 1105
rect 29382 1116 29416 1322
rect 31142 1320 31177 1327
rect 29450 1295 30035 1301
rect 29450 1275 29466 1295
rect 29486 1294 30035 1295
rect 29486 1275 30006 1294
rect 29450 1274 30006 1275
rect 30026 1274 30035 1294
rect 29450 1266 30035 1274
rect 31142 1300 31150 1320
rect 31170 1300 31177 1320
rect 31142 1227 31177 1300
rect 31356 1322 31412 1327
rect 31356 1302 31363 1322
rect 31383 1302 31412 1322
rect 31356 1295 31412 1302
rect 31447 1429 31477 1431
rect 32176 1429 32209 1430
rect 31447 1403 32210 1429
rect 31356 1294 31391 1295
rect 31447 1228 31477 1403
rect 32176 1382 32210 1403
rect 32175 1377 32210 1382
rect 32175 1357 32182 1377
rect 32202 1357 32210 1377
rect 32175 1349 32210 1357
rect 31442 1227 31477 1228
rect 31141 1200 31477 1227
rect 31447 1199 31477 1200
rect 31557 1191 32142 1199
rect 31557 1171 31566 1191
rect 31586 1190 32142 1191
rect 31586 1171 32106 1190
rect 31557 1170 32106 1171
rect 32126 1170 32142 1190
rect 31557 1164 32142 1170
rect 31381 1154 31413 1155
rect 31378 1149 31413 1154
rect 31378 1129 31385 1149
rect 31405 1129 31413 1149
rect 32176 1143 32210 1349
rect 32948 1313 32982 1519
rect 33745 1513 33753 1533
rect 33773 1513 33780 1533
rect 33745 1508 33780 1513
rect 33745 1507 33777 1508
rect 33016 1492 33601 1498
rect 33016 1472 33032 1492
rect 33052 1491 33601 1492
rect 33052 1472 33572 1491
rect 33016 1471 33572 1472
rect 33592 1471 33601 1491
rect 33016 1463 33601 1471
rect 33681 1462 33711 1463
rect 33681 1435 34017 1462
rect 33681 1434 33716 1435
rect 32948 1305 32983 1313
rect 32948 1285 32956 1305
rect 32976 1285 32983 1305
rect 32948 1280 32983 1285
rect 32948 1259 32982 1280
rect 33681 1259 33711 1434
rect 33767 1367 33802 1368
rect 32948 1233 33711 1259
rect 32949 1232 32982 1233
rect 33681 1231 33711 1233
rect 33746 1360 33802 1367
rect 33746 1340 33775 1360
rect 33795 1340 33802 1360
rect 33746 1335 33802 1340
rect 33981 1362 34016 1435
rect 33981 1342 33988 1362
rect 34008 1342 34016 1362
rect 33981 1335 34016 1342
rect 31378 1121 31413 1129
rect 29382 1108 29417 1116
rect 27790 1097 27825 1098
rect 27583 1065 27612 1095
rect 29382 1088 29390 1108
rect 29410 1088 29417 1108
rect 29382 1083 29417 1088
rect 29382 1082 29414 1083
rect 27583 1057 27965 1065
rect 27583 1038 27936 1057
rect 27957 1038 27965 1057
rect 27583 1033 27965 1038
rect 30760 963 31345 971
rect 30760 943 30769 963
rect 30789 962 31345 963
rect 30789 943 31309 962
rect 30760 942 31309 943
rect 31329 942 31345 962
rect 30760 936 31345 942
rect 26770 879 26778 899
rect 26798 879 26809 899
rect 22616 857 22651 858
rect 23851 810 23902 841
rect 23156 797 23195 810
rect 23156 792 23161 797
rect 22393 775 23161 792
rect 23185 792 23195 797
rect 23185 775 23196 792
rect 22393 767 23196 775
rect 23851 784 23868 810
rect 23896 784 23902 810
rect 22395 766 22681 767
rect 23851 761 23902 784
rect 23931 816 23977 847
rect 25775 845 25818 853
rect 23931 785 23945 816
rect 23973 785 23977 816
rect 23931 778 23977 785
rect 25769 838 25824 845
rect 25769 813 25782 838
rect 25814 813 25824 838
rect 21405 676 21416 708
rect 21456 676 21460 708
rect 22233 750 22294 759
rect 22233 723 22241 750
rect 22277 744 22294 750
rect 22335 744 22410 748
rect 22277 742 22410 744
rect 22277 723 22341 742
rect 22233 706 22341 723
rect 22386 706 22410 742
rect 22233 704 22410 706
rect 21405 663 21460 676
rect 22335 674 22410 704
rect 23864 569 23895 761
rect 23850 548 23896 569
rect 23850 527 23857 548
rect 23878 527 23896 548
rect 23850 523 23896 527
rect 23850 520 23885 523
rect 21989 483 22020 488
rect 19569 421 19575 441
rect 19595 421 19603 441
rect 19569 415 19603 421
rect 21191 463 22025 483
rect 17624 285 17667 296
rect 19248 295 19291 299
rect 19248 271 19259 295
rect 19282 271 19291 295
rect 19248 267 19291 271
rect 19465 296 19521 301
rect 19465 276 19472 296
rect 19492 276 19521 296
rect 19465 269 19521 276
rect 19465 268 19500 269
rect 19255 203 19286 267
rect 21191 203 21217 463
rect 21975 461 22021 463
rect 21975 440 21982 461
rect 22003 440 22021 461
rect 22055 453 23148 486
rect 21975 436 22021 440
rect 21975 433 22010 436
rect 21357 275 21942 283
rect 21357 255 21366 275
rect 21386 274 21942 275
rect 21386 255 21906 274
rect 21357 254 21906 255
rect 21926 254 21942 274
rect 21357 248 21942 254
rect 21976 227 22010 433
rect 22057 367 22100 453
rect 22057 347 22064 367
rect 22084 347 22100 367
rect 22057 336 22100 347
rect 21954 222 22010 227
rect 21744 217 21776 222
rect 19255 180 21218 203
rect 19263 178 21218 180
rect 21744 196 21751 217
rect 21768 196 21776 217
rect 21744 189 21776 196
rect 21954 202 21961 222
rect 21981 202 22010 222
rect 21954 195 22010 202
rect 23117 210 23146 453
rect 23232 362 23817 370
rect 23232 342 23241 362
rect 23261 361 23817 362
rect 23261 342 23781 361
rect 23232 341 23781 342
rect 23801 341 23817 361
rect 23232 335 23817 341
rect 23614 315 23657 317
rect 23610 309 23661 315
rect 23851 314 23885 520
rect 23933 454 23967 778
rect 25769 721 25824 813
rect 26770 804 26809 879
rect 26993 897 27049 902
rect 26993 877 27000 897
rect 27020 877 27049 897
rect 26993 870 27049 877
rect 31134 912 31173 916
rect 31379 915 31413 1121
rect 31943 1133 31977 1141
rect 31943 1115 31950 1133
rect 31969 1115 31977 1133
rect 31943 1108 31977 1115
rect 32154 1138 32210 1143
rect 32154 1118 32161 1138
rect 32181 1118 32210 1138
rect 32154 1111 32210 1118
rect 33746 1129 33780 1335
rect 33814 1308 34399 1314
rect 33814 1288 33830 1308
rect 33850 1307 34399 1308
rect 33850 1288 34370 1307
rect 33814 1287 34370 1288
rect 34390 1287 34399 1307
rect 33814 1279 34399 1287
rect 33746 1121 33781 1129
rect 32154 1110 32189 1111
rect 31947 1078 31976 1108
rect 33746 1101 33754 1121
rect 33774 1101 33781 1121
rect 33746 1096 33781 1101
rect 33746 1095 33778 1096
rect 31947 1070 32329 1078
rect 31947 1051 32300 1070
rect 32321 1051 32329 1070
rect 31947 1046 32329 1051
rect 31134 892 31142 912
rect 31162 892 31173 912
rect 26993 869 27028 870
rect 28228 822 28279 853
rect 27533 809 27572 822
rect 27533 804 27538 809
rect 26770 787 27538 804
rect 27562 804 27572 809
rect 27562 787 27573 804
rect 26770 779 27573 787
rect 28228 796 28245 822
rect 28273 796 28279 822
rect 26772 778 27058 779
rect 28228 773 28279 796
rect 28308 828 28354 859
rect 30152 857 30195 865
rect 28308 797 28322 828
rect 28350 797 28354 828
rect 28308 790 28354 797
rect 30146 850 30201 857
rect 30146 825 30159 850
rect 30191 825 30201 850
rect 25769 689 25780 721
rect 25820 689 25824 721
rect 26610 762 26671 771
rect 26610 735 26618 762
rect 26654 756 26671 762
rect 26712 756 26787 760
rect 26654 754 26787 756
rect 26654 735 26718 754
rect 26610 718 26718 735
rect 26763 718 26787 754
rect 26610 716 26787 718
rect 25769 676 25824 689
rect 26712 686 26787 716
rect 28241 581 28272 773
rect 28227 560 28273 581
rect 28227 539 28234 560
rect 28255 539 28273 560
rect 28227 535 28273 539
rect 28227 532 28262 535
rect 26437 507 26468 512
rect 23933 434 23939 454
rect 23959 434 23967 454
rect 23933 428 23967 434
rect 25639 487 26473 507
rect 23610 285 23626 309
rect 23649 285 23661 309
rect 23610 276 23661 285
rect 23829 309 23885 314
rect 23829 289 23836 309
rect 23856 289 23885 309
rect 23829 282 23885 289
rect 23829 281 23864 282
rect 23614 210 23657 276
rect 21954 194 21989 195
rect 17521 171 17577 176
rect 17521 151 17528 171
rect 17548 151 17577 171
rect 17521 144 17577 151
rect 17521 143 17556 144
rect 16735 121 16788 130
rect 16735 95 16747 121
rect 16778 95 16788 121
rect 21744 129 21772 189
rect 23117 182 23657 210
rect 23120 180 23657 182
rect 23614 178 23657 180
rect 25639 129 25665 487
rect 26423 485 26469 487
rect 26423 464 26430 485
rect 26451 464 26469 485
rect 26503 477 27432 510
rect 26423 460 26469 464
rect 26423 457 26458 460
rect 25805 299 26390 307
rect 25805 279 25814 299
rect 25834 298 26390 299
rect 25834 279 26354 298
rect 25805 278 26354 279
rect 26374 278 26390 298
rect 25805 272 26390 278
rect 26187 242 26228 255
rect 26424 251 26458 457
rect 26505 391 26548 477
rect 26632 471 27432 477
rect 26505 371 26512 391
rect 26532 371 26548 391
rect 26505 360 26548 371
rect 26187 221 26195 242
rect 26218 221 26228 242
rect 21744 95 25670 129
rect 16735 85 16788 95
rect 26187 77 26228 221
rect 26402 246 26458 251
rect 26402 226 26409 246
rect 26429 226 26458 246
rect 26402 219 26458 226
rect 26402 218 26437 219
rect 10022 2 13157 46
rect 26185 60 26248 77
rect 26185 34 26197 60
rect 26226 34 26248 60
rect 26185 22 26248 34
rect 27393 58 27432 471
rect 27609 374 28194 382
rect 27609 354 27618 374
rect 27638 373 28194 374
rect 27638 354 28158 373
rect 27609 353 28158 354
rect 28178 353 28194 373
rect 27609 347 28194 353
rect 28228 326 28262 532
rect 28310 466 28344 790
rect 30146 733 30201 825
rect 31134 817 31173 892
rect 31357 910 31413 915
rect 31357 890 31364 910
rect 31384 890 31413 910
rect 31357 883 31413 890
rect 31357 882 31392 883
rect 32592 835 32643 866
rect 31897 822 31936 835
rect 31897 817 31902 822
rect 31134 800 31902 817
rect 31926 817 31936 822
rect 31926 800 31937 817
rect 31134 792 31937 800
rect 32592 809 32609 835
rect 32637 809 32643 835
rect 31136 791 31422 792
rect 32592 786 32643 809
rect 32672 841 32718 872
rect 34516 870 34559 878
rect 32672 810 32686 841
rect 32714 810 32718 841
rect 32672 803 32718 810
rect 34510 863 34565 870
rect 34510 838 34523 863
rect 34555 838 34565 863
rect 30146 701 30157 733
rect 30197 701 30201 733
rect 30974 775 31035 784
rect 30974 748 30982 775
rect 31018 769 31035 775
rect 31076 769 31151 773
rect 31018 767 31151 769
rect 31018 748 31082 767
rect 30974 731 31082 748
rect 31127 731 31151 767
rect 30974 729 31151 731
rect 30146 688 30201 701
rect 31076 699 31151 729
rect 32605 594 32636 786
rect 32591 573 32637 594
rect 32591 552 32598 573
rect 32619 552 32637 573
rect 32591 548 32637 552
rect 32591 545 32626 548
rect 30730 508 30761 513
rect 28310 446 28316 466
rect 28336 446 28344 466
rect 28310 440 28344 446
rect 29932 488 30766 508
rect 27989 320 28032 324
rect 27989 296 28000 320
rect 28023 296 28032 320
rect 27989 292 28032 296
rect 28206 321 28262 326
rect 28206 301 28213 321
rect 28233 301 28262 321
rect 28206 294 28262 301
rect 28206 293 28241 294
rect 27996 228 28027 292
rect 29932 228 29958 488
rect 30716 486 30762 488
rect 30716 465 30723 486
rect 30744 465 30762 486
rect 30796 478 31889 511
rect 30716 461 30762 465
rect 30716 458 30751 461
rect 30098 300 30683 308
rect 30098 280 30107 300
rect 30127 299 30683 300
rect 30127 280 30647 299
rect 30098 279 30647 280
rect 30667 279 30683 299
rect 30098 273 30683 279
rect 30717 252 30751 458
rect 30798 392 30841 478
rect 30798 372 30805 392
rect 30825 372 30841 392
rect 30798 361 30841 372
rect 30476 245 30528 251
rect 27996 205 29959 228
rect 28004 203 29959 205
rect 30476 223 30488 245
rect 30509 223 30528 245
rect 30476 58 30528 223
rect 30695 247 30751 252
rect 30695 227 30702 247
rect 30722 227 30751 247
rect 30695 220 30751 227
rect 31858 235 31887 478
rect 31973 387 32558 395
rect 31973 367 31982 387
rect 32002 386 32558 387
rect 32002 367 32522 386
rect 31973 366 32522 367
rect 32542 366 32558 386
rect 31973 360 32558 366
rect 32355 340 32398 342
rect 32351 334 32402 340
rect 32592 339 32626 545
rect 32674 479 32708 803
rect 34510 746 34565 838
rect 34510 714 34521 746
rect 34561 714 34565 746
rect 34510 701 34565 714
rect 32674 459 32680 479
rect 32700 459 32708 479
rect 32674 453 32708 459
rect 32351 310 32367 334
rect 32390 310 32402 334
rect 32351 301 32402 310
rect 32570 334 32626 339
rect 32570 314 32577 334
rect 32597 314 32626 334
rect 32570 307 32626 314
rect 32570 306 32605 307
rect 32355 235 32398 301
rect 30695 219 30730 220
rect 31858 207 32398 235
rect 31861 205 32398 207
rect 32355 203 32398 205
rect 27393 17 30528 58
rect 10022 0 13102 2
<< via1 >>
rect 2200 5207 2227 5234
rect 2118 4388 2149 4414
rect 6564 5220 6591 5247
rect 6482 4401 6513 4427
rect 10941 5232 10968 5259
rect 10859 4413 10890 4439
rect 15305 5245 15332 5272
rect 15223 4426 15254 4452
rect 19571 5219 19598 5246
rect 19489 4400 19520 4426
rect 23935 5232 23962 5259
rect 23853 4413 23884 4439
rect 2133 759 2161 785
rect 2210 760 2238 791
rect 606 681 651 717
rect 6497 772 6525 798
rect 6574 773 6602 804
rect 4045 664 4085 696
rect 4970 694 5015 730
rect 28312 5244 28339 5271
rect 28230 4425 28261 4451
rect 32676 5257 32703 5284
rect 32594 4438 32625 4464
rect 10874 784 10902 810
rect 10951 785 10979 816
rect 8409 677 8449 709
rect 9347 706 9392 742
rect 8824 97 8853 128
rect 15238 797 15266 823
rect 15315 798 15343 829
rect 12786 689 12826 721
rect 13711 719 13756 755
rect 19504 771 19532 797
rect 19581 772 19609 803
rect 17150 702 17190 734
rect 17977 693 18022 729
rect 17903 386 17943 427
rect 23868 784 23896 810
rect 23945 785 23973 816
rect 21416 676 21456 708
rect 22341 706 22386 742
rect 28245 796 28273 822
rect 28322 797 28350 828
rect 25780 689 25820 721
rect 26718 718 26763 754
rect 16747 95 16778 121
rect 26197 34 26226 60
rect 32609 809 32637 835
rect 32686 810 32714 841
rect 30157 701 30197 733
rect 31082 731 31127 767
rect 34521 714 34561 746
<< metal2 >>
rect 32671 5284 32708 5288
rect 15300 5272 15337 5276
rect 10936 5259 10973 5263
rect 6559 5247 6596 5251
rect 2195 5234 2232 5238
rect 2195 5207 2200 5234
rect 2227 5207 2232 5234
rect 6559 5220 6564 5247
rect 6591 5220 6596 5247
rect 10936 5232 10941 5259
rect 10968 5232 10973 5259
rect 15300 5245 15305 5272
rect 15332 5245 15337 5272
rect 28307 5271 28344 5275
rect 23930 5259 23967 5263
rect 15300 5235 15337 5245
rect 19566 5246 19603 5250
rect 10936 5222 10973 5232
rect 6559 5210 6596 5220
rect 2195 5197 2232 5207
rect 2110 4414 2158 4432
rect 2110 4388 2118 4414
rect 2149 4388 2158 4414
rect 2110 4356 2158 4388
rect 2118 810 2158 4356
rect 2199 2460 2225 5197
rect 6474 4427 6522 4445
rect 6474 4401 6482 4427
rect 6513 4401 6522 4427
rect 6474 4369 6522 4401
rect 2197 822 2225 2460
rect 6482 823 6522 4369
rect 6563 2473 6589 5210
rect 10851 4439 10899 4457
rect 10851 4413 10859 4439
rect 10890 4413 10899 4439
rect 10851 4381 10899 4413
rect 6561 835 6589 2473
rect 10859 835 10899 4381
rect 10940 2485 10966 5222
rect 15215 4452 15263 4470
rect 15215 4426 15223 4452
rect 15254 4426 15263 4452
rect 15215 4394 15263 4426
rect 10938 847 10966 2485
rect 15223 848 15263 4394
rect 15304 2498 15330 5235
rect 19566 5219 19571 5246
rect 19598 5219 19603 5246
rect 23930 5232 23935 5259
rect 23962 5232 23967 5259
rect 28307 5244 28312 5271
rect 28339 5244 28344 5271
rect 32671 5257 32676 5284
rect 32703 5257 32708 5284
rect 32671 5247 32708 5257
rect 28307 5234 28344 5244
rect 23930 5222 23967 5232
rect 19566 5209 19603 5219
rect 19481 4426 19529 4444
rect 19481 4400 19489 4426
rect 19520 4400 19529 4426
rect 19481 4368 19529 4400
rect 15302 860 15330 2498
rect 2118 785 2164 810
rect 2118 759 2133 785
rect 2161 759 2164 785
rect 2118 740 2164 759
rect 2196 791 2242 822
rect 2196 760 2210 791
rect 2238 760 2242 791
rect 2196 753 2242 760
rect 6482 798 6528 823
rect 6482 772 6497 798
rect 6525 772 6528 798
rect 6482 753 6528 772
rect 6560 804 6606 835
rect 6560 773 6574 804
rect 6602 773 6606 804
rect 6560 766 6606 773
rect 10859 810 10905 835
rect 10859 784 10874 810
rect 10902 784 10905 810
rect 10859 765 10905 784
rect 10937 816 10983 847
rect 10937 785 10951 816
rect 10979 785 10983 816
rect 10937 778 10983 785
rect 15223 823 15269 848
rect 15223 797 15238 823
rect 15266 797 15269 823
rect 15223 778 15269 797
rect 15301 829 15347 860
rect 15301 798 15315 829
rect 15343 798 15347 829
rect 15301 791 15347 798
rect 19489 822 19529 4368
rect 19570 2472 19596 5209
rect 23845 4439 23893 4457
rect 23845 4413 23853 4439
rect 23884 4413 23893 4439
rect 23845 4381 23893 4413
rect 19568 834 19596 2472
rect 23853 835 23893 4381
rect 23934 2485 23960 5222
rect 28222 4451 28270 4469
rect 28222 4425 28230 4451
rect 28261 4425 28270 4451
rect 28222 4393 28270 4425
rect 23932 847 23960 2485
rect 28230 847 28270 4393
rect 28311 2497 28337 5234
rect 32586 4464 32634 4482
rect 32586 4438 32594 4464
rect 32625 4438 32634 4464
rect 32586 4406 32634 4438
rect 28309 859 28337 2497
rect 32594 860 32634 4406
rect 32675 2510 32701 5247
rect 32673 872 32701 2510
rect 19489 797 19535 822
rect 15227 774 15269 778
rect 19489 771 19504 797
rect 19532 771 19535 797
rect 10863 761 10905 765
rect 13697 755 13772 767
rect 6486 749 6528 753
rect 9333 742 9408 754
rect 2122 736 2164 740
rect 4956 730 5031 742
rect 592 717 667 729
rect 592 681 606 717
rect 651 704 667 717
rect 2109 704 2203 709
rect 651 696 4089 704
rect 651 681 4045 696
rect 592 664 4045 681
rect 4085 664 4089 696
rect 4956 694 4970 730
rect 5015 717 5031 730
rect 6473 717 6567 722
rect 5015 709 8453 717
rect 5015 694 8409 709
rect 4956 677 8409 694
rect 8449 677 8453 709
rect 9333 706 9347 742
rect 9392 729 9408 742
rect 10850 729 10944 734
rect 9392 721 12830 729
rect 9392 706 12786 721
rect 9333 689 12786 706
rect 12826 689 12830 721
rect 13697 719 13711 755
rect 13756 742 13772 755
rect 19489 752 19535 771
rect 19567 803 19613 834
rect 19567 772 19581 803
rect 19609 772 19613 803
rect 19567 765 19613 772
rect 23853 810 23899 835
rect 23853 784 23868 810
rect 23896 784 23899 810
rect 23853 765 23899 784
rect 23931 816 23977 847
rect 23931 785 23945 816
rect 23973 785 23977 816
rect 23931 778 23977 785
rect 28230 822 28276 847
rect 28230 796 28245 822
rect 28273 796 28276 822
rect 28230 777 28276 796
rect 28308 828 28354 859
rect 28308 797 28322 828
rect 28350 797 28354 828
rect 28308 790 28354 797
rect 32594 835 32640 860
rect 32594 809 32609 835
rect 32637 809 32640 835
rect 32594 790 32640 809
rect 32672 841 32718 872
rect 32672 810 32686 841
rect 32714 810 32718 841
rect 32672 803 32718 810
rect 32598 786 32640 790
rect 28234 773 28276 777
rect 31068 767 31143 779
rect 23857 761 23899 765
rect 26704 754 26779 766
rect 19493 748 19535 752
rect 15214 742 15308 747
rect 22327 742 22402 754
rect 13756 734 17194 742
rect 13756 719 17150 734
rect 13697 702 17150 719
rect 17190 702 17194 734
rect 13697 693 17194 702
rect 17963 729 18038 741
rect 17963 693 17977 729
rect 18022 716 18038 729
rect 19480 716 19574 721
rect 18022 708 21460 716
rect 18022 693 21416 708
rect 15214 690 15308 693
rect 9333 680 12830 689
rect 10850 677 10944 680
rect 4956 668 8453 677
rect 17963 676 21416 693
rect 21456 676 21460 708
rect 22327 706 22341 742
rect 22386 729 22402 742
rect 23844 729 23938 734
rect 22386 721 25824 729
rect 22386 706 25780 721
rect 22327 689 25780 706
rect 25820 689 25824 721
rect 26704 718 26718 754
rect 26763 741 26779 754
rect 28221 741 28315 746
rect 26763 733 30201 741
rect 26763 718 30157 733
rect 26704 701 30157 718
rect 30197 701 30201 733
rect 31068 731 31082 767
rect 31127 754 31143 767
rect 32585 754 32679 759
rect 31127 746 34565 754
rect 31127 731 34521 746
rect 31068 714 34521 731
rect 34561 714 34565 746
rect 31068 705 34565 714
rect 32585 702 32679 705
rect 26704 692 30201 701
rect 28221 689 28315 692
rect 22327 680 25824 689
rect 23844 677 23938 680
rect 6473 665 6567 668
rect 17963 667 21460 676
rect 19480 664 19574 667
rect 592 655 4089 664
rect 2109 652 2203 655
rect 17893 427 17957 434
rect 17893 386 17903 427
rect 17943 386 17957 427
rect 8817 130 8868 139
rect 8815 128 8868 130
rect 8815 97 8824 128
rect 8853 124 8868 128
rect 8853 121 16788 124
rect 8853 97 16747 121
rect 8815 95 16747 97
rect 16778 95 16788 121
rect 8815 93 16788 95
rect 8817 86 16788 93
rect 8817 85 8868 86
rect 17893 60 17957 386
rect 26185 60 26248 77
rect 17890 34 26197 60
rect 26226 34 26248 60
rect 17890 28 26248 34
rect 26185 22 26248 28
<< labels >>
rlabel locali 3939 243 3962 259 1 d6
rlabel locali 4003 433 4032 439 1 vdd
rlabel locali 4000 134 4029 140 1 gnd
rlabel space 4106 152 4135 161 1 gnd
rlabel nwell 4138 410 4161 413 1 vdd
rlabel locali 5820 333 5835 346 1 d5
rlabel locali 5878 520 5907 526 1 vdd
rlabel locali 5875 221 5904 227 1 gnd
rlabel space 5981 239 6010 248 1 gnd
rlabel nwell 6013 497 6036 500 1 vdd
rlabel locali 8302 1253 8324 1268 5 d0
rlabel locali 8241 1074 8270 1080 5 vdd
rlabel locali 8244 1373 8273 1379 5 gnd
rlabel space 8138 1352 8167 1361 5 gnd
rlabel nwell 8112 1100 8135 1103 5 vdd
rlabel locali 8301 1665 8323 1680 5 d0
rlabel locali 8240 1486 8269 1492 5 vdd
rlabel locali 8243 1785 8272 1791 5 gnd
rlabel space 8137 1764 8166 1773 5 gnd
rlabel nwell 8111 1512 8134 1515 5 vdd
rlabel locali 8319 2271 8341 2286 5 d0
rlabel locali 8258 2092 8287 2098 5 vdd
rlabel locali 8261 2391 8290 2397 5 gnd
rlabel space 8155 2370 8184 2379 5 gnd
rlabel nwell 8129 2118 8152 2121 5 vdd
rlabel locali 8318 2683 8340 2698 5 d0
rlabel locali 8257 2504 8286 2510 5 vdd
rlabel locali 8260 2803 8289 2809 5 gnd
rlabel space 8154 2782 8183 2791 5 gnd
rlabel nwell 8128 2530 8151 2533 5 vdd
rlabel locali 7443 1258 7472 1264 5 vdd
rlabel locali 7446 1557 7475 1563 5 gnd
rlabel space 7340 1536 7369 1545 5 gnd
rlabel nwell 7314 1284 7337 1287 5 vdd
rlabel locali 7510 1439 7532 1456 5 d1
rlabel locali 7460 2276 7489 2282 5 vdd
rlabel locali 7463 2575 7492 2581 5 gnd
rlabel space 7357 2554 7386 2563 5 gnd
rlabel nwell 7331 2302 7354 2305 5 vdd
rlabel locali 7527 2457 7549 2474 5 d1
rlabel locali 7361 1866 7390 1872 5 vdd
rlabel locali 7364 2165 7393 2171 5 gnd
rlabel space 7258 2144 7287 2153 5 gnd
rlabel nwell 7232 1892 7255 1895 5 vdd
rlabel locali 7428 2040 7448 2064 5 d2
rlabel locali 8339 3289 8361 3304 5 d0
rlabel locali 8278 3110 8307 3116 5 vdd
rlabel locali 8281 3409 8310 3415 5 gnd
rlabel space 8175 3388 8204 3397 5 gnd
rlabel nwell 8149 3136 8172 3139 5 vdd
rlabel locali 8338 3701 8360 3716 5 d0
rlabel locali 8277 3522 8306 3528 5 vdd
rlabel locali 8280 3821 8309 3827 5 gnd
rlabel space 8174 3800 8203 3809 5 gnd
rlabel nwell 8148 3548 8171 3551 5 vdd
rlabel locali 8356 4307 8378 4322 5 d0
rlabel locali 8295 4128 8324 4134 5 vdd
rlabel locali 8298 4427 8327 4433 5 gnd
rlabel space 8192 4406 8221 4415 5 gnd
rlabel nwell 8166 4154 8189 4157 5 vdd
rlabel locali 8355 4719 8377 4734 5 d0
rlabel locali 8294 4540 8323 4546 5 vdd
rlabel locali 8297 4839 8326 4845 5 gnd
rlabel space 8191 4818 8220 4827 5 gnd
rlabel nwell 8165 4566 8188 4569 5 vdd
rlabel locali 7480 3294 7509 3300 5 vdd
rlabel locali 7483 3593 7512 3599 5 gnd
rlabel space 7377 3572 7406 3581 5 gnd
rlabel nwell 7351 3320 7374 3323 5 vdd
rlabel locali 7547 3475 7569 3492 5 d1
rlabel locali 7497 4312 7526 4318 5 vdd
rlabel locali 7500 4611 7529 4617 5 gnd
rlabel space 7394 4590 7423 4599 5 gnd
rlabel nwell 7368 4338 7391 4341 5 vdd
rlabel locali 7564 4493 7586 4510 5 d1
rlabel locali 7398 3902 7427 3908 5 vdd
rlabel locali 7401 4201 7430 4207 5 gnd
rlabel space 7295 4180 7324 4189 5 gnd
rlabel nwell 7269 3928 7292 3931 5 vdd
rlabel locali 7465 4076 7485 4100 5 d2
rlabel locali 7315 2886 7344 2892 5 vdd
rlabel locali 7318 3185 7347 3191 5 gnd
rlabel space 7212 3164 7241 3173 5 gnd
rlabel nwell 7186 2912 7209 2915 5 vdd
rlabel locali 7380 3065 7400 3078 5 d3
rlabel locali 8375 5325 8397 5340 5 d0
rlabel locali 8314 5146 8343 5152 5 vdd
rlabel locali 8317 5445 8346 5451 5 gnd
rlabel space 8211 5424 8240 5433 5 gnd
rlabel nwell 8185 5172 8208 5175 5 vdd
rlabel locali 8374 5737 8396 5752 5 d0
rlabel locali 8313 5558 8342 5564 5 vdd
rlabel locali 8316 5857 8345 5863 5 gnd
rlabel space 8210 5836 8239 5845 5 gnd
rlabel nwell 8184 5584 8207 5587 5 vdd
rlabel locali 8392 6343 8414 6358 5 d0
rlabel locali 8331 6164 8360 6170 5 vdd
rlabel locali 8334 6463 8363 6469 5 gnd
rlabel space 8228 6442 8257 6451 5 gnd
rlabel nwell 8202 6190 8225 6193 5 vdd
rlabel locali 8391 6755 8413 6770 5 d0
rlabel locali 8330 6576 8359 6582 5 vdd
rlabel locali 8333 6875 8362 6881 5 gnd
rlabel space 8227 6854 8256 6863 5 gnd
rlabel nwell 8201 6602 8224 6605 5 vdd
rlabel locali 7516 5330 7545 5336 5 vdd
rlabel locali 7519 5629 7548 5635 5 gnd
rlabel space 7413 5608 7442 5617 5 gnd
rlabel nwell 7387 5356 7410 5359 5 vdd
rlabel locali 7583 5511 7605 5528 5 d1
rlabel locali 7533 6348 7562 6354 5 vdd
rlabel locali 7536 6647 7565 6653 5 gnd
rlabel space 7430 6626 7459 6635 5 gnd
rlabel nwell 7404 6374 7427 6377 5 vdd
rlabel locali 7600 6529 7622 6546 5 d1
rlabel locali 7434 5938 7463 5944 5 vdd
rlabel locali 7437 6237 7466 6243 5 gnd
rlabel space 7331 6216 7360 6225 5 gnd
rlabel nwell 7305 5964 7328 5967 5 vdd
rlabel locali 7501 6112 7521 6136 5 d2
rlabel locali 8412 7361 8434 7376 5 d0
rlabel locali 8351 7182 8380 7188 5 vdd
rlabel locali 8354 7481 8383 7487 5 gnd
rlabel space 8248 7460 8277 7469 5 gnd
rlabel nwell 8222 7208 8245 7211 5 vdd
rlabel locali 8411 7773 8433 7788 5 d0
rlabel locali 8350 7594 8379 7600 5 vdd
rlabel locali 8353 7893 8382 7899 5 gnd
rlabel space 8247 7872 8276 7881 5 gnd
rlabel nwell 8221 7620 8244 7623 5 vdd
rlabel locali 8429 8379 8451 8394 5 d0
rlabel locali 8368 8200 8397 8206 5 vdd
rlabel locali 8371 8499 8400 8505 5 gnd
rlabel space 8265 8478 8294 8487 5 gnd
rlabel nwell 8239 8226 8262 8229 5 vdd
rlabel locali 8428 8791 8450 8806 5 d0
rlabel locali 8367 8612 8396 8618 5 vdd
rlabel locali 8370 8911 8399 8917 5 gnd
rlabel space 8264 8890 8293 8899 5 gnd
rlabel nwell 8238 8638 8261 8641 5 vdd
rlabel locali 7553 7366 7582 7372 5 vdd
rlabel locali 7556 7665 7585 7671 5 gnd
rlabel space 7450 7644 7479 7653 5 gnd
rlabel nwell 7424 7392 7447 7395 5 vdd
rlabel locali 7620 7547 7642 7564 5 d1
rlabel locali 7570 8384 7599 8390 5 vdd
rlabel locali 7573 8683 7602 8689 5 gnd
rlabel space 7467 8662 7496 8671 5 gnd
rlabel nwell 7441 8410 7464 8413 5 vdd
rlabel locali 7637 8565 7659 8582 5 d1
rlabel locali 7471 7974 7500 7980 5 vdd
rlabel locali 7474 8273 7503 8279 5 gnd
rlabel space 7368 8252 7397 8261 5 gnd
rlabel nwell 7342 8000 7365 8003 5 vdd
rlabel locali 7538 8148 7558 8172 5 d2
rlabel locali 7388 6958 7417 6964 5 vdd
rlabel locali 7391 7257 7420 7263 5 gnd
rlabel space 7285 7236 7314 7245 5 gnd
rlabel nwell 7259 6984 7282 6987 5 vdd
rlabel locali 7453 7137 7473 7150 5 d3
rlabel locali 7212 4924 7241 4930 5 vdd
rlabel locali 7215 5223 7244 5229 5 gnd
rlabel space 7109 5202 7138 5211 5 gnd
rlabel nwell 7083 4950 7106 4953 5 vdd
rlabel locali 7276 5103 7295 5120 5 d4
rlabel locali 5766 4594 5785 4611 1 d4
rlabel nwell 5955 4761 5978 4764 1 vdd
rlabel space 5923 4503 5952 4512 1 gnd
rlabel locali 5817 4485 5846 4491 1 gnd
rlabel locali 5820 4784 5849 4790 1 vdd
rlabel locali 5588 2564 5608 2577 1 d3
rlabel nwell 5779 2727 5802 2730 1 vdd
rlabel space 5747 2469 5776 2478 1 gnd
rlabel locali 5641 2451 5670 2457 1 gnd
rlabel locali 5644 2750 5673 2756 1 vdd
rlabel locali 5503 1542 5523 1566 1 d2
rlabel nwell 5696 1711 5719 1714 1 vdd
rlabel space 5664 1453 5693 1462 1 gnd
rlabel locali 5558 1435 5587 1441 1 gnd
rlabel locali 5561 1734 5590 1740 1 vdd
rlabel locali 5402 1132 5424 1149 1 d1
rlabel nwell 5597 1301 5620 1304 1 vdd
rlabel space 5565 1043 5594 1052 1 gnd
rlabel locali 5459 1025 5488 1031 1 gnd
rlabel locali 5462 1324 5491 1330 1 vdd
rlabel locali 5419 2150 5441 2167 1 d1
rlabel nwell 5614 2319 5637 2322 1 vdd
rlabel space 5582 2061 5611 2070 1 gnd
rlabel locali 5476 2043 5505 2049 1 gnd
rlabel locali 5479 2342 5508 2348 1 vdd
rlabel nwell 4800 1073 4823 1076 1 vdd
rlabel space 4768 815 4797 824 1 gnd
rlabel locali 4662 797 4691 803 1 gnd
rlabel locali 4665 1096 4694 1102 1 vdd
rlabel locali 4611 908 4633 923 1 d0
rlabel nwell 4799 1485 4822 1488 1 vdd
rlabel space 4767 1227 4796 1236 1 gnd
rlabel locali 4661 1209 4690 1215 1 gnd
rlabel locali 4664 1508 4693 1514 1 vdd
rlabel locali 4610 1320 4632 1335 1 d0
rlabel nwell 4817 2091 4840 2094 1 vdd
rlabel space 4785 1833 4814 1842 1 gnd
rlabel locali 4679 1815 4708 1821 1 gnd
rlabel locali 4682 2114 4711 2120 1 vdd
rlabel locali 4628 1926 4650 1941 1 d0
rlabel nwell 4816 2503 4839 2506 1 vdd
rlabel space 4784 2245 4813 2254 1 gnd
rlabel locali 4678 2227 4707 2233 1 gnd
rlabel locali 4681 2526 4710 2532 1 vdd
rlabel locali 4627 2338 4649 2353 1 d0
rlabel locali 5540 3578 5560 3602 1 d2
rlabel nwell 5733 3747 5756 3750 1 vdd
rlabel space 5701 3489 5730 3498 1 gnd
rlabel locali 5595 3471 5624 3477 1 gnd
rlabel locali 5598 3770 5627 3776 1 vdd
rlabel locali 5439 3168 5461 3185 1 d1
rlabel nwell 5634 3337 5657 3340 1 vdd
rlabel space 5602 3079 5631 3088 1 gnd
rlabel locali 5496 3061 5525 3067 1 gnd
rlabel locali 5499 3360 5528 3366 1 vdd
rlabel locali 5456 4186 5478 4203 1 d1
rlabel nwell 5651 4355 5674 4358 1 vdd
rlabel space 5619 4097 5648 4106 1 gnd
rlabel locali 5513 4079 5542 4085 1 gnd
rlabel locali 5516 4378 5545 4384 1 vdd
rlabel nwell 4837 3109 4860 3112 1 vdd
rlabel space 4805 2851 4834 2860 1 gnd
rlabel locali 4699 2833 4728 2839 1 gnd
rlabel locali 4702 3132 4731 3138 1 vdd
rlabel locali 4648 2944 4670 2959 1 d0
rlabel nwell 4836 3521 4859 3524 1 vdd
rlabel space 4804 3263 4833 3272 1 gnd
rlabel locali 4698 3245 4727 3251 1 gnd
rlabel locali 4701 3544 4730 3550 1 vdd
rlabel locali 4647 3356 4669 3371 1 d0
rlabel nwell 4854 4127 4877 4130 1 vdd
rlabel space 4822 3869 4851 3878 1 gnd
rlabel locali 4716 3851 4745 3857 1 gnd
rlabel locali 4719 4150 4748 4156 1 vdd
rlabel locali 4665 3962 4687 3977 1 d0
rlabel nwell 4853 4539 4876 4542 1 vdd
rlabel space 4821 4281 4850 4290 1 gnd
rlabel locali 4715 4263 4744 4269 1 gnd
rlabel locali 4718 4562 4747 4568 1 vdd
rlabel locali 4664 4374 4686 4389 1 d0
rlabel locali 5661 6636 5681 6649 1 d3
rlabel nwell 5852 6799 5875 6802 1 vdd
rlabel space 5820 6541 5849 6550 1 gnd
rlabel locali 5714 6523 5743 6529 1 gnd
rlabel locali 5717 6822 5746 6828 1 vdd
rlabel locali 5576 5614 5596 5638 1 d2
rlabel nwell 5769 5783 5792 5786 1 vdd
rlabel space 5737 5525 5766 5534 1 gnd
rlabel locali 5631 5507 5660 5513 1 gnd
rlabel locali 5634 5806 5663 5812 1 vdd
rlabel locali 5475 5204 5497 5221 1 d1
rlabel nwell 5670 5373 5693 5376 1 vdd
rlabel space 5638 5115 5667 5124 1 gnd
rlabel locali 5532 5097 5561 5103 1 gnd
rlabel locali 5535 5396 5564 5402 1 vdd
rlabel locali 5492 6222 5514 6239 1 d1
rlabel nwell 5687 6391 5710 6394 1 vdd
rlabel space 5655 6133 5684 6142 1 gnd
rlabel locali 5549 6115 5578 6121 1 gnd
rlabel locali 5552 6414 5581 6420 1 vdd
rlabel nwell 4873 5145 4896 5148 1 vdd
rlabel space 4841 4887 4870 4896 1 gnd
rlabel locali 4735 4869 4764 4875 1 gnd
rlabel locali 4738 5168 4767 5174 1 vdd
rlabel locali 4684 4980 4706 4995 1 d0
rlabel nwell 4872 5557 4895 5560 1 vdd
rlabel space 4840 5299 4869 5308 1 gnd
rlabel locali 4734 5281 4763 5287 1 gnd
rlabel locali 4737 5580 4766 5586 1 vdd
rlabel locali 4683 5392 4705 5407 1 d0
rlabel nwell 4890 6163 4913 6166 1 vdd
rlabel space 4858 5905 4887 5914 1 gnd
rlabel locali 4752 5887 4781 5893 1 gnd
rlabel locali 4755 6186 4784 6192 1 vdd
rlabel locali 4701 5998 4723 6013 1 d0
rlabel nwell 4889 6575 4912 6578 1 vdd
rlabel space 4857 6317 4886 6326 1 gnd
rlabel locali 4751 6299 4780 6305 1 gnd
rlabel locali 4754 6598 4783 6604 1 vdd
rlabel locali 4700 6410 4722 6425 1 d0
rlabel locali 5613 7650 5633 7674 1 d2
rlabel nwell 5806 7819 5829 7822 1 vdd
rlabel space 5774 7561 5803 7570 1 gnd
rlabel locali 5668 7543 5697 7549 1 gnd
rlabel locali 5671 7842 5700 7848 1 vdd
rlabel locali 5512 7240 5534 7257 1 d1
rlabel nwell 5707 7409 5730 7412 1 vdd
rlabel space 5675 7151 5704 7160 1 gnd
rlabel locali 5569 7133 5598 7139 1 gnd
rlabel locali 5572 7432 5601 7438 1 vdd
rlabel locali 5529 8258 5551 8275 1 d1
rlabel nwell 5724 8427 5747 8430 1 vdd
rlabel space 5692 8169 5721 8178 1 gnd
rlabel locali 5586 8151 5615 8157 1 gnd
rlabel locali 5589 8450 5618 8456 1 vdd
rlabel nwell 4910 7181 4933 7184 1 vdd
rlabel space 4878 6923 4907 6932 1 gnd
rlabel locali 4772 6905 4801 6911 1 gnd
rlabel locali 4775 7204 4804 7210 1 vdd
rlabel locali 4721 7016 4743 7031 1 d0
rlabel nwell 4909 7593 4932 7596 1 vdd
rlabel space 4877 7335 4906 7344 1 gnd
rlabel locali 4771 7317 4800 7323 1 gnd
rlabel locali 4774 7616 4803 7622 1 vdd
rlabel locali 4720 7428 4742 7443 1 d0
rlabel nwell 4927 8199 4950 8202 1 vdd
rlabel space 4895 7941 4924 7950 1 gnd
rlabel locali 4789 7923 4818 7929 1 gnd
rlabel locali 4792 8222 4821 8228 1 vdd
rlabel locali 4738 8034 4760 8049 1 d0
rlabel nwell 4926 8611 4949 8614 1 vdd
rlabel space 4894 8353 4923 8362 1 gnd
rlabel locali 4788 8335 4817 8341 1 gnd
rlabel locali 4791 8634 4820 8640 1 vdd
rlabel locali 4737 8446 4759 8461 1 d0
rlabel locali 1456 320 1471 333 1 d5
rlabel locali 1514 507 1543 513 1 vdd
rlabel locali 1511 208 1540 214 1 gnd
rlabel space 1617 226 1646 235 1 gnd
rlabel nwell 1649 484 1672 487 1 vdd
rlabel locali 3938 1240 3960 1255 5 d0
rlabel locali 3877 1061 3906 1067 5 vdd
rlabel locali 3880 1360 3909 1366 5 gnd
rlabel space 3774 1339 3803 1348 5 gnd
rlabel nwell 3748 1087 3771 1090 5 vdd
rlabel locali 3937 1652 3959 1667 5 d0
rlabel locali 3876 1473 3905 1479 5 vdd
rlabel locali 3879 1772 3908 1778 5 gnd
rlabel space 3773 1751 3802 1760 5 gnd
rlabel nwell 3747 1499 3770 1502 5 vdd
rlabel locali 3955 2258 3977 2273 5 d0
rlabel locali 3894 2079 3923 2085 5 vdd
rlabel locali 3897 2378 3926 2384 5 gnd
rlabel space 3791 2357 3820 2366 5 gnd
rlabel nwell 3765 2105 3788 2108 5 vdd
rlabel locali 3954 2670 3976 2685 5 d0
rlabel locali 3893 2491 3922 2497 5 vdd
rlabel locali 3896 2790 3925 2796 5 gnd
rlabel space 3790 2769 3819 2778 5 gnd
rlabel nwell 3764 2517 3787 2520 5 vdd
rlabel locali 3079 1245 3108 1251 5 vdd
rlabel locali 3082 1544 3111 1550 5 gnd
rlabel space 2976 1523 3005 1532 5 gnd
rlabel nwell 2950 1271 2973 1274 5 vdd
rlabel locali 3146 1426 3168 1443 5 d1
rlabel locali 3096 2263 3125 2269 5 vdd
rlabel locali 3099 2562 3128 2568 5 gnd
rlabel space 2993 2541 3022 2550 5 gnd
rlabel nwell 2967 2289 2990 2292 5 vdd
rlabel locali 3163 2444 3185 2461 5 d1
rlabel locali 2997 1853 3026 1859 5 vdd
rlabel locali 3000 2152 3029 2158 5 gnd
rlabel space 2894 2131 2923 2140 5 gnd
rlabel nwell 2868 1879 2891 1882 5 vdd
rlabel locali 3064 2027 3084 2051 5 d2
rlabel locali 3975 3276 3997 3291 5 d0
rlabel locali 3914 3097 3943 3103 5 vdd
rlabel locali 3917 3396 3946 3402 5 gnd
rlabel space 3811 3375 3840 3384 5 gnd
rlabel nwell 3785 3123 3808 3126 5 vdd
rlabel locali 3974 3688 3996 3703 5 d0
rlabel locali 3913 3509 3942 3515 5 vdd
rlabel locali 3916 3808 3945 3814 5 gnd
rlabel space 3810 3787 3839 3796 5 gnd
rlabel nwell 3784 3535 3807 3538 5 vdd
rlabel locali 3992 4294 4014 4309 5 d0
rlabel locali 3931 4115 3960 4121 5 vdd
rlabel locali 3934 4414 3963 4420 5 gnd
rlabel space 3828 4393 3857 4402 5 gnd
rlabel nwell 3802 4141 3825 4144 5 vdd
rlabel locali 3991 4706 4013 4721 5 d0
rlabel locali 3930 4527 3959 4533 5 vdd
rlabel locali 3933 4826 3962 4832 5 gnd
rlabel space 3827 4805 3856 4814 5 gnd
rlabel nwell 3801 4553 3824 4556 5 vdd
rlabel locali 3116 3281 3145 3287 5 vdd
rlabel locali 3119 3580 3148 3586 5 gnd
rlabel space 3013 3559 3042 3568 5 gnd
rlabel nwell 2987 3307 3010 3310 5 vdd
rlabel locali 3183 3462 3205 3479 5 d1
rlabel locali 3133 4299 3162 4305 5 vdd
rlabel locali 3136 4598 3165 4604 5 gnd
rlabel space 3030 4577 3059 4586 5 gnd
rlabel nwell 3004 4325 3027 4328 5 vdd
rlabel locali 3200 4480 3222 4497 5 d1
rlabel locali 3034 3889 3063 3895 5 vdd
rlabel locali 3037 4188 3066 4194 5 gnd
rlabel space 2931 4167 2960 4176 5 gnd
rlabel nwell 2905 3915 2928 3918 5 vdd
rlabel locali 3101 4063 3121 4087 5 d2
rlabel locali 2951 2873 2980 2879 5 vdd
rlabel locali 2954 3172 2983 3178 5 gnd
rlabel space 2848 3151 2877 3160 5 gnd
rlabel nwell 2822 2899 2845 2902 5 vdd
rlabel locali 3016 3052 3036 3065 5 d3
rlabel locali 4011 5312 4033 5327 5 d0
rlabel locali 3950 5133 3979 5139 5 vdd
rlabel locali 3953 5432 3982 5438 5 gnd
rlabel space 3847 5411 3876 5420 5 gnd
rlabel nwell 3821 5159 3844 5162 5 vdd
rlabel locali 4010 5724 4032 5739 5 d0
rlabel locali 3949 5545 3978 5551 5 vdd
rlabel locali 3952 5844 3981 5850 5 gnd
rlabel space 3846 5823 3875 5832 5 gnd
rlabel nwell 3820 5571 3843 5574 5 vdd
rlabel locali 4028 6330 4050 6345 5 d0
rlabel locali 3967 6151 3996 6157 5 vdd
rlabel locali 3970 6450 3999 6456 5 gnd
rlabel space 3864 6429 3893 6438 5 gnd
rlabel nwell 3838 6177 3861 6180 5 vdd
rlabel locali 4027 6742 4049 6757 5 d0
rlabel locali 3966 6563 3995 6569 5 vdd
rlabel locali 3969 6862 3998 6868 5 gnd
rlabel space 3863 6841 3892 6850 5 gnd
rlabel nwell 3837 6589 3860 6592 5 vdd
rlabel locali 3152 5317 3181 5323 5 vdd
rlabel locali 3155 5616 3184 5622 5 gnd
rlabel space 3049 5595 3078 5604 5 gnd
rlabel nwell 3023 5343 3046 5346 5 vdd
rlabel locali 3219 5498 3241 5515 5 d1
rlabel locali 3169 6335 3198 6341 5 vdd
rlabel locali 3172 6634 3201 6640 5 gnd
rlabel space 3066 6613 3095 6622 5 gnd
rlabel nwell 3040 6361 3063 6364 5 vdd
rlabel locali 3236 6516 3258 6533 5 d1
rlabel locali 3070 5925 3099 5931 5 vdd
rlabel locali 3073 6224 3102 6230 5 gnd
rlabel space 2967 6203 2996 6212 5 gnd
rlabel nwell 2941 5951 2964 5954 5 vdd
rlabel locali 3137 6099 3157 6123 5 d2
rlabel locali 4048 7348 4070 7363 5 d0
rlabel locali 3987 7169 4016 7175 5 vdd
rlabel locali 3990 7468 4019 7474 5 gnd
rlabel space 3884 7447 3913 7456 5 gnd
rlabel nwell 3858 7195 3881 7198 5 vdd
rlabel locali 4047 7760 4069 7775 5 d0
rlabel locali 3986 7581 4015 7587 5 vdd
rlabel locali 3989 7880 4018 7886 5 gnd
rlabel space 3883 7859 3912 7868 5 gnd
rlabel nwell 3857 7607 3880 7610 5 vdd
rlabel locali 4065 8366 4087 8381 5 d0
rlabel locali 4004 8187 4033 8193 5 vdd
rlabel locali 4007 8486 4036 8492 5 gnd
rlabel space 3901 8465 3930 8474 5 gnd
rlabel nwell 3875 8213 3898 8216 5 vdd
rlabel locali 4064 8778 4086 8793 5 d0
rlabel locali 4003 8599 4032 8605 5 vdd
rlabel locali 4006 8898 4035 8904 5 gnd
rlabel space 3900 8877 3929 8886 5 gnd
rlabel nwell 3874 8625 3897 8628 5 vdd
rlabel locali 3189 7353 3218 7359 5 vdd
rlabel locali 3192 7652 3221 7658 5 gnd
rlabel space 3086 7631 3115 7640 5 gnd
rlabel nwell 3060 7379 3083 7382 5 vdd
rlabel locali 3256 7534 3278 7551 5 d1
rlabel locali 3206 8371 3235 8377 5 vdd
rlabel locali 3209 8670 3238 8676 5 gnd
rlabel space 3103 8649 3132 8658 5 gnd
rlabel nwell 3077 8397 3100 8400 5 vdd
rlabel locali 3273 8552 3295 8569 5 d1
rlabel locali 3107 7961 3136 7967 5 vdd
rlabel locali 3110 8260 3139 8266 5 gnd
rlabel space 3004 8239 3033 8248 5 gnd
rlabel nwell 2978 7987 3001 7990 5 vdd
rlabel locali 3174 8135 3194 8159 5 d2
rlabel locali 3024 6945 3053 6951 5 vdd
rlabel locali 3027 7244 3056 7250 5 gnd
rlabel space 2921 7223 2950 7232 5 gnd
rlabel nwell 2895 6971 2918 6974 5 vdd
rlabel locali 3089 7124 3109 7137 5 d3
rlabel locali 2848 4911 2877 4917 5 vdd
rlabel locali 2851 5210 2880 5216 5 gnd
rlabel space 2745 5189 2774 5198 5 gnd
rlabel nwell 2719 4937 2742 4940 5 vdd
rlabel locali 2912 5090 2931 5107 5 d4
rlabel locali 1402 4581 1421 4598 1 d4
rlabel nwell 1591 4748 1614 4751 1 vdd
rlabel space 1559 4490 1588 4499 1 gnd
rlabel locali 1453 4472 1482 4478 1 gnd
rlabel locali 1456 4771 1485 4777 1 vdd
rlabel locali 1224 2551 1244 2564 1 d3
rlabel nwell 1415 2714 1438 2717 1 vdd
rlabel space 1383 2456 1412 2465 1 gnd
rlabel locali 1277 2438 1306 2444 1 gnd
rlabel locali 1280 2737 1309 2743 1 vdd
rlabel locali 1139 1529 1159 1553 1 d2
rlabel nwell 1332 1698 1355 1701 1 vdd
rlabel space 1300 1440 1329 1449 1 gnd
rlabel locali 1194 1422 1223 1428 1 gnd
rlabel locali 1197 1721 1226 1727 1 vdd
rlabel locali 1038 1119 1060 1136 1 d1
rlabel nwell 1233 1288 1256 1291 1 vdd
rlabel space 1201 1030 1230 1039 1 gnd
rlabel locali 1095 1012 1124 1018 1 gnd
rlabel locali 1098 1311 1127 1317 1 vdd
rlabel locali 1055 2137 1077 2154 1 d1
rlabel nwell 1250 2306 1273 2309 1 vdd
rlabel space 1218 2048 1247 2057 1 gnd
rlabel locali 1112 2030 1141 2036 1 gnd
rlabel locali 1115 2329 1144 2335 1 vdd
rlabel nwell 436 1060 459 1063 1 vdd
rlabel space 404 802 433 811 1 gnd
rlabel locali 298 784 327 790 1 gnd
rlabel locali 301 1083 330 1089 1 vdd
rlabel locali 247 895 269 910 1 d0
rlabel nwell 435 1472 458 1475 1 vdd
rlabel space 403 1214 432 1223 1 gnd
rlabel locali 297 1196 326 1202 1 gnd
rlabel locali 300 1495 329 1501 1 vdd
rlabel locali 246 1307 268 1322 1 d0
rlabel nwell 453 2078 476 2081 1 vdd
rlabel space 421 1820 450 1829 1 gnd
rlabel locali 315 1802 344 1808 1 gnd
rlabel locali 318 2101 347 2107 1 vdd
rlabel locali 264 1913 286 1928 1 d0
rlabel nwell 452 2490 475 2493 1 vdd
rlabel space 420 2232 449 2241 1 gnd
rlabel locali 314 2214 343 2220 1 gnd
rlabel locali 317 2513 346 2519 1 vdd
rlabel locali 263 2325 285 2340 1 d0
rlabel locali 1176 3565 1196 3589 1 d2
rlabel nwell 1369 3734 1392 3737 1 vdd
rlabel space 1337 3476 1366 3485 1 gnd
rlabel locali 1231 3458 1260 3464 1 gnd
rlabel locali 1234 3757 1263 3763 1 vdd
rlabel locali 1075 3155 1097 3172 1 d1
rlabel nwell 1270 3324 1293 3327 1 vdd
rlabel space 1238 3066 1267 3075 1 gnd
rlabel locali 1132 3048 1161 3054 1 gnd
rlabel locali 1135 3347 1164 3353 1 vdd
rlabel locali 1092 4173 1114 4190 1 d1
rlabel nwell 1287 4342 1310 4345 1 vdd
rlabel space 1255 4084 1284 4093 1 gnd
rlabel locali 1149 4066 1178 4072 1 gnd
rlabel locali 1152 4365 1181 4371 1 vdd
rlabel nwell 473 3096 496 3099 1 vdd
rlabel space 441 2838 470 2847 1 gnd
rlabel locali 335 2820 364 2826 1 gnd
rlabel locali 338 3119 367 3125 1 vdd
rlabel locali 284 2931 306 2946 1 d0
rlabel nwell 472 3508 495 3511 1 vdd
rlabel space 440 3250 469 3259 1 gnd
rlabel locali 334 3232 363 3238 1 gnd
rlabel locali 337 3531 366 3537 1 vdd
rlabel locali 283 3343 305 3358 1 d0
rlabel nwell 490 4114 513 4117 1 vdd
rlabel space 458 3856 487 3865 1 gnd
rlabel locali 352 3838 381 3844 1 gnd
rlabel locali 355 4137 384 4143 1 vdd
rlabel locali 301 3949 323 3964 1 d0
rlabel nwell 489 4526 512 4529 1 vdd
rlabel space 457 4268 486 4277 1 gnd
rlabel locali 351 4250 380 4256 1 gnd
rlabel locali 354 4549 383 4555 1 vdd
rlabel locali 300 4361 322 4376 1 d0
rlabel locali 1297 6623 1317 6636 1 d3
rlabel nwell 1488 6786 1511 6789 1 vdd
rlabel space 1456 6528 1485 6537 1 gnd
rlabel locali 1350 6510 1379 6516 1 gnd
rlabel locali 1353 6809 1382 6815 1 vdd
rlabel locali 1212 5601 1232 5625 1 d2
rlabel nwell 1405 5770 1428 5773 1 vdd
rlabel space 1373 5512 1402 5521 1 gnd
rlabel locali 1267 5494 1296 5500 1 gnd
rlabel locali 1270 5793 1299 5799 1 vdd
rlabel locali 1111 5191 1133 5208 1 d1
rlabel nwell 1306 5360 1329 5363 1 vdd
rlabel space 1274 5102 1303 5111 1 gnd
rlabel locali 1168 5084 1197 5090 1 gnd
rlabel locali 1171 5383 1200 5389 1 vdd
rlabel locali 1128 6209 1150 6226 1 d1
rlabel nwell 1323 6378 1346 6381 1 vdd
rlabel space 1291 6120 1320 6129 1 gnd
rlabel locali 1185 6102 1214 6108 1 gnd
rlabel locali 1188 6401 1217 6407 1 vdd
rlabel nwell 509 5132 532 5135 1 vdd
rlabel space 477 4874 506 4883 1 gnd
rlabel locali 371 4856 400 4862 1 gnd
rlabel locali 374 5155 403 5161 1 vdd
rlabel locali 320 4967 342 4982 1 d0
rlabel nwell 508 5544 531 5547 1 vdd
rlabel space 476 5286 505 5295 1 gnd
rlabel locali 370 5268 399 5274 1 gnd
rlabel locali 373 5567 402 5573 1 vdd
rlabel locali 319 5379 341 5394 1 d0
rlabel nwell 526 6150 549 6153 1 vdd
rlabel space 494 5892 523 5901 1 gnd
rlabel locali 388 5874 417 5880 1 gnd
rlabel locali 391 6173 420 6179 1 vdd
rlabel locali 337 5985 359 6000 1 d0
rlabel nwell 525 6562 548 6565 1 vdd
rlabel space 493 6304 522 6313 1 gnd
rlabel locali 387 6286 416 6292 1 gnd
rlabel locali 390 6585 419 6591 1 vdd
rlabel locali 336 6397 358 6412 1 d0
rlabel locali 1249 7637 1269 7661 1 d2
rlabel nwell 1442 7806 1465 7809 1 vdd
rlabel space 1410 7548 1439 7557 1 gnd
rlabel locali 1304 7530 1333 7536 1 gnd
rlabel locali 1307 7829 1336 7835 1 vdd
rlabel locali 1148 7227 1170 7244 1 d1
rlabel nwell 1343 7396 1366 7399 1 vdd
rlabel space 1311 7138 1340 7147 1 gnd
rlabel locali 1205 7120 1234 7126 1 gnd
rlabel locali 1208 7419 1237 7425 1 vdd
rlabel locali 1165 8245 1187 8262 1 d1
rlabel nwell 1360 8414 1383 8417 1 vdd
rlabel space 1328 8156 1357 8165 1 gnd
rlabel locali 1222 8138 1251 8144 1 gnd
rlabel locali 1225 8437 1254 8443 1 vdd
rlabel nwell 546 7168 569 7171 1 vdd
rlabel space 514 6910 543 6919 1 gnd
rlabel locali 408 6892 437 6898 1 gnd
rlabel locali 411 7191 440 7197 1 vdd
rlabel locali 357 7003 379 7018 1 d0
rlabel nwell 545 7580 568 7583 1 vdd
rlabel space 513 7322 542 7331 1 gnd
rlabel locali 407 7304 436 7310 1 gnd
rlabel locali 410 7603 439 7609 1 vdd
rlabel locali 356 7415 378 7430 1 d0
rlabel locali 264 8866 288 8896 1 vref
rlabel nwell 563 8186 586 8189 1 vdd
rlabel space 531 7928 560 7937 1 gnd
rlabel locali 425 7910 454 7916 1 gnd
rlabel locali 428 8209 457 8215 1 vdd
rlabel locali 374 8021 396 8036 1 d0
rlabel nwell 562 8598 585 8601 1 vdd
rlabel space 530 8340 559 8349 1 gnd
rlabel locali 424 8322 453 8328 1 gnd
rlabel locali 427 8621 456 8627 1 vdd
rlabel locali 373 8433 395 8448 1 d0
rlabel locali 12680 268 12703 284 1 d6
rlabel locali 12744 458 12773 464 1 vdd
rlabel locali 12741 159 12770 165 1 gnd
rlabel space 12847 177 12876 186 1 gnd
rlabel nwell 12879 435 12902 438 1 vdd
rlabel locali 14561 358 14576 371 1 d5
rlabel locali 14619 545 14648 551 1 vdd
rlabel locali 14616 246 14645 252 1 gnd
rlabel space 14722 264 14751 273 1 gnd
rlabel nwell 14754 522 14777 525 1 vdd
rlabel locali 17043 1278 17065 1293 5 d0
rlabel locali 16982 1099 17011 1105 5 vdd
rlabel locali 16985 1398 17014 1404 5 gnd
rlabel space 16879 1377 16908 1386 5 gnd
rlabel nwell 16853 1125 16876 1128 5 vdd
rlabel locali 17042 1690 17064 1705 5 d0
rlabel locali 16981 1511 17010 1517 5 vdd
rlabel locali 16984 1810 17013 1816 5 gnd
rlabel space 16878 1789 16907 1798 5 gnd
rlabel nwell 16852 1537 16875 1540 5 vdd
rlabel locali 17060 2296 17082 2311 5 d0
rlabel locali 16999 2117 17028 2123 5 vdd
rlabel locali 17002 2416 17031 2422 5 gnd
rlabel space 16896 2395 16925 2404 5 gnd
rlabel nwell 16870 2143 16893 2146 5 vdd
rlabel locali 17059 2708 17081 2723 5 d0
rlabel locali 16998 2529 17027 2535 5 vdd
rlabel locali 17001 2828 17030 2834 5 gnd
rlabel space 16895 2807 16924 2816 5 gnd
rlabel nwell 16869 2555 16892 2558 5 vdd
rlabel locali 16184 1283 16213 1289 5 vdd
rlabel locali 16187 1582 16216 1588 5 gnd
rlabel space 16081 1561 16110 1570 5 gnd
rlabel nwell 16055 1309 16078 1312 5 vdd
rlabel locali 16251 1464 16273 1481 5 d1
rlabel locali 16201 2301 16230 2307 5 vdd
rlabel locali 16204 2600 16233 2606 5 gnd
rlabel space 16098 2579 16127 2588 5 gnd
rlabel nwell 16072 2327 16095 2330 5 vdd
rlabel locali 16268 2482 16290 2499 5 d1
rlabel locali 16102 1891 16131 1897 5 vdd
rlabel locali 16105 2190 16134 2196 5 gnd
rlabel space 15999 2169 16028 2178 5 gnd
rlabel nwell 15973 1917 15996 1920 5 vdd
rlabel locali 16169 2065 16189 2089 5 d2
rlabel locali 17080 3314 17102 3329 5 d0
rlabel locali 17019 3135 17048 3141 5 vdd
rlabel locali 17022 3434 17051 3440 5 gnd
rlabel space 16916 3413 16945 3422 5 gnd
rlabel nwell 16890 3161 16913 3164 5 vdd
rlabel locali 17079 3726 17101 3741 5 d0
rlabel locali 17018 3547 17047 3553 5 vdd
rlabel locali 17021 3846 17050 3852 5 gnd
rlabel space 16915 3825 16944 3834 5 gnd
rlabel nwell 16889 3573 16912 3576 5 vdd
rlabel locali 17097 4332 17119 4347 5 d0
rlabel locali 17036 4153 17065 4159 5 vdd
rlabel locali 17039 4452 17068 4458 5 gnd
rlabel space 16933 4431 16962 4440 5 gnd
rlabel nwell 16907 4179 16930 4182 5 vdd
rlabel locali 17096 4744 17118 4759 5 d0
rlabel locali 17035 4565 17064 4571 5 vdd
rlabel locali 17038 4864 17067 4870 5 gnd
rlabel space 16932 4843 16961 4852 5 gnd
rlabel nwell 16906 4591 16929 4594 5 vdd
rlabel locali 16221 3319 16250 3325 5 vdd
rlabel locali 16224 3618 16253 3624 5 gnd
rlabel space 16118 3597 16147 3606 5 gnd
rlabel nwell 16092 3345 16115 3348 5 vdd
rlabel locali 16288 3500 16310 3517 5 d1
rlabel locali 16238 4337 16267 4343 5 vdd
rlabel locali 16241 4636 16270 4642 5 gnd
rlabel space 16135 4615 16164 4624 5 gnd
rlabel nwell 16109 4363 16132 4366 5 vdd
rlabel locali 16305 4518 16327 4535 5 d1
rlabel locali 16139 3927 16168 3933 5 vdd
rlabel locali 16142 4226 16171 4232 5 gnd
rlabel space 16036 4205 16065 4214 5 gnd
rlabel nwell 16010 3953 16033 3956 5 vdd
rlabel locali 16206 4101 16226 4125 5 d2
rlabel locali 16056 2911 16085 2917 5 vdd
rlabel locali 16059 3210 16088 3216 5 gnd
rlabel space 15953 3189 15982 3198 5 gnd
rlabel nwell 15927 2937 15950 2940 5 vdd
rlabel locali 16121 3090 16141 3103 5 d3
rlabel locali 17116 5350 17138 5365 5 d0
rlabel locali 17055 5171 17084 5177 5 vdd
rlabel locali 17058 5470 17087 5476 5 gnd
rlabel space 16952 5449 16981 5458 5 gnd
rlabel nwell 16926 5197 16949 5200 5 vdd
rlabel locali 17115 5762 17137 5777 5 d0
rlabel locali 17054 5583 17083 5589 5 vdd
rlabel locali 17057 5882 17086 5888 5 gnd
rlabel space 16951 5861 16980 5870 5 gnd
rlabel nwell 16925 5609 16948 5612 5 vdd
rlabel locali 17133 6368 17155 6383 5 d0
rlabel locali 17072 6189 17101 6195 5 vdd
rlabel locali 17075 6488 17104 6494 5 gnd
rlabel space 16969 6467 16998 6476 5 gnd
rlabel nwell 16943 6215 16966 6218 5 vdd
rlabel locali 17132 6780 17154 6795 5 d0
rlabel locali 17071 6601 17100 6607 5 vdd
rlabel locali 17074 6900 17103 6906 5 gnd
rlabel space 16968 6879 16997 6888 5 gnd
rlabel nwell 16942 6627 16965 6630 5 vdd
rlabel locali 16257 5355 16286 5361 5 vdd
rlabel locali 16260 5654 16289 5660 5 gnd
rlabel space 16154 5633 16183 5642 5 gnd
rlabel nwell 16128 5381 16151 5384 5 vdd
rlabel locali 16324 5536 16346 5553 5 d1
rlabel locali 16274 6373 16303 6379 5 vdd
rlabel locali 16277 6672 16306 6678 5 gnd
rlabel space 16171 6651 16200 6660 5 gnd
rlabel nwell 16145 6399 16168 6402 5 vdd
rlabel locali 16341 6554 16363 6571 5 d1
rlabel locali 16175 5963 16204 5969 5 vdd
rlabel locali 16178 6262 16207 6268 5 gnd
rlabel space 16072 6241 16101 6250 5 gnd
rlabel nwell 16046 5989 16069 5992 5 vdd
rlabel locali 16242 6137 16262 6161 5 d2
rlabel locali 17153 7386 17175 7401 5 d0
rlabel locali 17092 7207 17121 7213 5 vdd
rlabel locali 17095 7506 17124 7512 5 gnd
rlabel space 16989 7485 17018 7494 5 gnd
rlabel nwell 16963 7233 16986 7236 5 vdd
rlabel locali 17152 7798 17174 7813 5 d0
rlabel locali 17091 7619 17120 7625 5 vdd
rlabel locali 17094 7918 17123 7924 5 gnd
rlabel space 16988 7897 17017 7906 5 gnd
rlabel nwell 16962 7645 16985 7648 5 vdd
rlabel locali 17170 8404 17192 8419 5 d0
rlabel locali 17109 8225 17138 8231 5 vdd
rlabel locali 17112 8524 17141 8530 5 gnd
rlabel space 17006 8503 17035 8512 5 gnd
rlabel nwell 16980 8251 17003 8254 5 vdd
rlabel locali 17169 8816 17191 8831 5 d0
rlabel locali 17108 8637 17137 8643 5 vdd
rlabel locali 17111 8936 17140 8942 5 gnd
rlabel space 17005 8915 17034 8924 5 gnd
rlabel nwell 16979 8663 17002 8666 5 vdd
rlabel locali 16294 7391 16323 7397 5 vdd
rlabel locali 16297 7690 16326 7696 5 gnd
rlabel space 16191 7669 16220 7678 5 gnd
rlabel nwell 16165 7417 16188 7420 5 vdd
rlabel locali 16361 7572 16383 7589 5 d1
rlabel locali 16311 8409 16340 8415 5 vdd
rlabel locali 16314 8708 16343 8714 5 gnd
rlabel space 16208 8687 16237 8696 5 gnd
rlabel nwell 16182 8435 16205 8438 5 vdd
rlabel locali 16378 8590 16400 8607 5 d1
rlabel locali 16212 7999 16241 8005 5 vdd
rlabel locali 16215 8298 16244 8304 5 gnd
rlabel space 16109 8277 16138 8286 5 gnd
rlabel nwell 16083 8025 16106 8028 5 vdd
rlabel locali 16279 8173 16299 8197 5 d2
rlabel locali 16129 6983 16158 6989 5 vdd
rlabel locali 16132 7282 16161 7288 5 gnd
rlabel space 16026 7261 16055 7270 5 gnd
rlabel nwell 16000 7009 16023 7012 5 vdd
rlabel locali 16194 7162 16214 7175 5 d3
rlabel locali 15953 4949 15982 4955 5 vdd
rlabel locali 15956 5248 15985 5254 5 gnd
rlabel space 15850 5227 15879 5236 5 gnd
rlabel nwell 15824 4975 15847 4978 5 vdd
rlabel locali 16017 5128 16036 5145 5 d4
rlabel locali 14507 4619 14526 4636 1 d4
rlabel nwell 14696 4786 14719 4789 1 vdd
rlabel space 14664 4528 14693 4537 1 gnd
rlabel locali 14558 4510 14587 4516 1 gnd
rlabel locali 14561 4809 14590 4815 1 vdd
rlabel locali 14329 2589 14349 2602 1 d3
rlabel nwell 14520 2752 14543 2755 1 vdd
rlabel space 14488 2494 14517 2503 1 gnd
rlabel locali 14382 2476 14411 2482 1 gnd
rlabel locali 14385 2775 14414 2781 1 vdd
rlabel locali 14244 1567 14264 1591 1 d2
rlabel nwell 14437 1736 14460 1739 1 vdd
rlabel space 14405 1478 14434 1487 1 gnd
rlabel locali 14299 1460 14328 1466 1 gnd
rlabel locali 14302 1759 14331 1765 1 vdd
rlabel locali 14143 1157 14165 1174 1 d1
rlabel nwell 14338 1326 14361 1329 1 vdd
rlabel space 14306 1068 14335 1077 1 gnd
rlabel locali 14200 1050 14229 1056 1 gnd
rlabel locali 14203 1349 14232 1355 1 vdd
rlabel locali 14160 2175 14182 2192 1 d1
rlabel nwell 14355 2344 14378 2347 1 vdd
rlabel space 14323 2086 14352 2095 1 gnd
rlabel locali 14217 2068 14246 2074 1 gnd
rlabel locali 14220 2367 14249 2373 1 vdd
rlabel nwell 13541 1098 13564 1101 1 vdd
rlabel space 13509 840 13538 849 1 gnd
rlabel locali 13403 822 13432 828 1 gnd
rlabel locali 13406 1121 13435 1127 1 vdd
rlabel locali 13352 933 13374 948 1 d0
rlabel nwell 13540 1510 13563 1513 1 vdd
rlabel space 13508 1252 13537 1261 1 gnd
rlabel locali 13402 1234 13431 1240 1 gnd
rlabel locali 13405 1533 13434 1539 1 vdd
rlabel locali 13351 1345 13373 1360 1 d0
rlabel nwell 13558 2116 13581 2119 1 vdd
rlabel space 13526 1858 13555 1867 1 gnd
rlabel locali 13420 1840 13449 1846 1 gnd
rlabel locali 13423 2139 13452 2145 1 vdd
rlabel locali 13369 1951 13391 1966 1 d0
rlabel nwell 13557 2528 13580 2531 1 vdd
rlabel space 13525 2270 13554 2279 1 gnd
rlabel locali 13419 2252 13448 2258 1 gnd
rlabel locali 13422 2551 13451 2557 1 vdd
rlabel locali 13368 2363 13390 2378 1 d0
rlabel locali 14281 3603 14301 3627 1 d2
rlabel nwell 14474 3772 14497 3775 1 vdd
rlabel space 14442 3514 14471 3523 1 gnd
rlabel locali 14336 3496 14365 3502 1 gnd
rlabel locali 14339 3795 14368 3801 1 vdd
rlabel locali 14180 3193 14202 3210 1 d1
rlabel nwell 14375 3362 14398 3365 1 vdd
rlabel space 14343 3104 14372 3113 1 gnd
rlabel locali 14237 3086 14266 3092 1 gnd
rlabel locali 14240 3385 14269 3391 1 vdd
rlabel locali 14197 4211 14219 4228 1 d1
rlabel nwell 14392 4380 14415 4383 1 vdd
rlabel space 14360 4122 14389 4131 1 gnd
rlabel locali 14254 4104 14283 4110 1 gnd
rlabel locali 14257 4403 14286 4409 1 vdd
rlabel nwell 13578 3134 13601 3137 1 vdd
rlabel space 13546 2876 13575 2885 1 gnd
rlabel locali 13440 2858 13469 2864 1 gnd
rlabel locali 13443 3157 13472 3163 1 vdd
rlabel locali 13389 2969 13411 2984 1 d0
rlabel nwell 13577 3546 13600 3549 1 vdd
rlabel space 13545 3288 13574 3297 1 gnd
rlabel locali 13439 3270 13468 3276 1 gnd
rlabel locali 13442 3569 13471 3575 1 vdd
rlabel locali 13388 3381 13410 3396 1 d0
rlabel nwell 13595 4152 13618 4155 1 vdd
rlabel space 13563 3894 13592 3903 1 gnd
rlabel locali 13457 3876 13486 3882 1 gnd
rlabel locali 13460 4175 13489 4181 1 vdd
rlabel locali 13406 3987 13428 4002 1 d0
rlabel nwell 13594 4564 13617 4567 1 vdd
rlabel space 13562 4306 13591 4315 1 gnd
rlabel locali 13456 4288 13485 4294 1 gnd
rlabel locali 13459 4587 13488 4593 1 vdd
rlabel locali 13405 4399 13427 4414 1 d0
rlabel locali 14402 6661 14422 6674 1 d3
rlabel nwell 14593 6824 14616 6827 1 vdd
rlabel space 14561 6566 14590 6575 1 gnd
rlabel locali 14455 6548 14484 6554 1 gnd
rlabel locali 14458 6847 14487 6853 1 vdd
rlabel locali 14317 5639 14337 5663 1 d2
rlabel nwell 14510 5808 14533 5811 1 vdd
rlabel space 14478 5550 14507 5559 1 gnd
rlabel locali 14372 5532 14401 5538 1 gnd
rlabel locali 14375 5831 14404 5837 1 vdd
rlabel locali 14216 5229 14238 5246 1 d1
rlabel nwell 14411 5398 14434 5401 1 vdd
rlabel space 14379 5140 14408 5149 1 gnd
rlabel locali 14273 5122 14302 5128 1 gnd
rlabel locali 14276 5421 14305 5427 1 vdd
rlabel locali 14233 6247 14255 6264 1 d1
rlabel nwell 14428 6416 14451 6419 1 vdd
rlabel space 14396 6158 14425 6167 1 gnd
rlabel locali 14290 6140 14319 6146 1 gnd
rlabel locali 14293 6439 14322 6445 1 vdd
rlabel nwell 13614 5170 13637 5173 1 vdd
rlabel space 13582 4912 13611 4921 1 gnd
rlabel locali 13476 4894 13505 4900 1 gnd
rlabel locali 13479 5193 13508 5199 1 vdd
rlabel locali 13425 5005 13447 5020 1 d0
rlabel nwell 13613 5582 13636 5585 1 vdd
rlabel space 13581 5324 13610 5333 1 gnd
rlabel locali 13475 5306 13504 5312 1 gnd
rlabel locali 13478 5605 13507 5611 1 vdd
rlabel locali 13424 5417 13446 5432 1 d0
rlabel nwell 13631 6188 13654 6191 1 vdd
rlabel space 13599 5930 13628 5939 1 gnd
rlabel locali 13493 5912 13522 5918 1 gnd
rlabel locali 13496 6211 13525 6217 1 vdd
rlabel locali 13442 6023 13464 6038 1 d0
rlabel nwell 13630 6600 13653 6603 1 vdd
rlabel space 13598 6342 13627 6351 1 gnd
rlabel locali 13492 6324 13521 6330 1 gnd
rlabel locali 13495 6623 13524 6629 1 vdd
rlabel locali 13441 6435 13463 6450 1 d0
rlabel locali 14354 7675 14374 7699 1 d2
rlabel nwell 14547 7844 14570 7847 1 vdd
rlabel space 14515 7586 14544 7595 1 gnd
rlabel locali 14409 7568 14438 7574 1 gnd
rlabel locali 14412 7867 14441 7873 1 vdd
rlabel locali 14253 7265 14275 7282 1 d1
rlabel nwell 14448 7434 14471 7437 1 vdd
rlabel space 14416 7176 14445 7185 1 gnd
rlabel locali 14310 7158 14339 7164 1 gnd
rlabel locali 14313 7457 14342 7463 1 vdd
rlabel locali 14270 8283 14292 8300 1 d1
rlabel nwell 14465 8452 14488 8455 1 vdd
rlabel space 14433 8194 14462 8203 1 gnd
rlabel locali 14327 8176 14356 8182 1 gnd
rlabel locali 14330 8475 14359 8481 1 vdd
rlabel nwell 13651 7206 13674 7209 1 vdd
rlabel space 13619 6948 13648 6957 1 gnd
rlabel locali 13513 6930 13542 6936 1 gnd
rlabel locali 13516 7229 13545 7235 1 vdd
rlabel locali 13462 7041 13484 7056 1 d0
rlabel nwell 13650 7618 13673 7621 1 vdd
rlabel space 13618 7360 13647 7369 1 gnd
rlabel locali 13512 7342 13541 7348 1 gnd
rlabel locali 13515 7641 13544 7647 1 vdd
rlabel locali 13461 7453 13483 7468 1 d0
rlabel nwell 13668 8224 13691 8227 1 vdd
rlabel space 13636 7966 13665 7975 1 gnd
rlabel locali 13530 7948 13559 7954 1 gnd
rlabel locali 13533 8247 13562 8253 1 vdd
rlabel locali 13479 8059 13501 8074 1 d0
rlabel nwell 13667 8636 13690 8639 1 vdd
rlabel space 13635 8378 13664 8387 1 gnd
rlabel locali 13529 8360 13558 8366 1 gnd
rlabel locali 13532 8659 13561 8665 1 vdd
rlabel locali 13478 8471 13500 8486 1 d0
rlabel locali 10197 345 10212 358 1 d5
rlabel locali 10255 532 10284 538 1 vdd
rlabel locali 10252 233 10281 239 1 gnd
rlabel space 10358 251 10387 260 1 gnd
rlabel nwell 10390 509 10413 512 1 vdd
rlabel locali 12679 1265 12701 1280 5 d0
rlabel locali 12618 1086 12647 1092 5 vdd
rlabel locali 12621 1385 12650 1391 5 gnd
rlabel space 12515 1364 12544 1373 5 gnd
rlabel nwell 12489 1112 12512 1115 5 vdd
rlabel locali 12678 1677 12700 1692 5 d0
rlabel locali 12617 1498 12646 1504 5 vdd
rlabel locali 12620 1797 12649 1803 5 gnd
rlabel space 12514 1776 12543 1785 5 gnd
rlabel nwell 12488 1524 12511 1527 5 vdd
rlabel locali 12696 2283 12718 2298 5 d0
rlabel locali 12635 2104 12664 2110 5 vdd
rlabel locali 12638 2403 12667 2409 5 gnd
rlabel space 12532 2382 12561 2391 5 gnd
rlabel nwell 12506 2130 12529 2133 5 vdd
rlabel locali 12695 2695 12717 2710 5 d0
rlabel locali 12634 2516 12663 2522 5 vdd
rlabel locali 12637 2815 12666 2821 5 gnd
rlabel space 12531 2794 12560 2803 5 gnd
rlabel nwell 12505 2542 12528 2545 5 vdd
rlabel locali 11820 1270 11849 1276 5 vdd
rlabel locali 11823 1569 11852 1575 5 gnd
rlabel space 11717 1548 11746 1557 5 gnd
rlabel nwell 11691 1296 11714 1299 5 vdd
rlabel locali 11887 1451 11909 1468 5 d1
rlabel locali 11837 2288 11866 2294 5 vdd
rlabel locali 11840 2587 11869 2593 5 gnd
rlabel space 11734 2566 11763 2575 5 gnd
rlabel nwell 11708 2314 11731 2317 5 vdd
rlabel locali 11904 2469 11926 2486 5 d1
rlabel locali 11738 1878 11767 1884 5 vdd
rlabel locali 11741 2177 11770 2183 5 gnd
rlabel space 11635 2156 11664 2165 5 gnd
rlabel nwell 11609 1904 11632 1907 5 vdd
rlabel locali 11805 2052 11825 2076 5 d2
rlabel locali 12716 3301 12738 3316 5 d0
rlabel locali 12655 3122 12684 3128 5 vdd
rlabel locali 12658 3421 12687 3427 5 gnd
rlabel space 12552 3400 12581 3409 5 gnd
rlabel nwell 12526 3148 12549 3151 5 vdd
rlabel locali 12715 3713 12737 3728 5 d0
rlabel locali 12654 3534 12683 3540 5 vdd
rlabel locali 12657 3833 12686 3839 5 gnd
rlabel space 12551 3812 12580 3821 5 gnd
rlabel nwell 12525 3560 12548 3563 5 vdd
rlabel locali 12733 4319 12755 4334 5 d0
rlabel locali 12672 4140 12701 4146 5 vdd
rlabel locali 12675 4439 12704 4445 5 gnd
rlabel space 12569 4418 12598 4427 5 gnd
rlabel nwell 12543 4166 12566 4169 5 vdd
rlabel locali 12732 4731 12754 4746 5 d0
rlabel locali 12671 4552 12700 4558 5 vdd
rlabel locali 12674 4851 12703 4857 5 gnd
rlabel space 12568 4830 12597 4839 5 gnd
rlabel nwell 12542 4578 12565 4581 5 vdd
rlabel locali 11857 3306 11886 3312 5 vdd
rlabel locali 11860 3605 11889 3611 5 gnd
rlabel space 11754 3584 11783 3593 5 gnd
rlabel nwell 11728 3332 11751 3335 5 vdd
rlabel locali 11924 3487 11946 3504 5 d1
rlabel locali 11874 4324 11903 4330 5 vdd
rlabel locali 11877 4623 11906 4629 5 gnd
rlabel space 11771 4602 11800 4611 5 gnd
rlabel nwell 11745 4350 11768 4353 5 vdd
rlabel locali 11941 4505 11963 4522 5 d1
rlabel locali 11775 3914 11804 3920 5 vdd
rlabel locali 11778 4213 11807 4219 5 gnd
rlabel space 11672 4192 11701 4201 5 gnd
rlabel nwell 11646 3940 11669 3943 5 vdd
rlabel locali 11842 4088 11862 4112 5 d2
rlabel locali 11692 2898 11721 2904 5 vdd
rlabel locali 11695 3197 11724 3203 5 gnd
rlabel space 11589 3176 11618 3185 5 gnd
rlabel nwell 11563 2924 11586 2927 5 vdd
rlabel locali 11757 3077 11777 3090 5 d3
rlabel locali 12752 5337 12774 5352 5 d0
rlabel locali 12691 5158 12720 5164 5 vdd
rlabel locali 12694 5457 12723 5463 5 gnd
rlabel space 12588 5436 12617 5445 5 gnd
rlabel nwell 12562 5184 12585 5187 5 vdd
rlabel locali 12751 5749 12773 5764 5 d0
rlabel locali 12690 5570 12719 5576 5 vdd
rlabel locali 12693 5869 12722 5875 5 gnd
rlabel space 12587 5848 12616 5857 5 gnd
rlabel nwell 12561 5596 12584 5599 5 vdd
rlabel locali 12769 6355 12791 6370 5 d0
rlabel locali 12708 6176 12737 6182 5 vdd
rlabel locali 12711 6475 12740 6481 5 gnd
rlabel space 12605 6454 12634 6463 5 gnd
rlabel nwell 12579 6202 12602 6205 5 vdd
rlabel locali 12768 6767 12790 6782 5 d0
rlabel locali 12707 6588 12736 6594 5 vdd
rlabel locali 12710 6887 12739 6893 5 gnd
rlabel space 12604 6866 12633 6875 5 gnd
rlabel nwell 12578 6614 12601 6617 5 vdd
rlabel locali 11893 5342 11922 5348 5 vdd
rlabel locali 11896 5641 11925 5647 5 gnd
rlabel space 11790 5620 11819 5629 5 gnd
rlabel nwell 11764 5368 11787 5371 5 vdd
rlabel locali 11960 5523 11982 5540 5 d1
rlabel locali 11910 6360 11939 6366 5 vdd
rlabel locali 11913 6659 11942 6665 5 gnd
rlabel space 11807 6638 11836 6647 5 gnd
rlabel nwell 11781 6386 11804 6389 5 vdd
rlabel locali 11977 6541 11999 6558 5 d1
rlabel locali 11811 5950 11840 5956 5 vdd
rlabel locali 11814 6249 11843 6255 5 gnd
rlabel space 11708 6228 11737 6237 5 gnd
rlabel nwell 11682 5976 11705 5979 5 vdd
rlabel locali 11878 6124 11898 6148 5 d2
rlabel locali 12789 7373 12811 7388 5 d0
rlabel locali 12728 7194 12757 7200 5 vdd
rlabel locali 12731 7493 12760 7499 5 gnd
rlabel space 12625 7472 12654 7481 5 gnd
rlabel nwell 12599 7220 12622 7223 5 vdd
rlabel locali 12788 7785 12810 7800 5 d0
rlabel locali 12727 7606 12756 7612 5 vdd
rlabel locali 12730 7905 12759 7911 5 gnd
rlabel space 12624 7884 12653 7893 5 gnd
rlabel nwell 12598 7632 12621 7635 5 vdd
rlabel locali 12806 8391 12828 8406 5 d0
rlabel locali 12745 8212 12774 8218 5 vdd
rlabel locali 12748 8511 12777 8517 5 gnd
rlabel space 12642 8490 12671 8499 5 gnd
rlabel nwell 12616 8238 12639 8241 5 vdd
rlabel locali 12805 8803 12827 8818 5 d0
rlabel locali 12744 8624 12773 8630 5 vdd
rlabel locali 12747 8923 12776 8929 5 gnd
rlabel space 12641 8902 12670 8911 5 gnd
rlabel nwell 12615 8650 12638 8653 5 vdd
rlabel locali 11930 7378 11959 7384 5 vdd
rlabel locali 11933 7677 11962 7683 5 gnd
rlabel space 11827 7656 11856 7665 5 gnd
rlabel nwell 11801 7404 11824 7407 5 vdd
rlabel locali 11997 7559 12019 7576 5 d1
rlabel locali 11947 8396 11976 8402 5 vdd
rlabel locali 11950 8695 11979 8701 5 gnd
rlabel space 11844 8674 11873 8683 5 gnd
rlabel nwell 11818 8422 11841 8425 5 vdd
rlabel locali 12014 8577 12036 8594 5 d1
rlabel locali 11848 7986 11877 7992 5 vdd
rlabel locali 11851 8285 11880 8291 5 gnd
rlabel space 11745 8264 11774 8273 5 gnd
rlabel nwell 11719 8012 11742 8015 5 vdd
rlabel locali 11915 8160 11935 8184 5 d2
rlabel locali 11765 6970 11794 6976 5 vdd
rlabel locali 11768 7269 11797 7275 5 gnd
rlabel space 11662 7248 11691 7257 5 gnd
rlabel nwell 11636 6996 11659 6999 5 vdd
rlabel locali 11830 7149 11850 7162 5 d3
rlabel locali 11589 4936 11618 4942 5 vdd
rlabel locali 11592 5235 11621 5241 5 gnd
rlabel space 11486 5214 11515 5223 5 gnd
rlabel nwell 11460 4962 11483 4965 5 vdd
rlabel locali 11653 5115 11672 5132 5 d4
rlabel locali 10143 4606 10162 4623 1 d4
rlabel nwell 10332 4773 10355 4776 1 vdd
rlabel space 10300 4515 10329 4524 1 gnd
rlabel locali 10194 4497 10223 4503 1 gnd
rlabel locali 10197 4796 10226 4802 1 vdd
rlabel locali 9965 2576 9985 2589 1 d3
rlabel nwell 10156 2739 10179 2742 1 vdd
rlabel space 10124 2481 10153 2490 1 gnd
rlabel locali 10018 2463 10047 2469 1 gnd
rlabel locali 10021 2762 10050 2768 1 vdd
rlabel locali 9880 1554 9900 1578 1 d2
rlabel nwell 10073 1723 10096 1726 1 vdd
rlabel space 10041 1465 10070 1474 1 gnd
rlabel locali 9935 1447 9964 1453 1 gnd
rlabel locali 9938 1746 9967 1752 1 vdd
rlabel locali 9779 1144 9801 1161 1 d1
rlabel nwell 9974 1313 9997 1316 1 vdd
rlabel space 9942 1055 9971 1064 1 gnd
rlabel locali 9836 1037 9865 1043 1 gnd
rlabel locali 9839 1336 9868 1342 1 vdd
rlabel locali 9796 2162 9818 2179 1 d1
rlabel nwell 9991 2331 10014 2334 1 vdd
rlabel space 9959 2073 9988 2082 1 gnd
rlabel locali 9853 2055 9882 2061 1 gnd
rlabel locali 9856 2354 9885 2360 1 vdd
rlabel nwell 9177 1085 9200 1088 1 vdd
rlabel space 9145 827 9174 836 1 gnd
rlabel locali 9039 809 9068 815 1 gnd
rlabel locali 9042 1108 9071 1114 1 vdd
rlabel locali 8988 920 9010 935 1 d0
rlabel nwell 9176 1497 9199 1500 1 vdd
rlabel space 9144 1239 9173 1248 1 gnd
rlabel locali 9038 1221 9067 1227 1 gnd
rlabel locali 9041 1520 9070 1526 1 vdd
rlabel locali 8987 1332 9009 1347 1 d0
rlabel nwell 9194 2103 9217 2106 1 vdd
rlabel space 9162 1845 9191 1854 1 gnd
rlabel locali 9056 1827 9085 1833 1 gnd
rlabel locali 9059 2126 9088 2132 1 vdd
rlabel locali 9005 1938 9027 1953 1 d0
rlabel nwell 9193 2515 9216 2518 1 vdd
rlabel space 9161 2257 9190 2266 1 gnd
rlabel locali 9055 2239 9084 2245 1 gnd
rlabel locali 9058 2538 9087 2544 1 vdd
rlabel locali 9004 2350 9026 2365 1 d0
rlabel locali 9917 3590 9937 3614 1 d2
rlabel nwell 10110 3759 10133 3762 1 vdd
rlabel space 10078 3501 10107 3510 1 gnd
rlabel locali 9972 3483 10001 3489 1 gnd
rlabel locali 9975 3782 10004 3788 1 vdd
rlabel locali 9816 3180 9838 3197 1 d1
rlabel nwell 10011 3349 10034 3352 1 vdd
rlabel space 9979 3091 10008 3100 1 gnd
rlabel locali 9873 3073 9902 3079 1 gnd
rlabel locali 9876 3372 9905 3378 1 vdd
rlabel locali 9833 4198 9855 4215 1 d1
rlabel nwell 10028 4367 10051 4370 1 vdd
rlabel space 9996 4109 10025 4118 1 gnd
rlabel locali 9890 4091 9919 4097 1 gnd
rlabel locali 9893 4390 9922 4396 1 vdd
rlabel nwell 9214 3121 9237 3124 1 vdd
rlabel space 9182 2863 9211 2872 1 gnd
rlabel locali 9076 2845 9105 2851 1 gnd
rlabel locali 9079 3144 9108 3150 1 vdd
rlabel locali 9025 2956 9047 2971 1 d0
rlabel nwell 9213 3533 9236 3536 1 vdd
rlabel space 9181 3275 9210 3284 1 gnd
rlabel locali 9075 3257 9104 3263 1 gnd
rlabel locali 9078 3556 9107 3562 1 vdd
rlabel locali 9024 3368 9046 3383 1 d0
rlabel nwell 9231 4139 9254 4142 1 vdd
rlabel space 9199 3881 9228 3890 1 gnd
rlabel locali 9093 3863 9122 3869 1 gnd
rlabel locali 9096 4162 9125 4168 1 vdd
rlabel locali 9042 3974 9064 3989 1 d0
rlabel nwell 9230 4551 9253 4554 1 vdd
rlabel space 9198 4293 9227 4302 1 gnd
rlabel locali 9092 4275 9121 4281 1 gnd
rlabel locali 9095 4574 9124 4580 1 vdd
rlabel locali 9041 4386 9063 4401 1 d0
rlabel locali 10038 6648 10058 6661 1 d3
rlabel nwell 10229 6811 10252 6814 1 vdd
rlabel space 10197 6553 10226 6562 1 gnd
rlabel locali 10091 6535 10120 6541 1 gnd
rlabel locali 10094 6834 10123 6840 1 vdd
rlabel locali 9953 5626 9973 5650 1 d2
rlabel nwell 10146 5795 10169 5798 1 vdd
rlabel space 10114 5537 10143 5546 1 gnd
rlabel locali 10008 5519 10037 5525 1 gnd
rlabel locali 10011 5818 10040 5824 1 vdd
rlabel locali 9852 5216 9874 5233 1 d1
rlabel nwell 10047 5385 10070 5388 1 vdd
rlabel space 10015 5127 10044 5136 1 gnd
rlabel locali 9909 5109 9938 5115 1 gnd
rlabel locali 9912 5408 9941 5414 1 vdd
rlabel locali 9869 6234 9891 6251 1 d1
rlabel nwell 10064 6403 10087 6406 1 vdd
rlabel space 10032 6145 10061 6154 1 gnd
rlabel locali 9926 6127 9955 6133 1 gnd
rlabel locali 9929 6426 9958 6432 1 vdd
rlabel nwell 9250 5157 9273 5160 1 vdd
rlabel space 9218 4899 9247 4908 1 gnd
rlabel locali 9112 4881 9141 4887 1 gnd
rlabel locali 9115 5180 9144 5186 1 vdd
rlabel locali 9061 4992 9083 5007 1 d0
rlabel nwell 9249 5569 9272 5572 1 vdd
rlabel space 9217 5311 9246 5320 1 gnd
rlabel locali 9111 5293 9140 5299 1 gnd
rlabel locali 9114 5592 9143 5598 1 vdd
rlabel locali 9060 5404 9082 5419 1 d0
rlabel nwell 9267 6175 9290 6178 1 vdd
rlabel space 9235 5917 9264 5926 1 gnd
rlabel locali 9129 5899 9158 5905 1 gnd
rlabel locali 9132 6198 9161 6204 1 vdd
rlabel locali 9078 6010 9100 6025 1 d0
rlabel nwell 9266 6587 9289 6590 1 vdd
rlabel space 9234 6329 9263 6338 1 gnd
rlabel locali 9128 6311 9157 6317 1 gnd
rlabel locali 9131 6610 9160 6616 1 vdd
rlabel locali 9077 6422 9099 6437 1 d0
rlabel locali 9990 7662 10010 7686 1 d2
rlabel nwell 10183 7831 10206 7834 1 vdd
rlabel space 10151 7573 10180 7582 1 gnd
rlabel locali 10045 7555 10074 7561 1 gnd
rlabel locali 10048 7854 10077 7860 1 vdd
rlabel locali 9889 7252 9911 7269 1 d1
rlabel nwell 10084 7421 10107 7424 1 vdd
rlabel space 10052 7163 10081 7172 1 gnd
rlabel locali 9946 7145 9975 7151 1 gnd
rlabel locali 9949 7444 9978 7450 1 vdd
rlabel locali 9906 8270 9928 8287 1 d1
rlabel nwell 10101 8439 10124 8442 1 vdd
rlabel space 10069 8181 10098 8190 1 gnd
rlabel locali 9963 8163 9992 8169 1 gnd
rlabel locali 9966 8462 9995 8468 1 vdd
rlabel nwell 9287 7193 9310 7196 1 vdd
rlabel space 9255 6935 9284 6944 1 gnd
rlabel locali 9149 6917 9178 6923 1 gnd
rlabel locali 9152 7216 9181 7222 1 vdd
rlabel locali 9098 7028 9120 7043 1 d0
rlabel nwell 9286 7605 9309 7608 1 vdd
rlabel space 9254 7347 9283 7356 1 gnd
rlabel locali 9148 7329 9177 7335 1 gnd
rlabel locali 9151 7628 9180 7634 1 vdd
rlabel locali 9097 7440 9119 7455 1 d0
rlabel nwell 9304 8211 9327 8214 1 vdd
rlabel space 9272 7953 9301 7962 1 gnd
rlabel locali 9166 7935 9195 7941 1 gnd
rlabel locali 9169 8234 9198 8240 1 vdd
rlabel locali 9115 8046 9137 8061 1 d0
rlabel nwell 9303 8623 9326 8626 1 vdd
rlabel space 9271 8365 9300 8374 1 gnd
rlabel locali 9165 8347 9194 8353 1 gnd
rlabel locali 9168 8646 9197 8652 1 vdd
rlabel locali 9114 8458 9136 8473 1 d0
rlabel locali 8451 457 8480 463 1 vdd
rlabel locali 8448 158 8477 164 1 gnd
rlabel space 8554 176 8583 185 1 gnd
rlabel nwell 8586 434 8609 437 1 vdd
rlabel locali 8390 270 8412 285 1 d7
rlabel locali 21310 255 21333 271 1 d6
rlabel locali 21374 445 21403 451 1 vdd
rlabel locali 21371 146 21400 152 1 gnd
rlabel space 21477 164 21506 173 1 gnd
rlabel nwell 21509 422 21532 425 1 vdd
rlabel locali 23191 345 23206 358 1 d5
rlabel locali 23249 532 23278 538 1 vdd
rlabel locali 23246 233 23275 239 1 gnd
rlabel space 23352 251 23381 260 1 gnd
rlabel nwell 23384 509 23407 512 1 vdd
rlabel locali 25673 1265 25695 1280 5 d0
rlabel locali 25612 1086 25641 1092 5 vdd
rlabel locali 25615 1385 25644 1391 5 gnd
rlabel space 25509 1364 25538 1373 5 gnd
rlabel nwell 25483 1112 25506 1115 5 vdd
rlabel locali 25672 1677 25694 1692 5 d0
rlabel locali 25611 1498 25640 1504 5 vdd
rlabel locali 25614 1797 25643 1803 5 gnd
rlabel space 25508 1776 25537 1785 5 gnd
rlabel nwell 25482 1524 25505 1527 5 vdd
rlabel locali 25690 2283 25712 2298 5 d0
rlabel locali 25629 2104 25658 2110 5 vdd
rlabel locali 25632 2403 25661 2409 5 gnd
rlabel space 25526 2382 25555 2391 5 gnd
rlabel nwell 25500 2130 25523 2133 5 vdd
rlabel locali 25689 2695 25711 2710 5 d0
rlabel locali 25628 2516 25657 2522 5 vdd
rlabel locali 25631 2815 25660 2821 5 gnd
rlabel space 25525 2794 25554 2803 5 gnd
rlabel nwell 25499 2542 25522 2545 5 vdd
rlabel locali 24814 1270 24843 1276 5 vdd
rlabel locali 24817 1569 24846 1575 5 gnd
rlabel space 24711 1548 24740 1557 5 gnd
rlabel nwell 24685 1296 24708 1299 5 vdd
rlabel locali 24881 1451 24903 1468 5 d1
rlabel locali 24831 2288 24860 2294 5 vdd
rlabel locali 24834 2587 24863 2593 5 gnd
rlabel space 24728 2566 24757 2575 5 gnd
rlabel nwell 24702 2314 24725 2317 5 vdd
rlabel locali 24898 2469 24920 2486 5 d1
rlabel locali 24732 1878 24761 1884 5 vdd
rlabel locali 24735 2177 24764 2183 5 gnd
rlabel space 24629 2156 24658 2165 5 gnd
rlabel nwell 24603 1904 24626 1907 5 vdd
rlabel locali 24799 2052 24819 2076 5 d2
rlabel locali 25710 3301 25732 3316 5 d0
rlabel locali 25649 3122 25678 3128 5 vdd
rlabel locali 25652 3421 25681 3427 5 gnd
rlabel space 25546 3400 25575 3409 5 gnd
rlabel nwell 25520 3148 25543 3151 5 vdd
rlabel locali 25709 3713 25731 3728 5 d0
rlabel locali 25648 3534 25677 3540 5 vdd
rlabel locali 25651 3833 25680 3839 5 gnd
rlabel space 25545 3812 25574 3821 5 gnd
rlabel nwell 25519 3560 25542 3563 5 vdd
rlabel locali 25727 4319 25749 4334 5 d0
rlabel locali 25666 4140 25695 4146 5 vdd
rlabel locali 25669 4439 25698 4445 5 gnd
rlabel space 25563 4418 25592 4427 5 gnd
rlabel nwell 25537 4166 25560 4169 5 vdd
rlabel locali 25726 4731 25748 4746 5 d0
rlabel locali 25665 4552 25694 4558 5 vdd
rlabel locali 25668 4851 25697 4857 5 gnd
rlabel space 25562 4830 25591 4839 5 gnd
rlabel nwell 25536 4578 25559 4581 5 vdd
rlabel locali 24851 3306 24880 3312 5 vdd
rlabel locali 24854 3605 24883 3611 5 gnd
rlabel space 24748 3584 24777 3593 5 gnd
rlabel nwell 24722 3332 24745 3335 5 vdd
rlabel locali 24918 3487 24940 3504 5 d1
rlabel locali 24868 4324 24897 4330 5 vdd
rlabel locali 24871 4623 24900 4629 5 gnd
rlabel space 24765 4602 24794 4611 5 gnd
rlabel nwell 24739 4350 24762 4353 5 vdd
rlabel locali 24935 4505 24957 4522 5 d1
rlabel locali 24769 3914 24798 3920 5 vdd
rlabel locali 24772 4213 24801 4219 5 gnd
rlabel space 24666 4192 24695 4201 5 gnd
rlabel nwell 24640 3940 24663 3943 5 vdd
rlabel locali 24836 4088 24856 4112 5 d2
rlabel locali 24686 2898 24715 2904 5 vdd
rlabel locali 24689 3197 24718 3203 5 gnd
rlabel space 24583 3176 24612 3185 5 gnd
rlabel nwell 24557 2924 24580 2927 5 vdd
rlabel locali 24751 3077 24771 3090 5 d3
rlabel locali 25746 5337 25768 5352 5 d0
rlabel locali 25685 5158 25714 5164 5 vdd
rlabel locali 25688 5457 25717 5463 5 gnd
rlabel space 25582 5436 25611 5445 5 gnd
rlabel nwell 25556 5184 25579 5187 5 vdd
rlabel locali 25745 5749 25767 5764 5 d0
rlabel locali 25684 5570 25713 5576 5 vdd
rlabel locali 25687 5869 25716 5875 5 gnd
rlabel space 25581 5848 25610 5857 5 gnd
rlabel nwell 25555 5596 25578 5599 5 vdd
rlabel locali 25763 6355 25785 6370 5 d0
rlabel locali 25702 6176 25731 6182 5 vdd
rlabel locali 25705 6475 25734 6481 5 gnd
rlabel space 25599 6454 25628 6463 5 gnd
rlabel nwell 25573 6202 25596 6205 5 vdd
rlabel locali 25762 6767 25784 6782 5 d0
rlabel locali 25701 6588 25730 6594 5 vdd
rlabel locali 25704 6887 25733 6893 5 gnd
rlabel space 25598 6866 25627 6875 5 gnd
rlabel nwell 25572 6614 25595 6617 5 vdd
rlabel locali 24887 5342 24916 5348 5 vdd
rlabel locali 24890 5641 24919 5647 5 gnd
rlabel space 24784 5620 24813 5629 5 gnd
rlabel nwell 24758 5368 24781 5371 5 vdd
rlabel locali 24954 5523 24976 5540 5 d1
rlabel locali 24904 6360 24933 6366 5 vdd
rlabel locali 24907 6659 24936 6665 5 gnd
rlabel space 24801 6638 24830 6647 5 gnd
rlabel nwell 24775 6386 24798 6389 5 vdd
rlabel locali 24971 6541 24993 6558 5 d1
rlabel locali 24805 5950 24834 5956 5 vdd
rlabel locali 24808 6249 24837 6255 5 gnd
rlabel space 24702 6228 24731 6237 5 gnd
rlabel nwell 24676 5976 24699 5979 5 vdd
rlabel locali 24872 6124 24892 6148 5 d2
rlabel locali 25783 7373 25805 7388 5 d0
rlabel locali 25722 7194 25751 7200 5 vdd
rlabel locali 25725 7493 25754 7499 5 gnd
rlabel space 25619 7472 25648 7481 5 gnd
rlabel nwell 25593 7220 25616 7223 5 vdd
rlabel locali 25782 7785 25804 7800 5 d0
rlabel locali 25721 7606 25750 7612 5 vdd
rlabel locali 25724 7905 25753 7911 5 gnd
rlabel space 25618 7884 25647 7893 5 gnd
rlabel nwell 25592 7632 25615 7635 5 vdd
rlabel locali 25800 8391 25822 8406 5 d0
rlabel locali 25739 8212 25768 8218 5 vdd
rlabel locali 25742 8511 25771 8517 5 gnd
rlabel space 25636 8490 25665 8499 5 gnd
rlabel nwell 25610 8238 25633 8241 5 vdd
rlabel locali 25799 8803 25821 8818 5 d0
rlabel locali 25738 8624 25767 8630 5 vdd
rlabel locali 25741 8923 25770 8929 5 gnd
rlabel space 25635 8902 25664 8911 5 gnd
rlabel nwell 25609 8650 25632 8653 5 vdd
rlabel locali 24924 7378 24953 7384 5 vdd
rlabel locali 24927 7677 24956 7683 5 gnd
rlabel space 24821 7656 24850 7665 5 gnd
rlabel nwell 24795 7404 24818 7407 5 vdd
rlabel locali 24991 7559 25013 7576 5 d1
rlabel locali 24941 8396 24970 8402 5 vdd
rlabel locali 24944 8695 24973 8701 5 gnd
rlabel space 24838 8674 24867 8683 5 gnd
rlabel nwell 24812 8422 24835 8425 5 vdd
rlabel locali 25008 8577 25030 8594 5 d1
rlabel locali 24842 7986 24871 7992 5 vdd
rlabel locali 24845 8285 24874 8291 5 gnd
rlabel space 24739 8264 24768 8273 5 gnd
rlabel nwell 24713 8012 24736 8015 5 vdd
rlabel locali 24909 8160 24929 8184 5 d2
rlabel locali 24759 6970 24788 6976 5 vdd
rlabel locali 24762 7269 24791 7275 5 gnd
rlabel space 24656 7248 24685 7257 5 gnd
rlabel nwell 24630 6996 24653 6999 5 vdd
rlabel locali 24824 7149 24844 7162 5 d3
rlabel locali 24583 4936 24612 4942 5 vdd
rlabel locali 24586 5235 24615 5241 5 gnd
rlabel space 24480 5214 24509 5223 5 gnd
rlabel nwell 24454 4962 24477 4965 5 vdd
rlabel locali 24647 5115 24666 5132 5 d4
rlabel locali 23137 4606 23156 4623 1 d4
rlabel nwell 23326 4773 23349 4776 1 vdd
rlabel space 23294 4515 23323 4524 1 gnd
rlabel locali 23188 4497 23217 4503 1 gnd
rlabel locali 23191 4796 23220 4802 1 vdd
rlabel locali 22959 2576 22979 2589 1 d3
rlabel nwell 23150 2739 23173 2742 1 vdd
rlabel space 23118 2481 23147 2490 1 gnd
rlabel locali 23012 2463 23041 2469 1 gnd
rlabel locali 23015 2762 23044 2768 1 vdd
rlabel locali 22874 1554 22894 1578 1 d2
rlabel nwell 23067 1723 23090 1726 1 vdd
rlabel space 23035 1465 23064 1474 1 gnd
rlabel locali 22929 1447 22958 1453 1 gnd
rlabel locali 22932 1746 22961 1752 1 vdd
rlabel locali 22773 1144 22795 1161 1 d1
rlabel nwell 22968 1313 22991 1316 1 vdd
rlabel space 22936 1055 22965 1064 1 gnd
rlabel locali 22830 1037 22859 1043 1 gnd
rlabel locali 22833 1336 22862 1342 1 vdd
rlabel locali 22790 2162 22812 2179 1 d1
rlabel nwell 22985 2331 23008 2334 1 vdd
rlabel space 22953 2073 22982 2082 1 gnd
rlabel locali 22847 2055 22876 2061 1 gnd
rlabel locali 22850 2354 22879 2360 1 vdd
rlabel nwell 22171 1085 22194 1088 1 vdd
rlabel space 22139 827 22168 836 1 gnd
rlabel locali 22033 809 22062 815 1 gnd
rlabel locali 22036 1108 22065 1114 1 vdd
rlabel locali 21982 920 22004 935 1 d0
rlabel nwell 22170 1497 22193 1500 1 vdd
rlabel space 22138 1239 22167 1248 1 gnd
rlabel locali 22032 1221 22061 1227 1 gnd
rlabel locali 22035 1520 22064 1526 1 vdd
rlabel locali 21981 1332 22003 1347 1 d0
rlabel nwell 22188 2103 22211 2106 1 vdd
rlabel space 22156 1845 22185 1854 1 gnd
rlabel locali 22050 1827 22079 1833 1 gnd
rlabel locali 22053 2126 22082 2132 1 vdd
rlabel locali 21999 1938 22021 1953 1 d0
rlabel nwell 22187 2515 22210 2518 1 vdd
rlabel space 22155 2257 22184 2266 1 gnd
rlabel locali 22049 2239 22078 2245 1 gnd
rlabel locali 22052 2538 22081 2544 1 vdd
rlabel locali 21998 2350 22020 2365 1 d0
rlabel locali 22911 3590 22931 3614 1 d2
rlabel nwell 23104 3759 23127 3762 1 vdd
rlabel space 23072 3501 23101 3510 1 gnd
rlabel locali 22966 3483 22995 3489 1 gnd
rlabel locali 22969 3782 22998 3788 1 vdd
rlabel locali 22810 3180 22832 3197 1 d1
rlabel nwell 23005 3349 23028 3352 1 vdd
rlabel space 22973 3091 23002 3100 1 gnd
rlabel locali 22867 3073 22896 3079 1 gnd
rlabel locali 22870 3372 22899 3378 1 vdd
rlabel locali 22827 4198 22849 4215 1 d1
rlabel nwell 23022 4367 23045 4370 1 vdd
rlabel space 22990 4109 23019 4118 1 gnd
rlabel locali 22884 4091 22913 4097 1 gnd
rlabel locali 22887 4390 22916 4396 1 vdd
rlabel nwell 22208 3121 22231 3124 1 vdd
rlabel space 22176 2863 22205 2872 1 gnd
rlabel locali 22070 2845 22099 2851 1 gnd
rlabel locali 22073 3144 22102 3150 1 vdd
rlabel locali 22019 2956 22041 2971 1 d0
rlabel nwell 22207 3533 22230 3536 1 vdd
rlabel space 22175 3275 22204 3284 1 gnd
rlabel locali 22069 3257 22098 3263 1 gnd
rlabel locali 22072 3556 22101 3562 1 vdd
rlabel locali 22018 3368 22040 3383 1 d0
rlabel nwell 22225 4139 22248 4142 1 vdd
rlabel space 22193 3881 22222 3890 1 gnd
rlabel locali 22087 3863 22116 3869 1 gnd
rlabel locali 22090 4162 22119 4168 1 vdd
rlabel locali 22036 3974 22058 3989 1 d0
rlabel nwell 22224 4551 22247 4554 1 vdd
rlabel space 22192 4293 22221 4302 1 gnd
rlabel locali 22086 4275 22115 4281 1 gnd
rlabel locali 22089 4574 22118 4580 1 vdd
rlabel locali 22035 4386 22057 4401 1 d0
rlabel locali 23032 6648 23052 6661 1 d3
rlabel nwell 23223 6811 23246 6814 1 vdd
rlabel space 23191 6553 23220 6562 1 gnd
rlabel locali 23085 6535 23114 6541 1 gnd
rlabel locali 23088 6834 23117 6840 1 vdd
rlabel locali 22947 5626 22967 5650 1 d2
rlabel nwell 23140 5795 23163 5798 1 vdd
rlabel space 23108 5537 23137 5546 1 gnd
rlabel locali 23002 5519 23031 5525 1 gnd
rlabel locali 23005 5818 23034 5824 1 vdd
rlabel locali 22846 5216 22868 5233 1 d1
rlabel nwell 23041 5385 23064 5388 1 vdd
rlabel space 23009 5127 23038 5136 1 gnd
rlabel locali 22903 5109 22932 5115 1 gnd
rlabel locali 22906 5408 22935 5414 1 vdd
rlabel locali 22863 6234 22885 6251 1 d1
rlabel nwell 23058 6403 23081 6406 1 vdd
rlabel space 23026 6145 23055 6154 1 gnd
rlabel locali 22920 6127 22949 6133 1 gnd
rlabel locali 22923 6426 22952 6432 1 vdd
rlabel nwell 22244 5157 22267 5160 1 vdd
rlabel space 22212 4899 22241 4908 1 gnd
rlabel locali 22106 4881 22135 4887 1 gnd
rlabel locali 22109 5180 22138 5186 1 vdd
rlabel locali 22055 4992 22077 5007 1 d0
rlabel nwell 22243 5569 22266 5572 1 vdd
rlabel space 22211 5311 22240 5320 1 gnd
rlabel locali 22105 5293 22134 5299 1 gnd
rlabel locali 22108 5592 22137 5598 1 vdd
rlabel locali 22054 5404 22076 5419 1 d0
rlabel nwell 22261 6175 22284 6178 1 vdd
rlabel space 22229 5917 22258 5926 1 gnd
rlabel locali 22123 5899 22152 5905 1 gnd
rlabel locali 22126 6198 22155 6204 1 vdd
rlabel locali 22072 6010 22094 6025 1 d0
rlabel nwell 22260 6587 22283 6590 1 vdd
rlabel space 22228 6329 22257 6338 1 gnd
rlabel locali 22122 6311 22151 6317 1 gnd
rlabel locali 22125 6610 22154 6616 1 vdd
rlabel locali 22071 6422 22093 6437 1 d0
rlabel locali 22984 7662 23004 7686 1 d2
rlabel nwell 23177 7831 23200 7834 1 vdd
rlabel space 23145 7573 23174 7582 1 gnd
rlabel locali 23039 7555 23068 7561 1 gnd
rlabel locali 23042 7854 23071 7860 1 vdd
rlabel locali 22883 7252 22905 7269 1 d1
rlabel nwell 23078 7421 23101 7424 1 vdd
rlabel space 23046 7163 23075 7172 1 gnd
rlabel locali 22940 7145 22969 7151 1 gnd
rlabel locali 22943 7444 22972 7450 1 vdd
rlabel locali 22900 8270 22922 8287 1 d1
rlabel nwell 23095 8439 23118 8442 1 vdd
rlabel space 23063 8181 23092 8190 1 gnd
rlabel locali 22957 8163 22986 8169 1 gnd
rlabel locali 22960 8462 22989 8468 1 vdd
rlabel nwell 22281 7193 22304 7196 1 vdd
rlabel space 22249 6935 22278 6944 1 gnd
rlabel locali 22143 6917 22172 6923 1 gnd
rlabel locali 22146 7216 22175 7222 1 vdd
rlabel locali 22092 7028 22114 7043 1 d0
rlabel nwell 22280 7605 22303 7608 1 vdd
rlabel space 22248 7347 22277 7356 1 gnd
rlabel locali 22142 7329 22171 7335 1 gnd
rlabel locali 22145 7628 22174 7634 1 vdd
rlabel locali 22091 7440 22113 7455 1 d0
rlabel nwell 22298 8211 22321 8214 1 vdd
rlabel space 22266 7953 22295 7962 1 gnd
rlabel locali 22160 7935 22189 7941 1 gnd
rlabel locali 22163 8234 22192 8240 1 vdd
rlabel locali 22109 8046 22131 8061 1 d0
rlabel nwell 22297 8623 22320 8626 1 vdd
rlabel space 22265 8365 22294 8374 1 gnd
rlabel locali 22159 8347 22188 8353 1 gnd
rlabel locali 22162 8646 22191 8652 1 vdd
rlabel locali 22108 8458 22130 8473 1 d0
rlabel locali 18827 332 18842 345 1 d5
rlabel locali 18885 519 18914 525 1 vdd
rlabel locali 18882 220 18911 226 1 gnd
rlabel space 18988 238 19017 247 1 gnd
rlabel nwell 19020 496 19043 499 1 vdd
rlabel locali 21309 1252 21331 1267 5 d0
rlabel locali 21248 1073 21277 1079 5 vdd
rlabel locali 21251 1372 21280 1378 5 gnd
rlabel space 21145 1351 21174 1360 5 gnd
rlabel nwell 21119 1099 21142 1102 5 vdd
rlabel locali 21308 1664 21330 1679 5 d0
rlabel locali 21247 1485 21276 1491 5 vdd
rlabel locali 21250 1784 21279 1790 5 gnd
rlabel space 21144 1763 21173 1772 5 gnd
rlabel nwell 21118 1511 21141 1514 5 vdd
rlabel locali 21326 2270 21348 2285 5 d0
rlabel locali 21265 2091 21294 2097 5 vdd
rlabel locali 21268 2390 21297 2396 5 gnd
rlabel space 21162 2369 21191 2378 5 gnd
rlabel nwell 21136 2117 21159 2120 5 vdd
rlabel locali 21325 2682 21347 2697 5 d0
rlabel locali 21264 2503 21293 2509 5 vdd
rlabel locali 21267 2802 21296 2808 5 gnd
rlabel space 21161 2781 21190 2790 5 gnd
rlabel nwell 21135 2529 21158 2532 5 vdd
rlabel locali 20450 1257 20479 1263 5 vdd
rlabel locali 20453 1556 20482 1562 5 gnd
rlabel space 20347 1535 20376 1544 5 gnd
rlabel nwell 20321 1283 20344 1286 5 vdd
rlabel locali 20517 1438 20539 1455 5 d1
rlabel locali 20467 2275 20496 2281 5 vdd
rlabel locali 20470 2574 20499 2580 5 gnd
rlabel space 20364 2553 20393 2562 5 gnd
rlabel nwell 20338 2301 20361 2304 5 vdd
rlabel locali 20534 2456 20556 2473 5 d1
rlabel locali 20368 1865 20397 1871 5 vdd
rlabel locali 20371 2164 20400 2170 5 gnd
rlabel space 20265 2143 20294 2152 5 gnd
rlabel nwell 20239 1891 20262 1894 5 vdd
rlabel locali 20435 2039 20455 2063 5 d2
rlabel locali 21346 3288 21368 3303 5 d0
rlabel locali 21285 3109 21314 3115 5 vdd
rlabel locali 21288 3408 21317 3414 5 gnd
rlabel space 21182 3387 21211 3396 5 gnd
rlabel nwell 21156 3135 21179 3138 5 vdd
rlabel locali 21345 3700 21367 3715 5 d0
rlabel locali 21284 3521 21313 3527 5 vdd
rlabel locali 21287 3820 21316 3826 5 gnd
rlabel space 21181 3799 21210 3808 5 gnd
rlabel nwell 21155 3547 21178 3550 5 vdd
rlabel locali 21363 4306 21385 4321 5 d0
rlabel locali 21302 4127 21331 4133 5 vdd
rlabel locali 21305 4426 21334 4432 5 gnd
rlabel space 21199 4405 21228 4414 5 gnd
rlabel nwell 21173 4153 21196 4156 5 vdd
rlabel locali 21362 4718 21384 4733 5 d0
rlabel locali 21301 4539 21330 4545 5 vdd
rlabel locali 21304 4838 21333 4844 5 gnd
rlabel space 21198 4817 21227 4826 5 gnd
rlabel nwell 21172 4565 21195 4568 5 vdd
rlabel locali 20487 3293 20516 3299 5 vdd
rlabel locali 20490 3592 20519 3598 5 gnd
rlabel space 20384 3571 20413 3580 5 gnd
rlabel nwell 20358 3319 20381 3322 5 vdd
rlabel locali 20554 3474 20576 3491 5 d1
rlabel locali 20504 4311 20533 4317 5 vdd
rlabel locali 20507 4610 20536 4616 5 gnd
rlabel space 20401 4589 20430 4598 5 gnd
rlabel nwell 20375 4337 20398 4340 5 vdd
rlabel locali 20571 4492 20593 4509 5 d1
rlabel locali 20405 3901 20434 3907 5 vdd
rlabel locali 20408 4200 20437 4206 5 gnd
rlabel space 20302 4179 20331 4188 5 gnd
rlabel nwell 20276 3927 20299 3930 5 vdd
rlabel locali 20472 4075 20492 4099 5 d2
rlabel locali 20322 2885 20351 2891 5 vdd
rlabel locali 20325 3184 20354 3190 5 gnd
rlabel space 20219 3163 20248 3172 5 gnd
rlabel nwell 20193 2911 20216 2914 5 vdd
rlabel locali 20387 3064 20407 3077 5 d3
rlabel locali 21382 5324 21404 5339 5 d0
rlabel locali 21321 5145 21350 5151 5 vdd
rlabel locali 21324 5444 21353 5450 5 gnd
rlabel space 21218 5423 21247 5432 5 gnd
rlabel nwell 21192 5171 21215 5174 5 vdd
rlabel locali 21381 5736 21403 5751 5 d0
rlabel locali 21320 5557 21349 5563 5 vdd
rlabel locali 21323 5856 21352 5862 5 gnd
rlabel space 21217 5835 21246 5844 5 gnd
rlabel nwell 21191 5583 21214 5586 5 vdd
rlabel locali 21399 6342 21421 6357 5 d0
rlabel locali 21338 6163 21367 6169 5 vdd
rlabel locali 21341 6462 21370 6468 5 gnd
rlabel space 21235 6441 21264 6450 5 gnd
rlabel nwell 21209 6189 21232 6192 5 vdd
rlabel locali 21398 6754 21420 6769 5 d0
rlabel locali 21337 6575 21366 6581 5 vdd
rlabel locali 21340 6874 21369 6880 5 gnd
rlabel space 21234 6853 21263 6862 5 gnd
rlabel nwell 21208 6601 21231 6604 5 vdd
rlabel locali 20523 5329 20552 5335 5 vdd
rlabel locali 20526 5628 20555 5634 5 gnd
rlabel space 20420 5607 20449 5616 5 gnd
rlabel nwell 20394 5355 20417 5358 5 vdd
rlabel locali 20590 5510 20612 5527 5 d1
rlabel locali 20540 6347 20569 6353 5 vdd
rlabel locali 20543 6646 20572 6652 5 gnd
rlabel space 20437 6625 20466 6634 5 gnd
rlabel nwell 20411 6373 20434 6376 5 vdd
rlabel locali 20607 6528 20629 6545 5 d1
rlabel locali 20441 5937 20470 5943 5 vdd
rlabel locali 20444 6236 20473 6242 5 gnd
rlabel space 20338 6215 20367 6224 5 gnd
rlabel nwell 20312 5963 20335 5966 5 vdd
rlabel locali 20508 6111 20528 6135 5 d2
rlabel locali 21419 7360 21441 7375 5 d0
rlabel locali 21358 7181 21387 7187 5 vdd
rlabel locali 21361 7480 21390 7486 5 gnd
rlabel space 21255 7459 21284 7468 5 gnd
rlabel nwell 21229 7207 21252 7210 5 vdd
rlabel locali 21418 7772 21440 7787 5 d0
rlabel locali 21357 7593 21386 7599 5 vdd
rlabel locali 21360 7892 21389 7898 5 gnd
rlabel space 21254 7871 21283 7880 5 gnd
rlabel nwell 21228 7619 21251 7622 5 vdd
rlabel locali 21436 8378 21458 8393 5 d0
rlabel locali 21375 8199 21404 8205 5 vdd
rlabel locali 21378 8498 21407 8504 5 gnd
rlabel space 21272 8477 21301 8486 5 gnd
rlabel nwell 21246 8225 21269 8228 5 vdd
rlabel locali 21435 8790 21457 8805 5 d0
rlabel locali 21374 8611 21403 8617 5 vdd
rlabel locali 21377 8910 21406 8916 5 gnd
rlabel space 21271 8889 21300 8898 5 gnd
rlabel nwell 21245 8637 21268 8640 5 vdd
rlabel locali 20560 7365 20589 7371 5 vdd
rlabel locali 20563 7664 20592 7670 5 gnd
rlabel space 20457 7643 20486 7652 5 gnd
rlabel nwell 20431 7391 20454 7394 5 vdd
rlabel locali 20627 7546 20649 7563 5 d1
rlabel locali 20577 8383 20606 8389 5 vdd
rlabel locali 20580 8682 20609 8688 5 gnd
rlabel space 20474 8661 20503 8670 5 gnd
rlabel nwell 20448 8409 20471 8412 5 vdd
rlabel locali 20644 8564 20666 8581 5 d1
rlabel locali 20478 7973 20507 7979 5 vdd
rlabel locali 20481 8272 20510 8278 5 gnd
rlabel space 20375 8251 20404 8260 5 gnd
rlabel nwell 20349 7999 20372 8002 5 vdd
rlabel locali 20545 8147 20565 8171 5 d2
rlabel locali 20395 6957 20424 6963 5 vdd
rlabel locali 20398 7256 20427 7262 5 gnd
rlabel space 20292 7235 20321 7244 5 gnd
rlabel nwell 20266 6983 20289 6986 5 vdd
rlabel locali 20460 7136 20480 7149 5 d3
rlabel locali 20219 4923 20248 4929 5 vdd
rlabel locali 20222 5222 20251 5228 5 gnd
rlabel space 20116 5201 20145 5210 5 gnd
rlabel nwell 20090 4949 20113 4952 5 vdd
rlabel locali 20283 5102 20302 5119 5 d4
rlabel locali 18773 4593 18792 4610 1 d4
rlabel nwell 18962 4760 18985 4763 1 vdd
rlabel space 18930 4502 18959 4511 1 gnd
rlabel locali 18824 4484 18853 4490 1 gnd
rlabel locali 18827 4783 18856 4789 1 vdd
rlabel locali 18595 2563 18615 2576 1 d3
rlabel nwell 18786 2726 18809 2729 1 vdd
rlabel space 18754 2468 18783 2477 1 gnd
rlabel locali 18648 2450 18677 2456 1 gnd
rlabel locali 18651 2749 18680 2755 1 vdd
rlabel locali 18510 1541 18530 1565 1 d2
rlabel nwell 18703 1710 18726 1713 1 vdd
rlabel space 18671 1452 18700 1461 1 gnd
rlabel locali 18565 1434 18594 1440 1 gnd
rlabel locali 18568 1733 18597 1739 1 vdd
rlabel locali 18409 1131 18431 1148 1 d1
rlabel nwell 18604 1300 18627 1303 1 vdd
rlabel space 18572 1042 18601 1051 1 gnd
rlabel locali 18466 1024 18495 1030 1 gnd
rlabel locali 18469 1323 18498 1329 1 vdd
rlabel locali 18426 2149 18448 2166 1 d1
rlabel nwell 18621 2318 18644 2321 1 vdd
rlabel space 18589 2060 18618 2069 1 gnd
rlabel locali 18483 2042 18512 2048 1 gnd
rlabel locali 18486 2341 18515 2347 1 vdd
rlabel nwell 17807 1072 17830 1075 1 vdd
rlabel space 17775 814 17804 823 1 gnd
rlabel locali 17669 796 17698 802 1 gnd
rlabel locali 17672 1095 17701 1101 1 vdd
rlabel locali 17618 907 17640 922 1 d0
rlabel nwell 17806 1484 17829 1487 1 vdd
rlabel space 17774 1226 17803 1235 1 gnd
rlabel locali 17668 1208 17697 1214 1 gnd
rlabel locali 17671 1507 17700 1513 1 vdd
rlabel locali 17617 1319 17639 1334 1 d0
rlabel nwell 17824 2090 17847 2093 1 vdd
rlabel space 17792 1832 17821 1841 1 gnd
rlabel locali 17686 1814 17715 1820 1 gnd
rlabel locali 17689 2113 17718 2119 1 vdd
rlabel locali 17635 1925 17657 1940 1 d0
rlabel nwell 17823 2502 17846 2505 1 vdd
rlabel space 17791 2244 17820 2253 1 gnd
rlabel locali 17685 2226 17714 2232 1 gnd
rlabel locali 17688 2525 17717 2531 1 vdd
rlabel locali 17634 2337 17656 2352 1 d0
rlabel locali 18547 3577 18567 3601 1 d2
rlabel nwell 18740 3746 18763 3749 1 vdd
rlabel space 18708 3488 18737 3497 1 gnd
rlabel locali 18602 3470 18631 3476 1 gnd
rlabel locali 18605 3769 18634 3775 1 vdd
rlabel locali 18446 3167 18468 3184 1 d1
rlabel nwell 18641 3336 18664 3339 1 vdd
rlabel space 18609 3078 18638 3087 1 gnd
rlabel locali 18503 3060 18532 3066 1 gnd
rlabel locali 18506 3359 18535 3365 1 vdd
rlabel locali 18463 4185 18485 4202 1 d1
rlabel nwell 18658 4354 18681 4357 1 vdd
rlabel space 18626 4096 18655 4105 1 gnd
rlabel locali 18520 4078 18549 4084 1 gnd
rlabel locali 18523 4377 18552 4383 1 vdd
rlabel nwell 17844 3108 17867 3111 1 vdd
rlabel space 17812 2850 17841 2859 1 gnd
rlabel locali 17706 2832 17735 2838 1 gnd
rlabel locali 17709 3131 17738 3137 1 vdd
rlabel locali 17655 2943 17677 2958 1 d0
rlabel nwell 17843 3520 17866 3523 1 vdd
rlabel space 17811 3262 17840 3271 1 gnd
rlabel locali 17705 3244 17734 3250 1 gnd
rlabel locali 17708 3543 17737 3549 1 vdd
rlabel locali 17654 3355 17676 3370 1 d0
rlabel nwell 17861 4126 17884 4129 1 vdd
rlabel space 17829 3868 17858 3877 1 gnd
rlabel locali 17723 3850 17752 3856 1 gnd
rlabel locali 17726 4149 17755 4155 1 vdd
rlabel locali 17672 3961 17694 3976 1 d0
rlabel nwell 17860 4538 17883 4541 1 vdd
rlabel space 17828 4280 17857 4289 1 gnd
rlabel locali 17722 4262 17751 4268 1 gnd
rlabel locali 17725 4561 17754 4567 1 vdd
rlabel locali 17671 4373 17693 4388 1 d0
rlabel locali 18668 6635 18688 6648 1 d3
rlabel nwell 18859 6798 18882 6801 1 vdd
rlabel space 18827 6540 18856 6549 1 gnd
rlabel locali 18721 6522 18750 6528 1 gnd
rlabel locali 18724 6821 18753 6827 1 vdd
rlabel locali 18583 5613 18603 5637 1 d2
rlabel nwell 18776 5782 18799 5785 1 vdd
rlabel space 18744 5524 18773 5533 1 gnd
rlabel locali 18638 5506 18667 5512 1 gnd
rlabel locali 18641 5805 18670 5811 1 vdd
rlabel locali 18482 5203 18504 5220 1 d1
rlabel nwell 18677 5372 18700 5375 1 vdd
rlabel space 18645 5114 18674 5123 1 gnd
rlabel locali 18539 5096 18568 5102 1 gnd
rlabel locali 18542 5395 18571 5401 1 vdd
rlabel locali 18499 6221 18521 6238 1 d1
rlabel nwell 18694 6390 18717 6393 1 vdd
rlabel space 18662 6132 18691 6141 1 gnd
rlabel locali 18556 6114 18585 6120 1 gnd
rlabel locali 18559 6413 18588 6419 1 vdd
rlabel nwell 17880 5144 17903 5147 1 vdd
rlabel space 17848 4886 17877 4895 1 gnd
rlabel locali 17742 4868 17771 4874 1 gnd
rlabel locali 17745 5167 17774 5173 1 vdd
rlabel locali 17691 4979 17713 4994 1 d0
rlabel nwell 17879 5556 17902 5559 1 vdd
rlabel space 17847 5298 17876 5307 1 gnd
rlabel locali 17741 5280 17770 5286 1 gnd
rlabel locali 17744 5579 17773 5585 1 vdd
rlabel locali 17690 5391 17712 5406 1 d0
rlabel nwell 17897 6162 17920 6165 1 vdd
rlabel space 17865 5904 17894 5913 1 gnd
rlabel locali 17759 5886 17788 5892 1 gnd
rlabel locali 17762 6185 17791 6191 1 vdd
rlabel locali 17708 5997 17730 6012 1 d0
rlabel nwell 17896 6574 17919 6577 1 vdd
rlabel space 17864 6316 17893 6325 1 gnd
rlabel locali 17758 6298 17787 6304 1 gnd
rlabel locali 17761 6597 17790 6603 1 vdd
rlabel locali 17707 6409 17729 6424 1 d0
rlabel locali 18620 7649 18640 7673 1 d2
rlabel nwell 18813 7818 18836 7821 1 vdd
rlabel space 18781 7560 18810 7569 1 gnd
rlabel locali 18675 7542 18704 7548 1 gnd
rlabel locali 18678 7841 18707 7847 1 vdd
rlabel locali 18519 7239 18541 7256 1 d1
rlabel nwell 18714 7408 18737 7411 1 vdd
rlabel space 18682 7150 18711 7159 1 gnd
rlabel locali 18576 7132 18605 7138 1 gnd
rlabel locali 18579 7431 18608 7437 1 vdd
rlabel locali 18536 8257 18558 8274 1 d1
rlabel nwell 18731 8426 18754 8429 1 vdd
rlabel space 18699 8168 18728 8177 1 gnd
rlabel locali 18593 8150 18622 8156 1 gnd
rlabel locali 18596 8449 18625 8455 1 vdd
rlabel nwell 17917 7180 17940 7183 1 vdd
rlabel space 17885 6922 17914 6931 1 gnd
rlabel locali 17779 6904 17808 6910 1 gnd
rlabel locali 17782 7203 17811 7209 1 vdd
rlabel locali 17728 7015 17750 7030 1 d0
rlabel nwell 17916 7592 17939 7595 1 vdd
rlabel space 17884 7334 17913 7343 1 gnd
rlabel locali 17778 7316 17807 7322 1 gnd
rlabel locali 17781 7615 17810 7621 1 vdd
rlabel locali 17727 7427 17749 7442 1 d0
rlabel nwell 17934 8198 17957 8201 1 vdd
rlabel space 17902 7940 17931 7949 1 gnd
rlabel locali 17796 7922 17825 7928 1 gnd
rlabel locali 17799 8221 17828 8227 1 vdd
rlabel locali 17745 8033 17767 8048 1 d0
rlabel nwell 17933 8610 17956 8613 1 vdd
rlabel space 17901 8352 17930 8361 1 gnd
rlabel locali 17795 8334 17824 8340 1 gnd
rlabel locali 17798 8633 17827 8639 1 vdd
rlabel locali 17744 8445 17766 8460 1 d0
rlabel locali 30051 280 30074 296 1 d6
rlabel locali 30115 470 30144 476 1 vdd
rlabel locali 30112 171 30141 177 1 gnd
rlabel space 30218 189 30247 198 1 gnd
rlabel nwell 30250 447 30273 450 1 vdd
rlabel locali 31932 370 31947 383 1 d5
rlabel locali 31990 557 32019 563 1 vdd
rlabel locali 31987 258 32016 264 1 gnd
rlabel space 32093 276 32122 285 1 gnd
rlabel nwell 32125 534 32148 537 1 vdd
rlabel locali 34414 1290 34436 1305 5 d0
rlabel locali 34353 1111 34382 1117 5 vdd
rlabel locali 34356 1410 34385 1416 5 gnd
rlabel space 34250 1389 34279 1398 5 gnd
rlabel nwell 34224 1137 34247 1140 5 vdd
rlabel locali 34413 1702 34435 1717 5 d0
rlabel locali 34352 1523 34381 1529 5 vdd
rlabel locali 34355 1822 34384 1828 5 gnd
rlabel space 34249 1801 34278 1810 5 gnd
rlabel nwell 34223 1549 34246 1552 5 vdd
rlabel locali 34431 2308 34453 2323 5 d0
rlabel locali 34370 2129 34399 2135 5 vdd
rlabel locali 34373 2428 34402 2434 5 gnd
rlabel space 34267 2407 34296 2416 5 gnd
rlabel nwell 34241 2155 34264 2158 5 vdd
rlabel locali 34430 2720 34452 2735 5 d0
rlabel locali 34369 2541 34398 2547 5 vdd
rlabel locali 34372 2840 34401 2846 5 gnd
rlabel space 34266 2819 34295 2828 5 gnd
rlabel nwell 34240 2567 34263 2570 5 vdd
rlabel locali 33555 1295 33584 1301 5 vdd
rlabel locali 33558 1594 33587 1600 5 gnd
rlabel space 33452 1573 33481 1582 5 gnd
rlabel nwell 33426 1321 33449 1324 5 vdd
rlabel locali 33622 1476 33644 1493 5 d1
rlabel locali 33572 2313 33601 2319 5 vdd
rlabel locali 33575 2612 33604 2618 5 gnd
rlabel space 33469 2591 33498 2600 5 gnd
rlabel nwell 33443 2339 33466 2342 5 vdd
rlabel locali 33639 2494 33661 2511 5 d1
rlabel locali 33473 1903 33502 1909 5 vdd
rlabel locali 33476 2202 33505 2208 5 gnd
rlabel space 33370 2181 33399 2190 5 gnd
rlabel nwell 33344 1929 33367 1932 5 vdd
rlabel locali 33540 2077 33560 2101 5 d2
rlabel locali 34451 3326 34473 3341 5 d0
rlabel locali 34390 3147 34419 3153 5 vdd
rlabel locali 34393 3446 34422 3452 5 gnd
rlabel space 34287 3425 34316 3434 5 gnd
rlabel nwell 34261 3173 34284 3176 5 vdd
rlabel locali 34450 3738 34472 3753 5 d0
rlabel locali 34389 3559 34418 3565 5 vdd
rlabel locali 34392 3858 34421 3864 5 gnd
rlabel space 34286 3837 34315 3846 5 gnd
rlabel nwell 34260 3585 34283 3588 5 vdd
rlabel locali 34468 4344 34490 4359 5 d0
rlabel locali 34407 4165 34436 4171 5 vdd
rlabel locali 34410 4464 34439 4470 5 gnd
rlabel space 34304 4443 34333 4452 5 gnd
rlabel nwell 34278 4191 34301 4194 5 vdd
rlabel locali 34467 4756 34489 4771 5 d0
rlabel locali 34406 4577 34435 4583 5 vdd
rlabel locali 34409 4876 34438 4882 5 gnd
rlabel space 34303 4855 34332 4864 5 gnd
rlabel nwell 34277 4603 34300 4606 5 vdd
rlabel locali 33592 3331 33621 3337 5 vdd
rlabel locali 33595 3630 33624 3636 5 gnd
rlabel space 33489 3609 33518 3618 5 gnd
rlabel nwell 33463 3357 33486 3360 5 vdd
rlabel locali 33659 3512 33681 3529 5 d1
rlabel locali 33609 4349 33638 4355 5 vdd
rlabel locali 33612 4648 33641 4654 5 gnd
rlabel space 33506 4627 33535 4636 5 gnd
rlabel nwell 33480 4375 33503 4378 5 vdd
rlabel locali 33676 4530 33698 4547 5 d1
rlabel locali 33510 3939 33539 3945 5 vdd
rlabel locali 33513 4238 33542 4244 5 gnd
rlabel space 33407 4217 33436 4226 5 gnd
rlabel nwell 33381 3965 33404 3968 5 vdd
rlabel locali 33577 4113 33597 4137 5 d2
rlabel locali 33427 2923 33456 2929 5 vdd
rlabel locali 33430 3222 33459 3228 5 gnd
rlabel space 33324 3201 33353 3210 5 gnd
rlabel nwell 33298 2949 33321 2952 5 vdd
rlabel locali 33492 3102 33512 3115 5 d3
rlabel locali 34487 5362 34509 5377 5 d0
rlabel locali 34426 5183 34455 5189 5 vdd
rlabel locali 34429 5482 34458 5488 5 gnd
rlabel space 34323 5461 34352 5470 5 gnd
rlabel nwell 34297 5209 34320 5212 5 vdd
rlabel locali 34486 5774 34508 5789 5 d0
rlabel locali 34425 5595 34454 5601 5 vdd
rlabel locali 34428 5894 34457 5900 5 gnd
rlabel space 34322 5873 34351 5882 5 gnd
rlabel nwell 34296 5621 34319 5624 5 vdd
rlabel locali 34504 6380 34526 6395 5 d0
rlabel locali 34443 6201 34472 6207 5 vdd
rlabel locali 34446 6500 34475 6506 5 gnd
rlabel space 34340 6479 34369 6488 5 gnd
rlabel nwell 34314 6227 34337 6230 5 vdd
rlabel locali 34503 6792 34525 6807 5 d0
rlabel locali 34442 6613 34471 6619 5 vdd
rlabel locali 34445 6912 34474 6918 5 gnd
rlabel space 34339 6891 34368 6900 5 gnd
rlabel nwell 34313 6639 34336 6642 5 vdd
rlabel locali 33628 5367 33657 5373 5 vdd
rlabel locali 33631 5666 33660 5672 5 gnd
rlabel space 33525 5645 33554 5654 5 gnd
rlabel nwell 33499 5393 33522 5396 5 vdd
rlabel locali 33695 5548 33717 5565 5 d1
rlabel locali 33645 6385 33674 6391 5 vdd
rlabel locali 33648 6684 33677 6690 5 gnd
rlabel space 33542 6663 33571 6672 5 gnd
rlabel nwell 33516 6411 33539 6414 5 vdd
rlabel locali 33712 6566 33734 6583 5 d1
rlabel locali 33546 5975 33575 5981 5 vdd
rlabel locali 33549 6274 33578 6280 5 gnd
rlabel space 33443 6253 33472 6262 5 gnd
rlabel nwell 33417 6001 33440 6004 5 vdd
rlabel locali 33613 6149 33633 6173 5 d2
rlabel locali 34524 7398 34546 7413 5 d0
rlabel locali 34463 7219 34492 7225 5 vdd
rlabel locali 34466 7518 34495 7524 5 gnd
rlabel space 34360 7497 34389 7506 5 gnd
rlabel nwell 34334 7245 34357 7248 5 vdd
rlabel locali 34523 7810 34545 7825 5 d0
rlabel locali 34462 7631 34491 7637 5 vdd
rlabel locali 34465 7930 34494 7936 5 gnd
rlabel space 34359 7909 34388 7918 5 gnd
rlabel nwell 34333 7657 34356 7660 5 vdd
rlabel locali 34541 8416 34563 8431 5 d0
rlabel locali 34480 8237 34509 8243 5 vdd
rlabel locali 34483 8536 34512 8542 5 gnd
rlabel space 34377 8515 34406 8524 5 gnd
rlabel nwell 34351 8263 34374 8266 5 vdd
rlabel locali 34540 8828 34562 8843 5 d0
rlabel locali 34479 8649 34508 8655 5 vdd
rlabel locali 34482 8948 34511 8954 5 gnd
rlabel space 34376 8927 34405 8936 5 gnd
rlabel nwell 34350 8675 34373 8678 5 vdd
rlabel locali 34668 8937 34696 8955 5 gnd
rlabel locali 33665 7403 33694 7409 5 vdd
rlabel locali 33668 7702 33697 7708 5 gnd
rlabel space 33562 7681 33591 7690 5 gnd
rlabel nwell 33536 7429 33559 7432 5 vdd
rlabel locali 33732 7584 33754 7601 5 d1
rlabel locali 33682 8421 33711 8427 5 vdd
rlabel locali 33685 8720 33714 8726 5 gnd
rlabel space 33579 8699 33608 8708 5 gnd
rlabel nwell 33553 8447 33576 8450 5 vdd
rlabel locali 33749 8602 33771 8619 5 d1
rlabel locali 33583 8011 33612 8017 5 vdd
rlabel locali 33586 8310 33615 8316 5 gnd
rlabel space 33480 8289 33509 8298 5 gnd
rlabel nwell 33454 8037 33477 8040 5 vdd
rlabel locali 33650 8185 33670 8209 5 d2
rlabel locali 33500 6995 33529 7001 5 vdd
rlabel locali 33503 7294 33532 7300 5 gnd
rlabel space 33397 7273 33426 7282 5 gnd
rlabel nwell 33371 7021 33394 7024 5 vdd
rlabel locali 33565 7174 33585 7187 5 d3
rlabel locali 33324 4961 33353 4967 5 vdd
rlabel locali 33327 5260 33356 5266 5 gnd
rlabel space 33221 5239 33250 5248 5 gnd
rlabel nwell 33195 4987 33218 4990 5 vdd
rlabel locali 33388 5140 33407 5157 5 d4
rlabel locali 31878 4631 31897 4648 1 d4
rlabel nwell 32067 4798 32090 4801 1 vdd
rlabel space 32035 4540 32064 4549 1 gnd
rlabel locali 31929 4522 31958 4528 1 gnd
rlabel locali 31932 4821 31961 4827 1 vdd
rlabel locali 31700 2601 31720 2614 1 d3
rlabel nwell 31891 2764 31914 2767 1 vdd
rlabel space 31859 2506 31888 2515 1 gnd
rlabel locali 31753 2488 31782 2494 1 gnd
rlabel locali 31756 2787 31785 2793 1 vdd
rlabel locali 31615 1579 31635 1603 1 d2
rlabel nwell 31808 1748 31831 1751 1 vdd
rlabel space 31776 1490 31805 1499 1 gnd
rlabel locali 31670 1472 31699 1478 1 gnd
rlabel locali 31673 1771 31702 1777 1 vdd
rlabel locali 31514 1169 31536 1186 1 d1
rlabel nwell 31709 1338 31732 1341 1 vdd
rlabel space 31677 1080 31706 1089 1 gnd
rlabel locali 31571 1062 31600 1068 1 gnd
rlabel locali 31574 1361 31603 1367 1 vdd
rlabel locali 31531 2187 31553 2204 1 d1
rlabel nwell 31726 2356 31749 2359 1 vdd
rlabel space 31694 2098 31723 2107 1 gnd
rlabel locali 31588 2080 31617 2086 1 gnd
rlabel locali 31591 2379 31620 2385 1 vdd
rlabel nwell 30912 1110 30935 1113 1 vdd
rlabel space 30880 852 30909 861 1 gnd
rlabel locali 30774 834 30803 840 1 gnd
rlabel locali 30777 1133 30806 1139 1 vdd
rlabel locali 30723 945 30745 960 1 d0
rlabel nwell 30911 1522 30934 1525 1 vdd
rlabel space 30879 1264 30908 1273 1 gnd
rlabel locali 30773 1246 30802 1252 1 gnd
rlabel locali 30776 1545 30805 1551 1 vdd
rlabel locali 30722 1357 30744 1372 1 d0
rlabel nwell 30929 2128 30952 2131 1 vdd
rlabel space 30897 1870 30926 1879 1 gnd
rlabel locali 30791 1852 30820 1858 1 gnd
rlabel locali 30794 2151 30823 2157 1 vdd
rlabel locali 30740 1963 30762 1978 1 d0
rlabel nwell 30928 2540 30951 2543 1 vdd
rlabel space 30896 2282 30925 2291 1 gnd
rlabel locali 30790 2264 30819 2270 1 gnd
rlabel locali 30793 2563 30822 2569 1 vdd
rlabel locali 30739 2375 30761 2390 1 d0
rlabel locali 31652 3615 31672 3639 1 d2
rlabel nwell 31845 3784 31868 3787 1 vdd
rlabel space 31813 3526 31842 3535 1 gnd
rlabel locali 31707 3508 31736 3514 1 gnd
rlabel locali 31710 3807 31739 3813 1 vdd
rlabel locali 31551 3205 31573 3222 1 d1
rlabel nwell 31746 3374 31769 3377 1 vdd
rlabel space 31714 3116 31743 3125 1 gnd
rlabel locali 31608 3098 31637 3104 1 gnd
rlabel locali 31611 3397 31640 3403 1 vdd
rlabel locali 31568 4223 31590 4240 1 d1
rlabel nwell 31763 4392 31786 4395 1 vdd
rlabel space 31731 4134 31760 4143 1 gnd
rlabel locali 31625 4116 31654 4122 1 gnd
rlabel locali 31628 4415 31657 4421 1 vdd
rlabel nwell 30949 3146 30972 3149 1 vdd
rlabel space 30917 2888 30946 2897 1 gnd
rlabel locali 30811 2870 30840 2876 1 gnd
rlabel locali 30814 3169 30843 3175 1 vdd
rlabel locali 30760 2981 30782 2996 1 d0
rlabel nwell 30948 3558 30971 3561 1 vdd
rlabel space 30916 3300 30945 3309 1 gnd
rlabel locali 30810 3282 30839 3288 1 gnd
rlabel locali 30813 3581 30842 3587 1 vdd
rlabel locali 30759 3393 30781 3408 1 d0
rlabel nwell 30966 4164 30989 4167 1 vdd
rlabel space 30934 3906 30963 3915 1 gnd
rlabel locali 30828 3888 30857 3894 1 gnd
rlabel locali 30831 4187 30860 4193 1 vdd
rlabel locali 30777 3999 30799 4014 1 d0
rlabel nwell 30965 4576 30988 4579 1 vdd
rlabel space 30933 4318 30962 4327 1 gnd
rlabel locali 30827 4300 30856 4306 1 gnd
rlabel locali 30830 4599 30859 4605 1 vdd
rlabel locali 30776 4411 30798 4426 1 d0
rlabel locali 31773 6673 31793 6686 1 d3
rlabel nwell 31964 6836 31987 6839 1 vdd
rlabel space 31932 6578 31961 6587 1 gnd
rlabel locali 31826 6560 31855 6566 1 gnd
rlabel locali 31829 6859 31858 6865 1 vdd
rlabel locali 31688 5651 31708 5675 1 d2
rlabel nwell 31881 5820 31904 5823 1 vdd
rlabel space 31849 5562 31878 5571 1 gnd
rlabel locali 31743 5544 31772 5550 1 gnd
rlabel locali 31746 5843 31775 5849 1 vdd
rlabel locali 31587 5241 31609 5258 1 d1
rlabel nwell 31782 5410 31805 5413 1 vdd
rlabel space 31750 5152 31779 5161 1 gnd
rlabel locali 31644 5134 31673 5140 1 gnd
rlabel locali 31647 5433 31676 5439 1 vdd
rlabel locali 31604 6259 31626 6276 1 d1
rlabel nwell 31799 6428 31822 6431 1 vdd
rlabel space 31767 6170 31796 6179 1 gnd
rlabel locali 31661 6152 31690 6158 1 gnd
rlabel locali 31664 6451 31693 6457 1 vdd
rlabel nwell 30985 5182 31008 5185 1 vdd
rlabel space 30953 4924 30982 4933 1 gnd
rlabel locali 30847 4906 30876 4912 1 gnd
rlabel locali 30850 5205 30879 5211 1 vdd
rlabel locali 30796 5017 30818 5032 1 d0
rlabel nwell 30984 5594 31007 5597 1 vdd
rlabel space 30952 5336 30981 5345 1 gnd
rlabel locali 30846 5318 30875 5324 1 gnd
rlabel locali 30849 5617 30878 5623 1 vdd
rlabel locali 30795 5429 30817 5444 1 d0
rlabel nwell 31002 6200 31025 6203 1 vdd
rlabel space 30970 5942 30999 5951 1 gnd
rlabel locali 30864 5924 30893 5930 1 gnd
rlabel locali 30867 6223 30896 6229 1 vdd
rlabel locali 30813 6035 30835 6050 1 d0
rlabel nwell 31001 6612 31024 6615 1 vdd
rlabel space 30969 6354 30998 6363 1 gnd
rlabel locali 30863 6336 30892 6342 1 gnd
rlabel locali 30866 6635 30895 6641 1 vdd
rlabel locali 30812 6447 30834 6462 1 d0
rlabel locali 31725 7687 31745 7711 1 d2
rlabel nwell 31918 7856 31941 7859 1 vdd
rlabel space 31886 7598 31915 7607 1 gnd
rlabel locali 31780 7580 31809 7586 1 gnd
rlabel locali 31783 7879 31812 7885 1 vdd
rlabel locali 31624 7277 31646 7294 1 d1
rlabel nwell 31819 7446 31842 7449 1 vdd
rlabel space 31787 7188 31816 7197 1 gnd
rlabel locali 31681 7170 31710 7176 1 gnd
rlabel locali 31684 7469 31713 7475 1 vdd
rlabel locali 31641 8295 31663 8312 1 d1
rlabel nwell 31836 8464 31859 8467 1 vdd
rlabel space 31804 8206 31833 8215 1 gnd
rlabel locali 31698 8188 31727 8194 1 gnd
rlabel locali 31701 8487 31730 8493 1 vdd
rlabel nwell 31022 7218 31045 7221 1 vdd
rlabel space 30990 6960 31019 6969 1 gnd
rlabel locali 30884 6942 30913 6948 1 gnd
rlabel locali 30887 7241 30916 7247 1 vdd
rlabel locali 30833 7053 30855 7068 1 d0
rlabel nwell 31021 7630 31044 7633 1 vdd
rlabel space 30989 7372 31018 7381 1 gnd
rlabel locali 30883 7354 30912 7360 1 gnd
rlabel locali 30886 7653 30915 7659 1 vdd
rlabel locali 30832 7465 30854 7480 1 d0
rlabel nwell 31039 8236 31062 8239 1 vdd
rlabel space 31007 7978 31036 7987 1 gnd
rlabel locali 30901 7960 30930 7966 1 gnd
rlabel locali 30904 8259 30933 8265 1 vdd
rlabel locali 30850 8071 30872 8086 1 d0
rlabel nwell 31038 8648 31061 8651 1 vdd
rlabel space 31006 8390 31035 8399 1 gnd
rlabel locali 30900 8372 30929 8378 1 gnd
rlabel locali 30903 8671 30932 8677 1 vdd
rlabel locali 30849 8483 30871 8498 1 d0
rlabel locali 27568 357 27583 370 1 d5
rlabel locali 27626 544 27655 550 1 vdd
rlabel locali 27623 245 27652 251 1 gnd
rlabel space 27729 263 27758 272 1 gnd
rlabel nwell 27761 521 27784 524 1 vdd
rlabel locali 30050 1277 30072 1292 5 d0
rlabel locali 29989 1098 30018 1104 5 vdd
rlabel locali 29992 1397 30021 1403 5 gnd
rlabel space 29886 1376 29915 1385 5 gnd
rlabel nwell 29860 1124 29883 1127 5 vdd
rlabel locali 30049 1689 30071 1704 5 d0
rlabel locali 29988 1510 30017 1516 5 vdd
rlabel locali 29991 1809 30020 1815 5 gnd
rlabel space 29885 1788 29914 1797 5 gnd
rlabel nwell 29859 1536 29882 1539 5 vdd
rlabel locali 30067 2295 30089 2310 5 d0
rlabel locali 30006 2116 30035 2122 5 vdd
rlabel locali 30009 2415 30038 2421 5 gnd
rlabel space 29903 2394 29932 2403 5 gnd
rlabel nwell 29877 2142 29900 2145 5 vdd
rlabel locali 30066 2707 30088 2722 5 d0
rlabel locali 30005 2528 30034 2534 5 vdd
rlabel locali 30008 2827 30037 2833 5 gnd
rlabel space 29902 2806 29931 2815 5 gnd
rlabel nwell 29876 2554 29899 2557 5 vdd
rlabel locali 29191 1282 29220 1288 5 vdd
rlabel locali 29194 1581 29223 1587 5 gnd
rlabel space 29088 1560 29117 1569 5 gnd
rlabel nwell 29062 1308 29085 1311 5 vdd
rlabel locali 29258 1463 29280 1480 5 d1
rlabel locali 29208 2300 29237 2306 5 vdd
rlabel locali 29211 2599 29240 2605 5 gnd
rlabel space 29105 2578 29134 2587 5 gnd
rlabel nwell 29079 2326 29102 2329 5 vdd
rlabel locali 29275 2481 29297 2498 5 d1
rlabel locali 29109 1890 29138 1896 5 vdd
rlabel locali 29112 2189 29141 2195 5 gnd
rlabel space 29006 2168 29035 2177 5 gnd
rlabel nwell 28980 1916 29003 1919 5 vdd
rlabel locali 29176 2064 29196 2088 5 d2
rlabel locali 30087 3313 30109 3328 5 d0
rlabel locali 30026 3134 30055 3140 5 vdd
rlabel locali 30029 3433 30058 3439 5 gnd
rlabel space 29923 3412 29952 3421 5 gnd
rlabel nwell 29897 3160 29920 3163 5 vdd
rlabel locali 30086 3725 30108 3740 5 d0
rlabel locali 30025 3546 30054 3552 5 vdd
rlabel locali 30028 3845 30057 3851 5 gnd
rlabel space 29922 3824 29951 3833 5 gnd
rlabel nwell 29896 3572 29919 3575 5 vdd
rlabel locali 30104 4331 30126 4346 5 d0
rlabel locali 30043 4152 30072 4158 5 vdd
rlabel locali 30046 4451 30075 4457 5 gnd
rlabel space 29940 4430 29969 4439 5 gnd
rlabel nwell 29914 4178 29937 4181 5 vdd
rlabel locali 30103 4743 30125 4758 5 d0
rlabel locali 30042 4564 30071 4570 5 vdd
rlabel locali 30045 4863 30074 4869 5 gnd
rlabel space 29939 4842 29968 4851 5 gnd
rlabel nwell 29913 4590 29936 4593 5 vdd
rlabel locali 29228 3318 29257 3324 5 vdd
rlabel locali 29231 3617 29260 3623 5 gnd
rlabel space 29125 3596 29154 3605 5 gnd
rlabel nwell 29099 3344 29122 3347 5 vdd
rlabel locali 29295 3499 29317 3516 5 d1
rlabel locali 29245 4336 29274 4342 5 vdd
rlabel locali 29248 4635 29277 4641 5 gnd
rlabel space 29142 4614 29171 4623 5 gnd
rlabel nwell 29116 4362 29139 4365 5 vdd
rlabel locali 29312 4517 29334 4534 5 d1
rlabel locali 29146 3926 29175 3932 5 vdd
rlabel locali 29149 4225 29178 4231 5 gnd
rlabel space 29043 4204 29072 4213 5 gnd
rlabel nwell 29017 3952 29040 3955 5 vdd
rlabel locali 29213 4100 29233 4124 5 d2
rlabel locali 29063 2910 29092 2916 5 vdd
rlabel locali 29066 3209 29095 3215 5 gnd
rlabel space 28960 3188 28989 3197 5 gnd
rlabel nwell 28934 2936 28957 2939 5 vdd
rlabel locali 29128 3089 29148 3102 5 d3
rlabel locali 30123 5349 30145 5364 5 d0
rlabel locali 30062 5170 30091 5176 5 vdd
rlabel locali 30065 5469 30094 5475 5 gnd
rlabel space 29959 5448 29988 5457 5 gnd
rlabel nwell 29933 5196 29956 5199 5 vdd
rlabel locali 30122 5761 30144 5776 5 d0
rlabel locali 30061 5582 30090 5588 5 vdd
rlabel locali 30064 5881 30093 5887 5 gnd
rlabel space 29958 5860 29987 5869 5 gnd
rlabel nwell 29932 5608 29955 5611 5 vdd
rlabel locali 30140 6367 30162 6382 5 d0
rlabel locali 30079 6188 30108 6194 5 vdd
rlabel locali 30082 6487 30111 6493 5 gnd
rlabel space 29976 6466 30005 6475 5 gnd
rlabel nwell 29950 6214 29973 6217 5 vdd
rlabel locali 30139 6779 30161 6794 5 d0
rlabel locali 30078 6600 30107 6606 5 vdd
rlabel locali 30081 6899 30110 6905 5 gnd
rlabel space 29975 6878 30004 6887 5 gnd
rlabel nwell 29949 6626 29972 6629 5 vdd
rlabel locali 29264 5354 29293 5360 5 vdd
rlabel locali 29267 5653 29296 5659 5 gnd
rlabel space 29161 5632 29190 5641 5 gnd
rlabel nwell 29135 5380 29158 5383 5 vdd
rlabel locali 29331 5535 29353 5552 5 d1
rlabel locali 29281 6372 29310 6378 5 vdd
rlabel locali 29284 6671 29313 6677 5 gnd
rlabel space 29178 6650 29207 6659 5 gnd
rlabel nwell 29152 6398 29175 6401 5 vdd
rlabel locali 29348 6553 29370 6570 5 d1
rlabel locali 29182 5962 29211 5968 5 vdd
rlabel locali 29185 6261 29214 6267 5 gnd
rlabel space 29079 6240 29108 6249 5 gnd
rlabel nwell 29053 5988 29076 5991 5 vdd
rlabel locali 29249 6136 29269 6160 5 d2
rlabel locali 30160 7385 30182 7400 5 d0
rlabel locali 30099 7206 30128 7212 5 vdd
rlabel locali 30102 7505 30131 7511 5 gnd
rlabel space 29996 7484 30025 7493 5 gnd
rlabel nwell 29970 7232 29993 7235 5 vdd
rlabel locali 30159 7797 30181 7812 5 d0
rlabel locali 30098 7618 30127 7624 5 vdd
rlabel locali 30101 7917 30130 7923 5 gnd
rlabel space 29995 7896 30024 7905 5 gnd
rlabel nwell 29969 7644 29992 7647 5 vdd
rlabel locali 30177 8403 30199 8418 5 d0
rlabel locali 30116 8224 30145 8230 5 vdd
rlabel locali 30119 8523 30148 8529 5 gnd
rlabel space 30013 8502 30042 8511 5 gnd
rlabel nwell 29987 8250 30010 8253 5 vdd
rlabel locali 30176 8815 30198 8830 5 d0
rlabel locali 30115 8636 30144 8642 5 vdd
rlabel locali 30118 8935 30147 8941 5 gnd
rlabel space 30012 8914 30041 8923 5 gnd
rlabel nwell 29986 8662 30009 8665 5 vdd
rlabel locali 29301 7390 29330 7396 5 vdd
rlabel locali 29304 7689 29333 7695 5 gnd
rlabel space 29198 7668 29227 7677 5 gnd
rlabel nwell 29172 7416 29195 7419 5 vdd
rlabel locali 29368 7571 29390 7588 5 d1
rlabel locali 29318 8408 29347 8414 5 vdd
rlabel locali 29321 8707 29350 8713 5 gnd
rlabel space 29215 8686 29244 8695 5 gnd
rlabel nwell 29189 8434 29212 8437 5 vdd
rlabel locali 29385 8589 29407 8606 5 d1
rlabel locali 29219 7998 29248 8004 5 vdd
rlabel locali 29222 8297 29251 8303 5 gnd
rlabel space 29116 8276 29145 8285 5 gnd
rlabel nwell 29090 8024 29113 8027 5 vdd
rlabel locali 29286 8172 29306 8196 5 d2
rlabel locali 29136 6982 29165 6988 5 vdd
rlabel locali 29139 7281 29168 7287 5 gnd
rlabel space 29033 7260 29062 7269 5 gnd
rlabel nwell 29007 7008 29030 7011 5 vdd
rlabel locali 29201 7161 29221 7174 5 d3
rlabel locali 28960 4948 28989 4954 5 vdd
rlabel locali 28963 5247 28992 5253 5 gnd
rlabel space 28857 5226 28886 5235 5 gnd
rlabel nwell 28831 4974 28854 4977 5 vdd
rlabel locali 29024 5127 29043 5144 5 d4
rlabel locali 27514 4618 27533 4635 1 d4
rlabel nwell 27703 4785 27726 4788 1 vdd
rlabel space 27671 4527 27700 4536 1 gnd
rlabel locali 27565 4509 27594 4515 1 gnd
rlabel locali 27568 4808 27597 4814 1 vdd
rlabel locali 27336 2588 27356 2601 1 d3
rlabel nwell 27527 2751 27550 2754 1 vdd
rlabel space 27495 2493 27524 2502 1 gnd
rlabel locali 27389 2475 27418 2481 1 gnd
rlabel locali 27392 2774 27421 2780 1 vdd
rlabel locali 27251 1566 27271 1590 1 d2
rlabel nwell 27444 1735 27467 1738 1 vdd
rlabel space 27412 1477 27441 1486 1 gnd
rlabel locali 27306 1459 27335 1465 1 gnd
rlabel locali 27309 1758 27338 1764 1 vdd
rlabel locali 27150 1156 27172 1173 1 d1
rlabel nwell 27345 1325 27368 1328 1 vdd
rlabel space 27313 1067 27342 1076 1 gnd
rlabel locali 27207 1049 27236 1055 1 gnd
rlabel locali 27210 1348 27239 1354 1 vdd
rlabel locali 27167 2174 27189 2191 1 d1
rlabel nwell 27362 2343 27385 2346 1 vdd
rlabel space 27330 2085 27359 2094 1 gnd
rlabel locali 27224 2067 27253 2073 1 gnd
rlabel locali 27227 2366 27256 2372 1 vdd
rlabel nwell 26548 1097 26571 1100 1 vdd
rlabel space 26516 839 26545 848 1 gnd
rlabel locali 26410 821 26439 827 1 gnd
rlabel locali 26413 1120 26442 1126 1 vdd
rlabel locali 26359 932 26381 947 1 d0
rlabel nwell 26547 1509 26570 1512 1 vdd
rlabel space 26515 1251 26544 1260 1 gnd
rlabel locali 26409 1233 26438 1239 1 gnd
rlabel locali 26412 1532 26441 1538 1 vdd
rlabel locali 26358 1344 26380 1359 1 d0
rlabel nwell 26565 2115 26588 2118 1 vdd
rlabel space 26533 1857 26562 1866 1 gnd
rlabel locali 26427 1839 26456 1845 1 gnd
rlabel locali 26430 2138 26459 2144 1 vdd
rlabel locali 26376 1950 26398 1965 1 d0
rlabel nwell 26564 2527 26587 2530 1 vdd
rlabel space 26532 2269 26561 2278 1 gnd
rlabel locali 26426 2251 26455 2257 1 gnd
rlabel locali 26429 2550 26458 2556 1 vdd
rlabel locali 26375 2362 26397 2377 1 d0
rlabel locali 27288 3602 27308 3626 1 d2
rlabel nwell 27481 3771 27504 3774 1 vdd
rlabel space 27449 3513 27478 3522 1 gnd
rlabel locali 27343 3495 27372 3501 1 gnd
rlabel locali 27346 3794 27375 3800 1 vdd
rlabel locali 27187 3192 27209 3209 1 d1
rlabel nwell 27382 3361 27405 3364 1 vdd
rlabel space 27350 3103 27379 3112 1 gnd
rlabel locali 27244 3085 27273 3091 1 gnd
rlabel locali 27247 3384 27276 3390 1 vdd
rlabel locali 27204 4210 27226 4227 1 d1
rlabel nwell 27399 4379 27422 4382 1 vdd
rlabel space 27367 4121 27396 4130 1 gnd
rlabel locali 27261 4103 27290 4109 1 gnd
rlabel locali 27264 4402 27293 4408 1 vdd
rlabel nwell 26585 3133 26608 3136 1 vdd
rlabel space 26553 2875 26582 2884 1 gnd
rlabel locali 26447 2857 26476 2863 1 gnd
rlabel locali 26450 3156 26479 3162 1 vdd
rlabel locali 26396 2968 26418 2983 1 d0
rlabel nwell 26584 3545 26607 3548 1 vdd
rlabel space 26552 3287 26581 3296 1 gnd
rlabel locali 26446 3269 26475 3275 1 gnd
rlabel locali 26449 3568 26478 3574 1 vdd
rlabel locali 26395 3380 26417 3395 1 d0
rlabel nwell 26602 4151 26625 4154 1 vdd
rlabel space 26570 3893 26599 3902 1 gnd
rlabel locali 26464 3875 26493 3881 1 gnd
rlabel locali 26467 4174 26496 4180 1 vdd
rlabel locali 26413 3986 26435 4001 1 d0
rlabel nwell 26601 4563 26624 4566 1 vdd
rlabel space 26569 4305 26598 4314 1 gnd
rlabel locali 26463 4287 26492 4293 1 gnd
rlabel locali 26466 4586 26495 4592 1 vdd
rlabel locali 26412 4398 26434 4413 1 d0
rlabel locali 27409 6660 27429 6673 1 d3
rlabel nwell 27600 6823 27623 6826 1 vdd
rlabel space 27568 6565 27597 6574 1 gnd
rlabel locali 27462 6547 27491 6553 1 gnd
rlabel locali 27465 6846 27494 6852 1 vdd
rlabel locali 27324 5638 27344 5662 1 d2
rlabel nwell 27517 5807 27540 5810 1 vdd
rlabel space 27485 5549 27514 5558 1 gnd
rlabel locali 27379 5531 27408 5537 1 gnd
rlabel locali 27382 5830 27411 5836 1 vdd
rlabel locali 27223 5228 27245 5245 1 d1
rlabel nwell 27418 5397 27441 5400 1 vdd
rlabel space 27386 5139 27415 5148 1 gnd
rlabel locali 27280 5121 27309 5127 1 gnd
rlabel locali 27283 5420 27312 5426 1 vdd
rlabel locali 27240 6246 27262 6263 1 d1
rlabel nwell 27435 6415 27458 6418 1 vdd
rlabel space 27403 6157 27432 6166 1 gnd
rlabel locali 27297 6139 27326 6145 1 gnd
rlabel locali 27300 6438 27329 6444 1 vdd
rlabel nwell 26621 5169 26644 5172 1 vdd
rlabel space 26589 4911 26618 4920 1 gnd
rlabel locali 26483 4893 26512 4899 1 gnd
rlabel locali 26486 5192 26515 5198 1 vdd
rlabel locali 26432 5004 26454 5019 1 d0
rlabel nwell 26620 5581 26643 5584 1 vdd
rlabel space 26588 5323 26617 5332 1 gnd
rlabel locali 26482 5305 26511 5311 1 gnd
rlabel locali 26485 5604 26514 5610 1 vdd
rlabel locali 26431 5416 26453 5431 1 d0
rlabel nwell 26638 6187 26661 6190 1 vdd
rlabel space 26606 5929 26635 5938 1 gnd
rlabel locali 26500 5911 26529 5917 1 gnd
rlabel locali 26503 6210 26532 6216 1 vdd
rlabel locali 26449 6022 26471 6037 1 d0
rlabel nwell 26637 6599 26660 6602 1 vdd
rlabel space 26605 6341 26634 6350 1 gnd
rlabel locali 26499 6323 26528 6329 1 gnd
rlabel locali 26502 6622 26531 6628 1 vdd
rlabel locali 26448 6434 26470 6449 1 d0
rlabel locali 27361 7674 27381 7698 1 d2
rlabel nwell 27554 7843 27577 7846 1 vdd
rlabel space 27522 7585 27551 7594 1 gnd
rlabel locali 27416 7567 27445 7573 1 gnd
rlabel locali 27419 7866 27448 7872 1 vdd
rlabel locali 27260 7264 27282 7281 1 d1
rlabel nwell 27455 7433 27478 7436 1 vdd
rlabel space 27423 7175 27452 7184 1 gnd
rlabel locali 27317 7157 27346 7163 1 gnd
rlabel locali 27320 7456 27349 7462 1 vdd
rlabel locali 27277 8282 27299 8299 1 d1
rlabel nwell 27472 8451 27495 8454 1 vdd
rlabel space 27440 8193 27469 8202 1 gnd
rlabel locali 27334 8175 27363 8181 1 gnd
rlabel locali 27337 8474 27366 8480 1 vdd
rlabel nwell 26658 7205 26681 7208 1 vdd
rlabel space 26626 6947 26655 6956 1 gnd
rlabel locali 26520 6929 26549 6935 1 gnd
rlabel locali 26523 7228 26552 7234 1 vdd
rlabel locali 26469 7040 26491 7055 1 d0
rlabel nwell 26657 7617 26680 7620 1 vdd
rlabel space 26625 7359 26654 7368 1 gnd
rlabel locali 26519 7341 26548 7347 1 gnd
rlabel locali 26522 7640 26551 7646 1 vdd
rlabel locali 26468 7452 26490 7467 1 d0
rlabel nwell 26675 8223 26698 8226 1 vdd
rlabel space 26643 7965 26672 7974 1 gnd
rlabel locali 26537 7947 26566 7953 1 gnd
rlabel locali 26540 8246 26569 8252 1 vdd
rlabel locali 26486 8058 26508 8073 1 d0
rlabel nwell 26674 8635 26697 8638 1 vdd
rlabel space 26642 8377 26671 8386 1 gnd
rlabel locali 26536 8359 26565 8365 1 gnd
rlabel locali 26539 8658 26568 8664 1 vdd
rlabel locali 26485 8470 26507 8485 1 d0
rlabel locali 25822 469 25851 475 1 vdd
rlabel locali 25819 170 25848 176 1 gnd
rlabel space 25925 188 25954 197 1 gnd
rlabel nwell 25957 446 25980 449 1 vdd
rlabel locali 25761 282 25783 297 1 d7
rlabel locali 16941 394 16970 400 1 vdd
rlabel locali 16938 95 16967 101 1 gnd
rlabel space 17044 113 17073 122 1 gnd
rlabel nwell 17076 371 17099 374 1 vdd
rlabel locali 17314 241 17336 256 1 vout
rlabel locali 16878 207 16895 219 1 d8
<< end >>

* SPICE3 file created from 4bit_DAC1.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_142_1423# a_148_1606# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1 a_586_n525# d1 a_1372_n1198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_388_493# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3 a_94_n1448# d0 a_569_n1543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_105_n613# a_111_n430# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5 a_586_n525# a_368_n525# a_111_n430# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6 a_98_n831# d0 a_587_n937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7 a_96_n930# a_98_n831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8 a_1166_n709# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9 a_405_1511# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 a_1450_n301# d3 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X11 a_1285_719# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 a_125_405# d0 a_606_493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X13 gnd a_81_n1849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X14 a_1186_309# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 a_606_493# a_388_493# a_125_405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_125_405# a_131_588# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X17 a_624_1099# a_406_1099# a_135_1205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X18 a_1248_n1317# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 a_569_n1543# d1 a_1367_n1727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 a_94_n1448# a_96_n930# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X21 a_131_588# a_133_1106# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X22 a_118_187# d0 a_607_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X23 a_133_1106# a_135_1205# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X24 a_135_1205# a_142_1423# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X25 vout a_1331_n301# a_1450_n301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X26 a_81_n1849# a_88_n1631# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X27 a_368_n525# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X28 a_1409_838# a_1203_1327# a_624_1099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X29 a_587_n937# a_369_n937# a_98_n831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X30 a_1455_n182# a_1285_719# a_1404_309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X31 a_569_n1543# a_351_n1543# a_94_n1448# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X32 a_586_n525# a_368_n525# a_105_n613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X33 a_135_1205# d0 a_624_1099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X34 a_1404_309# a_1186_309# a_607_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X35 a_1285_719# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X36 a_148_1606# d0 a_623_1511# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X37 a_352_n1955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X38 a_1186_309# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X39 a_406_1099# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X40 a_623_1511# d1 a_1409_838# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X41 a_1331_n301# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X42 a_116_n106# d0 a_607_81# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X43 a_1372_n1198# a_1166_n709# a_587_n937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X44 a_1367_n1727# a_1149_n1727# a_569_n1543# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X45 a_1450_n301# a_1248_n1317# a_1372_n1198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X46 a_1203_1327# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X47 a_369_n937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X48 a_1409_838# a_1203_1327# a_623_1511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X49 a_1455_n182# a_1285_719# a_1409_838# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X50 a_368_n525# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_587_n937# a_369_n937# a_96_n930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_1372_n1198# d2 a_1450_n301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X53 a_607_81# a_389_81# a_116_n106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_569_n1543# a_351_n1543# a_88_n1631# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X55 a_1404_309# a_1186_309# a_606_493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X56 a_388_493# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X57 a_587_n937# d1 a_1372_n1198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X58 a_142_1423# d0 a_623_1511# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X59 gnd d0 a_570_n1955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X60 a_624_1099# d1 a_1409_838# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X61 a_352_n1955# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X62 a_116_n106# a_118_187# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X63 a_1166_n709# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X64 a_1455_n182# d3 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X65 a_1203_1327# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X66 a_351_n1543# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X67 a_148_1606# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X68 a_131_588# d0 a_606_493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X69 a_1367_n1727# a_1149_n1727# a_570_n1955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X70 a_606_493# a_388_493# a_131_588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X71 a_369_n937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_1248_n1317# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X73 a_1149_n1727# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X74 a_98_n831# a_105_n613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X75 a_105_n613# d0 a_586_n525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X76 a_624_1099# a_406_1099# a_133_1106# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X77 a_111_n430# a_116_n106# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X78 a_623_1511# a_405_1511# a_142_1423# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X79 a_1409_838# d2 a_1455_n182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X80 vout a_1331_n301# a_1455_n182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X81 a_81_n1849# d0 a_570_n1955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X82 a_133_1106# d0 a_624_1099# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X83 a_570_n1955# a_352_n1955# a_81_n1849# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X84 a_606_493# d1 a_1404_309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X85 a_389_81# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X86 a_118_187# a_125_405# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X87 a_88_n1631# d0 a_569_n1543# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X88 a_88_n1631# a_94_n1448# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X89 a_351_n1543# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X90 a_96_n930# d0 a_587_n937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X91 a_406_1099# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_111_n430# d0 a_586_n525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 a_1149_n1727# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 a_1331_n301# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X95 a_405_1511# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X96 a_1372_n1198# a_1166_n709# a_586_n525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X97 a_1404_309# d2 a_1455_n182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X98 a_623_1511# a_405_1511# a_148_1606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X99 a_389_81# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X100 a_1450_n301# a_1248_n1317# a_1367_n1727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_607_81# a_389_81# a_118_187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X102 a_607_81# d1 a_1404_309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X103 a_570_n1955# d1 a_1367_n1727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X104 a_1367_n1727# d2 a_1450_n301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X105 a_570_n1955# a_352_n1955# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
C0 gnd SUB 3.38fF
C1 vdd SUB 9.87fF
C2 d0 SUB 2.56fF
C3 a_570_n1955# SUB 2.21fF
C4 a_569_n1543# SUB 2.30fF
C5 a_587_n937# SUB 2.21fF
C6 a_586_n525# SUB 2.30fF
C7 a_607_81# SUB 2.21fF
C8 a_606_493# SUB 2.30fF
C9 a_624_1099# SUB 2.21fF
C10 a_623_1511# SUB 2.30fF


Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40ns 80ns)


.tran 1ns 80ns
.control
run
plot V(vout) V(d0) V(d1) V(d2) V(d3)
.endc
.end

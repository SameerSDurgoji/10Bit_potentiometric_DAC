* SPICE3 file created from 3bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_388_493# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 a_1233_n709# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_1456_n180# a_1250_309# a_607_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3 a_589_n525# a_371_n525# a_114_n430# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4 a_101_n831# a_108_n613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5 a_125_405# d0 a_606_493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6 a_1456_n180# d2 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7 a_101_n831# d0 a_590_n937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X8 a_114_n430# a_116_88# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X9 a_1451_n709# a_1233_n709# a_589_n525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 a_125_405# a_131_588# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X11 a_606_493# a_388_493# a_125_405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 a_372_n937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_1332_n299# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X14 a_131_588# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X15 a_118_187# d0 a_607_81# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 a_1456_n180# a_1250_309# a_606_493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X17 a_590_n937# d1 a_1451_n709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X18 a_589_n525# a_371_n525# a_108_n613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 a_108_n613# a_114_n430# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X20 gnd a_101_n831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X21 a_116_88# d0 a_607_81# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X22 a_1332_n299# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X23 a_1250_309# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_607_81# a_389_81# a_116_88# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X25 a_388_493# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X26 a_606_493# d1 a_1456_n180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_1233_n709# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X28 a_116_88# a_118_187# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X29 a_606_493# a_388_493# a_131_588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X30 a_131_588# d0 a_606_493# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X31 a_1451_n709# a_1233_n709# a_590_n937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X32 a_1250_309# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X33 a_108_n613# d0 a_589_n525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X34 a_607_81# d1 a_1456_n180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X35 vout a_1332_n299# a_1456_n180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X36 a_371_n525# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X37 a_589_n525# d1 a_1451_n709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_590_n937# a_372_n937# a_101_n831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X39 a_118_187# a_125_405# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X40 a_389_81# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X41 gnd d0 a_590_n937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X42 a_389_81# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X43 a_1451_n709# d2 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X44 a_114_n430# d0 a_589_n525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X45 a_607_81# a_389_81# a_118_187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X46 a_371_n525# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X47 a_372_n937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X48 vout a_1332_n299# a_1451_n709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X49 a_590_n937# a_372_n937# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
C0 vdd SUB 4.51fF
C1 a_590_n937# SUB 2.27fF
C2 a_589_n525# SUB 2.35fF
C3 a_607_81# SUB 2.27fF
C4 a_606_493# SUB 2.36fF


Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)

.tran 0.1ns 40ns
.control
run
plot V(vout) V(d0) V(d1) V(d2)
.endc
.end

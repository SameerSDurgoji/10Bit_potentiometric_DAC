* SPICE3 file created from 2bit_DAC3.ext - technology: sky130A

*.option scale=1.000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_42_n7# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1 vrefh d1 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_36_n190# a_42_n7# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3 a_299_n102# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 gnd a_29_n408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5 vrefl a_300_n514# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_1161_n286# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7 a_29_n408# a_36_n190# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X8 a_299_n102# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X9 gnd d0 vrefl vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 vout a_1161_n286# vrefh vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X11 a_300_n514# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X12 vout a_1161_n286# vrefl SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_36_n190# d0 vrefh vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X14 a_42_n7# d0 vrefh SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X15 vrefl a_300_n514# a_29_n408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X16 a_29_n408# d0 vrefl SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 vrefh a_299_n102# a_42_n7# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X18 a_300_n514# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X19 vrefl d1 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X20 vrefh a_299_n102# a_36_n190# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X21 a_1161_n286# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
C0 vdd SUB 2.32fF
C1 vrefl SUB 2.27fF
C2 vrefh SUB 2.36fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)

.tran 0.1ns 20ns
.control
run
plot V(vout) V(d0) V(d1)
.endc
.end

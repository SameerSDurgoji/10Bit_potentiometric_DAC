magic
tech sky130A
timestamp 1616093997
<< nwell >>
rect 3450 8426 4058 8576
rect 7814 8439 8422 8589
rect 401 8272 1009 8422
rect 1199 8088 1807 8238
rect 2653 8198 3261 8348
rect 4765 8285 5373 8435
rect 3451 8014 4059 8164
rect 5563 8101 6171 8251
rect 7017 8211 7625 8361
rect 7815 8027 8423 8177
rect 402 7860 1010 8010
rect 2554 7788 3162 7938
rect 4766 7873 5374 8023
rect 6918 7801 7526 7951
rect 1281 7480 1889 7630
rect 3433 7408 4041 7558
rect 5645 7493 6253 7643
rect 7797 7421 8405 7571
rect 384 7254 992 7404
rect 1182 7070 1790 7220
rect 2636 7180 3244 7330
rect 4748 7267 5356 7417
rect 3434 6996 4042 7146
rect 5546 7083 6154 7233
rect 7000 7193 7608 7343
rect 7798 7009 8406 7159
rect 385 6842 993 6992
rect 2471 6772 3079 6922
rect 4749 6855 5357 7005
rect 6835 6785 7443 6935
rect 1327 6460 1935 6610
rect 3413 6390 4021 6540
rect 5691 6473 6299 6623
rect 7777 6403 8385 6553
rect 364 6236 972 6386
rect 1162 6052 1770 6202
rect 2616 6162 3224 6312
rect 4728 6249 5336 6399
rect 3414 5978 4022 6128
rect 5526 6065 6134 6215
rect 6980 6175 7588 6325
rect 7778 5991 8386 6141
rect 365 5824 973 5974
rect 2517 5752 3125 5902
rect 4729 5837 5337 5987
rect 6881 5765 7489 5915
rect 1244 5444 1852 5594
rect 3396 5372 4004 5522
rect 5608 5457 6216 5607
rect 7760 5385 8368 5535
rect 347 5218 955 5368
rect 1145 5034 1753 5184
rect 2599 5144 3207 5294
rect 4711 5231 5319 5381
rect 3397 4960 4005 5110
rect 5509 5047 6117 5197
rect 6963 5157 7571 5307
rect 7761 4973 8369 5123
rect 348 4806 956 4956
rect 2295 4738 2903 4888
rect 4712 4819 5320 4969
rect 6659 4751 7267 4901
rect 1430 4422 2038 4572
rect 3377 4354 3985 4504
rect 5794 4435 6402 4585
rect 7741 4367 8349 4517
rect 328 4200 936 4350
rect 1126 4016 1734 4166
rect 2580 4126 3188 4276
rect 4692 4213 5300 4363
rect 3378 3942 3986 4092
rect 5490 4029 6098 4179
rect 6944 4139 7552 4289
rect 7742 3955 8350 4105
rect 329 3788 937 3938
rect 2481 3716 3089 3866
rect 4693 3801 5301 3951
rect 6845 3729 7453 3879
rect 1208 3408 1816 3558
rect 3360 3336 3968 3486
rect 5572 3421 6180 3571
rect 7724 3349 8332 3499
rect 311 3182 919 3332
rect 1109 2998 1717 3148
rect 2563 3108 3171 3258
rect 4675 3195 5283 3345
rect 3361 2924 3969 3074
rect 5473 3011 6081 3161
rect 6927 3121 7535 3271
rect 7725 2937 8333 3087
rect 312 2770 920 2920
rect 2398 2700 3006 2850
rect 4676 2783 5284 2933
rect 6762 2713 7370 2863
rect 1254 2388 1862 2538
rect 3340 2318 3948 2468
rect 5618 2401 6226 2551
rect 7704 2331 8312 2481
rect 291 2164 899 2314
rect 1089 1980 1697 2130
rect 2543 2090 3151 2240
rect 4655 2177 5263 2327
rect 3341 1906 3949 2056
rect 5453 1993 6061 2143
rect 6907 2103 7515 2253
rect 7705 1919 8313 2069
rect 292 1752 900 1902
rect 2444 1680 3052 1830
rect 4656 1765 5264 1915
rect 6808 1693 7416 1843
rect 1171 1372 1779 1522
rect 3323 1300 3931 1450
rect 5535 1385 6143 1535
rect 7687 1313 8295 1463
rect 274 1146 882 1296
rect 1072 962 1680 1112
rect 2526 1072 3134 1222
rect 4638 1159 5246 1309
rect 3324 888 3932 1038
rect 5436 975 6044 1125
rect 6890 1085 7498 1235
rect 7688 901 8296 1051
rect 275 734 883 884
rect 4639 747 5247 897
rect 1488 158 2096 308
rect 3977 84 4585 234
rect 5852 171 6460 321
<< nmos >>
rect 3518 8635 3568 8677
rect 3726 8635 3776 8677
rect 3944 8635 3994 8677
rect 7882 8648 7932 8690
rect 8090 8648 8140 8690
rect 8308 8648 8358 8690
rect 2721 8407 2771 8449
rect 2929 8407 2979 8449
rect 3147 8407 3197 8449
rect 7085 8420 7135 8462
rect 7293 8420 7343 8462
rect 7511 8420 7561 8462
rect 465 8171 515 8213
rect 683 8171 733 8213
rect 891 8171 941 8213
rect 3519 8223 3569 8265
rect 3727 8223 3777 8265
rect 3945 8223 3995 8265
rect 4829 8184 4879 8226
rect 5047 8184 5097 8226
rect 5255 8184 5305 8226
rect 7883 8236 7933 8278
rect 8091 8236 8141 8278
rect 8309 8236 8359 8278
rect 1263 7987 1313 8029
rect 1481 7987 1531 8029
rect 1689 7987 1739 8029
rect 2622 7997 2672 8039
rect 2830 7997 2880 8039
rect 3048 7997 3098 8039
rect 5627 8000 5677 8042
rect 5845 8000 5895 8042
rect 6053 8000 6103 8042
rect 6986 8010 7036 8052
rect 7194 8010 7244 8052
rect 7412 8010 7462 8052
rect 466 7759 516 7801
rect 684 7759 734 7801
rect 892 7759 942 7801
rect 4830 7772 4880 7814
rect 5048 7772 5098 7814
rect 5256 7772 5306 7814
rect 3501 7617 3551 7659
rect 3709 7617 3759 7659
rect 3927 7617 3977 7659
rect 7865 7630 7915 7672
rect 8073 7630 8123 7672
rect 8291 7630 8341 7672
rect 1345 7379 1395 7421
rect 1563 7379 1613 7421
rect 1771 7379 1821 7421
rect 2704 7389 2754 7431
rect 2912 7389 2962 7431
rect 3130 7389 3180 7431
rect 5709 7392 5759 7434
rect 5927 7392 5977 7434
rect 6135 7392 6185 7434
rect 7068 7402 7118 7444
rect 7276 7402 7326 7444
rect 7494 7402 7544 7444
rect 448 7153 498 7195
rect 666 7153 716 7195
rect 874 7153 924 7195
rect 3502 7205 3552 7247
rect 3710 7205 3760 7247
rect 3928 7205 3978 7247
rect 4812 7166 4862 7208
rect 5030 7166 5080 7208
rect 5238 7166 5288 7208
rect 7866 7218 7916 7260
rect 8074 7218 8124 7260
rect 8292 7218 8342 7260
rect 1246 6969 1296 7011
rect 1464 6969 1514 7011
rect 1672 6969 1722 7011
rect 2539 6981 2589 7023
rect 2747 6981 2797 7023
rect 2965 6981 3015 7023
rect 5610 6982 5660 7024
rect 5828 6982 5878 7024
rect 6036 6982 6086 7024
rect 6903 6994 6953 7036
rect 7111 6994 7161 7036
rect 7329 6994 7379 7036
rect 449 6741 499 6783
rect 667 6741 717 6783
rect 875 6741 925 6783
rect 4813 6754 4863 6796
rect 5031 6754 5081 6796
rect 5239 6754 5289 6796
rect 3481 6599 3531 6641
rect 3689 6599 3739 6641
rect 3907 6599 3957 6641
rect 7845 6612 7895 6654
rect 8053 6612 8103 6654
rect 8271 6612 8321 6654
rect 1391 6359 1441 6401
rect 1609 6359 1659 6401
rect 1817 6359 1867 6401
rect 2684 6371 2734 6413
rect 2892 6371 2942 6413
rect 3110 6371 3160 6413
rect 5755 6372 5805 6414
rect 5973 6372 6023 6414
rect 6181 6372 6231 6414
rect 7048 6384 7098 6426
rect 7256 6384 7306 6426
rect 7474 6384 7524 6426
rect 428 6135 478 6177
rect 646 6135 696 6177
rect 854 6135 904 6177
rect 3482 6187 3532 6229
rect 3690 6187 3740 6229
rect 3908 6187 3958 6229
rect 4792 6148 4842 6190
rect 5010 6148 5060 6190
rect 5218 6148 5268 6190
rect 7846 6200 7896 6242
rect 8054 6200 8104 6242
rect 8272 6200 8322 6242
rect 1226 5951 1276 5993
rect 1444 5951 1494 5993
rect 1652 5951 1702 5993
rect 2585 5961 2635 6003
rect 2793 5961 2843 6003
rect 3011 5961 3061 6003
rect 5590 5964 5640 6006
rect 5808 5964 5858 6006
rect 6016 5964 6066 6006
rect 6949 5974 6999 6016
rect 7157 5974 7207 6016
rect 7375 5974 7425 6016
rect 429 5723 479 5765
rect 647 5723 697 5765
rect 855 5723 905 5765
rect 4793 5736 4843 5778
rect 5011 5736 5061 5778
rect 5219 5736 5269 5778
rect 3464 5581 3514 5623
rect 3672 5581 3722 5623
rect 3890 5581 3940 5623
rect 7828 5594 7878 5636
rect 8036 5594 8086 5636
rect 8254 5594 8304 5636
rect 1308 5343 1358 5385
rect 1526 5343 1576 5385
rect 1734 5343 1784 5385
rect 2667 5353 2717 5395
rect 2875 5353 2925 5395
rect 3093 5353 3143 5395
rect 5672 5356 5722 5398
rect 5890 5356 5940 5398
rect 6098 5356 6148 5398
rect 7031 5366 7081 5408
rect 7239 5366 7289 5408
rect 7457 5366 7507 5408
rect 411 5117 461 5159
rect 629 5117 679 5159
rect 837 5117 887 5159
rect 3465 5169 3515 5211
rect 3673 5169 3723 5211
rect 3891 5169 3941 5211
rect 4775 5130 4825 5172
rect 4993 5130 5043 5172
rect 5201 5130 5251 5172
rect 7829 5182 7879 5224
rect 8037 5182 8087 5224
rect 8255 5182 8305 5224
rect 1209 4933 1259 4975
rect 1427 4933 1477 4975
rect 1635 4933 1685 4975
rect 2363 4947 2413 4989
rect 2571 4947 2621 4989
rect 2789 4947 2839 4989
rect 5573 4946 5623 4988
rect 5791 4946 5841 4988
rect 5999 4946 6049 4988
rect 6727 4960 6777 5002
rect 6935 4960 6985 5002
rect 7153 4960 7203 5002
rect 412 4705 462 4747
rect 630 4705 680 4747
rect 838 4705 888 4747
rect 4776 4718 4826 4760
rect 4994 4718 5044 4760
rect 5202 4718 5252 4760
rect 3445 4563 3495 4605
rect 3653 4563 3703 4605
rect 3871 4563 3921 4605
rect 7809 4576 7859 4618
rect 8017 4576 8067 4618
rect 8235 4576 8285 4618
rect 1494 4321 1544 4363
rect 1712 4321 1762 4363
rect 1920 4321 1970 4363
rect 2648 4335 2698 4377
rect 2856 4335 2906 4377
rect 3074 4335 3124 4377
rect 5858 4334 5908 4376
rect 6076 4334 6126 4376
rect 6284 4334 6334 4376
rect 7012 4348 7062 4390
rect 7220 4348 7270 4390
rect 7438 4348 7488 4390
rect 392 4099 442 4141
rect 610 4099 660 4141
rect 818 4099 868 4141
rect 3446 4151 3496 4193
rect 3654 4151 3704 4193
rect 3872 4151 3922 4193
rect 4756 4112 4806 4154
rect 4974 4112 5024 4154
rect 5182 4112 5232 4154
rect 7810 4164 7860 4206
rect 8018 4164 8068 4206
rect 8236 4164 8286 4206
rect 1190 3915 1240 3957
rect 1408 3915 1458 3957
rect 1616 3915 1666 3957
rect 2549 3925 2599 3967
rect 2757 3925 2807 3967
rect 2975 3925 3025 3967
rect 5554 3928 5604 3970
rect 5772 3928 5822 3970
rect 5980 3928 6030 3970
rect 6913 3938 6963 3980
rect 7121 3938 7171 3980
rect 7339 3938 7389 3980
rect 393 3687 443 3729
rect 611 3687 661 3729
rect 819 3687 869 3729
rect 4757 3700 4807 3742
rect 4975 3700 5025 3742
rect 5183 3700 5233 3742
rect 3428 3545 3478 3587
rect 3636 3545 3686 3587
rect 3854 3545 3904 3587
rect 7792 3558 7842 3600
rect 8000 3558 8050 3600
rect 8218 3558 8268 3600
rect 1272 3307 1322 3349
rect 1490 3307 1540 3349
rect 1698 3307 1748 3349
rect 2631 3317 2681 3359
rect 2839 3317 2889 3359
rect 3057 3317 3107 3359
rect 5636 3320 5686 3362
rect 5854 3320 5904 3362
rect 6062 3320 6112 3362
rect 6995 3330 7045 3372
rect 7203 3330 7253 3372
rect 7421 3330 7471 3372
rect 375 3081 425 3123
rect 593 3081 643 3123
rect 801 3081 851 3123
rect 3429 3133 3479 3175
rect 3637 3133 3687 3175
rect 3855 3133 3905 3175
rect 4739 3094 4789 3136
rect 4957 3094 5007 3136
rect 5165 3094 5215 3136
rect 7793 3146 7843 3188
rect 8001 3146 8051 3188
rect 8219 3146 8269 3188
rect 1173 2897 1223 2939
rect 1391 2897 1441 2939
rect 1599 2897 1649 2939
rect 2466 2909 2516 2951
rect 2674 2909 2724 2951
rect 2892 2909 2942 2951
rect 5537 2910 5587 2952
rect 5755 2910 5805 2952
rect 5963 2910 6013 2952
rect 6830 2922 6880 2964
rect 7038 2922 7088 2964
rect 7256 2922 7306 2964
rect 376 2669 426 2711
rect 594 2669 644 2711
rect 802 2669 852 2711
rect 4740 2682 4790 2724
rect 4958 2682 5008 2724
rect 5166 2682 5216 2724
rect 3408 2527 3458 2569
rect 3616 2527 3666 2569
rect 3834 2527 3884 2569
rect 7772 2540 7822 2582
rect 7980 2540 8030 2582
rect 8198 2540 8248 2582
rect 1318 2287 1368 2329
rect 1536 2287 1586 2329
rect 1744 2287 1794 2329
rect 2611 2299 2661 2341
rect 2819 2299 2869 2341
rect 3037 2299 3087 2341
rect 5682 2300 5732 2342
rect 5900 2300 5950 2342
rect 6108 2300 6158 2342
rect 6975 2312 7025 2354
rect 7183 2312 7233 2354
rect 7401 2312 7451 2354
rect 355 2063 405 2105
rect 573 2063 623 2105
rect 781 2063 831 2105
rect 3409 2115 3459 2157
rect 3617 2115 3667 2157
rect 3835 2115 3885 2157
rect 4719 2076 4769 2118
rect 4937 2076 4987 2118
rect 5145 2076 5195 2118
rect 7773 2128 7823 2170
rect 7981 2128 8031 2170
rect 8199 2128 8249 2170
rect 1153 1879 1203 1921
rect 1371 1879 1421 1921
rect 1579 1879 1629 1921
rect 2512 1889 2562 1931
rect 2720 1889 2770 1931
rect 2938 1889 2988 1931
rect 5517 1892 5567 1934
rect 5735 1892 5785 1934
rect 5943 1892 5993 1934
rect 6876 1902 6926 1944
rect 7084 1902 7134 1944
rect 7302 1902 7352 1944
rect 356 1651 406 1693
rect 574 1651 624 1693
rect 782 1651 832 1693
rect 4720 1664 4770 1706
rect 4938 1664 4988 1706
rect 5146 1664 5196 1706
rect 3391 1509 3441 1551
rect 3599 1509 3649 1551
rect 3817 1509 3867 1551
rect 7755 1522 7805 1564
rect 7963 1522 8013 1564
rect 8181 1522 8231 1564
rect 1235 1271 1285 1313
rect 1453 1271 1503 1313
rect 1661 1271 1711 1313
rect 2594 1281 2644 1323
rect 2802 1281 2852 1323
rect 3020 1281 3070 1323
rect 5599 1284 5649 1326
rect 5817 1284 5867 1326
rect 6025 1284 6075 1326
rect 6958 1294 7008 1336
rect 7166 1294 7216 1336
rect 7384 1294 7434 1336
rect 338 1045 388 1087
rect 556 1045 606 1087
rect 764 1045 814 1087
rect 3392 1097 3442 1139
rect 3600 1097 3650 1139
rect 3818 1097 3868 1139
rect 4702 1058 4752 1100
rect 4920 1058 4970 1100
rect 5128 1058 5178 1100
rect 7756 1110 7806 1152
rect 7964 1110 8014 1152
rect 8182 1110 8232 1152
rect 1136 861 1186 903
rect 1354 861 1404 903
rect 1562 861 1612 903
rect 5500 874 5550 916
rect 5718 874 5768 916
rect 5926 874 5976 916
rect 339 633 389 675
rect 557 633 607 675
rect 765 633 815 675
rect 4703 646 4753 688
rect 4921 646 4971 688
rect 5129 646 5179 688
rect 1552 57 1602 99
rect 1770 57 1820 99
rect 1978 57 2028 99
rect 5916 70 5966 112
rect 6134 70 6184 112
rect 6342 70 6392 112
rect 4041 -17 4091 25
rect 4259 -17 4309 25
rect 4467 -17 4517 25
<< pmos >>
rect 3518 8458 3568 8558
rect 3726 8458 3776 8558
rect 3944 8458 3994 8558
rect 7882 8471 7932 8571
rect 8090 8471 8140 8571
rect 8308 8471 8358 8571
rect 465 8290 515 8390
rect 683 8290 733 8390
rect 891 8290 941 8390
rect 2721 8230 2771 8330
rect 2929 8230 2979 8330
rect 3147 8230 3197 8330
rect 4829 8303 4879 8403
rect 5047 8303 5097 8403
rect 5255 8303 5305 8403
rect 1263 8106 1313 8206
rect 1481 8106 1531 8206
rect 1689 8106 1739 8206
rect 7085 8243 7135 8343
rect 7293 8243 7343 8343
rect 7511 8243 7561 8343
rect 3519 8046 3569 8146
rect 3727 8046 3777 8146
rect 3945 8046 3995 8146
rect 5627 8119 5677 8219
rect 5845 8119 5895 8219
rect 6053 8119 6103 8219
rect 7883 8059 7933 8159
rect 8091 8059 8141 8159
rect 8309 8059 8359 8159
rect 466 7878 516 7978
rect 684 7878 734 7978
rect 892 7878 942 7978
rect 2622 7820 2672 7920
rect 2830 7820 2880 7920
rect 3048 7820 3098 7920
rect 4830 7891 4880 7991
rect 5048 7891 5098 7991
rect 5256 7891 5306 7991
rect 6986 7833 7036 7933
rect 7194 7833 7244 7933
rect 7412 7833 7462 7933
rect 1345 7498 1395 7598
rect 1563 7498 1613 7598
rect 1771 7498 1821 7598
rect 3501 7440 3551 7540
rect 3709 7440 3759 7540
rect 3927 7440 3977 7540
rect 5709 7511 5759 7611
rect 5927 7511 5977 7611
rect 6135 7511 6185 7611
rect 7865 7453 7915 7553
rect 8073 7453 8123 7553
rect 8291 7453 8341 7553
rect 448 7272 498 7372
rect 666 7272 716 7372
rect 874 7272 924 7372
rect 2704 7212 2754 7312
rect 2912 7212 2962 7312
rect 3130 7212 3180 7312
rect 4812 7285 4862 7385
rect 5030 7285 5080 7385
rect 5238 7285 5288 7385
rect 1246 7088 1296 7188
rect 1464 7088 1514 7188
rect 1672 7088 1722 7188
rect 7068 7225 7118 7325
rect 7276 7225 7326 7325
rect 7494 7225 7544 7325
rect 3502 7028 3552 7128
rect 3710 7028 3760 7128
rect 3928 7028 3978 7128
rect 5610 7101 5660 7201
rect 5828 7101 5878 7201
rect 6036 7101 6086 7201
rect 7866 7041 7916 7141
rect 8074 7041 8124 7141
rect 8292 7041 8342 7141
rect 449 6860 499 6960
rect 667 6860 717 6960
rect 875 6860 925 6960
rect 2539 6804 2589 6904
rect 2747 6804 2797 6904
rect 2965 6804 3015 6904
rect 4813 6873 4863 6973
rect 5031 6873 5081 6973
rect 5239 6873 5289 6973
rect 6903 6817 6953 6917
rect 7111 6817 7161 6917
rect 7329 6817 7379 6917
rect 1391 6478 1441 6578
rect 1609 6478 1659 6578
rect 1817 6478 1867 6578
rect 3481 6422 3531 6522
rect 3689 6422 3739 6522
rect 3907 6422 3957 6522
rect 5755 6491 5805 6591
rect 5973 6491 6023 6591
rect 6181 6491 6231 6591
rect 7845 6435 7895 6535
rect 8053 6435 8103 6535
rect 8271 6435 8321 6535
rect 428 6254 478 6354
rect 646 6254 696 6354
rect 854 6254 904 6354
rect 2684 6194 2734 6294
rect 2892 6194 2942 6294
rect 3110 6194 3160 6294
rect 4792 6267 4842 6367
rect 5010 6267 5060 6367
rect 5218 6267 5268 6367
rect 1226 6070 1276 6170
rect 1444 6070 1494 6170
rect 1652 6070 1702 6170
rect 7048 6207 7098 6307
rect 7256 6207 7306 6307
rect 7474 6207 7524 6307
rect 3482 6010 3532 6110
rect 3690 6010 3740 6110
rect 3908 6010 3958 6110
rect 5590 6083 5640 6183
rect 5808 6083 5858 6183
rect 6016 6083 6066 6183
rect 7846 6023 7896 6123
rect 8054 6023 8104 6123
rect 8272 6023 8322 6123
rect 429 5842 479 5942
rect 647 5842 697 5942
rect 855 5842 905 5942
rect 2585 5784 2635 5884
rect 2793 5784 2843 5884
rect 3011 5784 3061 5884
rect 4793 5855 4843 5955
rect 5011 5855 5061 5955
rect 5219 5855 5269 5955
rect 6949 5797 6999 5897
rect 7157 5797 7207 5897
rect 7375 5797 7425 5897
rect 1308 5462 1358 5562
rect 1526 5462 1576 5562
rect 1734 5462 1784 5562
rect 3464 5404 3514 5504
rect 3672 5404 3722 5504
rect 3890 5404 3940 5504
rect 5672 5475 5722 5575
rect 5890 5475 5940 5575
rect 6098 5475 6148 5575
rect 7828 5417 7878 5517
rect 8036 5417 8086 5517
rect 8254 5417 8304 5517
rect 411 5236 461 5336
rect 629 5236 679 5336
rect 837 5236 887 5336
rect 2667 5176 2717 5276
rect 2875 5176 2925 5276
rect 3093 5176 3143 5276
rect 4775 5249 4825 5349
rect 4993 5249 5043 5349
rect 5201 5249 5251 5349
rect 1209 5052 1259 5152
rect 1427 5052 1477 5152
rect 1635 5052 1685 5152
rect 7031 5189 7081 5289
rect 7239 5189 7289 5289
rect 7457 5189 7507 5289
rect 3465 4992 3515 5092
rect 3673 4992 3723 5092
rect 3891 4992 3941 5092
rect 5573 5065 5623 5165
rect 5791 5065 5841 5165
rect 5999 5065 6049 5165
rect 7829 5005 7879 5105
rect 8037 5005 8087 5105
rect 8255 5005 8305 5105
rect 412 4824 462 4924
rect 630 4824 680 4924
rect 838 4824 888 4924
rect 2363 4770 2413 4870
rect 2571 4770 2621 4870
rect 2789 4770 2839 4870
rect 4776 4837 4826 4937
rect 4994 4837 5044 4937
rect 5202 4837 5252 4937
rect 6727 4783 6777 4883
rect 6935 4783 6985 4883
rect 7153 4783 7203 4883
rect 1494 4440 1544 4540
rect 1712 4440 1762 4540
rect 1920 4440 1970 4540
rect 3445 4386 3495 4486
rect 3653 4386 3703 4486
rect 3871 4386 3921 4486
rect 5858 4453 5908 4553
rect 6076 4453 6126 4553
rect 6284 4453 6334 4553
rect 7809 4399 7859 4499
rect 8017 4399 8067 4499
rect 8235 4399 8285 4499
rect 392 4218 442 4318
rect 610 4218 660 4318
rect 818 4218 868 4318
rect 2648 4158 2698 4258
rect 2856 4158 2906 4258
rect 3074 4158 3124 4258
rect 4756 4231 4806 4331
rect 4974 4231 5024 4331
rect 5182 4231 5232 4331
rect 1190 4034 1240 4134
rect 1408 4034 1458 4134
rect 1616 4034 1666 4134
rect 7012 4171 7062 4271
rect 7220 4171 7270 4271
rect 7438 4171 7488 4271
rect 3446 3974 3496 4074
rect 3654 3974 3704 4074
rect 3872 3974 3922 4074
rect 5554 4047 5604 4147
rect 5772 4047 5822 4147
rect 5980 4047 6030 4147
rect 7810 3987 7860 4087
rect 8018 3987 8068 4087
rect 8236 3987 8286 4087
rect 393 3806 443 3906
rect 611 3806 661 3906
rect 819 3806 869 3906
rect 2549 3748 2599 3848
rect 2757 3748 2807 3848
rect 2975 3748 3025 3848
rect 4757 3819 4807 3919
rect 4975 3819 5025 3919
rect 5183 3819 5233 3919
rect 6913 3761 6963 3861
rect 7121 3761 7171 3861
rect 7339 3761 7389 3861
rect 1272 3426 1322 3526
rect 1490 3426 1540 3526
rect 1698 3426 1748 3526
rect 3428 3368 3478 3468
rect 3636 3368 3686 3468
rect 3854 3368 3904 3468
rect 5636 3439 5686 3539
rect 5854 3439 5904 3539
rect 6062 3439 6112 3539
rect 7792 3381 7842 3481
rect 8000 3381 8050 3481
rect 8218 3381 8268 3481
rect 375 3200 425 3300
rect 593 3200 643 3300
rect 801 3200 851 3300
rect 2631 3140 2681 3240
rect 2839 3140 2889 3240
rect 3057 3140 3107 3240
rect 4739 3213 4789 3313
rect 4957 3213 5007 3313
rect 5165 3213 5215 3313
rect 1173 3016 1223 3116
rect 1391 3016 1441 3116
rect 1599 3016 1649 3116
rect 6995 3153 7045 3253
rect 7203 3153 7253 3253
rect 7421 3153 7471 3253
rect 3429 2956 3479 3056
rect 3637 2956 3687 3056
rect 3855 2956 3905 3056
rect 5537 3029 5587 3129
rect 5755 3029 5805 3129
rect 5963 3029 6013 3129
rect 7793 2969 7843 3069
rect 8001 2969 8051 3069
rect 8219 2969 8269 3069
rect 376 2788 426 2888
rect 594 2788 644 2888
rect 802 2788 852 2888
rect 2466 2732 2516 2832
rect 2674 2732 2724 2832
rect 2892 2732 2942 2832
rect 4740 2801 4790 2901
rect 4958 2801 5008 2901
rect 5166 2801 5216 2901
rect 6830 2745 6880 2845
rect 7038 2745 7088 2845
rect 7256 2745 7306 2845
rect 1318 2406 1368 2506
rect 1536 2406 1586 2506
rect 1744 2406 1794 2506
rect 3408 2350 3458 2450
rect 3616 2350 3666 2450
rect 3834 2350 3884 2450
rect 5682 2419 5732 2519
rect 5900 2419 5950 2519
rect 6108 2419 6158 2519
rect 7772 2363 7822 2463
rect 7980 2363 8030 2463
rect 8198 2363 8248 2463
rect 355 2182 405 2282
rect 573 2182 623 2282
rect 781 2182 831 2282
rect 2611 2122 2661 2222
rect 2819 2122 2869 2222
rect 3037 2122 3087 2222
rect 4719 2195 4769 2295
rect 4937 2195 4987 2295
rect 5145 2195 5195 2295
rect 1153 1998 1203 2098
rect 1371 1998 1421 2098
rect 1579 1998 1629 2098
rect 6975 2135 7025 2235
rect 7183 2135 7233 2235
rect 7401 2135 7451 2235
rect 3409 1938 3459 2038
rect 3617 1938 3667 2038
rect 3835 1938 3885 2038
rect 5517 2011 5567 2111
rect 5735 2011 5785 2111
rect 5943 2011 5993 2111
rect 7773 1951 7823 2051
rect 7981 1951 8031 2051
rect 8199 1951 8249 2051
rect 356 1770 406 1870
rect 574 1770 624 1870
rect 782 1770 832 1870
rect 2512 1712 2562 1812
rect 2720 1712 2770 1812
rect 2938 1712 2988 1812
rect 4720 1783 4770 1883
rect 4938 1783 4988 1883
rect 5146 1783 5196 1883
rect 6876 1725 6926 1825
rect 7084 1725 7134 1825
rect 7302 1725 7352 1825
rect 1235 1390 1285 1490
rect 1453 1390 1503 1490
rect 1661 1390 1711 1490
rect 3391 1332 3441 1432
rect 3599 1332 3649 1432
rect 3817 1332 3867 1432
rect 5599 1403 5649 1503
rect 5817 1403 5867 1503
rect 6025 1403 6075 1503
rect 7755 1345 7805 1445
rect 7963 1345 8013 1445
rect 8181 1345 8231 1445
rect 338 1164 388 1264
rect 556 1164 606 1264
rect 764 1164 814 1264
rect 2594 1104 2644 1204
rect 2802 1104 2852 1204
rect 3020 1104 3070 1204
rect 4702 1177 4752 1277
rect 4920 1177 4970 1277
rect 5128 1177 5178 1277
rect 1136 980 1186 1080
rect 1354 980 1404 1080
rect 1562 980 1612 1080
rect 6958 1117 7008 1217
rect 7166 1117 7216 1217
rect 7384 1117 7434 1217
rect 3392 920 3442 1020
rect 3600 920 3650 1020
rect 3818 920 3868 1020
rect 5500 993 5550 1093
rect 5718 993 5768 1093
rect 5926 993 5976 1093
rect 7756 933 7806 1033
rect 7964 933 8014 1033
rect 8182 933 8232 1033
rect 339 752 389 852
rect 557 752 607 852
rect 765 752 815 852
rect 4703 765 4753 865
rect 4921 765 4971 865
rect 5129 765 5179 865
rect 1552 176 1602 276
rect 1770 176 1820 276
rect 1978 176 2028 276
rect 4041 102 4091 202
rect 4259 102 4309 202
rect 4467 102 4517 202
rect 5916 189 5966 289
rect 6134 189 6184 289
rect 6342 189 6392 289
<< ndiff >>
rect 3469 8665 3518 8677
rect 3469 8645 3480 8665
rect 3500 8645 3518 8665
rect 3469 8635 3518 8645
rect 3568 8661 3612 8677
rect 3568 8641 3583 8661
rect 3603 8641 3612 8661
rect 3568 8635 3612 8641
rect 3682 8661 3726 8677
rect 3682 8641 3691 8661
rect 3711 8641 3726 8661
rect 3682 8635 3726 8641
rect 3776 8665 3825 8677
rect 3776 8645 3794 8665
rect 3814 8645 3825 8665
rect 3776 8635 3825 8645
rect 3900 8661 3944 8677
rect 3900 8641 3909 8661
rect 3929 8641 3944 8661
rect 3900 8635 3944 8641
rect 3994 8665 4043 8677
rect 3994 8645 4012 8665
rect 4032 8645 4043 8665
rect 3994 8635 4043 8645
rect 7833 8678 7882 8690
rect 7833 8658 7844 8678
rect 7864 8658 7882 8678
rect 7833 8648 7882 8658
rect 7932 8674 7976 8690
rect 7932 8654 7947 8674
rect 7967 8654 7976 8674
rect 7932 8648 7976 8654
rect 8046 8674 8090 8690
rect 8046 8654 8055 8674
rect 8075 8654 8090 8674
rect 8046 8648 8090 8654
rect 8140 8678 8189 8690
rect 8140 8658 8158 8678
rect 8178 8658 8189 8678
rect 8140 8648 8189 8658
rect 8264 8674 8308 8690
rect 8264 8654 8273 8674
rect 8293 8654 8308 8674
rect 8264 8648 8308 8654
rect 8358 8678 8407 8690
rect 8358 8658 8376 8678
rect 8396 8658 8407 8678
rect 8358 8648 8407 8658
rect 2672 8437 2721 8449
rect 2672 8417 2683 8437
rect 2703 8417 2721 8437
rect 2672 8407 2721 8417
rect 2771 8433 2815 8449
rect 2771 8413 2786 8433
rect 2806 8413 2815 8433
rect 2771 8407 2815 8413
rect 2885 8433 2929 8449
rect 2885 8413 2894 8433
rect 2914 8413 2929 8433
rect 2885 8407 2929 8413
rect 2979 8437 3028 8449
rect 2979 8417 2997 8437
rect 3017 8417 3028 8437
rect 2979 8407 3028 8417
rect 3103 8433 3147 8449
rect 3103 8413 3112 8433
rect 3132 8413 3147 8433
rect 3103 8407 3147 8413
rect 3197 8437 3246 8449
rect 3197 8417 3215 8437
rect 3235 8417 3246 8437
rect 3197 8407 3246 8417
rect 7036 8450 7085 8462
rect 7036 8430 7047 8450
rect 7067 8430 7085 8450
rect 7036 8420 7085 8430
rect 7135 8446 7179 8462
rect 7135 8426 7150 8446
rect 7170 8426 7179 8446
rect 7135 8420 7179 8426
rect 7249 8446 7293 8462
rect 7249 8426 7258 8446
rect 7278 8426 7293 8446
rect 7249 8420 7293 8426
rect 7343 8450 7392 8462
rect 7343 8430 7361 8450
rect 7381 8430 7392 8450
rect 7343 8420 7392 8430
rect 7467 8446 7511 8462
rect 7467 8426 7476 8446
rect 7496 8426 7511 8446
rect 7467 8420 7511 8426
rect 7561 8450 7610 8462
rect 7561 8430 7579 8450
rect 7599 8430 7610 8450
rect 7561 8420 7610 8430
rect 3470 8253 3519 8265
rect 3470 8233 3481 8253
rect 3501 8233 3519 8253
rect 416 8203 465 8213
rect 416 8183 427 8203
rect 447 8183 465 8203
rect 416 8171 465 8183
rect 515 8207 559 8213
rect 515 8187 530 8207
rect 550 8187 559 8207
rect 515 8171 559 8187
rect 634 8203 683 8213
rect 634 8183 645 8203
rect 665 8183 683 8203
rect 634 8171 683 8183
rect 733 8207 777 8213
rect 733 8187 748 8207
rect 768 8187 777 8207
rect 733 8171 777 8187
rect 847 8207 891 8213
rect 847 8187 856 8207
rect 876 8187 891 8207
rect 847 8171 891 8187
rect 941 8203 990 8213
rect 3470 8223 3519 8233
rect 3569 8249 3613 8265
rect 3569 8229 3584 8249
rect 3604 8229 3613 8249
rect 3569 8223 3613 8229
rect 3683 8249 3727 8265
rect 3683 8229 3692 8249
rect 3712 8229 3727 8249
rect 3683 8223 3727 8229
rect 3777 8253 3826 8265
rect 3777 8233 3795 8253
rect 3815 8233 3826 8253
rect 3777 8223 3826 8233
rect 3901 8249 3945 8265
rect 3901 8229 3910 8249
rect 3930 8229 3945 8249
rect 3901 8223 3945 8229
rect 3995 8253 4044 8265
rect 3995 8233 4013 8253
rect 4033 8233 4044 8253
rect 3995 8223 4044 8233
rect 941 8183 959 8203
rect 979 8183 990 8203
rect 941 8171 990 8183
rect 7834 8266 7883 8278
rect 7834 8246 7845 8266
rect 7865 8246 7883 8266
rect 4780 8216 4829 8226
rect 4780 8196 4791 8216
rect 4811 8196 4829 8216
rect 4780 8184 4829 8196
rect 4879 8220 4923 8226
rect 4879 8200 4894 8220
rect 4914 8200 4923 8220
rect 4879 8184 4923 8200
rect 4998 8216 5047 8226
rect 4998 8196 5009 8216
rect 5029 8196 5047 8216
rect 4998 8184 5047 8196
rect 5097 8220 5141 8226
rect 5097 8200 5112 8220
rect 5132 8200 5141 8220
rect 5097 8184 5141 8200
rect 5211 8220 5255 8226
rect 5211 8200 5220 8220
rect 5240 8200 5255 8220
rect 5211 8184 5255 8200
rect 5305 8216 5354 8226
rect 7834 8236 7883 8246
rect 7933 8262 7977 8278
rect 7933 8242 7948 8262
rect 7968 8242 7977 8262
rect 7933 8236 7977 8242
rect 8047 8262 8091 8278
rect 8047 8242 8056 8262
rect 8076 8242 8091 8262
rect 8047 8236 8091 8242
rect 8141 8266 8190 8278
rect 8141 8246 8159 8266
rect 8179 8246 8190 8266
rect 8141 8236 8190 8246
rect 8265 8262 8309 8278
rect 8265 8242 8274 8262
rect 8294 8242 8309 8262
rect 8265 8236 8309 8242
rect 8359 8266 8408 8278
rect 8359 8246 8377 8266
rect 8397 8246 8408 8266
rect 8359 8236 8408 8246
rect 5305 8196 5323 8216
rect 5343 8196 5354 8216
rect 5305 8184 5354 8196
rect 1214 8019 1263 8029
rect 1214 7999 1225 8019
rect 1245 7999 1263 8019
rect 1214 7987 1263 7999
rect 1313 8023 1357 8029
rect 1313 8003 1328 8023
rect 1348 8003 1357 8023
rect 1313 7987 1357 8003
rect 1432 8019 1481 8029
rect 1432 7999 1443 8019
rect 1463 7999 1481 8019
rect 1432 7987 1481 7999
rect 1531 8023 1575 8029
rect 1531 8003 1546 8023
rect 1566 8003 1575 8023
rect 1531 7987 1575 8003
rect 1645 8023 1689 8029
rect 1645 8003 1654 8023
rect 1674 8003 1689 8023
rect 1645 7987 1689 8003
rect 1739 8019 1788 8029
rect 1739 7999 1757 8019
rect 1777 7999 1788 8019
rect 1739 7987 1788 7999
rect 2573 8027 2622 8039
rect 2573 8007 2584 8027
rect 2604 8007 2622 8027
rect 2573 7997 2622 8007
rect 2672 8023 2716 8039
rect 2672 8003 2687 8023
rect 2707 8003 2716 8023
rect 2672 7997 2716 8003
rect 2786 8023 2830 8039
rect 2786 8003 2795 8023
rect 2815 8003 2830 8023
rect 2786 7997 2830 8003
rect 2880 8027 2929 8039
rect 2880 8007 2898 8027
rect 2918 8007 2929 8027
rect 2880 7997 2929 8007
rect 3004 8023 3048 8039
rect 3004 8003 3013 8023
rect 3033 8003 3048 8023
rect 3004 7997 3048 8003
rect 3098 8027 3147 8039
rect 3098 8007 3116 8027
rect 3136 8007 3147 8027
rect 3098 7997 3147 8007
rect 5578 8032 5627 8042
rect 5578 8012 5589 8032
rect 5609 8012 5627 8032
rect 5578 8000 5627 8012
rect 5677 8036 5721 8042
rect 5677 8016 5692 8036
rect 5712 8016 5721 8036
rect 5677 8000 5721 8016
rect 5796 8032 5845 8042
rect 5796 8012 5807 8032
rect 5827 8012 5845 8032
rect 5796 8000 5845 8012
rect 5895 8036 5939 8042
rect 5895 8016 5910 8036
rect 5930 8016 5939 8036
rect 5895 8000 5939 8016
rect 6009 8036 6053 8042
rect 6009 8016 6018 8036
rect 6038 8016 6053 8036
rect 6009 8000 6053 8016
rect 6103 8032 6152 8042
rect 6103 8012 6121 8032
rect 6141 8012 6152 8032
rect 6103 8000 6152 8012
rect 6937 8040 6986 8052
rect 6937 8020 6948 8040
rect 6968 8020 6986 8040
rect 6937 8010 6986 8020
rect 7036 8036 7080 8052
rect 7036 8016 7051 8036
rect 7071 8016 7080 8036
rect 7036 8010 7080 8016
rect 7150 8036 7194 8052
rect 7150 8016 7159 8036
rect 7179 8016 7194 8036
rect 7150 8010 7194 8016
rect 7244 8040 7293 8052
rect 7244 8020 7262 8040
rect 7282 8020 7293 8040
rect 7244 8010 7293 8020
rect 7368 8036 7412 8052
rect 7368 8016 7377 8036
rect 7397 8016 7412 8036
rect 7368 8010 7412 8016
rect 7462 8040 7511 8052
rect 7462 8020 7480 8040
rect 7500 8020 7511 8040
rect 7462 8010 7511 8020
rect 417 7791 466 7801
rect 417 7771 428 7791
rect 448 7771 466 7791
rect 417 7759 466 7771
rect 516 7795 560 7801
rect 516 7775 531 7795
rect 551 7775 560 7795
rect 516 7759 560 7775
rect 635 7791 684 7801
rect 635 7771 646 7791
rect 666 7771 684 7791
rect 635 7759 684 7771
rect 734 7795 778 7801
rect 734 7775 749 7795
rect 769 7775 778 7795
rect 734 7759 778 7775
rect 848 7795 892 7801
rect 848 7775 857 7795
rect 877 7775 892 7795
rect 848 7759 892 7775
rect 942 7791 991 7801
rect 942 7771 960 7791
rect 980 7771 991 7791
rect 942 7759 991 7771
rect 4781 7804 4830 7814
rect 4781 7784 4792 7804
rect 4812 7784 4830 7804
rect 4781 7772 4830 7784
rect 4880 7808 4924 7814
rect 4880 7788 4895 7808
rect 4915 7788 4924 7808
rect 4880 7772 4924 7788
rect 4999 7804 5048 7814
rect 4999 7784 5010 7804
rect 5030 7784 5048 7804
rect 4999 7772 5048 7784
rect 5098 7808 5142 7814
rect 5098 7788 5113 7808
rect 5133 7788 5142 7808
rect 5098 7772 5142 7788
rect 5212 7808 5256 7814
rect 5212 7788 5221 7808
rect 5241 7788 5256 7808
rect 5212 7772 5256 7788
rect 5306 7804 5355 7814
rect 5306 7784 5324 7804
rect 5344 7784 5355 7804
rect 5306 7772 5355 7784
rect 3452 7647 3501 7659
rect 3452 7627 3463 7647
rect 3483 7627 3501 7647
rect 3452 7617 3501 7627
rect 3551 7643 3595 7659
rect 3551 7623 3566 7643
rect 3586 7623 3595 7643
rect 3551 7617 3595 7623
rect 3665 7643 3709 7659
rect 3665 7623 3674 7643
rect 3694 7623 3709 7643
rect 3665 7617 3709 7623
rect 3759 7647 3808 7659
rect 3759 7627 3777 7647
rect 3797 7627 3808 7647
rect 3759 7617 3808 7627
rect 3883 7643 3927 7659
rect 3883 7623 3892 7643
rect 3912 7623 3927 7643
rect 3883 7617 3927 7623
rect 3977 7647 4026 7659
rect 3977 7627 3995 7647
rect 4015 7627 4026 7647
rect 3977 7617 4026 7627
rect 7816 7660 7865 7672
rect 7816 7640 7827 7660
rect 7847 7640 7865 7660
rect 7816 7630 7865 7640
rect 7915 7656 7959 7672
rect 7915 7636 7930 7656
rect 7950 7636 7959 7656
rect 7915 7630 7959 7636
rect 8029 7656 8073 7672
rect 8029 7636 8038 7656
rect 8058 7636 8073 7656
rect 8029 7630 8073 7636
rect 8123 7660 8172 7672
rect 8123 7640 8141 7660
rect 8161 7640 8172 7660
rect 8123 7630 8172 7640
rect 8247 7656 8291 7672
rect 8247 7636 8256 7656
rect 8276 7636 8291 7656
rect 8247 7630 8291 7636
rect 8341 7660 8390 7672
rect 8341 7640 8359 7660
rect 8379 7640 8390 7660
rect 8341 7630 8390 7640
rect 1296 7411 1345 7421
rect 1296 7391 1307 7411
rect 1327 7391 1345 7411
rect 1296 7379 1345 7391
rect 1395 7415 1439 7421
rect 1395 7395 1410 7415
rect 1430 7395 1439 7415
rect 1395 7379 1439 7395
rect 1514 7411 1563 7421
rect 1514 7391 1525 7411
rect 1545 7391 1563 7411
rect 1514 7379 1563 7391
rect 1613 7415 1657 7421
rect 1613 7395 1628 7415
rect 1648 7395 1657 7415
rect 1613 7379 1657 7395
rect 1727 7415 1771 7421
rect 1727 7395 1736 7415
rect 1756 7395 1771 7415
rect 1727 7379 1771 7395
rect 1821 7411 1870 7421
rect 1821 7391 1839 7411
rect 1859 7391 1870 7411
rect 1821 7379 1870 7391
rect 2655 7419 2704 7431
rect 2655 7399 2666 7419
rect 2686 7399 2704 7419
rect 2655 7389 2704 7399
rect 2754 7415 2798 7431
rect 2754 7395 2769 7415
rect 2789 7395 2798 7415
rect 2754 7389 2798 7395
rect 2868 7415 2912 7431
rect 2868 7395 2877 7415
rect 2897 7395 2912 7415
rect 2868 7389 2912 7395
rect 2962 7419 3011 7431
rect 2962 7399 2980 7419
rect 3000 7399 3011 7419
rect 2962 7389 3011 7399
rect 3086 7415 3130 7431
rect 3086 7395 3095 7415
rect 3115 7395 3130 7415
rect 3086 7389 3130 7395
rect 3180 7419 3229 7431
rect 3180 7399 3198 7419
rect 3218 7399 3229 7419
rect 3180 7389 3229 7399
rect 5660 7424 5709 7434
rect 5660 7404 5671 7424
rect 5691 7404 5709 7424
rect 5660 7392 5709 7404
rect 5759 7428 5803 7434
rect 5759 7408 5774 7428
rect 5794 7408 5803 7428
rect 5759 7392 5803 7408
rect 5878 7424 5927 7434
rect 5878 7404 5889 7424
rect 5909 7404 5927 7424
rect 5878 7392 5927 7404
rect 5977 7428 6021 7434
rect 5977 7408 5992 7428
rect 6012 7408 6021 7428
rect 5977 7392 6021 7408
rect 6091 7428 6135 7434
rect 6091 7408 6100 7428
rect 6120 7408 6135 7428
rect 6091 7392 6135 7408
rect 6185 7424 6234 7434
rect 6185 7404 6203 7424
rect 6223 7404 6234 7424
rect 6185 7392 6234 7404
rect 7019 7432 7068 7444
rect 7019 7412 7030 7432
rect 7050 7412 7068 7432
rect 7019 7402 7068 7412
rect 7118 7428 7162 7444
rect 7118 7408 7133 7428
rect 7153 7408 7162 7428
rect 7118 7402 7162 7408
rect 7232 7428 7276 7444
rect 7232 7408 7241 7428
rect 7261 7408 7276 7428
rect 7232 7402 7276 7408
rect 7326 7432 7375 7444
rect 7326 7412 7344 7432
rect 7364 7412 7375 7432
rect 7326 7402 7375 7412
rect 7450 7428 7494 7444
rect 7450 7408 7459 7428
rect 7479 7408 7494 7428
rect 7450 7402 7494 7408
rect 7544 7432 7593 7444
rect 7544 7412 7562 7432
rect 7582 7412 7593 7432
rect 7544 7402 7593 7412
rect 3453 7235 3502 7247
rect 3453 7215 3464 7235
rect 3484 7215 3502 7235
rect 399 7185 448 7195
rect 399 7165 410 7185
rect 430 7165 448 7185
rect 399 7153 448 7165
rect 498 7189 542 7195
rect 498 7169 513 7189
rect 533 7169 542 7189
rect 498 7153 542 7169
rect 617 7185 666 7195
rect 617 7165 628 7185
rect 648 7165 666 7185
rect 617 7153 666 7165
rect 716 7189 760 7195
rect 716 7169 731 7189
rect 751 7169 760 7189
rect 716 7153 760 7169
rect 830 7189 874 7195
rect 830 7169 839 7189
rect 859 7169 874 7189
rect 830 7153 874 7169
rect 924 7185 973 7195
rect 3453 7205 3502 7215
rect 3552 7231 3596 7247
rect 3552 7211 3567 7231
rect 3587 7211 3596 7231
rect 3552 7205 3596 7211
rect 3666 7231 3710 7247
rect 3666 7211 3675 7231
rect 3695 7211 3710 7231
rect 3666 7205 3710 7211
rect 3760 7235 3809 7247
rect 3760 7215 3778 7235
rect 3798 7215 3809 7235
rect 3760 7205 3809 7215
rect 3884 7231 3928 7247
rect 3884 7211 3893 7231
rect 3913 7211 3928 7231
rect 3884 7205 3928 7211
rect 3978 7235 4027 7247
rect 3978 7215 3996 7235
rect 4016 7215 4027 7235
rect 3978 7205 4027 7215
rect 924 7165 942 7185
rect 962 7165 973 7185
rect 924 7153 973 7165
rect 7817 7248 7866 7260
rect 7817 7228 7828 7248
rect 7848 7228 7866 7248
rect 4763 7198 4812 7208
rect 4763 7178 4774 7198
rect 4794 7178 4812 7198
rect 4763 7166 4812 7178
rect 4862 7202 4906 7208
rect 4862 7182 4877 7202
rect 4897 7182 4906 7202
rect 4862 7166 4906 7182
rect 4981 7198 5030 7208
rect 4981 7178 4992 7198
rect 5012 7178 5030 7198
rect 4981 7166 5030 7178
rect 5080 7202 5124 7208
rect 5080 7182 5095 7202
rect 5115 7182 5124 7202
rect 5080 7166 5124 7182
rect 5194 7202 5238 7208
rect 5194 7182 5203 7202
rect 5223 7182 5238 7202
rect 5194 7166 5238 7182
rect 5288 7198 5337 7208
rect 7817 7218 7866 7228
rect 7916 7244 7960 7260
rect 7916 7224 7931 7244
rect 7951 7224 7960 7244
rect 7916 7218 7960 7224
rect 8030 7244 8074 7260
rect 8030 7224 8039 7244
rect 8059 7224 8074 7244
rect 8030 7218 8074 7224
rect 8124 7248 8173 7260
rect 8124 7228 8142 7248
rect 8162 7228 8173 7248
rect 8124 7218 8173 7228
rect 8248 7244 8292 7260
rect 8248 7224 8257 7244
rect 8277 7224 8292 7244
rect 8248 7218 8292 7224
rect 8342 7248 8391 7260
rect 8342 7228 8360 7248
rect 8380 7228 8391 7248
rect 8342 7218 8391 7228
rect 5288 7178 5306 7198
rect 5326 7178 5337 7198
rect 5288 7166 5337 7178
rect 2490 7011 2539 7023
rect 1197 7001 1246 7011
rect 1197 6981 1208 7001
rect 1228 6981 1246 7001
rect 1197 6969 1246 6981
rect 1296 7005 1340 7011
rect 1296 6985 1311 7005
rect 1331 6985 1340 7005
rect 1296 6969 1340 6985
rect 1415 7001 1464 7011
rect 1415 6981 1426 7001
rect 1446 6981 1464 7001
rect 1415 6969 1464 6981
rect 1514 7005 1558 7011
rect 1514 6985 1529 7005
rect 1549 6985 1558 7005
rect 1514 6969 1558 6985
rect 1628 7005 1672 7011
rect 1628 6985 1637 7005
rect 1657 6985 1672 7005
rect 1628 6969 1672 6985
rect 1722 7001 1771 7011
rect 1722 6981 1740 7001
rect 1760 6981 1771 7001
rect 2490 6991 2501 7011
rect 2521 6991 2539 7011
rect 2490 6981 2539 6991
rect 2589 7007 2633 7023
rect 2589 6987 2604 7007
rect 2624 6987 2633 7007
rect 2589 6981 2633 6987
rect 2703 7007 2747 7023
rect 2703 6987 2712 7007
rect 2732 6987 2747 7007
rect 2703 6981 2747 6987
rect 2797 7011 2846 7023
rect 2797 6991 2815 7011
rect 2835 6991 2846 7011
rect 2797 6981 2846 6991
rect 2921 7007 2965 7023
rect 2921 6987 2930 7007
rect 2950 6987 2965 7007
rect 2921 6981 2965 6987
rect 3015 7011 3064 7023
rect 6854 7024 6903 7036
rect 3015 6991 3033 7011
rect 3053 6991 3064 7011
rect 3015 6981 3064 6991
rect 1722 6969 1771 6981
rect 5561 7014 5610 7024
rect 5561 6994 5572 7014
rect 5592 6994 5610 7014
rect 5561 6982 5610 6994
rect 5660 7018 5704 7024
rect 5660 6998 5675 7018
rect 5695 6998 5704 7018
rect 5660 6982 5704 6998
rect 5779 7014 5828 7024
rect 5779 6994 5790 7014
rect 5810 6994 5828 7014
rect 5779 6982 5828 6994
rect 5878 7018 5922 7024
rect 5878 6998 5893 7018
rect 5913 6998 5922 7018
rect 5878 6982 5922 6998
rect 5992 7018 6036 7024
rect 5992 6998 6001 7018
rect 6021 6998 6036 7018
rect 5992 6982 6036 6998
rect 6086 7014 6135 7024
rect 6086 6994 6104 7014
rect 6124 6994 6135 7014
rect 6854 7004 6865 7024
rect 6885 7004 6903 7024
rect 6854 6994 6903 7004
rect 6953 7020 6997 7036
rect 6953 7000 6968 7020
rect 6988 7000 6997 7020
rect 6953 6994 6997 7000
rect 7067 7020 7111 7036
rect 7067 7000 7076 7020
rect 7096 7000 7111 7020
rect 7067 6994 7111 7000
rect 7161 7024 7210 7036
rect 7161 7004 7179 7024
rect 7199 7004 7210 7024
rect 7161 6994 7210 7004
rect 7285 7020 7329 7036
rect 7285 7000 7294 7020
rect 7314 7000 7329 7020
rect 7285 6994 7329 7000
rect 7379 7024 7428 7036
rect 7379 7004 7397 7024
rect 7417 7004 7428 7024
rect 7379 6994 7428 7004
rect 6086 6982 6135 6994
rect 400 6773 449 6783
rect 400 6753 411 6773
rect 431 6753 449 6773
rect 400 6741 449 6753
rect 499 6777 543 6783
rect 499 6757 514 6777
rect 534 6757 543 6777
rect 499 6741 543 6757
rect 618 6773 667 6783
rect 618 6753 629 6773
rect 649 6753 667 6773
rect 618 6741 667 6753
rect 717 6777 761 6783
rect 717 6757 732 6777
rect 752 6757 761 6777
rect 717 6741 761 6757
rect 831 6777 875 6783
rect 831 6757 840 6777
rect 860 6757 875 6777
rect 831 6741 875 6757
rect 925 6773 974 6783
rect 925 6753 943 6773
rect 963 6753 974 6773
rect 925 6741 974 6753
rect 4764 6786 4813 6796
rect 4764 6766 4775 6786
rect 4795 6766 4813 6786
rect 4764 6754 4813 6766
rect 4863 6790 4907 6796
rect 4863 6770 4878 6790
rect 4898 6770 4907 6790
rect 4863 6754 4907 6770
rect 4982 6786 5031 6796
rect 4982 6766 4993 6786
rect 5013 6766 5031 6786
rect 4982 6754 5031 6766
rect 5081 6790 5125 6796
rect 5081 6770 5096 6790
rect 5116 6770 5125 6790
rect 5081 6754 5125 6770
rect 5195 6790 5239 6796
rect 5195 6770 5204 6790
rect 5224 6770 5239 6790
rect 5195 6754 5239 6770
rect 5289 6786 5338 6796
rect 5289 6766 5307 6786
rect 5327 6766 5338 6786
rect 5289 6754 5338 6766
rect 3432 6629 3481 6641
rect 3432 6609 3443 6629
rect 3463 6609 3481 6629
rect 3432 6599 3481 6609
rect 3531 6625 3575 6641
rect 3531 6605 3546 6625
rect 3566 6605 3575 6625
rect 3531 6599 3575 6605
rect 3645 6625 3689 6641
rect 3645 6605 3654 6625
rect 3674 6605 3689 6625
rect 3645 6599 3689 6605
rect 3739 6629 3788 6641
rect 3739 6609 3757 6629
rect 3777 6609 3788 6629
rect 3739 6599 3788 6609
rect 3863 6625 3907 6641
rect 3863 6605 3872 6625
rect 3892 6605 3907 6625
rect 3863 6599 3907 6605
rect 3957 6629 4006 6641
rect 3957 6609 3975 6629
rect 3995 6609 4006 6629
rect 3957 6599 4006 6609
rect 7796 6642 7845 6654
rect 7796 6622 7807 6642
rect 7827 6622 7845 6642
rect 7796 6612 7845 6622
rect 7895 6638 7939 6654
rect 7895 6618 7910 6638
rect 7930 6618 7939 6638
rect 7895 6612 7939 6618
rect 8009 6638 8053 6654
rect 8009 6618 8018 6638
rect 8038 6618 8053 6638
rect 8009 6612 8053 6618
rect 8103 6642 8152 6654
rect 8103 6622 8121 6642
rect 8141 6622 8152 6642
rect 8103 6612 8152 6622
rect 8227 6638 8271 6654
rect 8227 6618 8236 6638
rect 8256 6618 8271 6638
rect 8227 6612 8271 6618
rect 8321 6642 8370 6654
rect 8321 6622 8339 6642
rect 8359 6622 8370 6642
rect 8321 6612 8370 6622
rect 2635 6401 2684 6413
rect 1342 6391 1391 6401
rect 1342 6371 1353 6391
rect 1373 6371 1391 6391
rect 1342 6359 1391 6371
rect 1441 6395 1485 6401
rect 1441 6375 1456 6395
rect 1476 6375 1485 6395
rect 1441 6359 1485 6375
rect 1560 6391 1609 6401
rect 1560 6371 1571 6391
rect 1591 6371 1609 6391
rect 1560 6359 1609 6371
rect 1659 6395 1703 6401
rect 1659 6375 1674 6395
rect 1694 6375 1703 6395
rect 1659 6359 1703 6375
rect 1773 6395 1817 6401
rect 1773 6375 1782 6395
rect 1802 6375 1817 6395
rect 1773 6359 1817 6375
rect 1867 6391 1916 6401
rect 1867 6371 1885 6391
rect 1905 6371 1916 6391
rect 2635 6381 2646 6401
rect 2666 6381 2684 6401
rect 2635 6371 2684 6381
rect 2734 6397 2778 6413
rect 2734 6377 2749 6397
rect 2769 6377 2778 6397
rect 2734 6371 2778 6377
rect 2848 6397 2892 6413
rect 2848 6377 2857 6397
rect 2877 6377 2892 6397
rect 2848 6371 2892 6377
rect 2942 6401 2991 6413
rect 2942 6381 2960 6401
rect 2980 6381 2991 6401
rect 2942 6371 2991 6381
rect 3066 6397 3110 6413
rect 3066 6377 3075 6397
rect 3095 6377 3110 6397
rect 3066 6371 3110 6377
rect 3160 6401 3209 6413
rect 3160 6381 3178 6401
rect 3198 6381 3209 6401
rect 3160 6371 3209 6381
rect 6999 6414 7048 6426
rect 5706 6404 5755 6414
rect 5706 6384 5717 6404
rect 5737 6384 5755 6404
rect 1867 6359 1916 6371
rect 5706 6372 5755 6384
rect 5805 6408 5849 6414
rect 5805 6388 5820 6408
rect 5840 6388 5849 6408
rect 5805 6372 5849 6388
rect 5924 6404 5973 6414
rect 5924 6384 5935 6404
rect 5955 6384 5973 6404
rect 5924 6372 5973 6384
rect 6023 6408 6067 6414
rect 6023 6388 6038 6408
rect 6058 6388 6067 6408
rect 6023 6372 6067 6388
rect 6137 6408 6181 6414
rect 6137 6388 6146 6408
rect 6166 6388 6181 6408
rect 6137 6372 6181 6388
rect 6231 6404 6280 6414
rect 6231 6384 6249 6404
rect 6269 6384 6280 6404
rect 6999 6394 7010 6414
rect 7030 6394 7048 6414
rect 6999 6384 7048 6394
rect 7098 6410 7142 6426
rect 7098 6390 7113 6410
rect 7133 6390 7142 6410
rect 7098 6384 7142 6390
rect 7212 6410 7256 6426
rect 7212 6390 7221 6410
rect 7241 6390 7256 6410
rect 7212 6384 7256 6390
rect 7306 6414 7355 6426
rect 7306 6394 7324 6414
rect 7344 6394 7355 6414
rect 7306 6384 7355 6394
rect 7430 6410 7474 6426
rect 7430 6390 7439 6410
rect 7459 6390 7474 6410
rect 7430 6384 7474 6390
rect 7524 6414 7573 6426
rect 7524 6394 7542 6414
rect 7562 6394 7573 6414
rect 7524 6384 7573 6394
rect 6231 6372 6280 6384
rect 3433 6217 3482 6229
rect 3433 6197 3444 6217
rect 3464 6197 3482 6217
rect 379 6167 428 6177
rect 379 6147 390 6167
rect 410 6147 428 6167
rect 379 6135 428 6147
rect 478 6171 522 6177
rect 478 6151 493 6171
rect 513 6151 522 6171
rect 478 6135 522 6151
rect 597 6167 646 6177
rect 597 6147 608 6167
rect 628 6147 646 6167
rect 597 6135 646 6147
rect 696 6171 740 6177
rect 696 6151 711 6171
rect 731 6151 740 6171
rect 696 6135 740 6151
rect 810 6171 854 6177
rect 810 6151 819 6171
rect 839 6151 854 6171
rect 810 6135 854 6151
rect 904 6167 953 6177
rect 3433 6187 3482 6197
rect 3532 6213 3576 6229
rect 3532 6193 3547 6213
rect 3567 6193 3576 6213
rect 3532 6187 3576 6193
rect 3646 6213 3690 6229
rect 3646 6193 3655 6213
rect 3675 6193 3690 6213
rect 3646 6187 3690 6193
rect 3740 6217 3789 6229
rect 3740 6197 3758 6217
rect 3778 6197 3789 6217
rect 3740 6187 3789 6197
rect 3864 6213 3908 6229
rect 3864 6193 3873 6213
rect 3893 6193 3908 6213
rect 3864 6187 3908 6193
rect 3958 6217 4007 6229
rect 3958 6197 3976 6217
rect 3996 6197 4007 6217
rect 3958 6187 4007 6197
rect 904 6147 922 6167
rect 942 6147 953 6167
rect 904 6135 953 6147
rect 7797 6230 7846 6242
rect 7797 6210 7808 6230
rect 7828 6210 7846 6230
rect 4743 6180 4792 6190
rect 4743 6160 4754 6180
rect 4774 6160 4792 6180
rect 4743 6148 4792 6160
rect 4842 6184 4886 6190
rect 4842 6164 4857 6184
rect 4877 6164 4886 6184
rect 4842 6148 4886 6164
rect 4961 6180 5010 6190
rect 4961 6160 4972 6180
rect 4992 6160 5010 6180
rect 4961 6148 5010 6160
rect 5060 6184 5104 6190
rect 5060 6164 5075 6184
rect 5095 6164 5104 6184
rect 5060 6148 5104 6164
rect 5174 6184 5218 6190
rect 5174 6164 5183 6184
rect 5203 6164 5218 6184
rect 5174 6148 5218 6164
rect 5268 6180 5317 6190
rect 7797 6200 7846 6210
rect 7896 6226 7940 6242
rect 7896 6206 7911 6226
rect 7931 6206 7940 6226
rect 7896 6200 7940 6206
rect 8010 6226 8054 6242
rect 8010 6206 8019 6226
rect 8039 6206 8054 6226
rect 8010 6200 8054 6206
rect 8104 6230 8153 6242
rect 8104 6210 8122 6230
rect 8142 6210 8153 6230
rect 8104 6200 8153 6210
rect 8228 6226 8272 6242
rect 8228 6206 8237 6226
rect 8257 6206 8272 6226
rect 8228 6200 8272 6206
rect 8322 6230 8371 6242
rect 8322 6210 8340 6230
rect 8360 6210 8371 6230
rect 8322 6200 8371 6210
rect 5268 6160 5286 6180
rect 5306 6160 5317 6180
rect 5268 6148 5317 6160
rect 1177 5983 1226 5993
rect 1177 5963 1188 5983
rect 1208 5963 1226 5983
rect 1177 5951 1226 5963
rect 1276 5987 1320 5993
rect 1276 5967 1291 5987
rect 1311 5967 1320 5987
rect 1276 5951 1320 5967
rect 1395 5983 1444 5993
rect 1395 5963 1406 5983
rect 1426 5963 1444 5983
rect 1395 5951 1444 5963
rect 1494 5987 1538 5993
rect 1494 5967 1509 5987
rect 1529 5967 1538 5987
rect 1494 5951 1538 5967
rect 1608 5987 1652 5993
rect 1608 5967 1617 5987
rect 1637 5967 1652 5987
rect 1608 5951 1652 5967
rect 1702 5983 1751 5993
rect 1702 5963 1720 5983
rect 1740 5963 1751 5983
rect 1702 5951 1751 5963
rect 2536 5991 2585 6003
rect 2536 5971 2547 5991
rect 2567 5971 2585 5991
rect 2536 5961 2585 5971
rect 2635 5987 2679 6003
rect 2635 5967 2650 5987
rect 2670 5967 2679 5987
rect 2635 5961 2679 5967
rect 2749 5987 2793 6003
rect 2749 5967 2758 5987
rect 2778 5967 2793 5987
rect 2749 5961 2793 5967
rect 2843 5991 2892 6003
rect 2843 5971 2861 5991
rect 2881 5971 2892 5991
rect 2843 5961 2892 5971
rect 2967 5987 3011 6003
rect 2967 5967 2976 5987
rect 2996 5967 3011 5987
rect 2967 5961 3011 5967
rect 3061 5991 3110 6003
rect 3061 5971 3079 5991
rect 3099 5971 3110 5991
rect 3061 5961 3110 5971
rect 5541 5996 5590 6006
rect 5541 5976 5552 5996
rect 5572 5976 5590 5996
rect 5541 5964 5590 5976
rect 5640 6000 5684 6006
rect 5640 5980 5655 6000
rect 5675 5980 5684 6000
rect 5640 5964 5684 5980
rect 5759 5996 5808 6006
rect 5759 5976 5770 5996
rect 5790 5976 5808 5996
rect 5759 5964 5808 5976
rect 5858 6000 5902 6006
rect 5858 5980 5873 6000
rect 5893 5980 5902 6000
rect 5858 5964 5902 5980
rect 5972 6000 6016 6006
rect 5972 5980 5981 6000
rect 6001 5980 6016 6000
rect 5972 5964 6016 5980
rect 6066 5996 6115 6006
rect 6066 5976 6084 5996
rect 6104 5976 6115 5996
rect 6066 5964 6115 5976
rect 6900 6004 6949 6016
rect 6900 5984 6911 6004
rect 6931 5984 6949 6004
rect 6900 5974 6949 5984
rect 6999 6000 7043 6016
rect 6999 5980 7014 6000
rect 7034 5980 7043 6000
rect 6999 5974 7043 5980
rect 7113 6000 7157 6016
rect 7113 5980 7122 6000
rect 7142 5980 7157 6000
rect 7113 5974 7157 5980
rect 7207 6004 7256 6016
rect 7207 5984 7225 6004
rect 7245 5984 7256 6004
rect 7207 5974 7256 5984
rect 7331 6000 7375 6016
rect 7331 5980 7340 6000
rect 7360 5980 7375 6000
rect 7331 5974 7375 5980
rect 7425 6004 7474 6016
rect 7425 5984 7443 6004
rect 7463 5984 7474 6004
rect 7425 5974 7474 5984
rect 380 5755 429 5765
rect 380 5735 391 5755
rect 411 5735 429 5755
rect 380 5723 429 5735
rect 479 5759 523 5765
rect 479 5739 494 5759
rect 514 5739 523 5759
rect 479 5723 523 5739
rect 598 5755 647 5765
rect 598 5735 609 5755
rect 629 5735 647 5755
rect 598 5723 647 5735
rect 697 5759 741 5765
rect 697 5739 712 5759
rect 732 5739 741 5759
rect 697 5723 741 5739
rect 811 5759 855 5765
rect 811 5739 820 5759
rect 840 5739 855 5759
rect 811 5723 855 5739
rect 905 5755 954 5765
rect 905 5735 923 5755
rect 943 5735 954 5755
rect 905 5723 954 5735
rect 4744 5768 4793 5778
rect 4744 5748 4755 5768
rect 4775 5748 4793 5768
rect 4744 5736 4793 5748
rect 4843 5772 4887 5778
rect 4843 5752 4858 5772
rect 4878 5752 4887 5772
rect 4843 5736 4887 5752
rect 4962 5768 5011 5778
rect 4962 5748 4973 5768
rect 4993 5748 5011 5768
rect 4962 5736 5011 5748
rect 5061 5772 5105 5778
rect 5061 5752 5076 5772
rect 5096 5752 5105 5772
rect 5061 5736 5105 5752
rect 5175 5772 5219 5778
rect 5175 5752 5184 5772
rect 5204 5752 5219 5772
rect 5175 5736 5219 5752
rect 5269 5768 5318 5778
rect 5269 5748 5287 5768
rect 5307 5748 5318 5768
rect 5269 5736 5318 5748
rect 3415 5611 3464 5623
rect 3415 5591 3426 5611
rect 3446 5591 3464 5611
rect 3415 5581 3464 5591
rect 3514 5607 3558 5623
rect 3514 5587 3529 5607
rect 3549 5587 3558 5607
rect 3514 5581 3558 5587
rect 3628 5607 3672 5623
rect 3628 5587 3637 5607
rect 3657 5587 3672 5607
rect 3628 5581 3672 5587
rect 3722 5611 3771 5623
rect 3722 5591 3740 5611
rect 3760 5591 3771 5611
rect 3722 5581 3771 5591
rect 3846 5607 3890 5623
rect 3846 5587 3855 5607
rect 3875 5587 3890 5607
rect 3846 5581 3890 5587
rect 3940 5611 3989 5623
rect 3940 5591 3958 5611
rect 3978 5591 3989 5611
rect 3940 5581 3989 5591
rect 7779 5624 7828 5636
rect 7779 5604 7790 5624
rect 7810 5604 7828 5624
rect 7779 5594 7828 5604
rect 7878 5620 7922 5636
rect 7878 5600 7893 5620
rect 7913 5600 7922 5620
rect 7878 5594 7922 5600
rect 7992 5620 8036 5636
rect 7992 5600 8001 5620
rect 8021 5600 8036 5620
rect 7992 5594 8036 5600
rect 8086 5624 8135 5636
rect 8086 5604 8104 5624
rect 8124 5604 8135 5624
rect 8086 5594 8135 5604
rect 8210 5620 8254 5636
rect 8210 5600 8219 5620
rect 8239 5600 8254 5620
rect 8210 5594 8254 5600
rect 8304 5624 8353 5636
rect 8304 5604 8322 5624
rect 8342 5604 8353 5624
rect 8304 5594 8353 5604
rect 1259 5375 1308 5385
rect 1259 5355 1270 5375
rect 1290 5355 1308 5375
rect 1259 5343 1308 5355
rect 1358 5379 1402 5385
rect 1358 5359 1373 5379
rect 1393 5359 1402 5379
rect 1358 5343 1402 5359
rect 1477 5375 1526 5385
rect 1477 5355 1488 5375
rect 1508 5355 1526 5375
rect 1477 5343 1526 5355
rect 1576 5379 1620 5385
rect 1576 5359 1591 5379
rect 1611 5359 1620 5379
rect 1576 5343 1620 5359
rect 1690 5379 1734 5385
rect 1690 5359 1699 5379
rect 1719 5359 1734 5379
rect 1690 5343 1734 5359
rect 1784 5375 1833 5385
rect 1784 5355 1802 5375
rect 1822 5355 1833 5375
rect 1784 5343 1833 5355
rect 2618 5383 2667 5395
rect 2618 5363 2629 5383
rect 2649 5363 2667 5383
rect 2618 5353 2667 5363
rect 2717 5379 2761 5395
rect 2717 5359 2732 5379
rect 2752 5359 2761 5379
rect 2717 5353 2761 5359
rect 2831 5379 2875 5395
rect 2831 5359 2840 5379
rect 2860 5359 2875 5379
rect 2831 5353 2875 5359
rect 2925 5383 2974 5395
rect 2925 5363 2943 5383
rect 2963 5363 2974 5383
rect 2925 5353 2974 5363
rect 3049 5379 3093 5395
rect 3049 5359 3058 5379
rect 3078 5359 3093 5379
rect 3049 5353 3093 5359
rect 3143 5383 3192 5395
rect 3143 5363 3161 5383
rect 3181 5363 3192 5383
rect 3143 5353 3192 5363
rect 5623 5388 5672 5398
rect 5623 5368 5634 5388
rect 5654 5368 5672 5388
rect 5623 5356 5672 5368
rect 5722 5392 5766 5398
rect 5722 5372 5737 5392
rect 5757 5372 5766 5392
rect 5722 5356 5766 5372
rect 5841 5388 5890 5398
rect 5841 5368 5852 5388
rect 5872 5368 5890 5388
rect 5841 5356 5890 5368
rect 5940 5392 5984 5398
rect 5940 5372 5955 5392
rect 5975 5372 5984 5392
rect 5940 5356 5984 5372
rect 6054 5392 6098 5398
rect 6054 5372 6063 5392
rect 6083 5372 6098 5392
rect 6054 5356 6098 5372
rect 6148 5388 6197 5398
rect 6148 5368 6166 5388
rect 6186 5368 6197 5388
rect 6148 5356 6197 5368
rect 6982 5396 7031 5408
rect 6982 5376 6993 5396
rect 7013 5376 7031 5396
rect 6982 5366 7031 5376
rect 7081 5392 7125 5408
rect 7081 5372 7096 5392
rect 7116 5372 7125 5392
rect 7081 5366 7125 5372
rect 7195 5392 7239 5408
rect 7195 5372 7204 5392
rect 7224 5372 7239 5392
rect 7195 5366 7239 5372
rect 7289 5396 7338 5408
rect 7289 5376 7307 5396
rect 7327 5376 7338 5396
rect 7289 5366 7338 5376
rect 7413 5392 7457 5408
rect 7413 5372 7422 5392
rect 7442 5372 7457 5392
rect 7413 5366 7457 5372
rect 7507 5396 7556 5408
rect 7507 5376 7525 5396
rect 7545 5376 7556 5396
rect 7507 5366 7556 5376
rect 3416 5199 3465 5211
rect 3416 5179 3427 5199
rect 3447 5179 3465 5199
rect 362 5149 411 5159
rect 362 5129 373 5149
rect 393 5129 411 5149
rect 362 5117 411 5129
rect 461 5153 505 5159
rect 461 5133 476 5153
rect 496 5133 505 5153
rect 461 5117 505 5133
rect 580 5149 629 5159
rect 580 5129 591 5149
rect 611 5129 629 5149
rect 580 5117 629 5129
rect 679 5153 723 5159
rect 679 5133 694 5153
rect 714 5133 723 5153
rect 679 5117 723 5133
rect 793 5153 837 5159
rect 793 5133 802 5153
rect 822 5133 837 5153
rect 793 5117 837 5133
rect 887 5149 936 5159
rect 3416 5169 3465 5179
rect 3515 5195 3559 5211
rect 3515 5175 3530 5195
rect 3550 5175 3559 5195
rect 3515 5169 3559 5175
rect 3629 5195 3673 5211
rect 3629 5175 3638 5195
rect 3658 5175 3673 5195
rect 3629 5169 3673 5175
rect 3723 5199 3772 5211
rect 3723 5179 3741 5199
rect 3761 5179 3772 5199
rect 3723 5169 3772 5179
rect 3847 5195 3891 5211
rect 3847 5175 3856 5195
rect 3876 5175 3891 5195
rect 3847 5169 3891 5175
rect 3941 5199 3990 5211
rect 3941 5179 3959 5199
rect 3979 5179 3990 5199
rect 3941 5169 3990 5179
rect 887 5129 905 5149
rect 925 5129 936 5149
rect 887 5117 936 5129
rect 7780 5212 7829 5224
rect 7780 5192 7791 5212
rect 7811 5192 7829 5212
rect 4726 5162 4775 5172
rect 4726 5142 4737 5162
rect 4757 5142 4775 5162
rect 4726 5130 4775 5142
rect 4825 5166 4869 5172
rect 4825 5146 4840 5166
rect 4860 5146 4869 5166
rect 4825 5130 4869 5146
rect 4944 5162 4993 5172
rect 4944 5142 4955 5162
rect 4975 5142 4993 5162
rect 4944 5130 4993 5142
rect 5043 5166 5087 5172
rect 5043 5146 5058 5166
rect 5078 5146 5087 5166
rect 5043 5130 5087 5146
rect 5157 5166 5201 5172
rect 5157 5146 5166 5166
rect 5186 5146 5201 5166
rect 5157 5130 5201 5146
rect 5251 5162 5300 5172
rect 7780 5182 7829 5192
rect 7879 5208 7923 5224
rect 7879 5188 7894 5208
rect 7914 5188 7923 5208
rect 7879 5182 7923 5188
rect 7993 5208 8037 5224
rect 7993 5188 8002 5208
rect 8022 5188 8037 5208
rect 7993 5182 8037 5188
rect 8087 5212 8136 5224
rect 8087 5192 8105 5212
rect 8125 5192 8136 5212
rect 8087 5182 8136 5192
rect 8211 5208 8255 5224
rect 8211 5188 8220 5208
rect 8240 5188 8255 5208
rect 8211 5182 8255 5188
rect 8305 5212 8354 5224
rect 8305 5192 8323 5212
rect 8343 5192 8354 5212
rect 8305 5182 8354 5192
rect 5251 5142 5269 5162
rect 5289 5142 5300 5162
rect 5251 5130 5300 5142
rect 2314 4977 2363 4989
rect 1160 4965 1209 4975
rect 1160 4945 1171 4965
rect 1191 4945 1209 4965
rect 1160 4933 1209 4945
rect 1259 4969 1303 4975
rect 1259 4949 1274 4969
rect 1294 4949 1303 4969
rect 1259 4933 1303 4949
rect 1378 4965 1427 4975
rect 1378 4945 1389 4965
rect 1409 4945 1427 4965
rect 1378 4933 1427 4945
rect 1477 4969 1521 4975
rect 1477 4949 1492 4969
rect 1512 4949 1521 4969
rect 1477 4933 1521 4949
rect 1591 4969 1635 4975
rect 1591 4949 1600 4969
rect 1620 4949 1635 4969
rect 1591 4933 1635 4949
rect 1685 4965 1734 4975
rect 1685 4945 1703 4965
rect 1723 4945 1734 4965
rect 2314 4957 2325 4977
rect 2345 4957 2363 4977
rect 2314 4947 2363 4957
rect 2413 4973 2457 4989
rect 2413 4953 2428 4973
rect 2448 4953 2457 4973
rect 2413 4947 2457 4953
rect 2527 4973 2571 4989
rect 2527 4953 2536 4973
rect 2556 4953 2571 4973
rect 2527 4947 2571 4953
rect 2621 4977 2670 4989
rect 2621 4957 2639 4977
rect 2659 4957 2670 4977
rect 2621 4947 2670 4957
rect 2745 4973 2789 4989
rect 2745 4953 2754 4973
rect 2774 4953 2789 4973
rect 2745 4947 2789 4953
rect 2839 4977 2888 4989
rect 6678 4990 6727 5002
rect 2839 4957 2857 4977
rect 2877 4957 2888 4977
rect 2839 4947 2888 4957
rect 1685 4933 1734 4945
rect 5524 4978 5573 4988
rect 5524 4958 5535 4978
rect 5555 4958 5573 4978
rect 5524 4946 5573 4958
rect 5623 4982 5667 4988
rect 5623 4962 5638 4982
rect 5658 4962 5667 4982
rect 5623 4946 5667 4962
rect 5742 4978 5791 4988
rect 5742 4958 5753 4978
rect 5773 4958 5791 4978
rect 5742 4946 5791 4958
rect 5841 4982 5885 4988
rect 5841 4962 5856 4982
rect 5876 4962 5885 4982
rect 5841 4946 5885 4962
rect 5955 4982 5999 4988
rect 5955 4962 5964 4982
rect 5984 4962 5999 4982
rect 5955 4946 5999 4962
rect 6049 4978 6098 4988
rect 6049 4958 6067 4978
rect 6087 4958 6098 4978
rect 6678 4970 6689 4990
rect 6709 4970 6727 4990
rect 6678 4960 6727 4970
rect 6777 4986 6821 5002
rect 6777 4966 6792 4986
rect 6812 4966 6821 4986
rect 6777 4960 6821 4966
rect 6891 4986 6935 5002
rect 6891 4966 6900 4986
rect 6920 4966 6935 4986
rect 6891 4960 6935 4966
rect 6985 4990 7034 5002
rect 6985 4970 7003 4990
rect 7023 4970 7034 4990
rect 6985 4960 7034 4970
rect 7109 4986 7153 5002
rect 7109 4966 7118 4986
rect 7138 4966 7153 4986
rect 7109 4960 7153 4966
rect 7203 4990 7252 5002
rect 7203 4970 7221 4990
rect 7241 4970 7252 4990
rect 7203 4960 7252 4970
rect 6049 4946 6098 4958
rect 363 4737 412 4747
rect 363 4717 374 4737
rect 394 4717 412 4737
rect 363 4705 412 4717
rect 462 4741 506 4747
rect 462 4721 477 4741
rect 497 4721 506 4741
rect 462 4705 506 4721
rect 581 4737 630 4747
rect 581 4717 592 4737
rect 612 4717 630 4737
rect 581 4705 630 4717
rect 680 4741 724 4747
rect 680 4721 695 4741
rect 715 4721 724 4741
rect 680 4705 724 4721
rect 794 4741 838 4747
rect 794 4721 803 4741
rect 823 4721 838 4741
rect 794 4705 838 4721
rect 888 4737 937 4747
rect 888 4717 906 4737
rect 926 4717 937 4737
rect 888 4705 937 4717
rect 4727 4750 4776 4760
rect 4727 4730 4738 4750
rect 4758 4730 4776 4750
rect 4727 4718 4776 4730
rect 4826 4754 4870 4760
rect 4826 4734 4841 4754
rect 4861 4734 4870 4754
rect 4826 4718 4870 4734
rect 4945 4750 4994 4760
rect 4945 4730 4956 4750
rect 4976 4730 4994 4750
rect 4945 4718 4994 4730
rect 5044 4754 5088 4760
rect 5044 4734 5059 4754
rect 5079 4734 5088 4754
rect 5044 4718 5088 4734
rect 5158 4754 5202 4760
rect 5158 4734 5167 4754
rect 5187 4734 5202 4754
rect 5158 4718 5202 4734
rect 5252 4750 5301 4760
rect 5252 4730 5270 4750
rect 5290 4730 5301 4750
rect 5252 4718 5301 4730
rect 3396 4593 3445 4605
rect 3396 4573 3407 4593
rect 3427 4573 3445 4593
rect 3396 4563 3445 4573
rect 3495 4589 3539 4605
rect 3495 4569 3510 4589
rect 3530 4569 3539 4589
rect 3495 4563 3539 4569
rect 3609 4589 3653 4605
rect 3609 4569 3618 4589
rect 3638 4569 3653 4589
rect 3609 4563 3653 4569
rect 3703 4593 3752 4605
rect 3703 4573 3721 4593
rect 3741 4573 3752 4593
rect 3703 4563 3752 4573
rect 3827 4589 3871 4605
rect 3827 4569 3836 4589
rect 3856 4569 3871 4589
rect 3827 4563 3871 4569
rect 3921 4593 3970 4605
rect 3921 4573 3939 4593
rect 3959 4573 3970 4593
rect 3921 4563 3970 4573
rect 7760 4606 7809 4618
rect 7760 4586 7771 4606
rect 7791 4586 7809 4606
rect 7760 4576 7809 4586
rect 7859 4602 7903 4618
rect 7859 4582 7874 4602
rect 7894 4582 7903 4602
rect 7859 4576 7903 4582
rect 7973 4602 8017 4618
rect 7973 4582 7982 4602
rect 8002 4582 8017 4602
rect 7973 4576 8017 4582
rect 8067 4606 8116 4618
rect 8067 4586 8085 4606
rect 8105 4586 8116 4606
rect 8067 4576 8116 4586
rect 8191 4602 8235 4618
rect 8191 4582 8200 4602
rect 8220 4582 8235 4602
rect 8191 4576 8235 4582
rect 8285 4606 8334 4618
rect 8285 4586 8303 4606
rect 8323 4586 8334 4606
rect 8285 4576 8334 4586
rect 2599 4365 2648 4377
rect 1445 4353 1494 4363
rect 1445 4333 1456 4353
rect 1476 4333 1494 4353
rect 1445 4321 1494 4333
rect 1544 4357 1588 4363
rect 1544 4337 1559 4357
rect 1579 4337 1588 4357
rect 1544 4321 1588 4337
rect 1663 4353 1712 4363
rect 1663 4333 1674 4353
rect 1694 4333 1712 4353
rect 1663 4321 1712 4333
rect 1762 4357 1806 4363
rect 1762 4337 1777 4357
rect 1797 4337 1806 4357
rect 1762 4321 1806 4337
rect 1876 4357 1920 4363
rect 1876 4337 1885 4357
rect 1905 4337 1920 4357
rect 1876 4321 1920 4337
rect 1970 4353 2019 4363
rect 1970 4333 1988 4353
rect 2008 4333 2019 4353
rect 2599 4345 2610 4365
rect 2630 4345 2648 4365
rect 2599 4335 2648 4345
rect 2698 4361 2742 4377
rect 2698 4341 2713 4361
rect 2733 4341 2742 4361
rect 2698 4335 2742 4341
rect 2812 4361 2856 4377
rect 2812 4341 2821 4361
rect 2841 4341 2856 4361
rect 2812 4335 2856 4341
rect 2906 4365 2955 4377
rect 2906 4345 2924 4365
rect 2944 4345 2955 4365
rect 2906 4335 2955 4345
rect 3030 4361 3074 4377
rect 3030 4341 3039 4361
rect 3059 4341 3074 4361
rect 3030 4335 3074 4341
rect 3124 4365 3173 4377
rect 3124 4345 3142 4365
rect 3162 4345 3173 4365
rect 3124 4335 3173 4345
rect 6963 4378 7012 4390
rect 5809 4366 5858 4376
rect 5809 4346 5820 4366
rect 5840 4346 5858 4366
rect 1970 4321 2019 4333
rect 5809 4334 5858 4346
rect 5908 4370 5952 4376
rect 5908 4350 5923 4370
rect 5943 4350 5952 4370
rect 5908 4334 5952 4350
rect 6027 4366 6076 4376
rect 6027 4346 6038 4366
rect 6058 4346 6076 4366
rect 6027 4334 6076 4346
rect 6126 4370 6170 4376
rect 6126 4350 6141 4370
rect 6161 4350 6170 4370
rect 6126 4334 6170 4350
rect 6240 4370 6284 4376
rect 6240 4350 6249 4370
rect 6269 4350 6284 4370
rect 6240 4334 6284 4350
rect 6334 4366 6383 4376
rect 6334 4346 6352 4366
rect 6372 4346 6383 4366
rect 6963 4358 6974 4378
rect 6994 4358 7012 4378
rect 6963 4348 7012 4358
rect 7062 4374 7106 4390
rect 7062 4354 7077 4374
rect 7097 4354 7106 4374
rect 7062 4348 7106 4354
rect 7176 4374 7220 4390
rect 7176 4354 7185 4374
rect 7205 4354 7220 4374
rect 7176 4348 7220 4354
rect 7270 4378 7319 4390
rect 7270 4358 7288 4378
rect 7308 4358 7319 4378
rect 7270 4348 7319 4358
rect 7394 4374 7438 4390
rect 7394 4354 7403 4374
rect 7423 4354 7438 4374
rect 7394 4348 7438 4354
rect 7488 4378 7537 4390
rect 7488 4358 7506 4378
rect 7526 4358 7537 4378
rect 7488 4348 7537 4358
rect 6334 4334 6383 4346
rect 3397 4181 3446 4193
rect 3397 4161 3408 4181
rect 3428 4161 3446 4181
rect 343 4131 392 4141
rect 343 4111 354 4131
rect 374 4111 392 4131
rect 343 4099 392 4111
rect 442 4135 486 4141
rect 442 4115 457 4135
rect 477 4115 486 4135
rect 442 4099 486 4115
rect 561 4131 610 4141
rect 561 4111 572 4131
rect 592 4111 610 4131
rect 561 4099 610 4111
rect 660 4135 704 4141
rect 660 4115 675 4135
rect 695 4115 704 4135
rect 660 4099 704 4115
rect 774 4135 818 4141
rect 774 4115 783 4135
rect 803 4115 818 4135
rect 774 4099 818 4115
rect 868 4131 917 4141
rect 3397 4151 3446 4161
rect 3496 4177 3540 4193
rect 3496 4157 3511 4177
rect 3531 4157 3540 4177
rect 3496 4151 3540 4157
rect 3610 4177 3654 4193
rect 3610 4157 3619 4177
rect 3639 4157 3654 4177
rect 3610 4151 3654 4157
rect 3704 4181 3753 4193
rect 3704 4161 3722 4181
rect 3742 4161 3753 4181
rect 3704 4151 3753 4161
rect 3828 4177 3872 4193
rect 3828 4157 3837 4177
rect 3857 4157 3872 4177
rect 3828 4151 3872 4157
rect 3922 4181 3971 4193
rect 3922 4161 3940 4181
rect 3960 4161 3971 4181
rect 3922 4151 3971 4161
rect 868 4111 886 4131
rect 906 4111 917 4131
rect 868 4099 917 4111
rect 7761 4194 7810 4206
rect 7761 4174 7772 4194
rect 7792 4174 7810 4194
rect 4707 4144 4756 4154
rect 4707 4124 4718 4144
rect 4738 4124 4756 4144
rect 4707 4112 4756 4124
rect 4806 4148 4850 4154
rect 4806 4128 4821 4148
rect 4841 4128 4850 4148
rect 4806 4112 4850 4128
rect 4925 4144 4974 4154
rect 4925 4124 4936 4144
rect 4956 4124 4974 4144
rect 4925 4112 4974 4124
rect 5024 4148 5068 4154
rect 5024 4128 5039 4148
rect 5059 4128 5068 4148
rect 5024 4112 5068 4128
rect 5138 4148 5182 4154
rect 5138 4128 5147 4148
rect 5167 4128 5182 4148
rect 5138 4112 5182 4128
rect 5232 4144 5281 4154
rect 7761 4164 7810 4174
rect 7860 4190 7904 4206
rect 7860 4170 7875 4190
rect 7895 4170 7904 4190
rect 7860 4164 7904 4170
rect 7974 4190 8018 4206
rect 7974 4170 7983 4190
rect 8003 4170 8018 4190
rect 7974 4164 8018 4170
rect 8068 4194 8117 4206
rect 8068 4174 8086 4194
rect 8106 4174 8117 4194
rect 8068 4164 8117 4174
rect 8192 4190 8236 4206
rect 8192 4170 8201 4190
rect 8221 4170 8236 4190
rect 8192 4164 8236 4170
rect 8286 4194 8335 4206
rect 8286 4174 8304 4194
rect 8324 4174 8335 4194
rect 8286 4164 8335 4174
rect 5232 4124 5250 4144
rect 5270 4124 5281 4144
rect 5232 4112 5281 4124
rect 1141 3947 1190 3957
rect 1141 3927 1152 3947
rect 1172 3927 1190 3947
rect 1141 3915 1190 3927
rect 1240 3951 1284 3957
rect 1240 3931 1255 3951
rect 1275 3931 1284 3951
rect 1240 3915 1284 3931
rect 1359 3947 1408 3957
rect 1359 3927 1370 3947
rect 1390 3927 1408 3947
rect 1359 3915 1408 3927
rect 1458 3951 1502 3957
rect 1458 3931 1473 3951
rect 1493 3931 1502 3951
rect 1458 3915 1502 3931
rect 1572 3951 1616 3957
rect 1572 3931 1581 3951
rect 1601 3931 1616 3951
rect 1572 3915 1616 3931
rect 1666 3947 1715 3957
rect 1666 3927 1684 3947
rect 1704 3927 1715 3947
rect 1666 3915 1715 3927
rect 2500 3955 2549 3967
rect 2500 3935 2511 3955
rect 2531 3935 2549 3955
rect 2500 3925 2549 3935
rect 2599 3951 2643 3967
rect 2599 3931 2614 3951
rect 2634 3931 2643 3951
rect 2599 3925 2643 3931
rect 2713 3951 2757 3967
rect 2713 3931 2722 3951
rect 2742 3931 2757 3951
rect 2713 3925 2757 3931
rect 2807 3955 2856 3967
rect 2807 3935 2825 3955
rect 2845 3935 2856 3955
rect 2807 3925 2856 3935
rect 2931 3951 2975 3967
rect 2931 3931 2940 3951
rect 2960 3931 2975 3951
rect 2931 3925 2975 3931
rect 3025 3955 3074 3967
rect 3025 3935 3043 3955
rect 3063 3935 3074 3955
rect 3025 3925 3074 3935
rect 5505 3960 5554 3970
rect 5505 3940 5516 3960
rect 5536 3940 5554 3960
rect 5505 3928 5554 3940
rect 5604 3964 5648 3970
rect 5604 3944 5619 3964
rect 5639 3944 5648 3964
rect 5604 3928 5648 3944
rect 5723 3960 5772 3970
rect 5723 3940 5734 3960
rect 5754 3940 5772 3960
rect 5723 3928 5772 3940
rect 5822 3964 5866 3970
rect 5822 3944 5837 3964
rect 5857 3944 5866 3964
rect 5822 3928 5866 3944
rect 5936 3964 5980 3970
rect 5936 3944 5945 3964
rect 5965 3944 5980 3964
rect 5936 3928 5980 3944
rect 6030 3960 6079 3970
rect 6030 3940 6048 3960
rect 6068 3940 6079 3960
rect 6030 3928 6079 3940
rect 6864 3968 6913 3980
rect 6864 3948 6875 3968
rect 6895 3948 6913 3968
rect 6864 3938 6913 3948
rect 6963 3964 7007 3980
rect 6963 3944 6978 3964
rect 6998 3944 7007 3964
rect 6963 3938 7007 3944
rect 7077 3964 7121 3980
rect 7077 3944 7086 3964
rect 7106 3944 7121 3964
rect 7077 3938 7121 3944
rect 7171 3968 7220 3980
rect 7171 3948 7189 3968
rect 7209 3948 7220 3968
rect 7171 3938 7220 3948
rect 7295 3964 7339 3980
rect 7295 3944 7304 3964
rect 7324 3944 7339 3964
rect 7295 3938 7339 3944
rect 7389 3968 7438 3980
rect 7389 3948 7407 3968
rect 7427 3948 7438 3968
rect 7389 3938 7438 3948
rect 344 3719 393 3729
rect 344 3699 355 3719
rect 375 3699 393 3719
rect 344 3687 393 3699
rect 443 3723 487 3729
rect 443 3703 458 3723
rect 478 3703 487 3723
rect 443 3687 487 3703
rect 562 3719 611 3729
rect 562 3699 573 3719
rect 593 3699 611 3719
rect 562 3687 611 3699
rect 661 3723 705 3729
rect 661 3703 676 3723
rect 696 3703 705 3723
rect 661 3687 705 3703
rect 775 3723 819 3729
rect 775 3703 784 3723
rect 804 3703 819 3723
rect 775 3687 819 3703
rect 869 3719 918 3729
rect 869 3699 887 3719
rect 907 3699 918 3719
rect 869 3687 918 3699
rect 4708 3732 4757 3742
rect 4708 3712 4719 3732
rect 4739 3712 4757 3732
rect 4708 3700 4757 3712
rect 4807 3736 4851 3742
rect 4807 3716 4822 3736
rect 4842 3716 4851 3736
rect 4807 3700 4851 3716
rect 4926 3732 4975 3742
rect 4926 3712 4937 3732
rect 4957 3712 4975 3732
rect 4926 3700 4975 3712
rect 5025 3736 5069 3742
rect 5025 3716 5040 3736
rect 5060 3716 5069 3736
rect 5025 3700 5069 3716
rect 5139 3736 5183 3742
rect 5139 3716 5148 3736
rect 5168 3716 5183 3736
rect 5139 3700 5183 3716
rect 5233 3732 5282 3742
rect 5233 3712 5251 3732
rect 5271 3712 5282 3732
rect 5233 3700 5282 3712
rect 3379 3575 3428 3587
rect 3379 3555 3390 3575
rect 3410 3555 3428 3575
rect 3379 3545 3428 3555
rect 3478 3571 3522 3587
rect 3478 3551 3493 3571
rect 3513 3551 3522 3571
rect 3478 3545 3522 3551
rect 3592 3571 3636 3587
rect 3592 3551 3601 3571
rect 3621 3551 3636 3571
rect 3592 3545 3636 3551
rect 3686 3575 3735 3587
rect 3686 3555 3704 3575
rect 3724 3555 3735 3575
rect 3686 3545 3735 3555
rect 3810 3571 3854 3587
rect 3810 3551 3819 3571
rect 3839 3551 3854 3571
rect 3810 3545 3854 3551
rect 3904 3575 3953 3587
rect 3904 3555 3922 3575
rect 3942 3555 3953 3575
rect 3904 3545 3953 3555
rect 7743 3588 7792 3600
rect 7743 3568 7754 3588
rect 7774 3568 7792 3588
rect 7743 3558 7792 3568
rect 7842 3584 7886 3600
rect 7842 3564 7857 3584
rect 7877 3564 7886 3584
rect 7842 3558 7886 3564
rect 7956 3584 8000 3600
rect 7956 3564 7965 3584
rect 7985 3564 8000 3584
rect 7956 3558 8000 3564
rect 8050 3588 8099 3600
rect 8050 3568 8068 3588
rect 8088 3568 8099 3588
rect 8050 3558 8099 3568
rect 8174 3584 8218 3600
rect 8174 3564 8183 3584
rect 8203 3564 8218 3584
rect 8174 3558 8218 3564
rect 8268 3588 8317 3600
rect 8268 3568 8286 3588
rect 8306 3568 8317 3588
rect 8268 3558 8317 3568
rect 1223 3339 1272 3349
rect 1223 3319 1234 3339
rect 1254 3319 1272 3339
rect 1223 3307 1272 3319
rect 1322 3343 1366 3349
rect 1322 3323 1337 3343
rect 1357 3323 1366 3343
rect 1322 3307 1366 3323
rect 1441 3339 1490 3349
rect 1441 3319 1452 3339
rect 1472 3319 1490 3339
rect 1441 3307 1490 3319
rect 1540 3343 1584 3349
rect 1540 3323 1555 3343
rect 1575 3323 1584 3343
rect 1540 3307 1584 3323
rect 1654 3343 1698 3349
rect 1654 3323 1663 3343
rect 1683 3323 1698 3343
rect 1654 3307 1698 3323
rect 1748 3339 1797 3349
rect 1748 3319 1766 3339
rect 1786 3319 1797 3339
rect 1748 3307 1797 3319
rect 2582 3347 2631 3359
rect 2582 3327 2593 3347
rect 2613 3327 2631 3347
rect 2582 3317 2631 3327
rect 2681 3343 2725 3359
rect 2681 3323 2696 3343
rect 2716 3323 2725 3343
rect 2681 3317 2725 3323
rect 2795 3343 2839 3359
rect 2795 3323 2804 3343
rect 2824 3323 2839 3343
rect 2795 3317 2839 3323
rect 2889 3347 2938 3359
rect 2889 3327 2907 3347
rect 2927 3327 2938 3347
rect 2889 3317 2938 3327
rect 3013 3343 3057 3359
rect 3013 3323 3022 3343
rect 3042 3323 3057 3343
rect 3013 3317 3057 3323
rect 3107 3347 3156 3359
rect 3107 3327 3125 3347
rect 3145 3327 3156 3347
rect 3107 3317 3156 3327
rect 5587 3352 5636 3362
rect 5587 3332 5598 3352
rect 5618 3332 5636 3352
rect 5587 3320 5636 3332
rect 5686 3356 5730 3362
rect 5686 3336 5701 3356
rect 5721 3336 5730 3356
rect 5686 3320 5730 3336
rect 5805 3352 5854 3362
rect 5805 3332 5816 3352
rect 5836 3332 5854 3352
rect 5805 3320 5854 3332
rect 5904 3356 5948 3362
rect 5904 3336 5919 3356
rect 5939 3336 5948 3356
rect 5904 3320 5948 3336
rect 6018 3356 6062 3362
rect 6018 3336 6027 3356
rect 6047 3336 6062 3356
rect 6018 3320 6062 3336
rect 6112 3352 6161 3362
rect 6112 3332 6130 3352
rect 6150 3332 6161 3352
rect 6112 3320 6161 3332
rect 6946 3360 6995 3372
rect 6946 3340 6957 3360
rect 6977 3340 6995 3360
rect 6946 3330 6995 3340
rect 7045 3356 7089 3372
rect 7045 3336 7060 3356
rect 7080 3336 7089 3356
rect 7045 3330 7089 3336
rect 7159 3356 7203 3372
rect 7159 3336 7168 3356
rect 7188 3336 7203 3356
rect 7159 3330 7203 3336
rect 7253 3360 7302 3372
rect 7253 3340 7271 3360
rect 7291 3340 7302 3360
rect 7253 3330 7302 3340
rect 7377 3356 7421 3372
rect 7377 3336 7386 3356
rect 7406 3336 7421 3356
rect 7377 3330 7421 3336
rect 7471 3360 7520 3372
rect 7471 3340 7489 3360
rect 7509 3340 7520 3360
rect 7471 3330 7520 3340
rect 3380 3163 3429 3175
rect 3380 3143 3391 3163
rect 3411 3143 3429 3163
rect 326 3113 375 3123
rect 326 3093 337 3113
rect 357 3093 375 3113
rect 326 3081 375 3093
rect 425 3117 469 3123
rect 425 3097 440 3117
rect 460 3097 469 3117
rect 425 3081 469 3097
rect 544 3113 593 3123
rect 544 3093 555 3113
rect 575 3093 593 3113
rect 544 3081 593 3093
rect 643 3117 687 3123
rect 643 3097 658 3117
rect 678 3097 687 3117
rect 643 3081 687 3097
rect 757 3117 801 3123
rect 757 3097 766 3117
rect 786 3097 801 3117
rect 757 3081 801 3097
rect 851 3113 900 3123
rect 3380 3133 3429 3143
rect 3479 3159 3523 3175
rect 3479 3139 3494 3159
rect 3514 3139 3523 3159
rect 3479 3133 3523 3139
rect 3593 3159 3637 3175
rect 3593 3139 3602 3159
rect 3622 3139 3637 3159
rect 3593 3133 3637 3139
rect 3687 3163 3736 3175
rect 3687 3143 3705 3163
rect 3725 3143 3736 3163
rect 3687 3133 3736 3143
rect 3811 3159 3855 3175
rect 3811 3139 3820 3159
rect 3840 3139 3855 3159
rect 3811 3133 3855 3139
rect 3905 3163 3954 3175
rect 3905 3143 3923 3163
rect 3943 3143 3954 3163
rect 3905 3133 3954 3143
rect 851 3093 869 3113
rect 889 3093 900 3113
rect 851 3081 900 3093
rect 7744 3176 7793 3188
rect 7744 3156 7755 3176
rect 7775 3156 7793 3176
rect 4690 3126 4739 3136
rect 4690 3106 4701 3126
rect 4721 3106 4739 3126
rect 4690 3094 4739 3106
rect 4789 3130 4833 3136
rect 4789 3110 4804 3130
rect 4824 3110 4833 3130
rect 4789 3094 4833 3110
rect 4908 3126 4957 3136
rect 4908 3106 4919 3126
rect 4939 3106 4957 3126
rect 4908 3094 4957 3106
rect 5007 3130 5051 3136
rect 5007 3110 5022 3130
rect 5042 3110 5051 3130
rect 5007 3094 5051 3110
rect 5121 3130 5165 3136
rect 5121 3110 5130 3130
rect 5150 3110 5165 3130
rect 5121 3094 5165 3110
rect 5215 3126 5264 3136
rect 7744 3146 7793 3156
rect 7843 3172 7887 3188
rect 7843 3152 7858 3172
rect 7878 3152 7887 3172
rect 7843 3146 7887 3152
rect 7957 3172 8001 3188
rect 7957 3152 7966 3172
rect 7986 3152 8001 3172
rect 7957 3146 8001 3152
rect 8051 3176 8100 3188
rect 8051 3156 8069 3176
rect 8089 3156 8100 3176
rect 8051 3146 8100 3156
rect 8175 3172 8219 3188
rect 8175 3152 8184 3172
rect 8204 3152 8219 3172
rect 8175 3146 8219 3152
rect 8269 3176 8318 3188
rect 8269 3156 8287 3176
rect 8307 3156 8318 3176
rect 8269 3146 8318 3156
rect 5215 3106 5233 3126
rect 5253 3106 5264 3126
rect 5215 3094 5264 3106
rect 2417 2939 2466 2951
rect 1124 2929 1173 2939
rect 1124 2909 1135 2929
rect 1155 2909 1173 2929
rect 1124 2897 1173 2909
rect 1223 2933 1267 2939
rect 1223 2913 1238 2933
rect 1258 2913 1267 2933
rect 1223 2897 1267 2913
rect 1342 2929 1391 2939
rect 1342 2909 1353 2929
rect 1373 2909 1391 2929
rect 1342 2897 1391 2909
rect 1441 2933 1485 2939
rect 1441 2913 1456 2933
rect 1476 2913 1485 2933
rect 1441 2897 1485 2913
rect 1555 2933 1599 2939
rect 1555 2913 1564 2933
rect 1584 2913 1599 2933
rect 1555 2897 1599 2913
rect 1649 2929 1698 2939
rect 1649 2909 1667 2929
rect 1687 2909 1698 2929
rect 2417 2919 2428 2939
rect 2448 2919 2466 2939
rect 2417 2909 2466 2919
rect 2516 2935 2560 2951
rect 2516 2915 2531 2935
rect 2551 2915 2560 2935
rect 2516 2909 2560 2915
rect 2630 2935 2674 2951
rect 2630 2915 2639 2935
rect 2659 2915 2674 2935
rect 2630 2909 2674 2915
rect 2724 2939 2773 2951
rect 2724 2919 2742 2939
rect 2762 2919 2773 2939
rect 2724 2909 2773 2919
rect 2848 2935 2892 2951
rect 2848 2915 2857 2935
rect 2877 2915 2892 2935
rect 2848 2909 2892 2915
rect 2942 2939 2991 2951
rect 6781 2952 6830 2964
rect 2942 2919 2960 2939
rect 2980 2919 2991 2939
rect 2942 2909 2991 2919
rect 1649 2897 1698 2909
rect 5488 2942 5537 2952
rect 5488 2922 5499 2942
rect 5519 2922 5537 2942
rect 5488 2910 5537 2922
rect 5587 2946 5631 2952
rect 5587 2926 5602 2946
rect 5622 2926 5631 2946
rect 5587 2910 5631 2926
rect 5706 2942 5755 2952
rect 5706 2922 5717 2942
rect 5737 2922 5755 2942
rect 5706 2910 5755 2922
rect 5805 2946 5849 2952
rect 5805 2926 5820 2946
rect 5840 2926 5849 2946
rect 5805 2910 5849 2926
rect 5919 2946 5963 2952
rect 5919 2926 5928 2946
rect 5948 2926 5963 2946
rect 5919 2910 5963 2926
rect 6013 2942 6062 2952
rect 6013 2922 6031 2942
rect 6051 2922 6062 2942
rect 6781 2932 6792 2952
rect 6812 2932 6830 2952
rect 6781 2922 6830 2932
rect 6880 2948 6924 2964
rect 6880 2928 6895 2948
rect 6915 2928 6924 2948
rect 6880 2922 6924 2928
rect 6994 2948 7038 2964
rect 6994 2928 7003 2948
rect 7023 2928 7038 2948
rect 6994 2922 7038 2928
rect 7088 2952 7137 2964
rect 7088 2932 7106 2952
rect 7126 2932 7137 2952
rect 7088 2922 7137 2932
rect 7212 2948 7256 2964
rect 7212 2928 7221 2948
rect 7241 2928 7256 2948
rect 7212 2922 7256 2928
rect 7306 2952 7355 2964
rect 7306 2932 7324 2952
rect 7344 2932 7355 2952
rect 7306 2922 7355 2932
rect 6013 2910 6062 2922
rect 327 2701 376 2711
rect 327 2681 338 2701
rect 358 2681 376 2701
rect 327 2669 376 2681
rect 426 2705 470 2711
rect 426 2685 441 2705
rect 461 2685 470 2705
rect 426 2669 470 2685
rect 545 2701 594 2711
rect 545 2681 556 2701
rect 576 2681 594 2701
rect 545 2669 594 2681
rect 644 2705 688 2711
rect 644 2685 659 2705
rect 679 2685 688 2705
rect 644 2669 688 2685
rect 758 2705 802 2711
rect 758 2685 767 2705
rect 787 2685 802 2705
rect 758 2669 802 2685
rect 852 2701 901 2711
rect 852 2681 870 2701
rect 890 2681 901 2701
rect 852 2669 901 2681
rect 4691 2714 4740 2724
rect 4691 2694 4702 2714
rect 4722 2694 4740 2714
rect 4691 2682 4740 2694
rect 4790 2718 4834 2724
rect 4790 2698 4805 2718
rect 4825 2698 4834 2718
rect 4790 2682 4834 2698
rect 4909 2714 4958 2724
rect 4909 2694 4920 2714
rect 4940 2694 4958 2714
rect 4909 2682 4958 2694
rect 5008 2718 5052 2724
rect 5008 2698 5023 2718
rect 5043 2698 5052 2718
rect 5008 2682 5052 2698
rect 5122 2718 5166 2724
rect 5122 2698 5131 2718
rect 5151 2698 5166 2718
rect 5122 2682 5166 2698
rect 5216 2714 5265 2724
rect 5216 2694 5234 2714
rect 5254 2694 5265 2714
rect 5216 2682 5265 2694
rect 3359 2557 3408 2569
rect 3359 2537 3370 2557
rect 3390 2537 3408 2557
rect 3359 2527 3408 2537
rect 3458 2553 3502 2569
rect 3458 2533 3473 2553
rect 3493 2533 3502 2553
rect 3458 2527 3502 2533
rect 3572 2553 3616 2569
rect 3572 2533 3581 2553
rect 3601 2533 3616 2553
rect 3572 2527 3616 2533
rect 3666 2557 3715 2569
rect 3666 2537 3684 2557
rect 3704 2537 3715 2557
rect 3666 2527 3715 2537
rect 3790 2553 3834 2569
rect 3790 2533 3799 2553
rect 3819 2533 3834 2553
rect 3790 2527 3834 2533
rect 3884 2557 3933 2569
rect 3884 2537 3902 2557
rect 3922 2537 3933 2557
rect 3884 2527 3933 2537
rect 7723 2570 7772 2582
rect 7723 2550 7734 2570
rect 7754 2550 7772 2570
rect 7723 2540 7772 2550
rect 7822 2566 7866 2582
rect 7822 2546 7837 2566
rect 7857 2546 7866 2566
rect 7822 2540 7866 2546
rect 7936 2566 7980 2582
rect 7936 2546 7945 2566
rect 7965 2546 7980 2566
rect 7936 2540 7980 2546
rect 8030 2570 8079 2582
rect 8030 2550 8048 2570
rect 8068 2550 8079 2570
rect 8030 2540 8079 2550
rect 8154 2566 8198 2582
rect 8154 2546 8163 2566
rect 8183 2546 8198 2566
rect 8154 2540 8198 2546
rect 8248 2570 8297 2582
rect 8248 2550 8266 2570
rect 8286 2550 8297 2570
rect 8248 2540 8297 2550
rect 2562 2329 2611 2341
rect 1269 2319 1318 2329
rect 1269 2299 1280 2319
rect 1300 2299 1318 2319
rect 1269 2287 1318 2299
rect 1368 2323 1412 2329
rect 1368 2303 1383 2323
rect 1403 2303 1412 2323
rect 1368 2287 1412 2303
rect 1487 2319 1536 2329
rect 1487 2299 1498 2319
rect 1518 2299 1536 2319
rect 1487 2287 1536 2299
rect 1586 2323 1630 2329
rect 1586 2303 1601 2323
rect 1621 2303 1630 2323
rect 1586 2287 1630 2303
rect 1700 2323 1744 2329
rect 1700 2303 1709 2323
rect 1729 2303 1744 2323
rect 1700 2287 1744 2303
rect 1794 2319 1843 2329
rect 1794 2299 1812 2319
rect 1832 2299 1843 2319
rect 2562 2309 2573 2329
rect 2593 2309 2611 2329
rect 2562 2299 2611 2309
rect 2661 2325 2705 2341
rect 2661 2305 2676 2325
rect 2696 2305 2705 2325
rect 2661 2299 2705 2305
rect 2775 2325 2819 2341
rect 2775 2305 2784 2325
rect 2804 2305 2819 2325
rect 2775 2299 2819 2305
rect 2869 2329 2918 2341
rect 2869 2309 2887 2329
rect 2907 2309 2918 2329
rect 2869 2299 2918 2309
rect 2993 2325 3037 2341
rect 2993 2305 3002 2325
rect 3022 2305 3037 2325
rect 2993 2299 3037 2305
rect 3087 2329 3136 2341
rect 3087 2309 3105 2329
rect 3125 2309 3136 2329
rect 3087 2299 3136 2309
rect 6926 2342 6975 2354
rect 5633 2332 5682 2342
rect 5633 2312 5644 2332
rect 5664 2312 5682 2332
rect 1794 2287 1843 2299
rect 5633 2300 5682 2312
rect 5732 2336 5776 2342
rect 5732 2316 5747 2336
rect 5767 2316 5776 2336
rect 5732 2300 5776 2316
rect 5851 2332 5900 2342
rect 5851 2312 5862 2332
rect 5882 2312 5900 2332
rect 5851 2300 5900 2312
rect 5950 2336 5994 2342
rect 5950 2316 5965 2336
rect 5985 2316 5994 2336
rect 5950 2300 5994 2316
rect 6064 2336 6108 2342
rect 6064 2316 6073 2336
rect 6093 2316 6108 2336
rect 6064 2300 6108 2316
rect 6158 2332 6207 2342
rect 6158 2312 6176 2332
rect 6196 2312 6207 2332
rect 6926 2322 6937 2342
rect 6957 2322 6975 2342
rect 6926 2312 6975 2322
rect 7025 2338 7069 2354
rect 7025 2318 7040 2338
rect 7060 2318 7069 2338
rect 7025 2312 7069 2318
rect 7139 2338 7183 2354
rect 7139 2318 7148 2338
rect 7168 2318 7183 2338
rect 7139 2312 7183 2318
rect 7233 2342 7282 2354
rect 7233 2322 7251 2342
rect 7271 2322 7282 2342
rect 7233 2312 7282 2322
rect 7357 2338 7401 2354
rect 7357 2318 7366 2338
rect 7386 2318 7401 2338
rect 7357 2312 7401 2318
rect 7451 2342 7500 2354
rect 7451 2322 7469 2342
rect 7489 2322 7500 2342
rect 7451 2312 7500 2322
rect 6158 2300 6207 2312
rect 3360 2145 3409 2157
rect 3360 2125 3371 2145
rect 3391 2125 3409 2145
rect 306 2095 355 2105
rect 306 2075 317 2095
rect 337 2075 355 2095
rect 306 2063 355 2075
rect 405 2099 449 2105
rect 405 2079 420 2099
rect 440 2079 449 2099
rect 405 2063 449 2079
rect 524 2095 573 2105
rect 524 2075 535 2095
rect 555 2075 573 2095
rect 524 2063 573 2075
rect 623 2099 667 2105
rect 623 2079 638 2099
rect 658 2079 667 2099
rect 623 2063 667 2079
rect 737 2099 781 2105
rect 737 2079 746 2099
rect 766 2079 781 2099
rect 737 2063 781 2079
rect 831 2095 880 2105
rect 3360 2115 3409 2125
rect 3459 2141 3503 2157
rect 3459 2121 3474 2141
rect 3494 2121 3503 2141
rect 3459 2115 3503 2121
rect 3573 2141 3617 2157
rect 3573 2121 3582 2141
rect 3602 2121 3617 2141
rect 3573 2115 3617 2121
rect 3667 2145 3716 2157
rect 3667 2125 3685 2145
rect 3705 2125 3716 2145
rect 3667 2115 3716 2125
rect 3791 2141 3835 2157
rect 3791 2121 3800 2141
rect 3820 2121 3835 2141
rect 3791 2115 3835 2121
rect 3885 2145 3934 2157
rect 3885 2125 3903 2145
rect 3923 2125 3934 2145
rect 3885 2115 3934 2125
rect 831 2075 849 2095
rect 869 2075 880 2095
rect 831 2063 880 2075
rect 7724 2158 7773 2170
rect 7724 2138 7735 2158
rect 7755 2138 7773 2158
rect 4670 2108 4719 2118
rect 4670 2088 4681 2108
rect 4701 2088 4719 2108
rect 4670 2076 4719 2088
rect 4769 2112 4813 2118
rect 4769 2092 4784 2112
rect 4804 2092 4813 2112
rect 4769 2076 4813 2092
rect 4888 2108 4937 2118
rect 4888 2088 4899 2108
rect 4919 2088 4937 2108
rect 4888 2076 4937 2088
rect 4987 2112 5031 2118
rect 4987 2092 5002 2112
rect 5022 2092 5031 2112
rect 4987 2076 5031 2092
rect 5101 2112 5145 2118
rect 5101 2092 5110 2112
rect 5130 2092 5145 2112
rect 5101 2076 5145 2092
rect 5195 2108 5244 2118
rect 7724 2128 7773 2138
rect 7823 2154 7867 2170
rect 7823 2134 7838 2154
rect 7858 2134 7867 2154
rect 7823 2128 7867 2134
rect 7937 2154 7981 2170
rect 7937 2134 7946 2154
rect 7966 2134 7981 2154
rect 7937 2128 7981 2134
rect 8031 2158 8080 2170
rect 8031 2138 8049 2158
rect 8069 2138 8080 2158
rect 8031 2128 8080 2138
rect 8155 2154 8199 2170
rect 8155 2134 8164 2154
rect 8184 2134 8199 2154
rect 8155 2128 8199 2134
rect 8249 2158 8298 2170
rect 8249 2138 8267 2158
rect 8287 2138 8298 2158
rect 8249 2128 8298 2138
rect 5195 2088 5213 2108
rect 5233 2088 5244 2108
rect 5195 2076 5244 2088
rect 1104 1911 1153 1921
rect 1104 1891 1115 1911
rect 1135 1891 1153 1911
rect 1104 1879 1153 1891
rect 1203 1915 1247 1921
rect 1203 1895 1218 1915
rect 1238 1895 1247 1915
rect 1203 1879 1247 1895
rect 1322 1911 1371 1921
rect 1322 1891 1333 1911
rect 1353 1891 1371 1911
rect 1322 1879 1371 1891
rect 1421 1915 1465 1921
rect 1421 1895 1436 1915
rect 1456 1895 1465 1915
rect 1421 1879 1465 1895
rect 1535 1915 1579 1921
rect 1535 1895 1544 1915
rect 1564 1895 1579 1915
rect 1535 1879 1579 1895
rect 1629 1911 1678 1921
rect 1629 1891 1647 1911
rect 1667 1891 1678 1911
rect 1629 1879 1678 1891
rect 2463 1919 2512 1931
rect 2463 1899 2474 1919
rect 2494 1899 2512 1919
rect 2463 1889 2512 1899
rect 2562 1915 2606 1931
rect 2562 1895 2577 1915
rect 2597 1895 2606 1915
rect 2562 1889 2606 1895
rect 2676 1915 2720 1931
rect 2676 1895 2685 1915
rect 2705 1895 2720 1915
rect 2676 1889 2720 1895
rect 2770 1919 2819 1931
rect 2770 1899 2788 1919
rect 2808 1899 2819 1919
rect 2770 1889 2819 1899
rect 2894 1915 2938 1931
rect 2894 1895 2903 1915
rect 2923 1895 2938 1915
rect 2894 1889 2938 1895
rect 2988 1919 3037 1931
rect 2988 1899 3006 1919
rect 3026 1899 3037 1919
rect 2988 1889 3037 1899
rect 5468 1924 5517 1934
rect 5468 1904 5479 1924
rect 5499 1904 5517 1924
rect 5468 1892 5517 1904
rect 5567 1928 5611 1934
rect 5567 1908 5582 1928
rect 5602 1908 5611 1928
rect 5567 1892 5611 1908
rect 5686 1924 5735 1934
rect 5686 1904 5697 1924
rect 5717 1904 5735 1924
rect 5686 1892 5735 1904
rect 5785 1928 5829 1934
rect 5785 1908 5800 1928
rect 5820 1908 5829 1928
rect 5785 1892 5829 1908
rect 5899 1928 5943 1934
rect 5899 1908 5908 1928
rect 5928 1908 5943 1928
rect 5899 1892 5943 1908
rect 5993 1924 6042 1934
rect 5993 1904 6011 1924
rect 6031 1904 6042 1924
rect 5993 1892 6042 1904
rect 6827 1932 6876 1944
rect 6827 1912 6838 1932
rect 6858 1912 6876 1932
rect 6827 1902 6876 1912
rect 6926 1928 6970 1944
rect 6926 1908 6941 1928
rect 6961 1908 6970 1928
rect 6926 1902 6970 1908
rect 7040 1928 7084 1944
rect 7040 1908 7049 1928
rect 7069 1908 7084 1928
rect 7040 1902 7084 1908
rect 7134 1932 7183 1944
rect 7134 1912 7152 1932
rect 7172 1912 7183 1932
rect 7134 1902 7183 1912
rect 7258 1928 7302 1944
rect 7258 1908 7267 1928
rect 7287 1908 7302 1928
rect 7258 1902 7302 1908
rect 7352 1932 7401 1944
rect 7352 1912 7370 1932
rect 7390 1912 7401 1932
rect 7352 1902 7401 1912
rect 307 1683 356 1693
rect 307 1663 318 1683
rect 338 1663 356 1683
rect 307 1651 356 1663
rect 406 1687 450 1693
rect 406 1667 421 1687
rect 441 1667 450 1687
rect 406 1651 450 1667
rect 525 1683 574 1693
rect 525 1663 536 1683
rect 556 1663 574 1683
rect 525 1651 574 1663
rect 624 1687 668 1693
rect 624 1667 639 1687
rect 659 1667 668 1687
rect 624 1651 668 1667
rect 738 1687 782 1693
rect 738 1667 747 1687
rect 767 1667 782 1687
rect 738 1651 782 1667
rect 832 1683 881 1693
rect 832 1663 850 1683
rect 870 1663 881 1683
rect 832 1651 881 1663
rect 4671 1696 4720 1706
rect 4671 1676 4682 1696
rect 4702 1676 4720 1696
rect 4671 1664 4720 1676
rect 4770 1700 4814 1706
rect 4770 1680 4785 1700
rect 4805 1680 4814 1700
rect 4770 1664 4814 1680
rect 4889 1696 4938 1706
rect 4889 1676 4900 1696
rect 4920 1676 4938 1696
rect 4889 1664 4938 1676
rect 4988 1700 5032 1706
rect 4988 1680 5003 1700
rect 5023 1680 5032 1700
rect 4988 1664 5032 1680
rect 5102 1700 5146 1706
rect 5102 1680 5111 1700
rect 5131 1680 5146 1700
rect 5102 1664 5146 1680
rect 5196 1696 5245 1706
rect 5196 1676 5214 1696
rect 5234 1676 5245 1696
rect 5196 1664 5245 1676
rect 3342 1539 3391 1551
rect 3342 1519 3353 1539
rect 3373 1519 3391 1539
rect 3342 1509 3391 1519
rect 3441 1535 3485 1551
rect 3441 1515 3456 1535
rect 3476 1515 3485 1535
rect 3441 1509 3485 1515
rect 3555 1535 3599 1551
rect 3555 1515 3564 1535
rect 3584 1515 3599 1535
rect 3555 1509 3599 1515
rect 3649 1539 3698 1551
rect 3649 1519 3667 1539
rect 3687 1519 3698 1539
rect 3649 1509 3698 1519
rect 3773 1535 3817 1551
rect 3773 1515 3782 1535
rect 3802 1515 3817 1535
rect 3773 1509 3817 1515
rect 3867 1539 3916 1551
rect 3867 1519 3885 1539
rect 3905 1519 3916 1539
rect 3867 1509 3916 1519
rect 7706 1552 7755 1564
rect 7706 1532 7717 1552
rect 7737 1532 7755 1552
rect 7706 1522 7755 1532
rect 7805 1548 7849 1564
rect 7805 1528 7820 1548
rect 7840 1528 7849 1548
rect 7805 1522 7849 1528
rect 7919 1548 7963 1564
rect 7919 1528 7928 1548
rect 7948 1528 7963 1548
rect 7919 1522 7963 1528
rect 8013 1552 8062 1564
rect 8013 1532 8031 1552
rect 8051 1532 8062 1552
rect 8013 1522 8062 1532
rect 8137 1548 8181 1564
rect 8137 1528 8146 1548
rect 8166 1528 8181 1548
rect 8137 1522 8181 1528
rect 8231 1552 8280 1564
rect 8231 1532 8249 1552
rect 8269 1532 8280 1552
rect 8231 1522 8280 1532
rect 1186 1303 1235 1313
rect 1186 1283 1197 1303
rect 1217 1283 1235 1303
rect 1186 1271 1235 1283
rect 1285 1307 1329 1313
rect 1285 1287 1300 1307
rect 1320 1287 1329 1307
rect 1285 1271 1329 1287
rect 1404 1303 1453 1313
rect 1404 1283 1415 1303
rect 1435 1283 1453 1303
rect 1404 1271 1453 1283
rect 1503 1307 1547 1313
rect 1503 1287 1518 1307
rect 1538 1287 1547 1307
rect 1503 1271 1547 1287
rect 1617 1307 1661 1313
rect 1617 1287 1626 1307
rect 1646 1287 1661 1307
rect 1617 1271 1661 1287
rect 1711 1303 1760 1313
rect 1711 1283 1729 1303
rect 1749 1283 1760 1303
rect 1711 1271 1760 1283
rect 2545 1311 2594 1323
rect 2545 1291 2556 1311
rect 2576 1291 2594 1311
rect 2545 1281 2594 1291
rect 2644 1307 2688 1323
rect 2644 1287 2659 1307
rect 2679 1287 2688 1307
rect 2644 1281 2688 1287
rect 2758 1307 2802 1323
rect 2758 1287 2767 1307
rect 2787 1287 2802 1307
rect 2758 1281 2802 1287
rect 2852 1311 2901 1323
rect 2852 1291 2870 1311
rect 2890 1291 2901 1311
rect 2852 1281 2901 1291
rect 2976 1307 3020 1323
rect 2976 1287 2985 1307
rect 3005 1287 3020 1307
rect 2976 1281 3020 1287
rect 3070 1311 3119 1323
rect 3070 1291 3088 1311
rect 3108 1291 3119 1311
rect 3070 1281 3119 1291
rect 5550 1316 5599 1326
rect 5550 1296 5561 1316
rect 5581 1296 5599 1316
rect 5550 1284 5599 1296
rect 5649 1320 5693 1326
rect 5649 1300 5664 1320
rect 5684 1300 5693 1320
rect 5649 1284 5693 1300
rect 5768 1316 5817 1326
rect 5768 1296 5779 1316
rect 5799 1296 5817 1316
rect 5768 1284 5817 1296
rect 5867 1320 5911 1326
rect 5867 1300 5882 1320
rect 5902 1300 5911 1320
rect 5867 1284 5911 1300
rect 5981 1320 6025 1326
rect 5981 1300 5990 1320
rect 6010 1300 6025 1320
rect 5981 1284 6025 1300
rect 6075 1316 6124 1326
rect 6075 1296 6093 1316
rect 6113 1296 6124 1316
rect 6075 1284 6124 1296
rect 6909 1324 6958 1336
rect 6909 1304 6920 1324
rect 6940 1304 6958 1324
rect 6909 1294 6958 1304
rect 7008 1320 7052 1336
rect 7008 1300 7023 1320
rect 7043 1300 7052 1320
rect 7008 1294 7052 1300
rect 7122 1320 7166 1336
rect 7122 1300 7131 1320
rect 7151 1300 7166 1320
rect 7122 1294 7166 1300
rect 7216 1324 7265 1336
rect 7216 1304 7234 1324
rect 7254 1304 7265 1324
rect 7216 1294 7265 1304
rect 7340 1320 7384 1336
rect 7340 1300 7349 1320
rect 7369 1300 7384 1320
rect 7340 1294 7384 1300
rect 7434 1324 7483 1336
rect 7434 1304 7452 1324
rect 7472 1304 7483 1324
rect 7434 1294 7483 1304
rect 3343 1127 3392 1139
rect 3343 1107 3354 1127
rect 3374 1107 3392 1127
rect 289 1077 338 1087
rect 289 1057 300 1077
rect 320 1057 338 1077
rect 289 1045 338 1057
rect 388 1081 432 1087
rect 388 1061 403 1081
rect 423 1061 432 1081
rect 388 1045 432 1061
rect 507 1077 556 1087
rect 507 1057 518 1077
rect 538 1057 556 1077
rect 507 1045 556 1057
rect 606 1081 650 1087
rect 606 1061 621 1081
rect 641 1061 650 1081
rect 606 1045 650 1061
rect 720 1081 764 1087
rect 720 1061 729 1081
rect 749 1061 764 1081
rect 720 1045 764 1061
rect 814 1077 863 1087
rect 3343 1097 3392 1107
rect 3442 1123 3486 1139
rect 3442 1103 3457 1123
rect 3477 1103 3486 1123
rect 3442 1097 3486 1103
rect 3556 1123 3600 1139
rect 3556 1103 3565 1123
rect 3585 1103 3600 1123
rect 3556 1097 3600 1103
rect 3650 1127 3699 1139
rect 3650 1107 3668 1127
rect 3688 1107 3699 1127
rect 3650 1097 3699 1107
rect 3774 1123 3818 1139
rect 3774 1103 3783 1123
rect 3803 1103 3818 1123
rect 3774 1097 3818 1103
rect 3868 1127 3917 1139
rect 3868 1107 3886 1127
rect 3906 1107 3917 1127
rect 3868 1097 3917 1107
rect 814 1057 832 1077
rect 852 1057 863 1077
rect 814 1045 863 1057
rect 7707 1140 7756 1152
rect 7707 1120 7718 1140
rect 7738 1120 7756 1140
rect 4653 1090 4702 1100
rect 4653 1070 4664 1090
rect 4684 1070 4702 1090
rect 4653 1058 4702 1070
rect 4752 1094 4796 1100
rect 4752 1074 4767 1094
rect 4787 1074 4796 1094
rect 4752 1058 4796 1074
rect 4871 1090 4920 1100
rect 4871 1070 4882 1090
rect 4902 1070 4920 1090
rect 4871 1058 4920 1070
rect 4970 1094 5014 1100
rect 4970 1074 4985 1094
rect 5005 1074 5014 1094
rect 4970 1058 5014 1074
rect 5084 1094 5128 1100
rect 5084 1074 5093 1094
rect 5113 1074 5128 1094
rect 5084 1058 5128 1074
rect 5178 1090 5227 1100
rect 7707 1110 7756 1120
rect 7806 1136 7850 1152
rect 7806 1116 7821 1136
rect 7841 1116 7850 1136
rect 7806 1110 7850 1116
rect 7920 1136 7964 1152
rect 7920 1116 7929 1136
rect 7949 1116 7964 1136
rect 7920 1110 7964 1116
rect 8014 1140 8063 1152
rect 8014 1120 8032 1140
rect 8052 1120 8063 1140
rect 8014 1110 8063 1120
rect 8138 1136 8182 1152
rect 8138 1116 8147 1136
rect 8167 1116 8182 1136
rect 8138 1110 8182 1116
rect 8232 1140 8281 1152
rect 8232 1120 8250 1140
rect 8270 1120 8281 1140
rect 8232 1110 8281 1120
rect 5178 1070 5196 1090
rect 5216 1070 5227 1090
rect 5178 1058 5227 1070
rect 1087 893 1136 903
rect 1087 873 1098 893
rect 1118 873 1136 893
rect 1087 861 1136 873
rect 1186 897 1230 903
rect 1186 877 1201 897
rect 1221 877 1230 897
rect 1186 861 1230 877
rect 1305 893 1354 903
rect 1305 873 1316 893
rect 1336 873 1354 893
rect 1305 861 1354 873
rect 1404 897 1448 903
rect 1404 877 1419 897
rect 1439 877 1448 897
rect 1404 861 1448 877
rect 1518 897 1562 903
rect 1518 877 1527 897
rect 1547 877 1562 897
rect 1518 861 1562 877
rect 1612 893 1661 903
rect 1612 873 1630 893
rect 1650 873 1661 893
rect 1612 861 1661 873
rect 5451 906 5500 916
rect 5451 886 5462 906
rect 5482 886 5500 906
rect 5451 874 5500 886
rect 5550 910 5594 916
rect 5550 890 5565 910
rect 5585 890 5594 910
rect 5550 874 5594 890
rect 5669 906 5718 916
rect 5669 886 5680 906
rect 5700 886 5718 906
rect 5669 874 5718 886
rect 5768 910 5812 916
rect 5768 890 5783 910
rect 5803 890 5812 910
rect 5768 874 5812 890
rect 5882 910 5926 916
rect 5882 890 5891 910
rect 5911 890 5926 910
rect 5882 874 5926 890
rect 5976 906 6025 916
rect 5976 886 5994 906
rect 6014 886 6025 906
rect 5976 874 6025 886
rect 290 665 339 675
rect 290 645 301 665
rect 321 645 339 665
rect 290 633 339 645
rect 389 669 433 675
rect 389 649 404 669
rect 424 649 433 669
rect 389 633 433 649
rect 508 665 557 675
rect 508 645 519 665
rect 539 645 557 665
rect 508 633 557 645
rect 607 669 651 675
rect 607 649 622 669
rect 642 649 651 669
rect 607 633 651 649
rect 721 669 765 675
rect 721 649 730 669
rect 750 649 765 669
rect 721 633 765 649
rect 815 665 864 675
rect 815 645 833 665
rect 853 645 864 665
rect 815 633 864 645
rect 4654 678 4703 688
rect 4654 658 4665 678
rect 4685 658 4703 678
rect 4654 646 4703 658
rect 4753 682 4797 688
rect 4753 662 4768 682
rect 4788 662 4797 682
rect 4753 646 4797 662
rect 4872 678 4921 688
rect 4872 658 4883 678
rect 4903 658 4921 678
rect 4872 646 4921 658
rect 4971 682 5015 688
rect 4971 662 4986 682
rect 5006 662 5015 682
rect 4971 646 5015 662
rect 5085 682 5129 688
rect 5085 662 5094 682
rect 5114 662 5129 682
rect 5085 646 5129 662
rect 5179 678 5228 688
rect 5179 658 5197 678
rect 5217 658 5228 678
rect 5179 646 5228 658
rect 5867 102 5916 112
rect 1503 89 1552 99
rect 1503 69 1514 89
rect 1534 69 1552 89
rect 1503 57 1552 69
rect 1602 93 1646 99
rect 1602 73 1617 93
rect 1637 73 1646 93
rect 1602 57 1646 73
rect 1721 89 1770 99
rect 1721 69 1732 89
rect 1752 69 1770 89
rect 1721 57 1770 69
rect 1820 93 1864 99
rect 1820 73 1835 93
rect 1855 73 1864 93
rect 1820 57 1864 73
rect 1934 93 1978 99
rect 1934 73 1943 93
rect 1963 73 1978 93
rect 1934 57 1978 73
rect 2028 89 2077 99
rect 2028 69 2046 89
rect 2066 69 2077 89
rect 2028 57 2077 69
rect 5867 82 5878 102
rect 5898 82 5916 102
rect 5867 70 5916 82
rect 5966 106 6010 112
rect 5966 86 5981 106
rect 6001 86 6010 106
rect 5966 70 6010 86
rect 6085 102 6134 112
rect 6085 82 6096 102
rect 6116 82 6134 102
rect 6085 70 6134 82
rect 6184 106 6228 112
rect 6184 86 6199 106
rect 6219 86 6228 106
rect 6184 70 6228 86
rect 6298 106 6342 112
rect 6298 86 6307 106
rect 6327 86 6342 106
rect 6298 70 6342 86
rect 6392 102 6441 112
rect 6392 82 6410 102
rect 6430 82 6441 102
rect 6392 70 6441 82
rect 3992 15 4041 25
rect 3992 -5 4003 15
rect 4023 -5 4041 15
rect 3992 -17 4041 -5
rect 4091 19 4135 25
rect 4091 -1 4106 19
rect 4126 -1 4135 19
rect 4091 -17 4135 -1
rect 4210 15 4259 25
rect 4210 -5 4221 15
rect 4241 -5 4259 15
rect 4210 -17 4259 -5
rect 4309 19 4353 25
rect 4309 -1 4324 19
rect 4344 -1 4353 19
rect 4309 -17 4353 -1
rect 4423 19 4467 25
rect 4423 -1 4432 19
rect 4452 -1 4467 19
rect 4423 -17 4467 -1
rect 4517 15 4566 25
rect 4517 -5 4535 15
rect 4555 -5 4566 15
rect 4517 -17 4566 -5
<< pdiff >>
rect 3474 8516 3518 8558
rect 3474 8496 3486 8516
rect 3506 8496 3518 8516
rect 3474 8489 3518 8496
rect 3473 8458 3518 8489
rect 3568 8516 3610 8558
rect 3568 8496 3582 8516
rect 3602 8496 3610 8516
rect 3568 8458 3610 8496
rect 3684 8516 3726 8558
rect 3684 8496 3692 8516
rect 3712 8496 3726 8516
rect 3684 8458 3726 8496
rect 3776 8516 3820 8558
rect 3776 8496 3788 8516
rect 3808 8496 3820 8516
rect 3776 8458 3820 8496
rect 3902 8516 3944 8558
rect 3902 8496 3910 8516
rect 3930 8496 3944 8516
rect 3902 8458 3944 8496
rect 3994 8516 4038 8558
rect 3994 8496 4006 8516
rect 4026 8496 4038 8516
rect 3994 8458 4038 8496
rect 7838 8529 7882 8571
rect 7838 8509 7850 8529
rect 7870 8509 7882 8529
rect 7838 8502 7882 8509
rect 7837 8471 7882 8502
rect 7932 8529 7974 8571
rect 7932 8509 7946 8529
rect 7966 8509 7974 8529
rect 7932 8471 7974 8509
rect 8048 8529 8090 8571
rect 8048 8509 8056 8529
rect 8076 8509 8090 8529
rect 8048 8471 8090 8509
rect 8140 8529 8184 8571
rect 8140 8509 8152 8529
rect 8172 8509 8184 8529
rect 8140 8471 8184 8509
rect 8266 8529 8308 8571
rect 8266 8509 8274 8529
rect 8294 8509 8308 8529
rect 8266 8471 8308 8509
rect 8358 8529 8402 8571
rect 8358 8509 8370 8529
rect 8390 8509 8402 8529
rect 8358 8471 8402 8509
rect 421 8352 465 8390
rect 421 8332 433 8352
rect 453 8332 465 8352
rect 421 8290 465 8332
rect 515 8352 557 8390
rect 515 8332 529 8352
rect 549 8332 557 8352
rect 515 8290 557 8332
rect 639 8352 683 8390
rect 639 8332 651 8352
rect 671 8332 683 8352
rect 639 8290 683 8332
rect 733 8352 775 8390
rect 733 8332 747 8352
rect 767 8332 775 8352
rect 733 8290 775 8332
rect 849 8352 891 8390
rect 849 8332 857 8352
rect 877 8332 891 8352
rect 849 8290 891 8332
rect 941 8359 986 8390
rect 941 8352 985 8359
rect 941 8332 953 8352
rect 973 8332 985 8352
rect 941 8290 985 8332
rect 4785 8365 4829 8403
rect 4785 8345 4797 8365
rect 4817 8345 4829 8365
rect 2677 8288 2721 8330
rect 2677 8268 2689 8288
rect 2709 8268 2721 8288
rect 2677 8261 2721 8268
rect 2676 8230 2721 8261
rect 2771 8288 2813 8330
rect 2771 8268 2785 8288
rect 2805 8268 2813 8288
rect 2771 8230 2813 8268
rect 2887 8288 2929 8330
rect 2887 8268 2895 8288
rect 2915 8268 2929 8288
rect 2887 8230 2929 8268
rect 2979 8288 3023 8330
rect 2979 8268 2991 8288
rect 3011 8268 3023 8288
rect 2979 8230 3023 8268
rect 3105 8288 3147 8330
rect 3105 8268 3113 8288
rect 3133 8268 3147 8288
rect 3105 8230 3147 8268
rect 3197 8288 3241 8330
rect 4785 8303 4829 8345
rect 4879 8365 4921 8403
rect 4879 8345 4893 8365
rect 4913 8345 4921 8365
rect 4879 8303 4921 8345
rect 5003 8365 5047 8403
rect 5003 8345 5015 8365
rect 5035 8345 5047 8365
rect 5003 8303 5047 8345
rect 5097 8365 5139 8403
rect 5097 8345 5111 8365
rect 5131 8345 5139 8365
rect 5097 8303 5139 8345
rect 5213 8365 5255 8403
rect 5213 8345 5221 8365
rect 5241 8345 5255 8365
rect 5213 8303 5255 8345
rect 5305 8372 5350 8403
rect 5305 8365 5349 8372
rect 5305 8345 5317 8365
rect 5337 8345 5349 8365
rect 5305 8303 5349 8345
rect 3197 8268 3209 8288
rect 3229 8268 3241 8288
rect 3197 8230 3241 8268
rect 1219 8168 1263 8206
rect 1219 8148 1231 8168
rect 1251 8148 1263 8168
rect 1219 8106 1263 8148
rect 1313 8168 1355 8206
rect 1313 8148 1327 8168
rect 1347 8148 1355 8168
rect 1313 8106 1355 8148
rect 1437 8168 1481 8206
rect 1437 8148 1449 8168
rect 1469 8148 1481 8168
rect 1437 8106 1481 8148
rect 1531 8168 1573 8206
rect 1531 8148 1545 8168
rect 1565 8148 1573 8168
rect 1531 8106 1573 8148
rect 1647 8168 1689 8206
rect 1647 8148 1655 8168
rect 1675 8148 1689 8168
rect 1647 8106 1689 8148
rect 1739 8175 1784 8206
rect 1739 8168 1783 8175
rect 1739 8148 1751 8168
rect 1771 8148 1783 8168
rect 1739 8106 1783 8148
rect 7041 8301 7085 8343
rect 7041 8281 7053 8301
rect 7073 8281 7085 8301
rect 7041 8274 7085 8281
rect 7040 8243 7085 8274
rect 7135 8301 7177 8343
rect 7135 8281 7149 8301
rect 7169 8281 7177 8301
rect 7135 8243 7177 8281
rect 7251 8301 7293 8343
rect 7251 8281 7259 8301
rect 7279 8281 7293 8301
rect 7251 8243 7293 8281
rect 7343 8301 7387 8343
rect 7343 8281 7355 8301
rect 7375 8281 7387 8301
rect 7343 8243 7387 8281
rect 7469 8301 7511 8343
rect 7469 8281 7477 8301
rect 7497 8281 7511 8301
rect 7469 8243 7511 8281
rect 7561 8301 7605 8343
rect 7561 8281 7573 8301
rect 7593 8281 7605 8301
rect 7561 8243 7605 8281
rect 5583 8181 5627 8219
rect 5583 8161 5595 8181
rect 5615 8161 5627 8181
rect 3475 8104 3519 8146
rect 3475 8084 3487 8104
rect 3507 8084 3519 8104
rect 3475 8077 3519 8084
rect 3474 8046 3519 8077
rect 3569 8104 3611 8146
rect 3569 8084 3583 8104
rect 3603 8084 3611 8104
rect 3569 8046 3611 8084
rect 3685 8104 3727 8146
rect 3685 8084 3693 8104
rect 3713 8084 3727 8104
rect 3685 8046 3727 8084
rect 3777 8104 3821 8146
rect 3777 8084 3789 8104
rect 3809 8084 3821 8104
rect 3777 8046 3821 8084
rect 3903 8104 3945 8146
rect 3903 8084 3911 8104
rect 3931 8084 3945 8104
rect 3903 8046 3945 8084
rect 3995 8104 4039 8146
rect 5583 8119 5627 8161
rect 5677 8181 5719 8219
rect 5677 8161 5691 8181
rect 5711 8161 5719 8181
rect 5677 8119 5719 8161
rect 5801 8181 5845 8219
rect 5801 8161 5813 8181
rect 5833 8161 5845 8181
rect 5801 8119 5845 8161
rect 5895 8181 5937 8219
rect 5895 8161 5909 8181
rect 5929 8161 5937 8181
rect 5895 8119 5937 8161
rect 6011 8181 6053 8219
rect 6011 8161 6019 8181
rect 6039 8161 6053 8181
rect 6011 8119 6053 8161
rect 6103 8188 6148 8219
rect 6103 8181 6147 8188
rect 6103 8161 6115 8181
rect 6135 8161 6147 8181
rect 6103 8119 6147 8161
rect 3995 8084 4007 8104
rect 4027 8084 4039 8104
rect 3995 8046 4039 8084
rect 7839 8117 7883 8159
rect 7839 8097 7851 8117
rect 7871 8097 7883 8117
rect 7839 8090 7883 8097
rect 7838 8059 7883 8090
rect 7933 8117 7975 8159
rect 7933 8097 7947 8117
rect 7967 8097 7975 8117
rect 7933 8059 7975 8097
rect 8049 8117 8091 8159
rect 8049 8097 8057 8117
rect 8077 8097 8091 8117
rect 8049 8059 8091 8097
rect 8141 8117 8185 8159
rect 8141 8097 8153 8117
rect 8173 8097 8185 8117
rect 8141 8059 8185 8097
rect 8267 8117 8309 8159
rect 8267 8097 8275 8117
rect 8295 8097 8309 8117
rect 8267 8059 8309 8097
rect 8359 8117 8403 8159
rect 8359 8097 8371 8117
rect 8391 8097 8403 8117
rect 8359 8059 8403 8097
rect 422 7940 466 7978
rect 422 7920 434 7940
rect 454 7920 466 7940
rect 422 7878 466 7920
rect 516 7940 558 7978
rect 516 7920 530 7940
rect 550 7920 558 7940
rect 516 7878 558 7920
rect 640 7940 684 7978
rect 640 7920 652 7940
rect 672 7920 684 7940
rect 640 7878 684 7920
rect 734 7940 776 7978
rect 734 7920 748 7940
rect 768 7920 776 7940
rect 734 7878 776 7920
rect 850 7940 892 7978
rect 850 7920 858 7940
rect 878 7920 892 7940
rect 850 7878 892 7920
rect 942 7947 987 7978
rect 942 7940 986 7947
rect 942 7920 954 7940
rect 974 7920 986 7940
rect 4786 7953 4830 7991
rect 942 7878 986 7920
rect 2578 7878 2622 7920
rect 2578 7858 2590 7878
rect 2610 7858 2622 7878
rect 2578 7851 2622 7858
rect 2577 7820 2622 7851
rect 2672 7878 2714 7920
rect 2672 7858 2686 7878
rect 2706 7858 2714 7878
rect 2672 7820 2714 7858
rect 2788 7878 2830 7920
rect 2788 7858 2796 7878
rect 2816 7858 2830 7878
rect 2788 7820 2830 7858
rect 2880 7878 2924 7920
rect 2880 7858 2892 7878
rect 2912 7858 2924 7878
rect 2880 7820 2924 7858
rect 3006 7878 3048 7920
rect 3006 7858 3014 7878
rect 3034 7858 3048 7878
rect 3006 7820 3048 7858
rect 3098 7878 3142 7920
rect 4786 7933 4798 7953
rect 4818 7933 4830 7953
rect 3098 7858 3110 7878
rect 3130 7858 3142 7878
rect 4786 7891 4830 7933
rect 4880 7953 4922 7991
rect 4880 7933 4894 7953
rect 4914 7933 4922 7953
rect 4880 7891 4922 7933
rect 5004 7953 5048 7991
rect 5004 7933 5016 7953
rect 5036 7933 5048 7953
rect 5004 7891 5048 7933
rect 5098 7953 5140 7991
rect 5098 7933 5112 7953
rect 5132 7933 5140 7953
rect 5098 7891 5140 7933
rect 5214 7953 5256 7991
rect 5214 7933 5222 7953
rect 5242 7933 5256 7953
rect 5214 7891 5256 7933
rect 5306 7960 5351 7991
rect 5306 7953 5350 7960
rect 5306 7933 5318 7953
rect 5338 7933 5350 7953
rect 5306 7891 5350 7933
rect 6942 7891 6986 7933
rect 3098 7820 3142 7858
rect 6942 7871 6954 7891
rect 6974 7871 6986 7891
rect 6942 7864 6986 7871
rect 6941 7833 6986 7864
rect 7036 7891 7078 7933
rect 7036 7871 7050 7891
rect 7070 7871 7078 7891
rect 7036 7833 7078 7871
rect 7152 7891 7194 7933
rect 7152 7871 7160 7891
rect 7180 7871 7194 7891
rect 7152 7833 7194 7871
rect 7244 7891 7288 7933
rect 7244 7871 7256 7891
rect 7276 7871 7288 7891
rect 7244 7833 7288 7871
rect 7370 7891 7412 7933
rect 7370 7871 7378 7891
rect 7398 7871 7412 7891
rect 7370 7833 7412 7871
rect 7462 7891 7506 7933
rect 7462 7871 7474 7891
rect 7494 7871 7506 7891
rect 7462 7833 7506 7871
rect 1301 7560 1345 7598
rect 1301 7540 1313 7560
rect 1333 7540 1345 7560
rect 1301 7498 1345 7540
rect 1395 7560 1437 7598
rect 1395 7540 1409 7560
rect 1429 7540 1437 7560
rect 1395 7498 1437 7540
rect 1519 7560 1563 7598
rect 1519 7540 1531 7560
rect 1551 7540 1563 7560
rect 1519 7498 1563 7540
rect 1613 7560 1655 7598
rect 1613 7540 1627 7560
rect 1647 7540 1655 7560
rect 1613 7498 1655 7540
rect 1729 7560 1771 7598
rect 1729 7540 1737 7560
rect 1757 7540 1771 7560
rect 1729 7498 1771 7540
rect 1821 7567 1866 7598
rect 1821 7560 1865 7567
rect 1821 7540 1833 7560
rect 1853 7540 1865 7560
rect 5665 7573 5709 7611
rect 1821 7498 1865 7540
rect 3457 7498 3501 7540
rect 3457 7478 3469 7498
rect 3489 7478 3501 7498
rect 3457 7471 3501 7478
rect 3456 7440 3501 7471
rect 3551 7498 3593 7540
rect 3551 7478 3565 7498
rect 3585 7478 3593 7498
rect 3551 7440 3593 7478
rect 3667 7498 3709 7540
rect 3667 7478 3675 7498
rect 3695 7478 3709 7498
rect 3667 7440 3709 7478
rect 3759 7498 3803 7540
rect 3759 7478 3771 7498
rect 3791 7478 3803 7498
rect 3759 7440 3803 7478
rect 3885 7498 3927 7540
rect 3885 7478 3893 7498
rect 3913 7478 3927 7498
rect 3885 7440 3927 7478
rect 3977 7498 4021 7540
rect 5665 7553 5677 7573
rect 5697 7553 5709 7573
rect 3977 7478 3989 7498
rect 4009 7478 4021 7498
rect 5665 7511 5709 7553
rect 5759 7573 5801 7611
rect 5759 7553 5773 7573
rect 5793 7553 5801 7573
rect 5759 7511 5801 7553
rect 5883 7573 5927 7611
rect 5883 7553 5895 7573
rect 5915 7553 5927 7573
rect 5883 7511 5927 7553
rect 5977 7573 6019 7611
rect 5977 7553 5991 7573
rect 6011 7553 6019 7573
rect 5977 7511 6019 7553
rect 6093 7573 6135 7611
rect 6093 7553 6101 7573
rect 6121 7553 6135 7573
rect 6093 7511 6135 7553
rect 6185 7580 6230 7611
rect 6185 7573 6229 7580
rect 6185 7553 6197 7573
rect 6217 7553 6229 7573
rect 6185 7511 6229 7553
rect 7821 7511 7865 7553
rect 3977 7440 4021 7478
rect 7821 7491 7833 7511
rect 7853 7491 7865 7511
rect 7821 7484 7865 7491
rect 7820 7453 7865 7484
rect 7915 7511 7957 7553
rect 7915 7491 7929 7511
rect 7949 7491 7957 7511
rect 7915 7453 7957 7491
rect 8031 7511 8073 7553
rect 8031 7491 8039 7511
rect 8059 7491 8073 7511
rect 8031 7453 8073 7491
rect 8123 7511 8167 7553
rect 8123 7491 8135 7511
rect 8155 7491 8167 7511
rect 8123 7453 8167 7491
rect 8249 7511 8291 7553
rect 8249 7491 8257 7511
rect 8277 7491 8291 7511
rect 8249 7453 8291 7491
rect 8341 7511 8385 7553
rect 8341 7491 8353 7511
rect 8373 7491 8385 7511
rect 8341 7453 8385 7491
rect 404 7334 448 7372
rect 404 7314 416 7334
rect 436 7314 448 7334
rect 404 7272 448 7314
rect 498 7334 540 7372
rect 498 7314 512 7334
rect 532 7314 540 7334
rect 498 7272 540 7314
rect 622 7334 666 7372
rect 622 7314 634 7334
rect 654 7314 666 7334
rect 622 7272 666 7314
rect 716 7334 758 7372
rect 716 7314 730 7334
rect 750 7314 758 7334
rect 716 7272 758 7314
rect 832 7334 874 7372
rect 832 7314 840 7334
rect 860 7314 874 7334
rect 832 7272 874 7314
rect 924 7341 969 7372
rect 924 7334 968 7341
rect 924 7314 936 7334
rect 956 7314 968 7334
rect 924 7272 968 7314
rect 4768 7347 4812 7385
rect 4768 7327 4780 7347
rect 4800 7327 4812 7347
rect 2660 7270 2704 7312
rect 2660 7250 2672 7270
rect 2692 7250 2704 7270
rect 2660 7243 2704 7250
rect 2659 7212 2704 7243
rect 2754 7270 2796 7312
rect 2754 7250 2768 7270
rect 2788 7250 2796 7270
rect 2754 7212 2796 7250
rect 2870 7270 2912 7312
rect 2870 7250 2878 7270
rect 2898 7250 2912 7270
rect 2870 7212 2912 7250
rect 2962 7270 3006 7312
rect 2962 7250 2974 7270
rect 2994 7250 3006 7270
rect 2962 7212 3006 7250
rect 3088 7270 3130 7312
rect 3088 7250 3096 7270
rect 3116 7250 3130 7270
rect 3088 7212 3130 7250
rect 3180 7270 3224 7312
rect 4768 7285 4812 7327
rect 4862 7347 4904 7385
rect 4862 7327 4876 7347
rect 4896 7327 4904 7347
rect 4862 7285 4904 7327
rect 4986 7347 5030 7385
rect 4986 7327 4998 7347
rect 5018 7327 5030 7347
rect 4986 7285 5030 7327
rect 5080 7347 5122 7385
rect 5080 7327 5094 7347
rect 5114 7327 5122 7347
rect 5080 7285 5122 7327
rect 5196 7347 5238 7385
rect 5196 7327 5204 7347
rect 5224 7327 5238 7347
rect 5196 7285 5238 7327
rect 5288 7354 5333 7385
rect 5288 7347 5332 7354
rect 5288 7327 5300 7347
rect 5320 7327 5332 7347
rect 5288 7285 5332 7327
rect 3180 7250 3192 7270
rect 3212 7250 3224 7270
rect 3180 7212 3224 7250
rect 1202 7150 1246 7188
rect 1202 7130 1214 7150
rect 1234 7130 1246 7150
rect 1202 7088 1246 7130
rect 1296 7150 1338 7188
rect 1296 7130 1310 7150
rect 1330 7130 1338 7150
rect 1296 7088 1338 7130
rect 1420 7150 1464 7188
rect 1420 7130 1432 7150
rect 1452 7130 1464 7150
rect 1420 7088 1464 7130
rect 1514 7150 1556 7188
rect 1514 7130 1528 7150
rect 1548 7130 1556 7150
rect 1514 7088 1556 7130
rect 1630 7150 1672 7188
rect 1630 7130 1638 7150
rect 1658 7130 1672 7150
rect 1630 7088 1672 7130
rect 1722 7157 1767 7188
rect 1722 7150 1766 7157
rect 1722 7130 1734 7150
rect 1754 7130 1766 7150
rect 1722 7088 1766 7130
rect 7024 7283 7068 7325
rect 7024 7263 7036 7283
rect 7056 7263 7068 7283
rect 7024 7256 7068 7263
rect 7023 7225 7068 7256
rect 7118 7283 7160 7325
rect 7118 7263 7132 7283
rect 7152 7263 7160 7283
rect 7118 7225 7160 7263
rect 7234 7283 7276 7325
rect 7234 7263 7242 7283
rect 7262 7263 7276 7283
rect 7234 7225 7276 7263
rect 7326 7283 7370 7325
rect 7326 7263 7338 7283
rect 7358 7263 7370 7283
rect 7326 7225 7370 7263
rect 7452 7283 7494 7325
rect 7452 7263 7460 7283
rect 7480 7263 7494 7283
rect 7452 7225 7494 7263
rect 7544 7283 7588 7325
rect 7544 7263 7556 7283
rect 7576 7263 7588 7283
rect 7544 7225 7588 7263
rect 5566 7163 5610 7201
rect 5566 7143 5578 7163
rect 5598 7143 5610 7163
rect 3458 7086 3502 7128
rect 3458 7066 3470 7086
rect 3490 7066 3502 7086
rect 3458 7059 3502 7066
rect 3457 7028 3502 7059
rect 3552 7086 3594 7128
rect 3552 7066 3566 7086
rect 3586 7066 3594 7086
rect 3552 7028 3594 7066
rect 3668 7086 3710 7128
rect 3668 7066 3676 7086
rect 3696 7066 3710 7086
rect 3668 7028 3710 7066
rect 3760 7086 3804 7128
rect 3760 7066 3772 7086
rect 3792 7066 3804 7086
rect 3760 7028 3804 7066
rect 3886 7086 3928 7128
rect 3886 7066 3894 7086
rect 3914 7066 3928 7086
rect 3886 7028 3928 7066
rect 3978 7086 4022 7128
rect 5566 7101 5610 7143
rect 5660 7163 5702 7201
rect 5660 7143 5674 7163
rect 5694 7143 5702 7163
rect 5660 7101 5702 7143
rect 5784 7163 5828 7201
rect 5784 7143 5796 7163
rect 5816 7143 5828 7163
rect 5784 7101 5828 7143
rect 5878 7163 5920 7201
rect 5878 7143 5892 7163
rect 5912 7143 5920 7163
rect 5878 7101 5920 7143
rect 5994 7163 6036 7201
rect 5994 7143 6002 7163
rect 6022 7143 6036 7163
rect 5994 7101 6036 7143
rect 6086 7170 6131 7201
rect 6086 7163 6130 7170
rect 6086 7143 6098 7163
rect 6118 7143 6130 7163
rect 6086 7101 6130 7143
rect 3978 7066 3990 7086
rect 4010 7066 4022 7086
rect 3978 7028 4022 7066
rect 7822 7099 7866 7141
rect 7822 7079 7834 7099
rect 7854 7079 7866 7099
rect 7822 7072 7866 7079
rect 7821 7041 7866 7072
rect 7916 7099 7958 7141
rect 7916 7079 7930 7099
rect 7950 7079 7958 7099
rect 7916 7041 7958 7079
rect 8032 7099 8074 7141
rect 8032 7079 8040 7099
rect 8060 7079 8074 7099
rect 8032 7041 8074 7079
rect 8124 7099 8168 7141
rect 8124 7079 8136 7099
rect 8156 7079 8168 7099
rect 8124 7041 8168 7079
rect 8250 7099 8292 7141
rect 8250 7079 8258 7099
rect 8278 7079 8292 7099
rect 8250 7041 8292 7079
rect 8342 7099 8386 7141
rect 8342 7079 8354 7099
rect 8374 7079 8386 7099
rect 8342 7041 8386 7079
rect 405 6922 449 6960
rect 405 6902 417 6922
rect 437 6902 449 6922
rect 405 6860 449 6902
rect 499 6922 541 6960
rect 499 6902 513 6922
rect 533 6902 541 6922
rect 499 6860 541 6902
rect 623 6922 667 6960
rect 623 6902 635 6922
rect 655 6902 667 6922
rect 623 6860 667 6902
rect 717 6922 759 6960
rect 717 6902 731 6922
rect 751 6902 759 6922
rect 717 6860 759 6902
rect 833 6922 875 6960
rect 833 6902 841 6922
rect 861 6902 875 6922
rect 833 6860 875 6902
rect 925 6929 970 6960
rect 925 6922 969 6929
rect 925 6902 937 6922
rect 957 6902 969 6922
rect 4769 6935 4813 6973
rect 925 6860 969 6902
rect 2495 6862 2539 6904
rect 2495 6842 2507 6862
rect 2527 6842 2539 6862
rect 2495 6835 2539 6842
rect 2494 6804 2539 6835
rect 2589 6862 2631 6904
rect 2589 6842 2603 6862
rect 2623 6842 2631 6862
rect 2589 6804 2631 6842
rect 2705 6862 2747 6904
rect 2705 6842 2713 6862
rect 2733 6842 2747 6862
rect 2705 6804 2747 6842
rect 2797 6862 2841 6904
rect 2797 6842 2809 6862
rect 2829 6842 2841 6862
rect 2797 6804 2841 6842
rect 2923 6862 2965 6904
rect 2923 6842 2931 6862
rect 2951 6842 2965 6862
rect 2923 6804 2965 6842
rect 3015 6862 3059 6904
rect 4769 6915 4781 6935
rect 4801 6915 4813 6935
rect 3015 6842 3027 6862
rect 3047 6842 3059 6862
rect 4769 6873 4813 6915
rect 4863 6935 4905 6973
rect 4863 6915 4877 6935
rect 4897 6915 4905 6935
rect 4863 6873 4905 6915
rect 4987 6935 5031 6973
rect 4987 6915 4999 6935
rect 5019 6915 5031 6935
rect 4987 6873 5031 6915
rect 5081 6935 5123 6973
rect 5081 6915 5095 6935
rect 5115 6915 5123 6935
rect 5081 6873 5123 6915
rect 5197 6935 5239 6973
rect 5197 6915 5205 6935
rect 5225 6915 5239 6935
rect 5197 6873 5239 6915
rect 5289 6942 5334 6973
rect 5289 6935 5333 6942
rect 5289 6915 5301 6935
rect 5321 6915 5333 6935
rect 5289 6873 5333 6915
rect 6859 6875 6903 6917
rect 3015 6804 3059 6842
rect 6859 6855 6871 6875
rect 6891 6855 6903 6875
rect 6859 6848 6903 6855
rect 6858 6817 6903 6848
rect 6953 6875 6995 6917
rect 6953 6855 6967 6875
rect 6987 6855 6995 6875
rect 6953 6817 6995 6855
rect 7069 6875 7111 6917
rect 7069 6855 7077 6875
rect 7097 6855 7111 6875
rect 7069 6817 7111 6855
rect 7161 6875 7205 6917
rect 7161 6855 7173 6875
rect 7193 6855 7205 6875
rect 7161 6817 7205 6855
rect 7287 6875 7329 6917
rect 7287 6855 7295 6875
rect 7315 6855 7329 6875
rect 7287 6817 7329 6855
rect 7379 6875 7423 6917
rect 7379 6855 7391 6875
rect 7411 6855 7423 6875
rect 7379 6817 7423 6855
rect 1347 6540 1391 6578
rect 1347 6520 1359 6540
rect 1379 6520 1391 6540
rect 1347 6478 1391 6520
rect 1441 6540 1483 6578
rect 1441 6520 1455 6540
rect 1475 6520 1483 6540
rect 1441 6478 1483 6520
rect 1565 6540 1609 6578
rect 1565 6520 1577 6540
rect 1597 6520 1609 6540
rect 1565 6478 1609 6520
rect 1659 6540 1701 6578
rect 1659 6520 1673 6540
rect 1693 6520 1701 6540
rect 1659 6478 1701 6520
rect 1775 6540 1817 6578
rect 1775 6520 1783 6540
rect 1803 6520 1817 6540
rect 1775 6478 1817 6520
rect 1867 6547 1912 6578
rect 1867 6540 1911 6547
rect 1867 6520 1879 6540
rect 1899 6520 1911 6540
rect 5711 6553 5755 6591
rect 1867 6478 1911 6520
rect 3437 6480 3481 6522
rect 3437 6460 3449 6480
rect 3469 6460 3481 6480
rect 3437 6453 3481 6460
rect 3436 6422 3481 6453
rect 3531 6480 3573 6522
rect 3531 6460 3545 6480
rect 3565 6460 3573 6480
rect 3531 6422 3573 6460
rect 3647 6480 3689 6522
rect 3647 6460 3655 6480
rect 3675 6460 3689 6480
rect 3647 6422 3689 6460
rect 3739 6480 3783 6522
rect 3739 6460 3751 6480
rect 3771 6460 3783 6480
rect 3739 6422 3783 6460
rect 3865 6480 3907 6522
rect 3865 6460 3873 6480
rect 3893 6460 3907 6480
rect 3865 6422 3907 6460
rect 3957 6480 4001 6522
rect 5711 6533 5723 6553
rect 5743 6533 5755 6553
rect 3957 6460 3969 6480
rect 3989 6460 4001 6480
rect 5711 6491 5755 6533
rect 5805 6553 5847 6591
rect 5805 6533 5819 6553
rect 5839 6533 5847 6553
rect 5805 6491 5847 6533
rect 5929 6553 5973 6591
rect 5929 6533 5941 6553
rect 5961 6533 5973 6553
rect 5929 6491 5973 6533
rect 6023 6553 6065 6591
rect 6023 6533 6037 6553
rect 6057 6533 6065 6553
rect 6023 6491 6065 6533
rect 6139 6553 6181 6591
rect 6139 6533 6147 6553
rect 6167 6533 6181 6553
rect 6139 6491 6181 6533
rect 6231 6560 6276 6591
rect 6231 6553 6275 6560
rect 6231 6533 6243 6553
rect 6263 6533 6275 6553
rect 6231 6491 6275 6533
rect 7801 6493 7845 6535
rect 3957 6422 4001 6460
rect 7801 6473 7813 6493
rect 7833 6473 7845 6493
rect 7801 6466 7845 6473
rect 7800 6435 7845 6466
rect 7895 6493 7937 6535
rect 7895 6473 7909 6493
rect 7929 6473 7937 6493
rect 7895 6435 7937 6473
rect 8011 6493 8053 6535
rect 8011 6473 8019 6493
rect 8039 6473 8053 6493
rect 8011 6435 8053 6473
rect 8103 6493 8147 6535
rect 8103 6473 8115 6493
rect 8135 6473 8147 6493
rect 8103 6435 8147 6473
rect 8229 6493 8271 6535
rect 8229 6473 8237 6493
rect 8257 6473 8271 6493
rect 8229 6435 8271 6473
rect 8321 6493 8365 6535
rect 8321 6473 8333 6493
rect 8353 6473 8365 6493
rect 8321 6435 8365 6473
rect 384 6316 428 6354
rect 384 6296 396 6316
rect 416 6296 428 6316
rect 384 6254 428 6296
rect 478 6316 520 6354
rect 478 6296 492 6316
rect 512 6296 520 6316
rect 478 6254 520 6296
rect 602 6316 646 6354
rect 602 6296 614 6316
rect 634 6296 646 6316
rect 602 6254 646 6296
rect 696 6316 738 6354
rect 696 6296 710 6316
rect 730 6296 738 6316
rect 696 6254 738 6296
rect 812 6316 854 6354
rect 812 6296 820 6316
rect 840 6296 854 6316
rect 812 6254 854 6296
rect 904 6323 949 6354
rect 904 6316 948 6323
rect 904 6296 916 6316
rect 936 6296 948 6316
rect 904 6254 948 6296
rect 4748 6329 4792 6367
rect 4748 6309 4760 6329
rect 4780 6309 4792 6329
rect 2640 6252 2684 6294
rect 2640 6232 2652 6252
rect 2672 6232 2684 6252
rect 2640 6225 2684 6232
rect 2639 6194 2684 6225
rect 2734 6252 2776 6294
rect 2734 6232 2748 6252
rect 2768 6232 2776 6252
rect 2734 6194 2776 6232
rect 2850 6252 2892 6294
rect 2850 6232 2858 6252
rect 2878 6232 2892 6252
rect 2850 6194 2892 6232
rect 2942 6252 2986 6294
rect 2942 6232 2954 6252
rect 2974 6232 2986 6252
rect 2942 6194 2986 6232
rect 3068 6252 3110 6294
rect 3068 6232 3076 6252
rect 3096 6232 3110 6252
rect 3068 6194 3110 6232
rect 3160 6252 3204 6294
rect 4748 6267 4792 6309
rect 4842 6329 4884 6367
rect 4842 6309 4856 6329
rect 4876 6309 4884 6329
rect 4842 6267 4884 6309
rect 4966 6329 5010 6367
rect 4966 6309 4978 6329
rect 4998 6309 5010 6329
rect 4966 6267 5010 6309
rect 5060 6329 5102 6367
rect 5060 6309 5074 6329
rect 5094 6309 5102 6329
rect 5060 6267 5102 6309
rect 5176 6329 5218 6367
rect 5176 6309 5184 6329
rect 5204 6309 5218 6329
rect 5176 6267 5218 6309
rect 5268 6336 5313 6367
rect 5268 6329 5312 6336
rect 5268 6309 5280 6329
rect 5300 6309 5312 6329
rect 5268 6267 5312 6309
rect 3160 6232 3172 6252
rect 3192 6232 3204 6252
rect 3160 6194 3204 6232
rect 1182 6132 1226 6170
rect 1182 6112 1194 6132
rect 1214 6112 1226 6132
rect 1182 6070 1226 6112
rect 1276 6132 1318 6170
rect 1276 6112 1290 6132
rect 1310 6112 1318 6132
rect 1276 6070 1318 6112
rect 1400 6132 1444 6170
rect 1400 6112 1412 6132
rect 1432 6112 1444 6132
rect 1400 6070 1444 6112
rect 1494 6132 1536 6170
rect 1494 6112 1508 6132
rect 1528 6112 1536 6132
rect 1494 6070 1536 6112
rect 1610 6132 1652 6170
rect 1610 6112 1618 6132
rect 1638 6112 1652 6132
rect 1610 6070 1652 6112
rect 1702 6139 1747 6170
rect 1702 6132 1746 6139
rect 1702 6112 1714 6132
rect 1734 6112 1746 6132
rect 1702 6070 1746 6112
rect 7004 6265 7048 6307
rect 7004 6245 7016 6265
rect 7036 6245 7048 6265
rect 7004 6238 7048 6245
rect 7003 6207 7048 6238
rect 7098 6265 7140 6307
rect 7098 6245 7112 6265
rect 7132 6245 7140 6265
rect 7098 6207 7140 6245
rect 7214 6265 7256 6307
rect 7214 6245 7222 6265
rect 7242 6245 7256 6265
rect 7214 6207 7256 6245
rect 7306 6265 7350 6307
rect 7306 6245 7318 6265
rect 7338 6245 7350 6265
rect 7306 6207 7350 6245
rect 7432 6265 7474 6307
rect 7432 6245 7440 6265
rect 7460 6245 7474 6265
rect 7432 6207 7474 6245
rect 7524 6265 7568 6307
rect 7524 6245 7536 6265
rect 7556 6245 7568 6265
rect 7524 6207 7568 6245
rect 5546 6145 5590 6183
rect 5546 6125 5558 6145
rect 5578 6125 5590 6145
rect 3438 6068 3482 6110
rect 3438 6048 3450 6068
rect 3470 6048 3482 6068
rect 3438 6041 3482 6048
rect 3437 6010 3482 6041
rect 3532 6068 3574 6110
rect 3532 6048 3546 6068
rect 3566 6048 3574 6068
rect 3532 6010 3574 6048
rect 3648 6068 3690 6110
rect 3648 6048 3656 6068
rect 3676 6048 3690 6068
rect 3648 6010 3690 6048
rect 3740 6068 3784 6110
rect 3740 6048 3752 6068
rect 3772 6048 3784 6068
rect 3740 6010 3784 6048
rect 3866 6068 3908 6110
rect 3866 6048 3874 6068
rect 3894 6048 3908 6068
rect 3866 6010 3908 6048
rect 3958 6068 4002 6110
rect 5546 6083 5590 6125
rect 5640 6145 5682 6183
rect 5640 6125 5654 6145
rect 5674 6125 5682 6145
rect 5640 6083 5682 6125
rect 5764 6145 5808 6183
rect 5764 6125 5776 6145
rect 5796 6125 5808 6145
rect 5764 6083 5808 6125
rect 5858 6145 5900 6183
rect 5858 6125 5872 6145
rect 5892 6125 5900 6145
rect 5858 6083 5900 6125
rect 5974 6145 6016 6183
rect 5974 6125 5982 6145
rect 6002 6125 6016 6145
rect 5974 6083 6016 6125
rect 6066 6152 6111 6183
rect 6066 6145 6110 6152
rect 6066 6125 6078 6145
rect 6098 6125 6110 6145
rect 6066 6083 6110 6125
rect 3958 6048 3970 6068
rect 3990 6048 4002 6068
rect 3958 6010 4002 6048
rect 7802 6081 7846 6123
rect 7802 6061 7814 6081
rect 7834 6061 7846 6081
rect 7802 6054 7846 6061
rect 7801 6023 7846 6054
rect 7896 6081 7938 6123
rect 7896 6061 7910 6081
rect 7930 6061 7938 6081
rect 7896 6023 7938 6061
rect 8012 6081 8054 6123
rect 8012 6061 8020 6081
rect 8040 6061 8054 6081
rect 8012 6023 8054 6061
rect 8104 6081 8148 6123
rect 8104 6061 8116 6081
rect 8136 6061 8148 6081
rect 8104 6023 8148 6061
rect 8230 6081 8272 6123
rect 8230 6061 8238 6081
rect 8258 6061 8272 6081
rect 8230 6023 8272 6061
rect 8322 6081 8366 6123
rect 8322 6061 8334 6081
rect 8354 6061 8366 6081
rect 8322 6023 8366 6061
rect 385 5904 429 5942
rect 385 5884 397 5904
rect 417 5884 429 5904
rect 385 5842 429 5884
rect 479 5904 521 5942
rect 479 5884 493 5904
rect 513 5884 521 5904
rect 479 5842 521 5884
rect 603 5904 647 5942
rect 603 5884 615 5904
rect 635 5884 647 5904
rect 603 5842 647 5884
rect 697 5904 739 5942
rect 697 5884 711 5904
rect 731 5884 739 5904
rect 697 5842 739 5884
rect 813 5904 855 5942
rect 813 5884 821 5904
rect 841 5884 855 5904
rect 813 5842 855 5884
rect 905 5911 950 5942
rect 905 5904 949 5911
rect 905 5884 917 5904
rect 937 5884 949 5904
rect 4749 5917 4793 5955
rect 905 5842 949 5884
rect 2541 5842 2585 5884
rect 2541 5822 2553 5842
rect 2573 5822 2585 5842
rect 2541 5815 2585 5822
rect 2540 5784 2585 5815
rect 2635 5842 2677 5884
rect 2635 5822 2649 5842
rect 2669 5822 2677 5842
rect 2635 5784 2677 5822
rect 2751 5842 2793 5884
rect 2751 5822 2759 5842
rect 2779 5822 2793 5842
rect 2751 5784 2793 5822
rect 2843 5842 2887 5884
rect 2843 5822 2855 5842
rect 2875 5822 2887 5842
rect 2843 5784 2887 5822
rect 2969 5842 3011 5884
rect 2969 5822 2977 5842
rect 2997 5822 3011 5842
rect 2969 5784 3011 5822
rect 3061 5842 3105 5884
rect 4749 5897 4761 5917
rect 4781 5897 4793 5917
rect 3061 5822 3073 5842
rect 3093 5822 3105 5842
rect 4749 5855 4793 5897
rect 4843 5917 4885 5955
rect 4843 5897 4857 5917
rect 4877 5897 4885 5917
rect 4843 5855 4885 5897
rect 4967 5917 5011 5955
rect 4967 5897 4979 5917
rect 4999 5897 5011 5917
rect 4967 5855 5011 5897
rect 5061 5917 5103 5955
rect 5061 5897 5075 5917
rect 5095 5897 5103 5917
rect 5061 5855 5103 5897
rect 5177 5917 5219 5955
rect 5177 5897 5185 5917
rect 5205 5897 5219 5917
rect 5177 5855 5219 5897
rect 5269 5924 5314 5955
rect 5269 5917 5313 5924
rect 5269 5897 5281 5917
rect 5301 5897 5313 5917
rect 5269 5855 5313 5897
rect 6905 5855 6949 5897
rect 3061 5784 3105 5822
rect 6905 5835 6917 5855
rect 6937 5835 6949 5855
rect 6905 5828 6949 5835
rect 6904 5797 6949 5828
rect 6999 5855 7041 5897
rect 6999 5835 7013 5855
rect 7033 5835 7041 5855
rect 6999 5797 7041 5835
rect 7115 5855 7157 5897
rect 7115 5835 7123 5855
rect 7143 5835 7157 5855
rect 7115 5797 7157 5835
rect 7207 5855 7251 5897
rect 7207 5835 7219 5855
rect 7239 5835 7251 5855
rect 7207 5797 7251 5835
rect 7333 5855 7375 5897
rect 7333 5835 7341 5855
rect 7361 5835 7375 5855
rect 7333 5797 7375 5835
rect 7425 5855 7469 5897
rect 7425 5835 7437 5855
rect 7457 5835 7469 5855
rect 7425 5797 7469 5835
rect 1264 5524 1308 5562
rect 1264 5504 1276 5524
rect 1296 5504 1308 5524
rect 1264 5462 1308 5504
rect 1358 5524 1400 5562
rect 1358 5504 1372 5524
rect 1392 5504 1400 5524
rect 1358 5462 1400 5504
rect 1482 5524 1526 5562
rect 1482 5504 1494 5524
rect 1514 5504 1526 5524
rect 1482 5462 1526 5504
rect 1576 5524 1618 5562
rect 1576 5504 1590 5524
rect 1610 5504 1618 5524
rect 1576 5462 1618 5504
rect 1692 5524 1734 5562
rect 1692 5504 1700 5524
rect 1720 5504 1734 5524
rect 1692 5462 1734 5504
rect 1784 5531 1829 5562
rect 1784 5524 1828 5531
rect 1784 5504 1796 5524
rect 1816 5504 1828 5524
rect 5628 5537 5672 5575
rect 1784 5462 1828 5504
rect 3420 5462 3464 5504
rect 3420 5442 3432 5462
rect 3452 5442 3464 5462
rect 3420 5435 3464 5442
rect 3419 5404 3464 5435
rect 3514 5462 3556 5504
rect 3514 5442 3528 5462
rect 3548 5442 3556 5462
rect 3514 5404 3556 5442
rect 3630 5462 3672 5504
rect 3630 5442 3638 5462
rect 3658 5442 3672 5462
rect 3630 5404 3672 5442
rect 3722 5462 3766 5504
rect 3722 5442 3734 5462
rect 3754 5442 3766 5462
rect 3722 5404 3766 5442
rect 3848 5462 3890 5504
rect 3848 5442 3856 5462
rect 3876 5442 3890 5462
rect 3848 5404 3890 5442
rect 3940 5462 3984 5504
rect 5628 5517 5640 5537
rect 5660 5517 5672 5537
rect 3940 5442 3952 5462
rect 3972 5442 3984 5462
rect 5628 5475 5672 5517
rect 5722 5537 5764 5575
rect 5722 5517 5736 5537
rect 5756 5517 5764 5537
rect 5722 5475 5764 5517
rect 5846 5537 5890 5575
rect 5846 5517 5858 5537
rect 5878 5517 5890 5537
rect 5846 5475 5890 5517
rect 5940 5537 5982 5575
rect 5940 5517 5954 5537
rect 5974 5517 5982 5537
rect 5940 5475 5982 5517
rect 6056 5537 6098 5575
rect 6056 5517 6064 5537
rect 6084 5517 6098 5537
rect 6056 5475 6098 5517
rect 6148 5544 6193 5575
rect 6148 5537 6192 5544
rect 6148 5517 6160 5537
rect 6180 5517 6192 5537
rect 6148 5475 6192 5517
rect 7784 5475 7828 5517
rect 3940 5404 3984 5442
rect 7784 5455 7796 5475
rect 7816 5455 7828 5475
rect 7784 5448 7828 5455
rect 7783 5417 7828 5448
rect 7878 5475 7920 5517
rect 7878 5455 7892 5475
rect 7912 5455 7920 5475
rect 7878 5417 7920 5455
rect 7994 5475 8036 5517
rect 7994 5455 8002 5475
rect 8022 5455 8036 5475
rect 7994 5417 8036 5455
rect 8086 5475 8130 5517
rect 8086 5455 8098 5475
rect 8118 5455 8130 5475
rect 8086 5417 8130 5455
rect 8212 5475 8254 5517
rect 8212 5455 8220 5475
rect 8240 5455 8254 5475
rect 8212 5417 8254 5455
rect 8304 5475 8348 5517
rect 8304 5455 8316 5475
rect 8336 5455 8348 5475
rect 8304 5417 8348 5455
rect 367 5298 411 5336
rect 367 5278 379 5298
rect 399 5278 411 5298
rect 367 5236 411 5278
rect 461 5298 503 5336
rect 461 5278 475 5298
rect 495 5278 503 5298
rect 461 5236 503 5278
rect 585 5298 629 5336
rect 585 5278 597 5298
rect 617 5278 629 5298
rect 585 5236 629 5278
rect 679 5298 721 5336
rect 679 5278 693 5298
rect 713 5278 721 5298
rect 679 5236 721 5278
rect 795 5298 837 5336
rect 795 5278 803 5298
rect 823 5278 837 5298
rect 795 5236 837 5278
rect 887 5305 932 5336
rect 887 5298 931 5305
rect 887 5278 899 5298
rect 919 5278 931 5298
rect 887 5236 931 5278
rect 4731 5311 4775 5349
rect 4731 5291 4743 5311
rect 4763 5291 4775 5311
rect 2623 5234 2667 5276
rect 2623 5214 2635 5234
rect 2655 5214 2667 5234
rect 2623 5207 2667 5214
rect 2622 5176 2667 5207
rect 2717 5234 2759 5276
rect 2717 5214 2731 5234
rect 2751 5214 2759 5234
rect 2717 5176 2759 5214
rect 2833 5234 2875 5276
rect 2833 5214 2841 5234
rect 2861 5214 2875 5234
rect 2833 5176 2875 5214
rect 2925 5234 2969 5276
rect 2925 5214 2937 5234
rect 2957 5214 2969 5234
rect 2925 5176 2969 5214
rect 3051 5234 3093 5276
rect 3051 5214 3059 5234
rect 3079 5214 3093 5234
rect 3051 5176 3093 5214
rect 3143 5234 3187 5276
rect 4731 5249 4775 5291
rect 4825 5311 4867 5349
rect 4825 5291 4839 5311
rect 4859 5291 4867 5311
rect 4825 5249 4867 5291
rect 4949 5311 4993 5349
rect 4949 5291 4961 5311
rect 4981 5291 4993 5311
rect 4949 5249 4993 5291
rect 5043 5311 5085 5349
rect 5043 5291 5057 5311
rect 5077 5291 5085 5311
rect 5043 5249 5085 5291
rect 5159 5311 5201 5349
rect 5159 5291 5167 5311
rect 5187 5291 5201 5311
rect 5159 5249 5201 5291
rect 5251 5318 5296 5349
rect 5251 5311 5295 5318
rect 5251 5291 5263 5311
rect 5283 5291 5295 5311
rect 5251 5249 5295 5291
rect 3143 5214 3155 5234
rect 3175 5214 3187 5234
rect 3143 5176 3187 5214
rect 1165 5114 1209 5152
rect 1165 5094 1177 5114
rect 1197 5094 1209 5114
rect 1165 5052 1209 5094
rect 1259 5114 1301 5152
rect 1259 5094 1273 5114
rect 1293 5094 1301 5114
rect 1259 5052 1301 5094
rect 1383 5114 1427 5152
rect 1383 5094 1395 5114
rect 1415 5094 1427 5114
rect 1383 5052 1427 5094
rect 1477 5114 1519 5152
rect 1477 5094 1491 5114
rect 1511 5094 1519 5114
rect 1477 5052 1519 5094
rect 1593 5114 1635 5152
rect 1593 5094 1601 5114
rect 1621 5094 1635 5114
rect 1593 5052 1635 5094
rect 1685 5121 1730 5152
rect 1685 5114 1729 5121
rect 1685 5094 1697 5114
rect 1717 5094 1729 5114
rect 1685 5052 1729 5094
rect 6987 5247 7031 5289
rect 6987 5227 6999 5247
rect 7019 5227 7031 5247
rect 6987 5220 7031 5227
rect 6986 5189 7031 5220
rect 7081 5247 7123 5289
rect 7081 5227 7095 5247
rect 7115 5227 7123 5247
rect 7081 5189 7123 5227
rect 7197 5247 7239 5289
rect 7197 5227 7205 5247
rect 7225 5227 7239 5247
rect 7197 5189 7239 5227
rect 7289 5247 7333 5289
rect 7289 5227 7301 5247
rect 7321 5227 7333 5247
rect 7289 5189 7333 5227
rect 7415 5247 7457 5289
rect 7415 5227 7423 5247
rect 7443 5227 7457 5247
rect 7415 5189 7457 5227
rect 7507 5247 7551 5289
rect 7507 5227 7519 5247
rect 7539 5227 7551 5247
rect 7507 5189 7551 5227
rect 5529 5127 5573 5165
rect 5529 5107 5541 5127
rect 5561 5107 5573 5127
rect 3421 5050 3465 5092
rect 3421 5030 3433 5050
rect 3453 5030 3465 5050
rect 3421 5023 3465 5030
rect 3420 4992 3465 5023
rect 3515 5050 3557 5092
rect 3515 5030 3529 5050
rect 3549 5030 3557 5050
rect 3515 4992 3557 5030
rect 3631 5050 3673 5092
rect 3631 5030 3639 5050
rect 3659 5030 3673 5050
rect 3631 4992 3673 5030
rect 3723 5050 3767 5092
rect 3723 5030 3735 5050
rect 3755 5030 3767 5050
rect 3723 4992 3767 5030
rect 3849 5050 3891 5092
rect 3849 5030 3857 5050
rect 3877 5030 3891 5050
rect 3849 4992 3891 5030
rect 3941 5050 3985 5092
rect 5529 5065 5573 5107
rect 5623 5127 5665 5165
rect 5623 5107 5637 5127
rect 5657 5107 5665 5127
rect 5623 5065 5665 5107
rect 5747 5127 5791 5165
rect 5747 5107 5759 5127
rect 5779 5107 5791 5127
rect 5747 5065 5791 5107
rect 5841 5127 5883 5165
rect 5841 5107 5855 5127
rect 5875 5107 5883 5127
rect 5841 5065 5883 5107
rect 5957 5127 5999 5165
rect 5957 5107 5965 5127
rect 5985 5107 5999 5127
rect 5957 5065 5999 5107
rect 6049 5134 6094 5165
rect 6049 5127 6093 5134
rect 6049 5107 6061 5127
rect 6081 5107 6093 5127
rect 6049 5065 6093 5107
rect 3941 5030 3953 5050
rect 3973 5030 3985 5050
rect 3941 4992 3985 5030
rect 7785 5063 7829 5105
rect 7785 5043 7797 5063
rect 7817 5043 7829 5063
rect 7785 5036 7829 5043
rect 7784 5005 7829 5036
rect 7879 5063 7921 5105
rect 7879 5043 7893 5063
rect 7913 5043 7921 5063
rect 7879 5005 7921 5043
rect 7995 5063 8037 5105
rect 7995 5043 8003 5063
rect 8023 5043 8037 5063
rect 7995 5005 8037 5043
rect 8087 5063 8131 5105
rect 8087 5043 8099 5063
rect 8119 5043 8131 5063
rect 8087 5005 8131 5043
rect 8213 5063 8255 5105
rect 8213 5043 8221 5063
rect 8241 5043 8255 5063
rect 8213 5005 8255 5043
rect 8305 5063 8349 5105
rect 8305 5043 8317 5063
rect 8337 5043 8349 5063
rect 8305 5005 8349 5043
rect 368 4886 412 4924
rect 368 4866 380 4886
rect 400 4866 412 4886
rect 368 4824 412 4866
rect 462 4886 504 4924
rect 462 4866 476 4886
rect 496 4866 504 4886
rect 462 4824 504 4866
rect 586 4886 630 4924
rect 586 4866 598 4886
rect 618 4866 630 4886
rect 586 4824 630 4866
rect 680 4886 722 4924
rect 680 4866 694 4886
rect 714 4866 722 4886
rect 680 4824 722 4866
rect 796 4886 838 4924
rect 796 4866 804 4886
rect 824 4866 838 4886
rect 796 4824 838 4866
rect 888 4893 933 4924
rect 888 4886 932 4893
rect 888 4866 900 4886
rect 920 4866 932 4886
rect 4732 4899 4776 4937
rect 888 4824 932 4866
rect 2319 4828 2363 4870
rect 2319 4808 2331 4828
rect 2351 4808 2363 4828
rect 2319 4801 2363 4808
rect 2318 4770 2363 4801
rect 2413 4828 2455 4870
rect 2413 4808 2427 4828
rect 2447 4808 2455 4828
rect 2413 4770 2455 4808
rect 2529 4828 2571 4870
rect 2529 4808 2537 4828
rect 2557 4808 2571 4828
rect 2529 4770 2571 4808
rect 2621 4828 2665 4870
rect 2621 4808 2633 4828
rect 2653 4808 2665 4828
rect 2621 4770 2665 4808
rect 2747 4828 2789 4870
rect 2747 4808 2755 4828
rect 2775 4808 2789 4828
rect 2747 4770 2789 4808
rect 2839 4828 2883 4870
rect 4732 4879 4744 4899
rect 4764 4879 4776 4899
rect 2839 4808 2851 4828
rect 2871 4808 2883 4828
rect 4732 4837 4776 4879
rect 4826 4899 4868 4937
rect 4826 4879 4840 4899
rect 4860 4879 4868 4899
rect 4826 4837 4868 4879
rect 4950 4899 4994 4937
rect 4950 4879 4962 4899
rect 4982 4879 4994 4899
rect 4950 4837 4994 4879
rect 5044 4899 5086 4937
rect 5044 4879 5058 4899
rect 5078 4879 5086 4899
rect 5044 4837 5086 4879
rect 5160 4899 5202 4937
rect 5160 4879 5168 4899
rect 5188 4879 5202 4899
rect 5160 4837 5202 4879
rect 5252 4906 5297 4937
rect 5252 4899 5296 4906
rect 5252 4879 5264 4899
rect 5284 4879 5296 4899
rect 5252 4837 5296 4879
rect 6683 4841 6727 4883
rect 2839 4770 2883 4808
rect 6683 4821 6695 4841
rect 6715 4821 6727 4841
rect 6683 4814 6727 4821
rect 6682 4783 6727 4814
rect 6777 4841 6819 4883
rect 6777 4821 6791 4841
rect 6811 4821 6819 4841
rect 6777 4783 6819 4821
rect 6893 4841 6935 4883
rect 6893 4821 6901 4841
rect 6921 4821 6935 4841
rect 6893 4783 6935 4821
rect 6985 4841 7029 4883
rect 6985 4821 6997 4841
rect 7017 4821 7029 4841
rect 6985 4783 7029 4821
rect 7111 4841 7153 4883
rect 7111 4821 7119 4841
rect 7139 4821 7153 4841
rect 7111 4783 7153 4821
rect 7203 4841 7247 4883
rect 7203 4821 7215 4841
rect 7235 4821 7247 4841
rect 7203 4783 7247 4821
rect 1450 4502 1494 4540
rect 1450 4482 1462 4502
rect 1482 4482 1494 4502
rect 1450 4440 1494 4482
rect 1544 4502 1586 4540
rect 1544 4482 1558 4502
rect 1578 4482 1586 4502
rect 1544 4440 1586 4482
rect 1668 4502 1712 4540
rect 1668 4482 1680 4502
rect 1700 4482 1712 4502
rect 1668 4440 1712 4482
rect 1762 4502 1804 4540
rect 1762 4482 1776 4502
rect 1796 4482 1804 4502
rect 1762 4440 1804 4482
rect 1878 4502 1920 4540
rect 1878 4482 1886 4502
rect 1906 4482 1920 4502
rect 1878 4440 1920 4482
rect 1970 4509 2015 4540
rect 1970 4502 2014 4509
rect 1970 4482 1982 4502
rect 2002 4482 2014 4502
rect 5814 4515 5858 4553
rect 1970 4440 2014 4482
rect 3401 4444 3445 4486
rect 3401 4424 3413 4444
rect 3433 4424 3445 4444
rect 3401 4417 3445 4424
rect 3400 4386 3445 4417
rect 3495 4444 3537 4486
rect 3495 4424 3509 4444
rect 3529 4424 3537 4444
rect 3495 4386 3537 4424
rect 3611 4444 3653 4486
rect 3611 4424 3619 4444
rect 3639 4424 3653 4444
rect 3611 4386 3653 4424
rect 3703 4444 3747 4486
rect 3703 4424 3715 4444
rect 3735 4424 3747 4444
rect 3703 4386 3747 4424
rect 3829 4444 3871 4486
rect 3829 4424 3837 4444
rect 3857 4424 3871 4444
rect 3829 4386 3871 4424
rect 3921 4444 3965 4486
rect 5814 4495 5826 4515
rect 5846 4495 5858 4515
rect 3921 4424 3933 4444
rect 3953 4424 3965 4444
rect 5814 4453 5858 4495
rect 5908 4515 5950 4553
rect 5908 4495 5922 4515
rect 5942 4495 5950 4515
rect 5908 4453 5950 4495
rect 6032 4515 6076 4553
rect 6032 4495 6044 4515
rect 6064 4495 6076 4515
rect 6032 4453 6076 4495
rect 6126 4515 6168 4553
rect 6126 4495 6140 4515
rect 6160 4495 6168 4515
rect 6126 4453 6168 4495
rect 6242 4515 6284 4553
rect 6242 4495 6250 4515
rect 6270 4495 6284 4515
rect 6242 4453 6284 4495
rect 6334 4522 6379 4553
rect 6334 4515 6378 4522
rect 6334 4495 6346 4515
rect 6366 4495 6378 4515
rect 6334 4453 6378 4495
rect 7765 4457 7809 4499
rect 3921 4386 3965 4424
rect 7765 4437 7777 4457
rect 7797 4437 7809 4457
rect 7765 4430 7809 4437
rect 7764 4399 7809 4430
rect 7859 4457 7901 4499
rect 7859 4437 7873 4457
rect 7893 4437 7901 4457
rect 7859 4399 7901 4437
rect 7975 4457 8017 4499
rect 7975 4437 7983 4457
rect 8003 4437 8017 4457
rect 7975 4399 8017 4437
rect 8067 4457 8111 4499
rect 8067 4437 8079 4457
rect 8099 4437 8111 4457
rect 8067 4399 8111 4437
rect 8193 4457 8235 4499
rect 8193 4437 8201 4457
rect 8221 4437 8235 4457
rect 8193 4399 8235 4437
rect 8285 4457 8329 4499
rect 8285 4437 8297 4457
rect 8317 4437 8329 4457
rect 8285 4399 8329 4437
rect 348 4280 392 4318
rect 348 4260 360 4280
rect 380 4260 392 4280
rect 348 4218 392 4260
rect 442 4280 484 4318
rect 442 4260 456 4280
rect 476 4260 484 4280
rect 442 4218 484 4260
rect 566 4280 610 4318
rect 566 4260 578 4280
rect 598 4260 610 4280
rect 566 4218 610 4260
rect 660 4280 702 4318
rect 660 4260 674 4280
rect 694 4260 702 4280
rect 660 4218 702 4260
rect 776 4280 818 4318
rect 776 4260 784 4280
rect 804 4260 818 4280
rect 776 4218 818 4260
rect 868 4287 913 4318
rect 868 4280 912 4287
rect 868 4260 880 4280
rect 900 4260 912 4280
rect 868 4218 912 4260
rect 4712 4293 4756 4331
rect 4712 4273 4724 4293
rect 4744 4273 4756 4293
rect 2604 4216 2648 4258
rect 2604 4196 2616 4216
rect 2636 4196 2648 4216
rect 2604 4189 2648 4196
rect 2603 4158 2648 4189
rect 2698 4216 2740 4258
rect 2698 4196 2712 4216
rect 2732 4196 2740 4216
rect 2698 4158 2740 4196
rect 2814 4216 2856 4258
rect 2814 4196 2822 4216
rect 2842 4196 2856 4216
rect 2814 4158 2856 4196
rect 2906 4216 2950 4258
rect 2906 4196 2918 4216
rect 2938 4196 2950 4216
rect 2906 4158 2950 4196
rect 3032 4216 3074 4258
rect 3032 4196 3040 4216
rect 3060 4196 3074 4216
rect 3032 4158 3074 4196
rect 3124 4216 3168 4258
rect 4712 4231 4756 4273
rect 4806 4293 4848 4331
rect 4806 4273 4820 4293
rect 4840 4273 4848 4293
rect 4806 4231 4848 4273
rect 4930 4293 4974 4331
rect 4930 4273 4942 4293
rect 4962 4273 4974 4293
rect 4930 4231 4974 4273
rect 5024 4293 5066 4331
rect 5024 4273 5038 4293
rect 5058 4273 5066 4293
rect 5024 4231 5066 4273
rect 5140 4293 5182 4331
rect 5140 4273 5148 4293
rect 5168 4273 5182 4293
rect 5140 4231 5182 4273
rect 5232 4300 5277 4331
rect 5232 4293 5276 4300
rect 5232 4273 5244 4293
rect 5264 4273 5276 4293
rect 5232 4231 5276 4273
rect 3124 4196 3136 4216
rect 3156 4196 3168 4216
rect 3124 4158 3168 4196
rect 1146 4096 1190 4134
rect 1146 4076 1158 4096
rect 1178 4076 1190 4096
rect 1146 4034 1190 4076
rect 1240 4096 1282 4134
rect 1240 4076 1254 4096
rect 1274 4076 1282 4096
rect 1240 4034 1282 4076
rect 1364 4096 1408 4134
rect 1364 4076 1376 4096
rect 1396 4076 1408 4096
rect 1364 4034 1408 4076
rect 1458 4096 1500 4134
rect 1458 4076 1472 4096
rect 1492 4076 1500 4096
rect 1458 4034 1500 4076
rect 1574 4096 1616 4134
rect 1574 4076 1582 4096
rect 1602 4076 1616 4096
rect 1574 4034 1616 4076
rect 1666 4103 1711 4134
rect 1666 4096 1710 4103
rect 1666 4076 1678 4096
rect 1698 4076 1710 4096
rect 1666 4034 1710 4076
rect 6968 4229 7012 4271
rect 6968 4209 6980 4229
rect 7000 4209 7012 4229
rect 6968 4202 7012 4209
rect 6967 4171 7012 4202
rect 7062 4229 7104 4271
rect 7062 4209 7076 4229
rect 7096 4209 7104 4229
rect 7062 4171 7104 4209
rect 7178 4229 7220 4271
rect 7178 4209 7186 4229
rect 7206 4209 7220 4229
rect 7178 4171 7220 4209
rect 7270 4229 7314 4271
rect 7270 4209 7282 4229
rect 7302 4209 7314 4229
rect 7270 4171 7314 4209
rect 7396 4229 7438 4271
rect 7396 4209 7404 4229
rect 7424 4209 7438 4229
rect 7396 4171 7438 4209
rect 7488 4229 7532 4271
rect 7488 4209 7500 4229
rect 7520 4209 7532 4229
rect 7488 4171 7532 4209
rect 5510 4109 5554 4147
rect 5510 4089 5522 4109
rect 5542 4089 5554 4109
rect 3402 4032 3446 4074
rect 3402 4012 3414 4032
rect 3434 4012 3446 4032
rect 3402 4005 3446 4012
rect 3401 3974 3446 4005
rect 3496 4032 3538 4074
rect 3496 4012 3510 4032
rect 3530 4012 3538 4032
rect 3496 3974 3538 4012
rect 3612 4032 3654 4074
rect 3612 4012 3620 4032
rect 3640 4012 3654 4032
rect 3612 3974 3654 4012
rect 3704 4032 3748 4074
rect 3704 4012 3716 4032
rect 3736 4012 3748 4032
rect 3704 3974 3748 4012
rect 3830 4032 3872 4074
rect 3830 4012 3838 4032
rect 3858 4012 3872 4032
rect 3830 3974 3872 4012
rect 3922 4032 3966 4074
rect 5510 4047 5554 4089
rect 5604 4109 5646 4147
rect 5604 4089 5618 4109
rect 5638 4089 5646 4109
rect 5604 4047 5646 4089
rect 5728 4109 5772 4147
rect 5728 4089 5740 4109
rect 5760 4089 5772 4109
rect 5728 4047 5772 4089
rect 5822 4109 5864 4147
rect 5822 4089 5836 4109
rect 5856 4089 5864 4109
rect 5822 4047 5864 4089
rect 5938 4109 5980 4147
rect 5938 4089 5946 4109
rect 5966 4089 5980 4109
rect 5938 4047 5980 4089
rect 6030 4116 6075 4147
rect 6030 4109 6074 4116
rect 6030 4089 6042 4109
rect 6062 4089 6074 4109
rect 6030 4047 6074 4089
rect 3922 4012 3934 4032
rect 3954 4012 3966 4032
rect 3922 3974 3966 4012
rect 7766 4045 7810 4087
rect 7766 4025 7778 4045
rect 7798 4025 7810 4045
rect 7766 4018 7810 4025
rect 7765 3987 7810 4018
rect 7860 4045 7902 4087
rect 7860 4025 7874 4045
rect 7894 4025 7902 4045
rect 7860 3987 7902 4025
rect 7976 4045 8018 4087
rect 7976 4025 7984 4045
rect 8004 4025 8018 4045
rect 7976 3987 8018 4025
rect 8068 4045 8112 4087
rect 8068 4025 8080 4045
rect 8100 4025 8112 4045
rect 8068 3987 8112 4025
rect 8194 4045 8236 4087
rect 8194 4025 8202 4045
rect 8222 4025 8236 4045
rect 8194 3987 8236 4025
rect 8286 4045 8330 4087
rect 8286 4025 8298 4045
rect 8318 4025 8330 4045
rect 8286 3987 8330 4025
rect 349 3868 393 3906
rect 349 3848 361 3868
rect 381 3848 393 3868
rect 349 3806 393 3848
rect 443 3868 485 3906
rect 443 3848 457 3868
rect 477 3848 485 3868
rect 443 3806 485 3848
rect 567 3868 611 3906
rect 567 3848 579 3868
rect 599 3848 611 3868
rect 567 3806 611 3848
rect 661 3868 703 3906
rect 661 3848 675 3868
rect 695 3848 703 3868
rect 661 3806 703 3848
rect 777 3868 819 3906
rect 777 3848 785 3868
rect 805 3848 819 3868
rect 777 3806 819 3848
rect 869 3875 914 3906
rect 869 3868 913 3875
rect 869 3848 881 3868
rect 901 3848 913 3868
rect 4713 3881 4757 3919
rect 869 3806 913 3848
rect 2505 3806 2549 3848
rect 2505 3786 2517 3806
rect 2537 3786 2549 3806
rect 2505 3779 2549 3786
rect 2504 3748 2549 3779
rect 2599 3806 2641 3848
rect 2599 3786 2613 3806
rect 2633 3786 2641 3806
rect 2599 3748 2641 3786
rect 2715 3806 2757 3848
rect 2715 3786 2723 3806
rect 2743 3786 2757 3806
rect 2715 3748 2757 3786
rect 2807 3806 2851 3848
rect 2807 3786 2819 3806
rect 2839 3786 2851 3806
rect 2807 3748 2851 3786
rect 2933 3806 2975 3848
rect 2933 3786 2941 3806
rect 2961 3786 2975 3806
rect 2933 3748 2975 3786
rect 3025 3806 3069 3848
rect 4713 3861 4725 3881
rect 4745 3861 4757 3881
rect 3025 3786 3037 3806
rect 3057 3786 3069 3806
rect 4713 3819 4757 3861
rect 4807 3881 4849 3919
rect 4807 3861 4821 3881
rect 4841 3861 4849 3881
rect 4807 3819 4849 3861
rect 4931 3881 4975 3919
rect 4931 3861 4943 3881
rect 4963 3861 4975 3881
rect 4931 3819 4975 3861
rect 5025 3881 5067 3919
rect 5025 3861 5039 3881
rect 5059 3861 5067 3881
rect 5025 3819 5067 3861
rect 5141 3881 5183 3919
rect 5141 3861 5149 3881
rect 5169 3861 5183 3881
rect 5141 3819 5183 3861
rect 5233 3888 5278 3919
rect 5233 3881 5277 3888
rect 5233 3861 5245 3881
rect 5265 3861 5277 3881
rect 5233 3819 5277 3861
rect 6869 3819 6913 3861
rect 3025 3748 3069 3786
rect 6869 3799 6881 3819
rect 6901 3799 6913 3819
rect 6869 3792 6913 3799
rect 6868 3761 6913 3792
rect 6963 3819 7005 3861
rect 6963 3799 6977 3819
rect 6997 3799 7005 3819
rect 6963 3761 7005 3799
rect 7079 3819 7121 3861
rect 7079 3799 7087 3819
rect 7107 3799 7121 3819
rect 7079 3761 7121 3799
rect 7171 3819 7215 3861
rect 7171 3799 7183 3819
rect 7203 3799 7215 3819
rect 7171 3761 7215 3799
rect 7297 3819 7339 3861
rect 7297 3799 7305 3819
rect 7325 3799 7339 3819
rect 7297 3761 7339 3799
rect 7389 3819 7433 3861
rect 7389 3799 7401 3819
rect 7421 3799 7433 3819
rect 7389 3761 7433 3799
rect 1228 3488 1272 3526
rect 1228 3468 1240 3488
rect 1260 3468 1272 3488
rect 1228 3426 1272 3468
rect 1322 3488 1364 3526
rect 1322 3468 1336 3488
rect 1356 3468 1364 3488
rect 1322 3426 1364 3468
rect 1446 3488 1490 3526
rect 1446 3468 1458 3488
rect 1478 3468 1490 3488
rect 1446 3426 1490 3468
rect 1540 3488 1582 3526
rect 1540 3468 1554 3488
rect 1574 3468 1582 3488
rect 1540 3426 1582 3468
rect 1656 3488 1698 3526
rect 1656 3468 1664 3488
rect 1684 3468 1698 3488
rect 1656 3426 1698 3468
rect 1748 3495 1793 3526
rect 1748 3488 1792 3495
rect 1748 3468 1760 3488
rect 1780 3468 1792 3488
rect 5592 3501 5636 3539
rect 1748 3426 1792 3468
rect 3384 3426 3428 3468
rect 3384 3406 3396 3426
rect 3416 3406 3428 3426
rect 3384 3399 3428 3406
rect 3383 3368 3428 3399
rect 3478 3426 3520 3468
rect 3478 3406 3492 3426
rect 3512 3406 3520 3426
rect 3478 3368 3520 3406
rect 3594 3426 3636 3468
rect 3594 3406 3602 3426
rect 3622 3406 3636 3426
rect 3594 3368 3636 3406
rect 3686 3426 3730 3468
rect 3686 3406 3698 3426
rect 3718 3406 3730 3426
rect 3686 3368 3730 3406
rect 3812 3426 3854 3468
rect 3812 3406 3820 3426
rect 3840 3406 3854 3426
rect 3812 3368 3854 3406
rect 3904 3426 3948 3468
rect 5592 3481 5604 3501
rect 5624 3481 5636 3501
rect 3904 3406 3916 3426
rect 3936 3406 3948 3426
rect 5592 3439 5636 3481
rect 5686 3501 5728 3539
rect 5686 3481 5700 3501
rect 5720 3481 5728 3501
rect 5686 3439 5728 3481
rect 5810 3501 5854 3539
rect 5810 3481 5822 3501
rect 5842 3481 5854 3501
rect 5810 3439 5854 3481
rect 5904 3501 5946 3539
rect 5904 3481 5918 3501
rect 5938 3481 5946 3501
rect 5904 3439 5946 3481
rect 6020 3501 6062 3539
rect 6020 3481 6028 3501
rect 6048 3481 6062 3501
rect 6020 3439 6062 3481
rect 6112 3508 6157 3539
rect 6112 3501 6156 3508
rect 6112 3481 6124 3501
rect 6144 3481 6156 3501
rect 6112 3439 6156 3481
rect 7748 3439 7792 3481
rect 3904 3368 3948 3406
rect 7748 3419 7760 3439
rect 7780 3419 7792 3439
rect 7748 3412 7792 3419
rect 7747 3381 7792 3412
rect 7842 3439 7884 3481
rect 7842 3419 7856 3439
rect 7876 3419 7884 3439
rect 7842 3381 7884 3419
rect 7958 3439 8000 3481
rect 7958 3419 7966 3439
rect 7986 3419 8000 3439
rect 7958 3381 8000 3419
rect 8050 3439 8094 3481
rect 8050 3419 8062 3439
rect 8082 3419 8094 3439
rect 8050 3381 8094 3419
rect 8176 3439 8218 3481
rect 8176 3419 8184 3439
rect 8204 3419 8218 3439
rect 8176 3381 8218 3419
rect 8268 3439 8312 3481
rect 8268 3419 8280 3439
rect 8300 3419 8312 3439
rect 8268 3381 8312 3419
rect 331 3262 375 3300
rect 331 3242 343 3262
rect 363 3242 375 3262
rect 331 3200 375 3242
rect 425 3262 467 3300
rect 425 3242 439 3262
rect 459 3242 467 3262
rect 425 3200 467 3242
rect 549 3262 593 3300
rect 549 3242 561 3262
rect 581 3242 593 3262
rect 549 3200 593 3242
rect 643 3262 685 3300
rect 643 3242 657 3262
rect 677 3242 685 3262
rect 643 3200 685 3242
rect 759 3262 801 3300
rect 759 3242 767 3262
rect 787 3242 801 3262
rect 759 3200 801 3242
rect 851 3269 896 3300
rect 851 3262 895 3269
rect 851 3242 863 3262
rect 883 3242 895 3262
rect 851 3200 895 3242
rect 4695 3275 4739 3313
rect 4695 3255 4707 3275
rect 4727 3255 4739 3275
rect 2587 3198 2631 3240
rect 2587 3178 2599 3198
rect 2619 3178 2631 3198
rect 2587 3171 2631 3178
rect 2586 3140 2631 3171
rect 2681 3198 2723 3240
rect 2681 3178 2695 3198
rect 2715 3178 2723 3198
rect 2681 3140 2723 3178
rect 2797 3198 2839 3240
rect 2797 3178 2805 3198
rect 2825 3178 2839 3198
rect 2797 3140 2839 3178
rect 2889 3198 2933 3240
rect 2889 3178 2901 3198
rect 2921 3178 2933 3198
rect 2889 3140 2933 3178
rect 3015 3198 3057 3240
rect 3015 3178 3023 3198
rect 3043 3178 3057 3198
rect 3015 3140 3057 3178
rect 3107 3198 3151 3240
rect 4695 3213 4739 3255
rect 4789 3275 4831 3313
rect 4789 3255 4803 3275
rect 4823 3255 4831 3275
rect 4789 3213 4831 3255
rect 4913 3275 4957 3313
rect 4913 3255 4925 3275
rect 4945 3255 4957 3275
rect 4913 3213 4957 3255
rect 5007 3275 5049 3313
rect 5007 3255 5021 3275
rect 5041 3255 5049 3275
rect 5007 3213 5049 3255
rect 5123 3275 5165 3313
rect 5123 3255 5131 3275
rect 5151 3255 5165 3275
rect 5123 3213 5165 3255
rect 5215 3282 5260 3313
rect 5215 3275 5259 3282
rect 5215 3255 5227 3275
rect 5247 3255 5259 3275
rect 5215 3213 5259 3255
rect 3107 3178 3119 3198
rect 3139 3178 3151 3198
rect 3107 3140 3151 3178
rect 1129 3078 1173 3116
rect 1129 3058 1141 3078
rect 1161 3058 1173 3078
rect 1129 3016 1173 3058
rect 1223 3078 1265 3116
rect 1223 3058 1237 3078
rect 1257 3058 1265 3078
rect 1223 3016 1265 3058
rect 1347 3078 1391 3116
rect 1347 3058 1359 3078
rect 1379 3058 1391 3078
rect 1347 3016 1391 3058
rect 1441 3078 1483 3116
rect 1441 3058 1455 3078
rect 1475 3058 1483 3078
rect 1441 3016 1483 3058
rect 1557 3078 1599 3116
rect 1557 3058 1565 3078
rect 1585 3058 1599 3078
rect 1557 3016 1599 3058
rect 1649 3085 1694 3116
rect 1649 3078 1693 3085
rect 1649 3058 1661 3078
rect 1681 3058 1693 3078
rect 1649 3016 1693 3058
rect 6951 3211 6995 3253
rect 6951 3191 6963 3211
rect 6983 3191 6995 3211
rect 6951 3184 6995 3191
rect 6950 3153 6995 3184
rect 7045 3211 7087 3253
rect 7045 3191 7059 3211
rect 7079 3191 7087 3211
rect 7045 3153 7087 3191
rect 7161 3211 7203 3253
rect 7161 3191 7169 3211
rect 7189 3191 7203 3211
rect 7161 3153 7203 3191
rect 7253 3211 7297 3253
rect 7253 3191 7265 3211
rect 7285 3191 7297 3211
rect 7253 3153 7297 3191
rect 7379 3211 7421 3253
rect 7379 3191 7387 3211
rect 7407 3191 7421 3211
rect 7379 3153 7421 3191
rect 7471 3211 7515 3253
rect 7471 3191 7483 3211
rect 7503 3191 7515 3211
rect 7471 3153 7515 3191
rect 5493 3091 5537 3129
rect 5493 3071 5505 3091
rect 5525 3071 5537 3091
rect 3385 3014 3429 3056
rect 3385 2994 3397 3014
rect 3417 2994 3429 3014
rect 3385 2987 3429 2994
rect 3384 2956 3429 2987
rect 3479 3014 3521 3056
rect 3479 2994 3493 3014
rect 3513 2994 3521 3014
rect 3479 2956 3521 2994
rect 3595 3014 3637 3056
rect 3595 2994 3603 3014
rect 3623 2994 3637 3014
rect 3595 2956 3637 2994
rect 3687 3014 3731 3056
rect 3687 2994 3699 3014
rect 3719 2994 3731 3014
rect 3687 2956 3731 2994
rect 3813 3014 3855 3056
rect 3813 2994 3821 3014
rect 3841 2994 3855 3014
rect 3813 2956 3855 2994
rect 3905 3014 3949 3056
rect 5493 3029 5537 3071
rect 5587 3091 5629 3129
rect 5587 3071 5601 3091
rect 5621 3071 5629 3091
rect 5587 3029 5629 3071
rect 5711 3091 5755 3129
rect 5711 3071 5723 3091
rect 5743 3071 5755 3091
rect 5711 3029 5755 3071
rect 5805 3091 5847 3129
rect 5805 3071 5819 3091
rect 5839 3071 5847 3091
rect 5805 3029 5847 3071
rect 5921 3091 5963 3129
rect 5921 3071 5929 3091
rect 5949 3071 5963 3091
rect 5921 3029 5963 3071
rect 6013 3098 6058 3129
rect 6013 3091 6057 3098
rect 6013 3071 6025 3091
rect 6045 3071 6057 3091
rect 6013 3029 6057 3071
rect 3905 2994 3917 3014
rect 3937 2994 3949 3014
rect 3905 2956 3949 2994
rect 7749 3027 7793 3069
rect 7749 3007 7761 3027
rect 7781 3007 7793 3027
rect 7749 3000 7793 3007
rect 7748 2969 7793 3000
rect 7843 3027 7885 3069
rect 7843 3007 7857 3027
rect 7877 3007 7885 3027
rect 7843 2969 7885 3007
rect 7959 3027 8001 3069
rect 7959 3007 7967 3027
rect 7987 3007 8001 3027
rect 7959 2969 8001 3007
rect 8051 3027 8095 3069
rect 8051 3007 8063 3027
rect 8083 3007 8095 3027
rect 8051 2969 8095 3007
rect 8177 3027 8219 3069
rect 8177 3007 8185 3027
rect 8205 3007 8219 3027
rect 8177 2969 8219 3007
rect 8269 3027 8313 3069
rect 8269 3007 8281 3027
rect 8301 3007 8313 3027
rect 8269 2969 8313 3007
rect 332 2850 376 2888
rect 332 2830 344 2850
rect 364 2830 376 2850
rect 332 2788 376 2830
rect 426 2850 468 2888
rect 426 2830 440 2850
rect 460 2830 468 2850
rect 426 2788 468 2830
rect 550 2850 594 2888
rect 550 2830 562 2850
rect 582 2830 594 2850
rect 550 2788 594 2830
rect 644 2850 686 2888
rect 644 2830 658 2850
rect 678 2830 686 2850
rect 644 2788 686 2830
rect 760 2850 802 2888
rect 760 2830 768 2850
rect 788 2830 802 2850
rect 760 2788 802 2830
rect 852 2857 897 2888
rect 852 2850 896 2857
rect 852 2830 864 2850
rect 884 2830 896 2850
rect 4696 2863 4740 2901
rect 852 2788 896 2830
rect 2422 2790 2466 2832
rect 2422 2770 2434 2790
rect 2454 2770 2466 2790
rect 2422 2763 2466 2770
rect 2421 2732 2466 2763
rect 2516 2790 2558 2832
rect 2516 2770 2530 2790
rect 2550 2770 2558 2790
rect 2516 2732 2558 2770
rect 2632 2790 2674 2832
rect 2632 2770 2640 2790
rect 2660 2770 2674 2790
rect 2632 2732 2674 2770
rect 2724 2790 2768 2832
rect 2724 2770 2736 2790
rect 2756 2770 2768 2790
rect 2724 2732 2768 2770
rect 2850 2790 2892 2832
rect 2850 2770 2858 2790
rect 2878 2770 2892 2790
rect 2850 2732 2892 2770
rect 2942 2790 2986 2832
rect 4696 2843 4708 2863
rect 4728 2843 4740 2863
rect 2942 2770 2954 2790
rect 2974 2770 2986 2790
rect 4696 2801 4740 2843
rect 4790 2863 4832 2901
rect 4790 2843 4804 2863
rect 4824 2843 4832 2863
rect 4790 2801 4832 2843
rect 4914 2863 4958 2901
rect 4914 2843 4926 2863
rect 4946 2843 4958 2863
rect 4914 2801 4958 2843
rect 5008 2863 5050 2901
rect 5008 2843 5022 2863
rect 5042 2843 5050 2863
rect 5008 2801 5050 2843
rect 5124 2863 5166 2901
rect 5124 2843 5132 2863
rect 5152 2843 5166 2863
rect 5124 2801 5166 2843
rect 5216 2870 5261 2901
rect 5216 2863 5260 2870
rect 5216 2843 5228 2863
rect 5248 2843 5260 2863
rect 5216 2801 5260 2843
rect 6786 2803 6830 2845
rect 2942 2732 2986 2770
rect 6786 2783 6798 2803
rect 6818 2783 6830 2803
rect 6786 2776 6830 2783
rect 6785 2745 6830 2776
rect 6880 2803 6922 2845
rect 6880 2783 6894 2803
rect 6914 2783 6922 2803
rect 6880 2745 6922 2783
rect 6996 2803 7038 2845
rect 6996 2783 7004 2803
rect 7024 2783 7038 2803
rect 6996 2745 7038 2783
rect 7088 2803 7132 2845
rect 7088 2783 7100 2803
rect 7120 2783 7132 2803
rect 7088 2745 7132 2783
rect 7214 2803 7256 2845
rect 7214 2783 7222 2803
rect 7242 2783 7256 2803
rect 7214 2745 7256 2783
rect 7306 2803 7350 2845
rect 7306 2783 7318 2803
rect 7338 2783 7350 2803
rect 7306 2745 7350 2783
rect 1274 2468 1318 2506
rect 1274 2448 1286 2468
rect 1306 2448 1318 2468
rect 1274 2406 1318 2448
rect 1368 2468 1410 2506
rect 1368 2448 1382 2468
rect 1402 2448 1410 2468
rect 1368 2406 1410 2448
rect 1492 2468 1536 2506
rect 1492 2448 1504 2468
rect 1524 2448 1536 2468
rect 1492 2406 1536 2448
rect 1586 2468 1628 2506
rect 1586 2448 1600 2468
rect 1620 2448 1628 2468
rect 1586 2406 1628 2448
rect 1702 2468 1744 2506
rect 1702 2448 1710 2468
rect 1730 2448 1744 2468
rect 1702 2406 1744 2448
rect 1794 2475 1839 2506
rect 1794 2468 1838 2475
rect 1794 2448 1806 2468
rect 1826 2448 1838 2468
rect 5638 2481 5682 2519
rect 1794 2406 1838 2448
rect 3364 2408 3408 2450
rect 3364 2388 3376 2408
rect 3396 2388 3408 2408
rect 3364 2381 3408 2388
rect 3363 2350 3408 2381
rect 3458 2408 3500 2450
rect 3458 2388 3472 2408
rect 3492 2388 3500 2408
rect 3458 2350 3500 2388
rect 3574 2408 3616 2450
rect 3574 2388 3582 2408
rect 3602 2388 3616 2408
rect 3574 2350 3616 2388
rect 3666 2408 3710 2450
rect 3666 2388 3678 2408
rect 3698 2388 3710 2408
rect 3666 2350 3710 2388
rect 3792 2408 3834 2450
rect 3792 2388 3800 2408
rect 3820 2388 3834 2408
rect 3792 2350 3834 2388
rect 3884 2408 3928 2450
rect 5638 2461 5650 2481
rect 5670 2461 5682 2481
rect 3884 2388 3896 2408
rect 3916 2388 3928 2408
rect 5638 2419 5682 2461
rect 5732 2481 5774 2519
rect 5732 2461 5746 2481
rect 5766 2461 5774 2481
rect 5732 2419 5774 2461
rect 5856 2481 5900 2519
rect 5856 2461 5868 2481
rect 5888 2461 5900 2481
rect 5856 2419 5900 2461
rect 5950 2481 5992 2519
rect 5950 2461 5964 2481
rect 5984 2461 5992 2481
rect 5950 2419 5992 2461
rect 6066 2481 6108 2519
rect 6066 2461 6074 2481
rect 6094 2461 6108 2481
rect 6066 2419 6108 2461
rect 6158 2488 6203 2519
rect 6158 2481 6202 2488
rect 6158 2461 6170 2481
rect 6190 2461 6202 2481
rect 6158 2419 6202 2461
rect 7728 2421 7772 2463
rect 3884 2350 3928 2388
rect 7728 2401 7740 2421
rect 7760 2401 7772 2421
rect 7728 2394 7772 2401
rect 7727 2363 7772 2394
rect 7822 2421 7864 2463
rect 7822 2401 7836 2421
rect 7856 2401 7864 2421
rect 7822 2363 7864 2401
rect 7938 2421 7980 2463
rect 7938 2401 7946 2421
rect 7966 2401 7980 2421
rect 7938 2363 7980 2401
rect 8030 2421 8074 2463
rect 8030 2401 8042 2421
rect 8062 2401 8074 2421
rect 8030 2363 8074 2401
rect 8156 2421 8198 2463
rect 8156 2401 8164 2421
rect 8184 2401 8198 2421
rect 8156 2363 8198 2401
rect 8248 2421 8292 2463
rect 8248 2401 8260 2421
rect 8280 2401 8292 2421
rect 8248 2363 8292 2401
rect 311 2244 355 2282
rect 311 2224 323 2244
rect 343 2224 355 2244
rect 311 2182 355 2224
rect 405 2244 447 2282
rect 405 2224 419 2244
rect 439 2224 447 2244
rect 405 2182 447 2224
rect 529 2244 573 2282
rect 529 2224 541 2244
rect 561 2224 573 2244
rect 529 2182 573 2224
rect 623 2244 665 2282
rect 623 2224 637 2244
rect 657 2224 665 2244
rect 623 2182 665 2224
rect 739 2244 781 2282
rect 739 2224 747 2244
rect 767 2224 781 2244
rect 739 2182 781 2224
rect 831 2251 876 2282
rect 831 2244 875 2251
rect 831 2224 843 2244
rect 863 2224 875 2244
rect 831 2182 875 2224
rect 4675 2257 4719 2295
rect 4675 2237 4687 2257
rect 4707 2237 4719 2257
rect 2567 2180 2611 2222
rect 2567 2160 2579 2180
rect 2599 2160 2611 2180
rect 2567 2153 2611 2160
rect 2566 2122 2611 2153
rect 2661 2180 2703 2222
rect 2661 2160 2675 2180
rect 2695 2160 2703 2180
rect 2661 2122 2703 2160
rect 2777 2180 2819 2222
rect 2777 2160 2785 2180
rect 2805 2160 2819 2180
rect 2777 2122 2819 2160
rect 2869 2180 2913 2222
rect 2869 2160 2881 2180
rect 2901 2160 2913 2180
rect 2869 2122 2913 2160
rect 2995 2180 3037 2222
rect 2995 2160 3003 2180
rect 3023 2160 3037 2180
rect 2995 2122 3037 2160
rect 3087 2180 3131 2222
rect 4675 2195 4719 2237
rect 4769 2257 4811 2295
rect 4769 2237 4783 2257
rect 4803 2237 4811 2257
rect 4769 2195 4811 2237
rect 4893 2257 4937 2295
rect 4893 2237 4905 2257
rect 4925 2237 4937 2257
rect 4893 2195 4937 2237
rect 4987 2257 5029 2295
rect 4987 2237 5001 2257
rect 5021 2237 5029 2257
rect 4987 2195 5029 2237
rect 5103 2257 5145 2295
rect 5103 2237 5111 2257
rect 5131 2237 5145 2257
rect 5103 2195 5145 2237
rect 5195 2264 5240 2295
rect 5195 2257 5239 2264
rect 5195 2237 5207 2257
rect 5227 2237 5239 2257
rect 5195 2195 5239 2237
rect 3087 2160 3099 2180
rect 3119 2160 3131 2180
rect 3087 2122 3131 2160
rect 1109 2060 1153 2098
rect 1109 2040 1121 2060
rect 1141 2040 1153 2060
rect 1109 1998 1153 2040
rect 1203 2060 1245 2098
rect 1203 2040 1217 2060
rect 1237 2040 1245 2060
rect 1203 1998 1245 2040
rect 1327 2060 1371 2098
rect 1327 2040 1339 2060
rect 1359 2040 1371 2060
rect 1327 1998 1371 2040
rect 1421 2060 1463 2098
rect 1421 2040 1435 2060
rect 1455 2040 1463 2060
rect 1421 1998 1463 2040
rect 1537 2060 1579 2098
rect 1537 2040 1545 2060
rect 1565 2040 1579 2060
rect 1537 1998 1579 2040
rect 1629 2067 1674 2098
rect 1629 2060 1673 2067
rect 1629 2040 1641 2060
rect 1661 2040 1673 2060
rect 1629 1998 1673 2040
rect 6931 2193 6975 2235
rect 6931 2173 6943 2193
rect 6963 2173 6975 2193
rect 6931 2166 6975 2173
rect 6930 2135 6975 2166
rect 7025 2193 7067 2235
rect 7025 2173 7039 2193
rect 7059 2173 7067 2193
rect 7025 2135 7067 2173
rect 7141 2193 7183 2235
rect 7141 2173 7149 2193
rect 7169 2173 7183 2193
rect 7141 2135 7183 2173
rect 7233 2193 7277 2235
rect 7233 2173 7245 2193
rect 7265 2173 7277 2193
rect 7233 2135 7277 2173
rect 7359 2193 7401 2235
rect 7359 2173 7367 2193
rect 7387 2173 7401 2193
rect 7359 2135 7401 2173
rect 7451 2193 7495 2235
rect 7451 2173 7463 2193
rect 7483 2173 7495 2193
rect 7451 2135 7495 2173
rect 5473 2073 5517 2111
rect 5473 2053 5485 2073
rect 5505 2053 5517 2073
rect 3365 1996 3409 2038
rect 3365 1976 3377 1996
rect 3397 1976 3409 1996
rect 3365 1969 3409 1976
rect 3364 1938 3409 1969
rect 3459 1996 3501 2038
rect 3459 1976 3473 1996
rect 3493 1976 3501 1996
rect 3459 1938 3501 1976
rect 3575 1996 3617 2038
rect 3575 1976 3583 1996
rect 3603 1976 3617 1996
rect 3575 1938 3617 1976
rect 3667 1996 3711 2038
rect 3667 1976 3679 1996
rect 3699 1976 3711 1996
rect 3667 1938 3711 1976
rect 3793 1996 3835 2038
rect 3793 1976 3801 1996
rect 3821 1976 3835 1996
rect 3793 1938 3835 1976
rect 3885 1996 3929 2038
rect 5473 2011 5517 2053
rect 5567 2073 5609 2111
rect 5567 2053 5581 2073
rect 5601 2053 5609 2073
rect 5567 2011 5609 2053
rect 5691 2073 5735 2111
rect 5691 2053 5703 2073
rect 5723 2053 5735 2073
rect 5691 2011 5735 2053
rect 5785 2073 5827 2111
rect 5785 2053 5799 2073
rect 5819 2053 5827 2073
rect 5785 2011 5827 2053
rect 5901 2073 5943 2111
rect 5901 2053 5909 2073
rect 5929 2053 5943 2073
rect 5901 2011 5943 2053
rect 5993 2080 6038 2111
rect 5993 2073 6037 2080
rect 5993 2053 6005 2073
rect 6025 2053 6037 2073
rect 5993 2011 6037 2053
rect 3885 1976 3897 1996
rect 3917 1976 3929 1996
rect 3885 1938 3929 1976
rect 7729 2009 7773 2051
rect 7729 1989 7741 2009
rect 7761 1989 7773 2009
rect 7729 1982 7773 1989
rect 7728 1951 7773 1982
rect 7823 2009 7865 2051
rect 7823 1989 7837 2009
rect 7857 1989 7865 2009
rect 7823 1951 7865 1989
rect 7939 2009 7981 2051
rect 7939 1989 7947 2009
rect 7967 1989 7981 2009
rect 7939 1951 7981 1989
rect 8031 2009 8075 2051
rect 8031 1989 8043 2009
rect 8063 1989 8075 2009
rect 8031 1951 8075 1989
rect 8157 2009 8199 2051
rect 8157 1989 8165 2009
rect 8185 1989 8199 2009
rect 8157 1951 8199 1989
rect 8249 2009 8293 2051
rect 8249 1989 8261 2009
rect 8281 1989 8293 2009
rect 8249 1951 8293 1989
rect 312 1832 356 1870
rect 312 1812 324 1832
rect 344 1812 356 1832
rect 312 1770 356 1812
rect 406 1832 448 1870
rect 406 1812 420 1832
rect 440 1812 448 1832
rect 406 1770 448 1812
rect 530 1832 574 1870
rect 530 1812 542 1832
rect 562 1812 574 1832
rect 530 1770 574 1812
rect 624 1832 666 1870
rect 624 1812 638 1832
rect 658 1812 666 1832
rect 624 1770 666 1812
rect 740 1832 782 1870
rect 740 1812 748 1832
rect 768 1812 782 1832
rect 740 1770 782 1812
rect 832 1839 877 1870
rect 832 1832 876 1839
rect 832 1812 844 1832
rect 864 1812 876 1832
rect 4676 1845 4720 1883
rect 832 1770 876 1812
rect 2468 1770 2512 1812
rect 2468 1750 2480 1770
rect 2500 1750 2512 1770
rect 2468 1743 2512 1750
rect 2467 1712 2512 1743
rect 2562 1770 2604 1812
rect 2562 1750 2576 1770
rect 2596 1750 2604 1770
rect 2562 1712 2604 1750
rect 2678 1770 2720 1812
rect 2678 1750 2686 1770
rect 2706 1750 2720 1770
rect 2678 1712 2720 1750
rect 2770 1770 2814 1812
rect 2770 1750 2782 1770
rect 2802 1750 2814 1770
rect 2770 1712 2814 1750
rect 2896 1770 2938 1812
rect 2896 1750 2904 1770
rect 2924 1750 2938 1770
rect 2896 1712 2938 1750
rect 2988 1770 3032 1812
rect 4676 1825 4688 1845
rect 4708 1825 4720 1845
rect 2988 1750 3000 1770
rect 3020 1750 3032 1770
rect 4676 1783 4720 1825
rect 4770 1845 4812 1883
rect 4770 1825 4784 1845
rect 4804 1825 4812 1845
rect 4770 1783 4812 1825
rect 4894 1845 4938 1883
rect 4894 1825 4906 1845
rect 4926 1825 4938 1845
rect 4894 1783 4938 1825
rect 4988 1845 5030 1883
rect 4988 1825 5002 1845
rect 5022 1825 5030 1845
rect 4988 1783 5030 1825
rect 5104 1845 5146 1883
rect 5104 1825 5112 1845
rect 5132 1825 5146 1845
rect 5104 1783 5146 1825
rect 5196 1852 5241 1883
rect 5196 1845 5240 1852
rect 5196 1825 5208 1845
rect 5228 1825 5240 1845
rect 5196 1783 5240 1825
rect 6832 1783 6876 1825
rect 2988 1712 3032 1750
rect 6832 1763 6844 1783
rect 6864 1763 6876 1783
rect 6832 1756 6876 1763
rect 6831 1725 6876 1756
rect 6926 1783 6968 1825
rect 6926 1763 6940 1783
rect 6960 1763 6968 1783
rect 6926 1725 6968 1763
rect 7042 1783 7084 1825
rect 7042 1763 7050 1783
rect 7070 1763 7084 1783
rect 7042 1725 7084 1763
rect 7134 1783 7178 1825
rect 7134 1763 7146 1783
rect 7166 1763 7178 1783
rect 7134 1725 7178 1763
rect 7260 1783 7302 1825
rect 7260 1763 7268 1783
rect 7288 1763 7302 1783
rect 7260 1725 7302 1763
rect 7352 1783 7396 1825
rect 7352 1763 7364 1783
rect 7384 1763 7396 1783
rect 7352 1725 7396 1763
rect 1191 1452 1235 1490
rect 1191 1432 1203 1452
rect 1223 1432 1235 1452
rect 1191 1390 1235 1432
rect 1285 1452 1327 1490
rect 1285 1432 1299 1452
rect 1319 1432 1327 1452
rect 1285 1390 1327 1432
rect 1409 1452 1453 1490
rect 1409 1432 1421 1452
rect 1441 1432 1453 1452
rect 1409 1390 1453 1432
rect 1503 1452 1545 1490
rect 1503 1432 1517 1452
rect 1537 1432 1545 1452
rect 1503 1390 1545 1432
rect 1619 1452 1661 1490
rect 1619 1432 1627 1452
rect 1647 1432 1661 1452
rect 1619 1390 1661 1432
rect 1711 1459 1756 1490
rect 1711 1452 1755 1459
rect 1711 1432 1723 1452
rect 1743 1432 1755 1452
rect 5555 1465 5599 1503
rect 1711 1390 1755 1432
rect 3347 1390 3391 1432
rect 3347 1370 3359 1390
rect 3379 1370 3391 1390
rect 3347 1363 3391 1370
rect 3346 1332 3391 1363
rect 3441 1390 3483 1432
rect 3441 1370 3455 1390
rect 3475 1370 3483 1390
rect 3441 1332 3483 1370
rect 3557 1390 3599 1432
rect 3557 1370 3565 1390
rect 3585 1370 3599 1390
rect 3557 1332 3599 1370
rect 3649 1390 3693 1432
rect 3649 1370 3661 1390
rect 3681 1370 3693 1390
rect 3649 1332 3693 1370
rect 3775 1390 3817 1432
rect 3775 1370 3783 1390
rect 3803 1370 3817 1390
rect 3775 1332 3817 1370
rect 3867 1390 3911 1432
rect 5555 1445 5567 1465
rect 5587 1445 5599 1465
rect 3867 1370 3879 1390
rect 3899 1370 3911 1390
rect 5555 1403 5599 1445
rect 5649 1465 5691 1503
rect 5649 1445 5663 1465
rect 5683 1445 5691 1465
rect 5649 1403 5691 1445
rect 5773 1465 5817 1503
rect 5773 1445 5785 1465
rect 5805 1445 5817 1465
rect 5773 1403 5817 1445
rect 5867 1465 5909 1503
rect 5867 1445 5881 1465
rect 5901 1445 5909 1465
rect 5867 1403 5909 1445
rect 5983 1465 6025 1503
rect 5983 1445 5991 1465
rect 6011 1445 6025 1465
rect 5983 1403 6025 1445
rect 6075 1472 6120 1503
rect 6075 1465 6119 1472
rect 6075 1445 6087 1465
rect 6107 1445 6119 1465
rect 6075 1403 6119 1445
rect 7711 1403 7755 1445
rect 3867 1332 3911 1370
rect 7711 1383 7723 1403
rect 7743 1383 7755 1403
rect 7711 1376 7755 1383
rect 7710 1345 7755 1376
rect 7805 1403 7847 1445
rect 7805 1383 7819 1403
rect 7839 1383 7847 1403
rect 7805 1345 7847 1383
rect 7921 1403 7963 1445
rect 7921 1383 7929 1403
rect 7949 1383 7963 1403
rect 7921 1345 7963 1383
rect 8013 1403 8057 1445
rect 8013 1383 8025 1403
rect 8045 1383 8057 1403
rect 8013 1345 8057 1383
rect 8139 1403 8181 1445
rect 8139 1383 8147 1403
rect 8167 1383 8181 1403
rect 8139 1345 8181 1383
rect 8231 1403 8275 1445
rect 8231 1383 8243 1403
rect 8263 1383 8275 1403
rect 8231 1345 8275 1383
rect 294 1226 338 1264
rect 294 1206 306 1226
rect 326 1206 338 1226
rect 294 1164 338 1206
rect 388 1226 430 1264
rect 388 1206 402 1226
rect 422 1206 430 1226
rect 388 1164 430 1206
rect 512 1226 556 1264
rect 512 1206 524 1226
rect 544 1206 556 1226
rect 512 1164 556 1206
rect 606 1226 648 1264
rect 606 1206 620 1226
rect 640 1206 648 1226
rect 606 1164 648 1206
rect 722 1226 764 1264
rect 722 1206 730 1226
rect 750 1206 764 1226
rect 722 1164 764 1206
rect 814 1233 859 1264
rect 814 1226 858 1233
rect 814 1206 826 1226
rect 846 1206 858 1226
rect 814 1164 858 1206
rect 4658 1239 4702 1277
rect 4658 1219 4670 1239
rect 4690 1219 4702 1239
rect 2550 1162 2594 1204
rect 2550 1142 2562 1162
rect 2582 1142 2594 1162
rect 2550 1135 2594 1142
rect 2549 1104 2594 1135
rect 2644 1162 2686 1204
rect 2644 1142 2658 1162
rect 2678 1142 2686 1162
rect 2644 1104 2686 1142
rect 2760 1162 2802 1204
rect 2760 1142 2768 1162
rect 2788 1142 2802 1162
rect 2760 1104 2802 1142
rect 2852 1162 2896 1204
rect 2852 1142 2864 1162
rect 2884 1142 2896 1162
rect 2852 1104 2896 1142
rect 2978 1162 3020 1204
rect 2978 1142 2986 1162
rect 3006 1142 3020 1162
rect 2978 1104 3020 1142
rect 3070 1162 3114 1204
rect 4658 1177 4702 1219
rect 4752 1239 4794 1277
rect 4752 1219 4766 1239
rect 4786 1219 4794 1239
rect 4752 1177 4794 1219
rect 4876 1239 4920 1277
rect 4876 1219 4888 1239
rect 4908 1219 4920 1239
rect 4876 1177 4920 1219
rect 4970 1239 5012 1277
rect 4970 1219 4984 1239
rect 5004 1219 5012 1239
rect 4970 1177 5012 1219
rect 5086 1239 5128 1277
rect 5086 1219 5094 1239
rect 5114 1219 5128 1239
rect 5086 1177 5128 1219
rect 5178 1246 5223 1277
rect 5178 1239 5222 1246
rect 5178 1219 5190 1239
rect 5210 1219 5222 1239
rect 5178 1177 5222 1219
rect 3070 1142 3082 1162
rect 3102 1142 3114 1162
rect 3070 1104 3114 1142
rect 1092 1042 1136 1080
rect 1092 1022 1104 1042
rect 1124 1022 1136 1042
rect 1092 980 1136 1022
rect 1186 1042 1228 1080
rect 1186 1022 1200 1042
rect 1220 1022 1228 1042
rect 1186 980 1228 1022
rect 1310 1042 1354 1080
rect 1310 1022 1322 1042
rect 1342 1022 1354 1042
rect 1310 980 1354 1022
rect 1404 1042 1446 1080
rect 1404 1022 1418 1042
rect 1438 1022 1446 1042
rect 1404 980 1446 1022
rect 1520 1042 1562 1080
rect 1520 1022 1528 1042
rect 1548 1022 1562 1042
rect 1520 980 1562 1022
rect 1612 1049 1657 1080
rect 1612 1042 1656 1049
rect 1612 1022 1624 1042
rect 1644 1022 1656 1042
rect 1612 980 1656 1022
rect 6914 1175 6958 1217
rect 6914 1155 6926 1175
rect 6946 1155 6958 1175
rect 6914 1148 6958 1155
rect 6913 1117 6958 1148
rect 7008 1175 7050 1217
rect 7008 1155 7022 1175
rect 7042 1155 7050 1175
rect 7008 1117 7050 1155
rect 7124 1175 7166 1217
rect 7124 1155 7132 1175
rect 7152 1155 7166 1175
rect 7124 1117 7166 1155
rect 7216 1175 7260 1217
rect 7216 1155 7228 1175
rect 7248 1155 7260 1175
rect 7216 1117 7260 1155
rect 7342 1175 7384 1217
rect 7342 1155 7350 1175
rect 7370 1155 7384 1175
rect 7342 1117 7384 1155
rect 7434 1175 7478 1217
rect 7434 1155 7446 1175
rect 7466 1155 7478 1175
rect 7434 1117 7478 1155
rect 5456 1055 5500 1093
rect 5456 1035 5468 1055
rect 5488 1035 5500 1055
rect 3348 978 3392 1020
rect 3348 958 3360 978
rect 3380 958 3392 978
rect 3348 951 3392 958
rect 3347 920 3392 951
rect 3442 978 3484 1020
rect 3442 958 3456 978
rect 3476 958 3484 978
rect 3442 920 3484 958
rect 3558 978 3600 1020
rect 3558 958 3566 978
rect 3586 958 3600 978
rect 3558 920 3600 958
rect 3650 978 3694 1020
rect 3650 958 3662 978
rect 3682 958 3694 978
rect 3650 920 3694 958
rect 3776 978 3818 1020
rect 3776 958 3784 978
rect 3804 958 3818 978
rect 3776 920 3818 958
rect 3868 978 3912 1020
rect 5456 993 5500 1035
rect 5550 1055 5592 1093
rect 5550 1035 5564 1055
rect 5584 1035 5592 1055
rect 5550 993 5592 1035
rect 5674 1055 5718 1093
rect 5674 1035 5686 1055
rect 5706 1035 5718 1055
rect 5674 993 5718 1035
rect 5768 1055 5810 1093
rect 5768 1035 5782 1055
rect 5802 1035 5810 1055
rect 5768 993 5810 1035
rect 5884 1055 5926 1093
rect 5884 1035 5892 1055
rect 5912 1035 5926 1055
rect 5884 993 5926 1035
rect 5976 1062 6021 1093
rect 5976 1055 6020 1062
rect 5976 1035 5988 1055
rect 6008 1035 6020 1055
rect 5976 993 6020 1035
rect 3868 958 3880 978
rect 3900 958 3912 978
rect 3868 920 3912 958
rect 7712 991 7756 1033
rect 7712 971 7724 991
rect 7744 971 7756 991
rect 7712 964 7756 971
rect 7711 933 7756 964
rect 7806 991 7848 1033
rect 7806 971 7820 991
rect 7840 971 7848 991
rect 7806 933 7848 971
rect 7922 991 7964 1033
rect 7922 971 7930 991
rect 7950 971 7964 991
rect 7922 933 7964 971
rect 8014 991 8058 1033
rect 8014 971 8026 991
rect 8046 971 8058 991
rect 8014 933 8058 971
rect 8140 991 8182 1033
rect 8140 971 8148 991
rect 8168 971 8182 991
rect 8140 933 8182 971
rect 8232 991 8276 1033
rect 8232 971 8244 991
rect 8264 971 8276 991
rect 8232 933 8276 971
rect 295 814 339 852
rect 295 794 307 814
rect 327 794 339 814
rect 295 752 339 794
rect 389 814 431 852
rect 389 794 403 814
rect 423 794 431 814
rect 389 752 431 794
rect 513 814 557 852
rect 513 794 525 814
rect 545 794 557 814
rect 513 752 557 794
rect 607 814 649 852
rect 607 794 621 814
rect 641 794 649 814
rect 607 752 649 794
rect 723 814 765 852
rect 723 794 731 814
rect 751 794 765 814
rect 723 752 765 794
rect 815 821 860 852
rect 815 814 859 821
rect 815 794 827 814
rect 847 794 859 814
rect 815 752 859 794
rect 4659 827 4703 865
rect 4659 807 4671 827
rect 4691 807 4703 827
rect 4659 765 4703 807
rect 4753 827 4795 865
rect 4753 807 4767 827
rect 4787 807 4795 827
rect 4753 765 4795 807
rect 4877 827 4921 865
rect 4877 807 4889 827
rect 4909 807 4921 827
rect 4877 765 4921 807
rect 4971 827 5013 865
rect 4971 807 4985 827
rect 5005 807 5013 827
rect 4971 765 5013 807
rect 5087 827 5129 865
rect 5087 807 5095 827
rect 5115 807 5129 827
rect 5087 765 5129 807
rect 5179 834 5224 865
rect 5179 827 5223 834
rect 5179 807 5191 827
rect 5211 807 5223 827
rect 5179 765 5223 807
rect 1508 238 1552 276
rect 1508 218 1520 238
rect 1540 218 1552 238
rect 1508 176 1552 218
rect 1602 238 1644 276
rect 1602 218 1616 238
rect 1636 218 1644 238
rect 1602 176 1644 218
rect 1726 238 1770 276
rect 1726 218 1738 238
rect 1758 218 1770 238
rect 1726 176 1770 218
rect 1820 238 1862 276
rect 1820 218 1834 238
rect 1854 218 1862 238
rect 1820 176 1862 218
rect 1936 238 1978 276
rect 1936 218 1944 238
rect 1964 218 1978 238
rect 1936 176 1978 218
rect 2028 245 2073 276
rect 5872 251 5916 289
rect 2028 238 2072 245
rect 2028 218 2040 238
rect 2060 218 2072 238
rect 2028 176 2072 218
rect 5872 231 5884 251
rect 5904 231 5916 251
rect 3997 164 4041 202
rect 3997 144 4009 164
rect 4029 144 4041 164
rect 3997 102 4041 144
rect 4091 164 4133 202
rect 4091 144 4105 164
rect 4125 144 4133 164
rect 4091 102 4133 144
rect 4215 164 4259 202
rect 4215 144 4227 164
rect 4247 144 4259 164
rect 4215 102 4259 144
rect 4309 164 4351 202
rect 4309 144 4323 164
rect 4343 144 4351 164
rect 4309 102 4351 144
rect 4425 164 4467 202
rect 4425 144 4433 164
rect 4453 144 4467 164
rect 4425 102 4467 144
rect 4517 171 4562 202
rect 5872 189 5916 231
rect 5966 251 6008 289
rect 5966 231 5980 251
rect 6000 231 6008 251
rect 5966 189 6008 231
rect 6090 251 6134 289
rect 6090 231 6102 251
rect 6122 231 6134 251
rect 6090 189 6134 231
rect 6184 251 6226 289
rect 6184 231 6198 251
rect 6218 231 6226 251
rect 6184 189 6226 231
rect 6300 251 6342 289
rect 6300 231 6308 251
rect 6328 231 6342 251
rect 6300 189 6342 231
rect 6392 258 6437 289
rect 6392 251 6436 258
rect 6392 231 6404 251
rect 6424 231 6436 251
rect 6392 189 6436 231
rect 4517 164 4561 171
rect 4517 144 4529 164
rect 4549 144 4561 164
rect 4517 102 4561 144
<< ndiffc >>
rect 3480 8645 3500 8665
rect 3583 8641 3603 8661
rect 3691 8641 3711 8661
rect 3794 8645 3814 8665
rect 3909 8641 3929 8661
rect 4012 8645 4032 8665
rect 4199 8652 4217 8670
rect 263 8590 281 8608
rect 7844 8658 7864 8678
rect 7947 8654 7967 8674
rect 8055 8654 8075 8674
rect 8158 8658 8178 8678
rect 8273 8654 8293 8674
rect 8376 8658 8396 8678
rect 8563 8665 8581 8683
rect 4627 8603 4645 8621
rect 261 8491 279 8509
rect 4197 8553 4215 8571
rect 4625 8504 4643 8522
rect 2683 8417 2703 8437
rect 2786 8413 2806 8433
rect 2894 8413 2914 8433
rect 2997 8417 3017 8437
rect 3112 8413 3132 8433
rect 8561 8566 8579 8584
rect 3215 8417 3235 8437
rect 4192 8434 4210 8452
rect 7047 8430 7067 8450
rect 7150 8426 7170 8446
rect 7258 8426 7278 8446
rect 7361 8430 7381 8450
rect 7476 8426 7496 8446
rect 7579 8430 7599 8450
rect 8556 8447 8574 8465
rect 4190 8335 4208 8353
rect 258 8266 276 8284
rect 8554 8348 8572 8366
rect 3481 8233 3501 8253
rect 256 8167 274 8185
rect 427 8183 447 8203
rect 530 8187 550 8207
rect 645 8183 665 8203
rect 748 8187 768 8207
rect 856 8187 876 8207
rect 3584 8229 3604 8249
rect 3692 8229 3712 8249
rect 3795 8233 3815 8253
rect 3910 8229 3930 8249
rect 4013 8233 4033 8253
rect 4186 8251 4204 8269
rect 4622 8279 4640 8297
rect 959 8183 979 8203
rect 7845 8246 7865 8266
rect 4184 8152 4202 8170
rect 4620 8180 4638 8198
rect 4791 8196 4811 8216
rect 4894 8200 4914 8220
rect 5009 8196 5029 8216
rect 5112 8200 5132 8220
rect 5220 8200 5240 8220
rect 7948 8242 7968 8262
rect 8056 8242 8076 8262
rect 8159 8246 8179 8266
rect 8274 8242 8294 8262
rect 8377 8246 8397 8266
rect 8550 8264 8568 8282
rect 5323 8196 5343 8216
rect 252 8083 270 8101
rect 8548 8165 8566 8183
rect 4616 8096 4634 8114
rect 250 7984 268 8002
rect 1225 7999 1245 8019
rect 1328 8003 1348 8023
rect 1443 7999 1463 8019
rect 1546 8003 1566 8023
rect 1654 8003 1674 8023
rect 1757 7999 1777 8019
rect 2584 8007 2604 8027
rect 2687 8003 2707 8023
rect 2795 8003 2815 8023
rect 2898 8007 2918 8027
rect 3013 8003 3033 8023
rect 3116 8007 3136 8027
rect 4614 7997 4632 8015
rect 5589 8012 5609 8032
rect 245 7865 263 7883
rect 5692 8016 5712 8036
rect 5807 8012 5827 8032
rect 5910 8016 5930 8036
rect 6018 8016 6038 8036
rect 6121 8012 6141 8032
rect 6948 8020 6968 8040
rect 7051 8016 7071 8036
rect 7159 8016 7179 8036
rect 7262 8020 7282 8040
rect 7377 8016 7397 8036
rect 7480 8020 7500 8040
rect 4181 7927 4199 7945
rect 4609 7878 4627 7896
rect 8545 7940 8563 7958
rect 4179 7828 4197 7846
rect 243 7766 261 7784
rect 428 7771 448 7791
rect 531 7775 551 7795
rect 646 7771 666 7791
rect 749 7775 769 7795
rect 857 7775 877 7795
rect 960 7771 980 7791
rect 8543 7841 8561 7859
rect 4607 7779 4625 7797
rect 4792 7784 4812 7804
rect 4895 7788 4915 7808
rect 5010 7784 5030 7804
rect 5113 7788 5133 7808
rect 5221 7788 5241 7808
rect 5324 7784 5344 7804
rect 3463 7627 3483 7647
rect 3566 7623 3586 7643
rect 3674 7623 3694 7643
rect 3777 7627 3797 7647
rect 3892 7623 3912 7643
rect 3995 7627 4015 7647
rect 4182 7634 4200 7652
rect 246 7572 264 7590
rect 7827 7640 7847 7660
rect 7930 7636 7950 7656
rect 8038 7636 8058 7656
rect 8141 7640 8161 7660
rect 8256 7636 8276 7656
rect 8359 7640 8379 7660
rect 8546 7647 8564 7665
rect 4610 7585 4628 7603
rect 244 7473 262 7491
rect 4180 7535 4198 7553
rect 4608 7486 4626 7504
rect 1307 7391 1327 7411
rect 1410 7395 1430 7415
rect 1525 7391 1545 7411
rect 1628 7395 1648 7415
rect 1736 7395 1756 7415
rect 1839 7391 1859 7411
rect 2666 7399 2686 7419
rect 2769 7395 2789 7415
rect 2877 7395 2897 7415
rect 2980 7399 3000 7419
rect 3095 7395 3115 7415
rect 8544 7548 8562 7566
rect 3198 7399 3218 7419
rect 4175 7416 4193 7434
rect 5671 7404 5691 7424
rect 5774 7408 5794 7428
rect 5889 7404 5909 7424
rect 5992 7408 6012 7428
rect 6100 7408 6120 7428
rect 6203 7404 6223 7424
rect 7030 7412 7050 7432
rect 7133 7408 7153 7428
rect 7241 7408 7261 7428
rect 7344 7412 7364 7432
rect 7459 7408 7479 7428
rect 7562 7412 7582 7432
rect 8539 7429 8557 7447
rect 4173 7317 4191 7335
rect 241 7248 259 7266
rect 8537 7330 8555 7348
rect 3464 7215 3484 7235
rect 239 7149 257 7167
rect 410 7165 430 7185
rect 513 7169 533 7189
rect 628 7165 648 7185
rect 731 7169 751 7189
rect 839 7169 859 7189
rect 3567 7211 3587 7231
rect 3675 7211 3695 7231
rect 3778 7215 3798 7235
rect 3893 7211 3913 7231
rect 3996 7215 4016 7235
rect 4169 7233 4187 7251
rect 4605 7261 4623 7279
rect 942 7165 962 7185
rect 7828 7228 7848 7248
rect 4167 7134 4185 7152
rect 4603 7162 4621 7180
rect 4774 7178 4794 7198
rect 4877 7182 4897 7202
rect 4992 7178 5012 7198
rect 5095 7182 5115 7202
rect 5203 7182 5223 7202
rect 7931 7224 7951 7244
rect 8039 7224 8059 7244
rect 8142 7228 8162 7248
rect 8257 7224 8277 7244
rect 8360 7228 8380 7248
rect 8533 7246 8551 7264
rect 5306 7178 5326 7198
rect 235 7065 253 7083
rect 8531 7147 8549 7165
rect 4599 7078 4617 7096
rect 233 6966 251 6984
rect 1208 6981 1228 7001
rect 1311 6985 1331 7005
rect 1426 6981 1446 7001
rect 1529 6985 1549 7005
rect 1637 6985 1657 7005
rect 1740 6981 1760 7001
rect 2501 6991 2521 7011
rect 2604 6987 2624 7007
rect 2712 6987 2732 7007
rect 2815 6991 2835 7011
rect 2930 6987 2950 7007
rect 3033 6991 3053 7011
rect 228 6847 246 6865
rect 4597 6979 4615 6997
rect 5572 6994 5592 7014
rect 5675 6998 5695 7018
rect 5790 6994 5810 7014
rect 5893 6998 5913 7018
rect 6001 6998 6021 7018
rect 6104 6994 6124 7014
rect 6865 7004 6885 7024
rect 6968 7000 6988 7020
rect 7076 7000 7096 7020
rect 7179 7004 7199 7024
rect 7294 7000 7314 7020
rect 7397 7004 7417 7024
rect 4164 6909 4182 6927
rect 4592 6860 4610 6878
rect 8528 6922 8546 6940
rect 4162 6810 4180 6828
rect 226 6748 244 6766
rect 411 6753 431 6773
rect 514 6757 534 6777
rect 629 6753 649 6773
rect 732 6757 752 6777
rect 840 6757 860 6777
rect 943 6753 963 6773
rect 8526 6823 8544 6841
rect 4590 6761 4608 6779
rect 4775 6766 4795 6786
rect 4878 6770 4898 6790
rect 4993 6766 5013 6786
rect 5096 6770 5116 6790
rect 5204 6770 5224 6790
rect 5307 6766 5327 6786
rect 3443 6609 3463 6629
rect 3546 6605 3566 6625
rect 3654 6605 3674 6625
rect 3757 6609 3777 6629
rect 3872 6605 3892 6625
rect 3975 6609 3995 6629
rect 4162 6616 4180 6634
rect 226 6554 244 6572
rect 7807 6622 7827 6642
rect 7910 6618 7930 6638
rect 8018 6618 8038 6638
rect 8121 6622 8141 6642
rect 8236 6618 8256 6638
rect 8339 6622 8359 6642
rect 8526 6629 8544 6647
rect 4590 6567 4608 6585
rect 224 6455 242 6473
rect 4160 6517 4178 6535
rect 4588 6468 4606 6486
rect 1353 6371 1373 6391
rect 1456 6375 1476 6395
rect 1571 6371 1591 6391
rect 1674 6375 1694 6395
rect 1782 6375 1802 6395
rect 1885 6371 1905 6391
rect 2646 6381 2666 6401
rect 2749 6377 2769 6397
rect 2857 6377 2877 6397
rect 2960 6381 2980 6401
rect 3075 6377 3095 6397
rect 3178 6381 3198 6401
rect 4155 6398 4173 6416
rect 8524 6530 8542 6548
rect 5717 6384 5737 6404
rect 5820 6388 5840 6408
rect 5935 6384 5955 6404
rect 6038 6388 6058 6408
rect 6146 6388 6166 6408
rect 6249 6384 6269 6404
rect 7010 6394 7030 6414
rect 7113 6390 7133 6410
rect 7221 6390 7241 6410
rect 7324 6394 7344 6414
rect 7439 6390 7459 6410
rect 7542 6394 7562 6414
rect 8519 6411 8537 6429
rect 4153 6299 4171 6317
rect 221 6230 239 6248
rect 8517 6312 8535 6330
rect 3444 6197 3464 6217
rect 219 6131 237 6149
rect 390 6147 410 6167
rect 493 6151 513 6171
rect 608 6147 628 6167
rect 711 6151 731 6171
rect 819 6151 839 6171
rect 3547 6193 3567 6213
rect 3655 6193 3675 6213
rect 3758 6197 3778 6217
rect 3873 6193 3893 6213
rect 3976 6197 3996 6217
rect 4149 6215 4167 6233
rect 4585 6243 4603 6261
rect 922 6147 942 6167
rect 7808 6210 7828 6230
rect 4147 6116 4165 6134
rect 4583 6144 4601 6162
rect 4754 6160 4774 6180
rect 4857 6164 4877 6184
rect 4972 6160 4992 6180
rect 5075 6164 5095 6184
rect 5183 6164 5203 6184
rect 7911 6206 7931 6226
rect 8019 6206 8039 6226
rect 8122 6210 8142 6230
rect 8237 6206 8257 6226
rect 8340 6210 8360 6230
rect 8513 6228 8531 6246
rect 5286 6160 5306 6180
rect 215 6047 233 6065
rect 8511 6129 8529 6147
rect 4579 6060 4597 6078
rect 213 5948 231 5966
rect 1188 5963 1208 5983
rect 1291 5967 1311 5987
rect 1406 5963 1426 5983
rect 1509 5967 1529 5987
rect 1617 5967 1637 5987
rect 1720 5963 1740 5983
rect 2547 5971 2567 5991
rect 2650 5967 2670 5987
rect 2758 5967 2778 5987
rect 2861 5971 2881 5991
rect 2976 5967 2996 5987
rect 3079 5971 3099 5991
rect 4577 5961 4595 5979
rect 5552 5976 5572 5996
rect 208 5829 226 5847
rect 5655 5980 5675 6000
rect 5770 5976 5790 5996
rect 5873 5980 5893 6000
rect 5981 5980 6001 6000
rect 6084 5976 6104 5996
rect 6911 5984 6931 6004
rect 7014 5980 7034 6000
rect 7122 5980 7142 6000
rect 7225 5984 7245 6004
rect 7340 5980 7360 6000
rect 7443 5984 7463 6004
rect 4144 5891 4162 5909
rect 4572 5842 4590 5860
rect 8508 5904 8526 5922
rect 4142 5792 4160 5810
rect 206 5730 224 5748
rect 391 5735 411 5755
rect 494 5739 514 5759
rect 609 5735 629 5755
rect 712 5739 732 5759
rect 820 5739 840 5759
rect 923 5735 943 5755
rect 8506 5805 8524 5823
rect 4570 5743 4588 5761
rect 4755 5748 4775 5768
rect 4858 5752 4878 5772
rect 4973 5748 4993 5768
rect 5076 5752 5096 5772
rect 5184 5752 5204 5772
rect 5287 5748 5307 5768
rect 3426 5591 3446 5611
rect 3529 5587 3549 5607
rect 3637 5587 3657 5607
rect 3740 5591 3760 5611
rect 3855 5587 3875 5607
rect 3958 5591 3978 5611
rect 4145 5598 4163 5616
rect 209 5536 227 5554
rect 7790 5604 7810 5624
rect 7893 5600 7913 5620
rect 8001 5600 8021 5620
rect 8104 5604 8124 5624
rect 8219 5600 8239 5620
rect 8322 5604 8342 5624
rect 8509 5611 8527 5629
rect 4573 5549 4591 5567
rect 207 5437 225 5455
rect 4143 5499 4161 5517
rect 4571 5450 4589 5468
rect 1270 5355 1290 5375
rect 1373 5359 1393 5379
rect 1488 5355 1508 5375
rect 1591 5359 1611 5379
rect 1699 5359 1719 5379
rect 1802 5355 1822 5375
rect 2629 5363 2649 5383
rect 2732 5359 2752 5379
rect 2840 5359 2860 5379
rect 2943 5363 2963 5383
rect 3058 5359 3078 5379
rect 8507 5512 8525 5530
rect 3161 5363 3181 5383
rect 4138 5380 4156 5398
rect 5634 5368 5654 5388
rect 5737 5372 5757 5392
rect 5852 5368 5872 5388
rect 5955 5372 5975 5392
rect 6063 5372 6083 5392
rect 6166 5368 6186 5388
rect 6993 5376 7013 5396
rect 7096 5372 7116 5392
rect 7204 5372 7224 5392
rect 7307 5376 7327 5396
rect 7422 5372 7442 5392
rect 7525 5376 7545 5396
rect 8502 5393 8520 5411
rect 4136 5281 4154 5299
rect 204 5212 222 5230
rect 8500 5294 8518 5312
rect 3427 5179 3447 5199
rect 202 5113 220 5131
rect 373 5129 393 5149
rect 476 5133 496 5153
rect 591 5129 611 5149
rect 694 5133 714 5153
rect 802 5133 822 5153
rect 3530 5175 3550 5195
rect 3638 5175 3658 5195
rect 3741 5179 3761 5199
rect 3856 5175 3876 5195
rect 3959 5179 3979 5199
rect 4132 5197 4150 5215
rect 4568 5225 4586 5243
rect 905 5129 925 5149
rect 7791 5192 7811 5212
rect 4130 5098 4148 5116
rect 4566 5126 4584 5144
rect 4737 5142 4757 5162
rect 4840 5146 4860 5166
rect 4955 5142 4975 5162
rect 5058 5146 5078 5166
rect 5166 5146 5186 5166
rect 7894 5188 7914 5208
rect 8002 5188 8022 5208
rect 8105 5192 8125 5212
rect 8220 5188 8240 5208
rect 8323 5192 8343 5212
rect 8496 5210 8514 5228
rect 5269 5142 5289 5162
rect 198 5029 216 5047
rect 8494 5111 8512 5129
rect 4562 5042 4580 5060
rect 196 4930 214 4948
rect 1171 4945 1191 4965
rect 1274 4949 1294 4969
rect 1389 4945 1409 4965
rect 1492 4949 1512 4969
rect 1600 4949 1620 4969
rect 1703 4945 1723 4965
rect 2325 4957 2345 4977
rect 2428 4953 2448 4973
rect 2536 4953 2556 4973
rect 2639 4957 2659 4977
rect 2754 4953 2774 4973
rect 2857 4957 2877 4977
rect 191 4811 209 4829
rect 4560 4943 4578 4961
rect 5535 4958 5555 4978
rect 5638 4962 5658 4982
rect 5753 4958 5773 4978
rect 5856 4962 5876 4982
rect 5964 4962 5984 4982
rect 6067 4958 6087 4978
rect 6689 4970 6709 4990
rect 6792 4966 6812 4986
rect 6900 4966 6920 4986
rect 7003 4970 7023 4990
rect 7118 4966 7138 4986
rect 7221 4970 7241 4990
rect 4127 4873 4145 4891
rect 4555 4824 4573 4842
rect 8491 4886 8509 4904
rect 4125 4774 4143 4792
rect 189 4712 207 4730
rect 374 4717 394 4737
rect 477 4721 497 4741
rect 592 4717 612 4737
rect 695 4721 715 4741
rect 803 4721 823 4741
rect 906 4717 926 4737
rect 8489 4787 8507 4805
rect 4553 4725 4571 4743
rect 4738 4730 4758 4750
rect 4841 4734 4861 4754
rect 4956 4730 4976 4750
rect 5059 4734 5079 4754
rect 5167 4734 5187 4754
rect 5270 4730 5290 4750
rect 3407 4573 3427 4593
rect 3510 4569 3530 4589
rect 3618 4569 3638 4589
rect 3721 4573 3741 4593
rect 3836 4569 3856 4589
rect 3939 4573 3959 4593
rect 4126 4580 4144 4598
rect 190 4518 208 4536
rect 7771 4586 7791 4606
rect 7874 4582 7894 4602
rect 7982 4582 8002 4602
rect 8085 4586 8105 4606
rect 8200 4582 8220 4602
rect 8303 4586 8323 4606
rect 8490 4593 8508 4611
rect 4554 4531 4572 4549
rect 188 4419 206 4437
rect 4124 4481 4142 4499
rect 4552 4432 4570 4450
rect 1456 4333 1476 4353
rect 1559 4337 1579 4357
rect 1674 4333 1694 4353
rect 1777 4337 1797 4357
rect 1885 4337 1905 4357
rect 1988 4333 2008 4353
rect 2610 4345 2630 4365
rect 2713 4341 2733 4361
rect 2821 4341 2841 4361
rect 2924 4345 2944 4365
rect 3039 4341 3059 4361
rect 3142 4345 3162 4365
rect 4119 4362 4137 4380
rect 8488 4494 8506 4512
rect 5820 4346 5840 4366
rect 5923 4350 5943 4370
rect 6038 4346 6058 4366
rect 6141 4350 6161 4370
rect 6249 4350 6269 4370
rect 6352 4346 6372 4366
rect 6974 4358 6994 4378
rect 7077 4354 7097 4374
rect 7185 4354 7205 4374
rect 7288 4358 7308 4378
rect 7403 4354 7423 4374
rect 7506 4358 7526 4378
rect 8483 4375 8501 4393
rect 4117 4263 4135 4281
rect 185 4194 203 4212
rect 8481 4276 8499 4294
rect 3408 4161 3428 4181
rect 183 4095 201 4113
rect 354 4111 374 4131
rect 457 4115 477 4135
rect 572 4111 592 4131
rect 675 4115 695 4135
rect 783 4115 803 4135
rect 3511 4157 3531 4177
rect 3619 4157 3639 4177
rect 3722 4161 3742 4181
rect 3837 4157 3857 4177
rect 3940 4161 3960 4181
rect 4113 4179 4131 4197
rect 4549 4207 4567 4225
rect 886 4111 906 4131
rect 7772 4174 7792 4194
rect 4111 4080 4129 4098
rect 4547 4108 4565 4126
rect 4718 4124 4738 4144
rect 4821 4128 4841 4148
rect 4936 4124 4956 4144
rect 5039 4128 5059 4148
rect 5147 4128 5167 4148
rect 7875 4170 7895 4190
rect 7983 4170 8003 4190
rect 8086 4174 8106 4194
rect 8201 4170 8221 4190
rect 8304 4174 8324 4194
rect 8477 4192 8495 4210
rect 5250 4124 5270 4144
rect 179 4011 197 4029
rect 8475 4093 8493 4111
rect 4543 4024 4561 4042
rect 177 3912 195 3930
rect 1152 3927 1172 3947
rect 1255 3931 1275 3951
rect 1370 3927 1390 3947
rect 1473 3931 1493 3951
rect 1581 3931 1601 3951
rect 1684 3927 1704 3947
rect 2511 3935 2531 3955
rect 2614 3931 2634 3951
rect 2722 3931 2742 3951
rect 2825 3935 2845 3955
rect 2940 3931 2960 3951
rect 3043 3935 3063 3955
rect 4541 3925 4559 3943
rect 5516 3940 5536 3960
rect 172 3793 190 3811
rect 5619 3944 5639 3964
rect 5734 3940 5754 3960
rect 5837 3944 5857 3964
rect 5945 3944 5965 3964
rect 6048 3940 6068 3960
rect 6875 3948 6895 3968
rect 6978 3944 6998 3964
rect 7086 3944 7106 3964
rect 7189 3948 7209 3968
rect 7304 3944 7324 3964
rect 7407 3948 7427 3968
rect 4108 3855 4126 3873
rect 4536 3806 4554 3824
rect 8472 3868 8490 3886
rect 4106 3756 4124 3774
rect 170 3694 188 3712
rect 355 3699 375 3719
rect 458 3703 478 3723
rect 573 3699 593 3719
rect 676 3703 696 3723
rect 784 3703 804 3723
rect 887 3699 907 3719
rect 8470 3769 8488 3787
rect 4534 3707 4552 3725
rect 4719 3712 4739 3732
rect 4822 3716 4842 3736
rect 4937 3712 4957 3732
rect 5040 3716 5060 3736
rect 5148 3716 5168 3736
rect 5251 3712 5271 3732
rect 3390 3555 3410 3575
rect 3493 3551 3513 3571
rect 3601 3551 3621 3571
rect 3704 3555 3724 3575
rect 3819 3551 3839 3571
rect 3922 3555 3942 3575
rect 4109 3562 4127 3580
rect 173 3500 191 3518
rect 7754 3568 7774 3588
rect 7857 3564 7877 3584
rect 7965 3564 7985 3584
rect 8068 3568 8088 3588
rect 8183 3564 8203 3584
rect 8286 3568 8306 3588
rect 8473 3575 8491 3593
rect 4537 3513 4555 3531
rect 171 3401 189 3419
rect 4107 3463 4125 3481
rect 4535 3414 4553 3432
rect 1234 3319 1254 3339
rect 1337 3323 1357 3343
rect 1452 3319 1472 3339
rect 1555 3323 1575 3343
rect 1663 3323 1683 3343
rect 1766 3319 1786 3339
rect 2593 3327 2613 3347
rect 2696 3323 2716 3343
rect 2804 3323 2824 3343
rect 2907 3327 2927 3347
rect 3022 3323 3042 3343
rect 8471 3476 8489 3494
rect 3125 3327 3145 3347
rect 4102 3344 4120 3362
rect 5598 3332 5618 3352
rect 5701 3336 5721 3356
rect 5816 3332 5836 3352
rect 5919 3336 5939 3356
rect 6027 3336 6047 3356
rect 6130 3332 6150 3352
rect 6957 3340 6977 3360
rect 7060 3336 7080 3356
rect 7168 3336 7188 3356
rect 7271 3340 7291 3360
rect 7386 3336 7406 3356
rect 7489 3340 7509 3360
rect 8466 3357 8484 3375
rect 4100 3245 4118 3263
rect 168 3176 186 3194
rect 8464 3258 8482 3276
rect 3391 3143 3411 3163
rect 166 3077 184 3095
rect 337 3093 357 3113
rect 440 3097 460 3117
rect 555 3093 575 3113
rect 658 3097 678 3117
rect 766 3097 786 3117
rect 3494 3139 3514 3159
rect 3602 3139 3622 3159
rect 3705 3143 3725 3163
rect 3820 3139 3840 3159
rect 3923 3143 3943 3163
rect 4096 3161 4114 3179
rect 4532 3189 4550 3207
rect 869 3093 889 3113
rect 7755 3156 7775 3176
rect 4094 3062 4112 3080
rect 4530 3090 4548 3108
rect 4701 3106 4721 3126
rect 4804 3110 4824 3130
rect 4919 3106 4939 3126
rect 5022 3110 5042 3130
rect 5130 3110 5150 3130
rect 7858 3152 7878 3172
rect 7966 3152 7986 3172
rect 8069 3156 8089 3176
rect 8184 3152 8204 3172
rect 8287 3156 8307 3176
rect 8460 3174 8478 3192
rect 5233 3106 5253 3126
rect 162 2993 180 3011
rect 8458 3075 8476 3093
rect 4526 3006 4544 3024
rect 160 2894 178 2912
rect 1135 2909 1155 2929
rect 1238 2913 1258 2933
rect 1353 2909 1373 2929
rect 1456 2913 1476 2933
rect 1564 2913 1584 2933
rect 1667 2909 1687 2929
rect 2428 2919 2448 2939
rect 2531 2915 2551 2935
rect 2639 2915 2659 2935
rect 2742 2919 2762 2939
rect 2857 2915 2877 2935
rect 2960 2919 2980 2939
rect 155 2775 173 2793
rect 4524 2907 4542 2925
rect 5499 2922 5519 2942
rect 5602 2926 5622 2946
rect 5717 2922 5737 2942
rect 5820 2926 5840 2946
rect 5928 2926 5948 2946
rect 6031 2922 6051 2942
rect 6792 2932 6812 2952
rect 6895 2928 6915 2948
rect 7003 2928 7023 2948
rect 7106 2932 7126 2952
rect 7221 2928 7241 2948
rect 7324 2932 7344 2952
rect 4091 2837 4109 2855
rect 4519 2788 4537 2806
rect 8455 2850 8473 2868
rect 4089 2738 4107 2756
rect 153 2676 171 2694
rect 338 2681 358 2701
rect 441 2685 461 2705
rect 556 2681 576 2701
rect 659 2685 679 2705
rect 767 2685 787 2705
rect 870 2681 890 2701
rect 8453 2751 8471 2769
rect 4517 2689 4535 2707
rect 4702 2694 4722 2714
rect 4805 2698 4825 2718
rect 4920 2694 4940 2714
rect 5023 2698 5043 2718
rect 5131 2698 5151 2718
rect 5234 2694 5254 2714
rect 3370 2537 3390 2557
rect 3473 2533 3493 2553
rect 3581 2533 3601 2553
rect 3684 2537 3704 2557
rect 3799 2533 3819 2553
rect 3902 2537 3922 2557
rect 4089 2544 4107 2562
rect 153 2482 171 2500
rect 7734 2550 7754 2570
rect 7837 2546 7857 2566
rect 7945 2546 7965 2566
rect 8048 2550 8068 2570
rect 8163 2546 8183 2566
rect 8266 2550 8286 2570
rect 8453 2557 8471 2575
rect 4517 2495 4535 2513
rect 151 2383 169 2401
rect 4087 2445 4105 2463
rect 4515 2396 4533 2414
rect 1280 2299 1300 2319
rect 1383 2303 1403 2323
rect 1498 2299 1518 2319
rect 1601 2303 1621 2323
rect 1709 2303 1729 2323
rect 1812 2299 1832 2319
rect 2573 2309 2593 2329
rect 2676 2305 2696 2325
rect 2784 2305 2804 2325
rect 2887 2309 2907 2329
rect 3002 2305 3022 2325
rect 3105 2309 3125 2329
rect 4082 2326 4100 2344
rect 8451 2458 8469 2476
rect 5644 2312 5664 2332
rect 5747 2316 5767 2336
rect 5862 2312 5882 2332
rect 5965 2316 5985 2336
rect 6073 2316 6093 2336
rect 6176 2312 6196 2332
rect 6937 2322 6957 2342
rect 7040 2318 7060 2338
rect 7148 2318 7168 2338
rect 7251 2322 7271 2342
rect 7366 2318 7386 2338
rect 7469 2322 7489 2342
rect 8446 2339 8464 2357
rect 4080 2227 4098 2245
rect 148 2158 166 2176
rect 8444 2240 8462 2258
rect 3371 2125 3391 2145
rect 146 2059 164 2077
rect 317 2075 337 2095
rect 420 2079 440 2099
rect 535 2075 555 2095
rect 638 2079 658 2099
rect 746 2079 766 2099
rect 3474 2121 3494 2141
rect 3582 2121 3602 2141
rect 3685 2125 3705 2145
rect 3800 2121 3820 2141
rect 3903 2125 3923 2145
rect 4076 2143 4094 2161
rect 4512 2171 4530 2189
rect 849 2075 869 2095
rect 7735 2138 7755 2158
rect 4074 2044 4092 2062
rect 4510 2072 4528 2090
rect 4681 2088 4701 2108
rect 4784 2092 4804 2112
rect 4899 2088 4919 2108
rect 5002 2092 5022 2112
rect 5110 2092 5130 2112
rect 7838 2134 7858 2154
rect 7946 2134 7966 2154
rect 8049 2138 8069 2158
rect 8164 2134 8184 2154
rect 8267 2138 8287 2158
rect 8440 2156 8458 2174
rect 5213 2088 5233 2108
rect 142 1975 160 1993
rect 8438 2057 8456 2075
rect 4506 1988 4524 2006
rect 140 1876 158 1894
rect 1115 1891 1135 1911
rect 1218 1895 1238 1915
rect 1333 1891 1353 1911
rect 1436 1895 1456 1915
rect 1544 1895 1564 1915
rect 1647 1891 1667 1911
rect 2474 1899 2494 1919
rect 2577 1895 2597 1915
rect 2685 1895 2705 1915
rect 2788 1899 2808 1919
rect 2903 1895 2923 1915
rect 3006 1899 3026 1919
rect 4504 1889 4522 1907
rect 5479 1904 5499 1924
rect 135 1757 153 1775
rect 5582 1908 5602 1928
rect 5697 1904 5717 1924
rect 5800 1908 5820 1928
rect 5908 1908 5928 1928
rect 6011 1904 6031 1924
rect 6838 1912 6858 1932
rect 6941 1908 6961 1928
rect 7049 1908 7069 1928
rect 7152 1912 7172 1932
rect 7267 1908 7287 1928
rect 7370 1912 7390 1932
rect 4071 1819 4089 1837
rect 4499 1770 4517 1788
rect 8435 1832 8453 1850
rect 4069 1720 4087 1738
rect 133 1658 151 1676
rect 318 1663 338 1683
rect 421 1667 441 1687
rect 536 1663 556 1683
rect 639 1667 659 1687
rect 747 1667 767 1687
rect 850 1663 870 1683
rect 8433 1733 8451 1751
rect 4497 1671 4515 1689
rect 4682 1676 4702 1696
rect 4785 1680 4805 1700
rect 4900 1676 4920 1696
rect 5003 1680 5023 1700
rect 5111 1680 5131 1700
rect 5214 1676 5234 1696
rect 3353 1519 3373 1539
rect 3456 1515 3476 1535
rect 3564 1515 3584 1535
rect 3667 1519 3687 1539
rect 3782 1515 3802 1535
rect 3885 1519 3905 1539
rect 4072 1526 4090 1544
rect 136 1464 154 1482
rect 7717 1532 7737 1552
rect 7820 1528 7840 1548
rect 7928 1528 7948 1548
rect 8031 1532 8051 1552
rect 8146 1528 8166 1548
rect 8249 1532 8269 1552
rect 8436 1539 8454 1557
rect 4500 1477 4518 1495
rect 134 1365 152 1383
rect 4070 1427 4088 1445
rect 4498 1378 4516 1396
rect 1197 1283 1217 1303
rect 1300 1287 1320 1307
rect 1415 1283 1435 1303
rect 1518 1287 1538 1307
rect 1626 1287 1646 1307
rect 1729 1283 1749 1303
rect 2556 1291 2576 1311
rect 2659 1287 2679 1307
rect 2767 1287 2787 1307
rect 2870 1291 2890 1311
rect 2985 1287 3005 1307
rect 8434 1440 8452 1458
rect 3088 1291 3108 1311
rect 4065 1308 4083 1326
rect 5561 1296 5581 1316
rect 5664 1300 5684 1320
rect 5779 1296 5799 1316
rect 5882 1300 5902 1320
rect 5990 1300 6010 1320
rect 6093 1296 6113 1316
rect 6920 1304 6940 1324
rect 7023 1300 7043 1320
rect 7131 1300 7151 1320
rect 7234 1304 7254 1324
rect 7349 1300 7369 1320
rect 7452 1304 7472 1324
rect 8429 1321 8447 1339
rect 4063 1209 4081 1227
rect 131 1140 149 1158
rect 8427 1222 8445 1240
rect 3354 1107 3374 1127
rect 129 1041 147 1059
rect 300 1057 320 1077
rect 403 1061 423 1081
rect 518 1057 538 1077
rect 621 1061 641 1081
rect 729 1061 749 1081
rect 3457 1103 3477 1123
rect 3565 1103 3585 1123
rect 3668 1107 3688 1127
rect 3783 1103 3803 1123
rect 3886 1107 3906 1127
rect 4059 1125 4077 1143
rect 4495 1153 4513 1171
rect 832 1057 852 1077
rect 7718 1120 7738 1140
rect 4057 1026 4075 1044
rect 4493 1054 4511 1072
rect 4664 1070 4684 1090
rect 4767 1074 4787 1094
rect 4882 1070 4902 1090
rect 4985 1074 5005 1094
rect 5093 1074 5113 1094
rect 7821 1116 7841 1136
rect 7929 1116 7949 1136
rect 8032 1120 8052 1140
rect 8147 1116 8167 1136
rect 8250 1120 8270 1140
rect 8423 1138 8441 1156
rect 5196 1070 5216 1090
rect 125 957 143 975
rect 8421 1039 8439 1057
rect 4489 970 4507 988
rect 123 858 141 876
rect 1098 873 1118 893
rect 1201 877 1221 897
rect 1316 873 1336 893
rect 1419 877 1439 897
rect 1527 877 1547 897
rect 1630 873 1650 893
rect 4487 871 4505 889
rect 5462 886 5482 906
rect 118 739 136 757
rect 5565 890 5585 910
rect 5680 886 5700 906
rect 5783 890 5803 910
rect 5891 890 5911 910
rect 5994 886 6014 906
rect 4054 801 4072 819
rect 4482 752 4500 770
rect 8418 814 8436 832
rect 4052 702 4070 720
rect 116 640 134 658
rect 301 645 321 665
rect 404 649 424 669
rect 519 645 539 665
rect 622 649 642 669
rect 730 649 750 669
rect 833 645 853 665
rect 8416 715 8434 733
rect 4480 653 4498 671
rect 4665 658 4685 678
rect 4768 662 4788 682
rect 4883 658 4903 678
rect 4986 662 5006 682
rect 5094 662 5114 682
rect 5197 658 5217 678
rect 1514 69 1534 89
rect 1617 73 1637 93
rect 1732 69 1752 89
rect 1835 73 1855 93
rect 1943 73 1963 93
rect 2046 69 2066 89
rect 5878 82 5898 102
rect 5981 86 6001 106
rect 6096 82 6116 102
rect 6199 86 6219 106
rect 6307 86 6327 106
rect 6410 82 6430 102
rect 4003 -5 4023 15
rect 4106 -1 4126 19
rect 4221 -5 4241 15
rect 4324 -1 4344 19
rect 4432 -1 4452 19
rect 4535 -5 4555 15
<< pdiffc >>
rect 3486 8496 3506 8516
rect 3582 8496 3602 8516
rect 3692 8496 3712 8516
rect 3788 8496 3808 8516
rect 3910 8496 3930 8516
rect 4006 8496 4026 8516
rect 7850 8509 7870 8529
rect 7946 8509 7966 8529
rect 8056 8509 8076 8529
rect 8152 8509 8172 8529
rect 8274 8509 8294 8529
rect 8370 8509 8390 8529
rect 433 8332 453 8352
rect 529 8332 549 8352
rect 651 8332 671 8352
rect 747 8332 767 8352
rect 857 8332 877 8352
rect 953 8332 973 8352
rect 4797 8345 4817 8365
rect 2689 8268 2709 8288
rect 2785 8268 2805 8288
rect 2895 8268 2915 8288
rect 2991 8268 3011 8288
rect 3113 8268 3133 8288
rect 4893 8345 4913 8365
rect 5015 8345 5035 8365
rect 5111 8345 5131 8365
rect 5221 8345 5241 8365
rect 5317 8345 5337 8365
rect 3209 8268 3229 8288
rect 1231 8148 1251 8168
rect 1327 8148 1347 8168
rect 1449 8148 1469 8168
rect 1545 8148 1565 8168
rect 1655 8148 1675 8168
rect 1751 8148 1771 8168
rect 7053 8281 7073 8301
rect 7149 8281 7169 8301
rect 7259 8281 7279 8301
rect 7355 8281 7375 8301
rect 7477 8281 7497 8301
rect 7573 8281 7593 8301
rect 5595 8161 5615 8181
rect 3487 8084 3507 8104
rect 3583 8084 3603 8104
rect 3693 8084 3713 8104
rect 3789 8084 3809 8104
rect 3911 8084 3931 8104
rect 5691 8161 5711 8181
rect 5813 8161 5833 8181
rect 5909 8161 5929 8181
rect 6019 8161 6039 8181
rect 6115 8161 6135 8181
rect 4007 8084 4027 8104
rect 7851 8097 7871 8117
rect 7947 8097 7967 8117
rect 8057 8097 8077 8117
rect 8153 8097 8173 8117
rect 8275 8097 8295 8117
rect 8371 8097 8391 8117
rect 434 7920 454 7940
rect 530 7920 550 7940
rect 652 7920 672 7940
rect 748 7920 768 7940
rect 858 7920 878 7940
rect 954 7920 974 7940
rect 2590 7858 2610 7878
rect 2686 7858 2706 7878
rect 2796 7858 2816 7878
rect 2892 7858 2912 7878
rect 3014 7858 3034 7878
rect 4798 7933 4818 7953
rect 3110 7858 3130 7878
rect 4894 7933 4914 7953
rect 5016 7933 5036 7953
rect 5112 7933 5132 7953
rect 5222 7933 5242 7953
rect 5318 7933 5338 7953
rect 6954 7871 6974 7891
rect 7050 7871 7070 7891
rect 7160 7871 7180 7891
rect 7256 7871 7276 7891
rect 7378 7871 7398 7891
rect 7474 7871 7494 7891
rect 1313 7540 1333 7560
rect 1409 7540 1429 7560
rect 1531 7540 1551 7560
rect 1627 7540 1647 7560
rect 1737 7540 1757 7560
rect 1833 7540 1853 7560
rect 3469 7478 3489 7498
rect 3565 7478 3585 7498
rect 3675 7478 3695 7498
rect 3771 7478 3791 7498
rect 3893 7478 3913 7498
rect 5677 7553 5697 7573
rect 3989 7478 4009 7498
rect 5773 7553 5793 7573
rect 5895 7553 5915 7573
rect 5991 7553 6011 7573
rect 6101 7553 6121 7573
rect 6197 7553 6217 7573
rect 7833 7491 7853 7511
rect 7929 7491 7949 7511
rect 8039 7491 8059 7511
rect 8135 7491 8155 7511
rect 8257 7491 8277 7511
rect 8353 7491 8373 7511
rect 416 7314 436 7334
rect 512 7314 532 7334
rect 634 7314 654 7334
rect 730 7314 750 7334
rect 840 7314 860 7334
rect 936 7314 956 7334
rect 4780 7327 4800 7347
rect 2672 7250 2692 7270
rect 2768 7250 2788 7270
rect 2878 7250 2898 7270
rect 2974 7250 2994 7270
rect 3096 7250 3116 7270
rect 4876 7327 4896 7347
rect 4998 7327 5018 7347
rect 5094 7327 5114 7347
rect 5204 7327 5224 7347
rect 5300 7327 5320 7347
rect 3192 7250 3212 7270
rect 1214 7130 1234 7150
rect 1310 7130 1330 7150
rect 1432 7130 1452 7150
rect 1528 7130 1548 7150
rect 1638 7130 1658 7150
rect 1734 7130 1754 7150
rect 7036 7263 7056 7283
rect 7132 7263 7152 7283
rect 7242 7263 7262 7283
rect 7338 7263 7358 7283
rect 7460 7263 7480 7283
rect 7556 7263 7576 7283
rect 5578 7143 5598 7163
rect 3470 7066 3490 7086
rect 3566 7066 3586 7086
rect 3676 7066 3696 7086
rect 3772 7066 3792 7086
rect 3894 7066 3914 7086
rect 5674 7143 5694 7163
rect 5796 7143 5816 7163
rect 5892 7143 5912 7163
rect 6002 7143 6022 7163
rect 6098 7143 6118 7163
rect 3990 7066 4010 7086
rect 7834 7079 7854 7099
rect 7930 7079 7950 7099
rect 8040 7079 8060 7099
rect 8136 7079 8156 7099
rect 8258 7079 8278 7099
rect 8354 7079 8374 7099
rect 417 6902 437 6922
rect 513 6902 533 6922
rect 635 6902 655 6922
rect 731 6902 751 6922
rect 841 6902 861 6922
rect 937 6902 957 6922
rect 2507 6842 2527 6862
rect 2603 6842 2623 6862
rect 2713 6842 2733 6862
rect 2809 6842 2829 6862
rect 2931 6842 2951 6862
rect 4781 6915 4801 6935
rect 3027 6842 3047 6862
rect 4877 6915 4897 6935
rect 4999 6915 5019 6935
rect 5095 6915 5115 6935
rect 5205 6915 5225 6935
rect 5301 6915 5321 6935
rect 6871 6855 6891 6875
rect 6967 6855 6987 6875
rect 7077 6855 7097 6875
rect 7173 6855 7193 6875
rect 7295 6855 7315 6875
rect 7391 6855 7411 6875
rect 1359 6520 1379 6540
rect 1455 6520 1475 6540
rect 1577 6520 1597 6540
rect 1673 6520 1693 6540
rect 1783 6520 1803 6540
rect 1879 6520 1899 6540
rect 3449 6460 3469 6480
rect 3545 6460 3565 6480
rect 3655 6460 3675 6480
rect 3751 6460 3771 6480
rect 3873 6460 3893 6480
rect 5723 6533 5743 6553
rect 3969 6460 3989 6480
rect 5819 6533 5839 6553
rect 5941 6533 5961 6553
rect 6037 6533 6057 6553
rect 6147 6533 6167 6553
rect 6243 6533 6263 6553
rect 7813 6473 7833 6493
rect 7909 6473 7929 6493
rect 8019 6473 8039 6493
rect 8115 6473 8135 6493
rect 8237 6473 8257 6493
rect 8333 6473 8353 6493
rect 396 6296 416 6316
rect 492 6296 512 6316
rect 614 6296 634 6316
rect 710 6296 730 6316
rect 820 6296 840 6316
rect 916 6296 936 6316
rect 4760 6309 4780 6329
rect 2652 6232 2672 6252
rect 2748 6232 2768 6252
rect 2858 6232 2878 6252
rect 2954 6232 2974 6252
rect 3076 6232 3096 6252
rect 4856 6309 4876 6329
rect 4978 6309 4998 6329
rect 5074 6309 5094 6329
rect 5184 6309 5204 6329
rect 5280 6309 5300 6329
rect 3172 6232 3192 6252
rect 1194 6112 1214 6132
rect 1290 6112 1310 6132
rect 1412 6112 1432 6132
rect 1508 6112 1528 6132
rect 1618 6112 1638 6132
rect 1714 6112 1734 6132
rect 7016 6245 7036 6265
rect 7112 6245 7132 6265
rect 7222 6245 7242 6265
rect 7318 6245 7338 6265
rect 7440 6245 7460 6265
rect 7536 6245 7556 6265
rect 5558 6125 5578 6145
rect 3450 6048 3470 6068
rect 3546 6048 3566 6068
rect 3656 6048 3676 6068
rect 3752 6048 3772 6068
rect 3874 6048 3894 6068
rect 5654 6125 5674 6145
rect 5776 6125 5796 6145
rect 5872 6125 5892 6145
rect 5982 6125 6002 6145
rect 6078 6125 6098 6145
rect 3970 6048 3990 6068
rect 7814 6061 7834 6081
rect 7910 6061 7930 6081
rect 8020 6061 8040 6081
rect 8116 6061 8136 6081
rect 8238 6061 8258 6081
rect 8334 6061 8354 6081
rect 397 5884 417 5904
rect 493 5884 513 5904
rect 615 5884 635 5904
rect 711 5884 731 5904
rect 821 5884 841 5904
rect 917 5884 937 5904
rect 2553 5822 2573 5842
rect 2649 5822 2669 5842
rect 2759 5822 2779 5842
rect 2855 5822 2875 5842
rect 2977 5822 2997 5842
rect 4761 5897 4781 5917
rect 3073 5822 3093 5842
rect 4857 5897 4877 5917
rect 4979 5897 4999 5917
rect 5075 5897 5095 5917
rect 5185 5897 5205 5917
rect 5281 5897 5301 5917
rect 6917 5835 6937 5855
rect 7013 5835 7033 5855
rect 7123 5835 7143 5855
rect 7219 5835 7239 5855
rect 7341 5835 7361 5855
rect 7437 5835 7457 5855
rect 1276 5504 1296 5524
rect 1372 5504 1392 5524
rect 1494 5504 1514 5524
rect 1590 5504 1610 5524
rect 1700 5504 1720 5524
rect 1796 5504 1816 5524
rect 3432 5442 3452 5462
rect 3528 5442 3548 5462
rect 3638 5442 3658 5462
rect 3734 5442 3754 5462
rect 3856 5442 3876 5462
rect 5640 5517 5660 5537
rect 3952 5442 3972 5462
rect 5736 5517 5756 5537
rect 5858 5517 5878 5537
rect 5954 5517 5974 5537
rect 6064 5517 6084 5537
rect 6160 5517 6180 5537
rect 7796 5455 7816 5475
rect 7892 5455 7912 5475
rect 8002 5455 8022 5475
rect 8098 5455 8118 5475
rect 8220 5455 8240 5475
rect 8316 5455 8336 5475
rect 379 5278 399 5298
rect 475 5278 495 5298
rect 597 5278 617 5298
rect 693 5278 713 5298
rect 803 5278 823 5298
rect 899 5278 919 5298
rect 4743 5291 4763 5311
rect 2635 5214 2655 5234
rect 2731 5214 2751 5234
rect 2841 5214 2861 5234
rect 2937 5214 2957 5234
rect 3059 5214 3079 5234
rect 4839 5291 4859 5311
rect 4961 5291 4981 5311
rect 5057 5291 5077 5311
rect 5167 5291 5187 5311
rect 5263 5291 5283 5311
rect 3155 5214 3175 5234
rect 1177 5094 1197 5114
rect 1273 5094 1293 5114
rect 1395 5094 1415 5114
rect 1491 5094 1511 5114
rect 1601 5094 1621 5114
rect 1697 5094 1717 5114
rect 6999 5227 7019 5247
rect 7095 5227 7115 5247
rect 7205 5227 7225 5247
rect 7301 5227 7321 5247
rect 7423 5227 7443 5247
rect 7519 5227 7539 5247
rect 5541 5107 5561 5127
rect 3433 5030 3453 5050
rect 3529 5030 3549 5050
rect 3639 5030 3659 5050
rect 3735 5030 3755 5050
rect 3857 5030 3877 5050
rect 5637 5107 5657 5127
rect 5759 5107 5779 5127
rect 5855 5107 5875 5127
rect 5965 5107 5985 5127
rect 6061 5107 6081 5127
rect 3953 5030 3973 5050
rect 7797 5043 7817 5063
rect 7893 5043 7913 5063
rect 8003 5043 8023 5063
rect 8099 5043 8119 5063
rect 8221 5043 8241 5063
rect 8317 5043 8337 5063
rect 380 4866 400 4886
rect 476 4866 496 4886
rect 598 4866 618 4886
rect 694 4866 714 4886
rect 804 4866 824 4886
rect 900 4866 920 4886
rect 2331 4808 2351 4828
rect 2427 4808 2447 4828
rect 2537 4808 2557 4828
rect 2633 4808 2653 4828
rect 2755 4808 2775 4828
rect 4744 4879 4764 4899
rect 2851 4808 2871 4828
rect 4840 4879 4860 4899
rect 4962 4879 4982 4899
rect 5058 4879 5078 4899
rect 5168 4879 5188 4899
rect 5264 4879 5284 4899
rect 6695 4821 6715 4841
rect 6791 4821 6811 4841
rect 6901 4821 6921 4841
rect 6997 4821 7017 4841
rect 7119 4821 7139 4841
rect 7215 4821 7235 4841
rect 1462 4482 1482 4502
rect 1558 4482 1578 4502
rect 1680 4482 1700 4502
rect 1776 4482 1796 4502
rect 1886 4482 1906 4502
rect 1982 4482 2002 4502
rect 3413 4424 3433 4444
rect 3509 4424 3529 4444
rect 3619 4424 3639 4444
rect 3715 4424 3735 4444
rect 3837 4424 3857 4444
rect 5826 4495 5846 4515
rect 3933 4424 3953 4444
rect 5922 4495 5942 4515
rect 6044 4495 6064 4515
rect 6140 4495 6160 4515
rect 6250 4495 6270 4515
rect 6346 4495 6366 4515
rect 7777 4437 7797 4457
rect 7873 4437 7893 4457
rect 7983 4437 8003 4457
rect 8079 4437 8099 4457
rect 8201 4437 8221 4457
rect 8297 4437 8317 4457
rect 360 4260 380 4280
rect 456 4260 476 4280
rect 578 4260 598 4280
rect 674 4260 694 4280
rect 784 4260 804 4280
rect 880 4260 900 4280
rect 4724 4273 4744 4293
rect 2616 4196 2636 4216
rect 2712 4196 2732 4216
rect 2822 4196 2842 4216
rect 2918 4196 2938 4216
rect 3040 4196 3060 4216
rect 4820 4273 4840 4293
rect 4942 4273 4962 4293
rect 5038 4273 5058 4293
rect 5148 4273 5168 4293
rect 5244 4273 5264 4293
rect 3136 4196 3156 4216
rect 1158 4076 1178 4096
rect 1254 4076 1274 4096
rect 1376 4076 1396 4096
rect 1472 4076 1492 4096
rect 1582 4076 1602 4096
rect 1678 4076 1698 4096
rect 6980 4209 7000 4229
rect 7076 4209 7096 4229
rect 7186 4209 7206 4229
rect 7282 4209 7302 4229
rect 7404 4209 7424 4229
rect 7500 4209 7520 4229
rect 5522 4089 5542 4109
rect 3414 4012 3434 4032
rect 3510 4012 3530 4032
rect 3620 4012 3640 4032
rect 3716 4012 3736 4032
rect 3838 4012 3858 4032
rect 5618 4089 5638 4109
rect 5740 4089 5760 4109
rect 5836 4089 5856 4109
rect 5946 4089 5966 4109
rect 6042 4089 6062 4109
rect 3934 4012 3954 4032
rect 7778 4025 7798 4045
rect 7874 4025 7894 4045
rect 7984 4025 8004 4045
rect 8080 4025 8100 4045
rect 8202 4025 8222 4045
rect 8298 4025 8318 4045
rect 361 3848 381 3868
rect 457 3848 477 3868
rect 579 3848 599 3868
rect 675 3848 695 3868
rect 785 3848 805 3868
rect 881 3848 901 3868
rect 2517 3786 2537 3806
rect 2613 3786 2633 3806
rect 2723 3786 2743 3806
rect 2819 3786 2839 3806
rect 2941 3786 2961 3806
rect 4725 3861 4745 3881
rect 3037 3786 3057 3806
rect 4821 3861 4841 3881
rect 4943 3861 4963 3881
rect 5039 3861 5059 3881
rect 5149 3861 5169 3881
rect 5245 3861 5265 3881
rect 6881 3799 6901 3819
rect 6977 3799 6997 3819
rect 7087 3799 7107 3819
rect 7183 3799 7203 3819
rect 7305 3799 7325 3819
rect 7401 3799 7421 3819
rect 1240 3468 1260 3488
rect 1336 3468 1356 3488
rect 1458 3468 1478 3488
rect 1554 3468 1574 3488
rect 1664 3468 1684 3488
rect 1760 3468 1780 3488
rect 3396 3406 3416 3426
rect 3492 3406 3512 3426
rect 3602 3406 3622 3426
rect 3698 3406 3718 3426
rect 3820 3406 3840 3426
rect 5604 3481 5624 3501
rect 3916 3406 3936 3426
rect 5700 3481 5720 3501
rect 5822 3481 5842 3501
rect 5918 3481 5938 3501
rect 6028 3481 6048 3501
rect 6124 3481 6144 3501
rect 7760 3419 7780 3439
rect 7856 3419 7876 3439
rect 7966 3419 7986 3439
rect 8062 3419 8082 3439
rect 8184 3419 8204 3439
rect 8280 3419 8300 3439
rect 343 3242 363 3262
rect 439 3242 459 3262
rect 561 3242 581 3262
rect 657 3242 677 3262
rect 767 3242 787 3262
rect 863 3242 883 3262
rect 4707 3255 4727 3275
rect 2599 3178 2619 3198
rect 2695 3178 2715 3198
rect 2805 3178 2825 3198
rect 2901 3178 2921 3198
rect 3023 3178 3043 3198
rect 4803 3255 4823 3275
rect 4925 3255 4945 3275
rect 5021 3255 5041 3275
rect 5131 3255 5151 3275
rect 5227 3255 5247 3275
rect 3119 3178 3139 3198
rect 1141 3058 1161 3078
rect 1237 3058 1257 3078
rect 1359 3058 1379 3078
rect 1455 3058 1475 3078
rect 1565 3058 1585 3078
rect 1661 3058 1681 3078
rect 6963 3191 6983 3211
rect 7059 3191 7079 3211
rect 7169 3191 7189 3211
rect 7265 3191 7285 3211
rect 7387 3191 7407 3211
rect 7483 3191 7503 3211
rect 5505 3071 5525 3091
rect 3397 2994 3417 3014
rect 3493 2994 3513 3014
rect 3603 2994 3623 3014
rect 3699 2994 3719 3014
rect 3821 2994 3841 3014
rect 5601 3071 5621 3091
rect 5723 3071 5743 3091
rect 5819 3071 5839 3091
rect 5929 3071 5949 3091
rect 6025 3071 6045 3091
rect 3917 2994 3937 3014
rect 7761 3007 7781 3027
rect 7857 3007 7877 3027
rect 7967 3007 7987 3027
rect 8063 3007 8083 3027
rect 8185 3007 8205 3027
rect 8281 3007 8301 3027
rect 344 2830 364 2850
rect 440 2830 460 2850
rect 562 2830 582 2850
rect 658 2830 678 2850
rect 768 2830 788 2850
rect 864 2830 884 2850
rect 2434 2770 2454 2790
rect 2530 2770 2550 2790
rect 2640 2770 2660 2790
rect 2736 2770 2756 2790
rect 2858 2770 2878 2790
rect 4708 2843 4728 2863
rect 2954 2770 2974 2790
rect 4804 2843 4824 2863
rect 4926 2843 4946 2863
rect 5022 2843 5042 2863
rect 5132 2843 5152 2863
rect 5228 2843 5248 2863
rect 6798 2783 6818 2803
rect 6894 2783 6914 2803
rect 7004 2783 7024 2803
rect 7100 2783 7120 2803
rect 7222 2783 7242 2803
rect 7318 2783 7338 2803
rect 1286 2448 1306 2468
rect 1382 2448 1402 2468
rect 1504 2448 1524 2468
rect 1600 2448 1620 2468
rect 1710 2448 1730 2468
rect 1806 2448 1826 2468
rect 3376 2388 3396 2408
rect 3472 2388 3492 2408
rect 3582 2388 3602 2408
rect 3678 2388 3698 2408
rect 3800 2388 3820 2408
rect 5650 2461 5670 2481
rect 3896 2388 3916 2408
rect 5746 2461 5766 2481
rect 5868 2461 5888 2481
rect 5964 2461 5984 2481
rect 6074 2461 6094 2481
rect 6170 2461 6190 2481
rect 7740 2401 7760 2421
rect 7836 2401 7856 2421
rect 7946 2401 7966 2421
rect 8042 2401 8062 2421
rect 8164 2401 8184 2421
rect 8260 2401 8280 2421
rect 323 2224 343 2244
rect 419 2224 439 2244
rect 541 2224 561 2244
rect 637 2224 657 2244
rect 747 2224 767 2244
rect 843 2224 863 2244
rect 4687 2237 4707 2257
rect 2579 2160 2599 2180
rect 2675 2160 2695 2180
rect 2785 2160 2805 2180
rect 2881 2160 2901 2180
rect 3003 2160 3023 2180
rect 4783 2237 4803 2257
rect 4905 2237 4925 2257
rect 5001 2237 5021 2257
rect 5111 2237 5131 2257
rect 5207 2237 5227 2257
rect 3099 2160 3119 2180
rect 1121 2040 1141 2060
rect 1217 2040 1237 2060
rect 1339 2040 1359 2060
rect 1435 2040 1455 2060
rect 1545 2040 1565 2060
rect 1641 2040 1661 2060
rect 6943 2173 6963 2193
rect 7039 2173 7059 2193
rect 7149 2173 7169 2193
rect 7245 2173 7265 2193
rect 7367 2173 7387 2193
rect 7463 2173 7483 2193
rect 5485 2053 5505 2073
rect 3377 1976 3397 1996
rect 3473 1976 3493 1996
rect 3583 1976 3603 1996
rect 3679 1976 3699 1996
rect 3801 1976 3821 1996
rect 5581 2053 5601 2073
rect 5703 2053 5723 2073
rect 5799 2053 5819 2073
rect 5909 2053 5929 2073
rect 6005 2053 6025 2073
rect 3897 1976 3917 1996
rect 7741 1989 7761 2009
rect 7837 1989 7857 2009
rect 7947 1989 7967 2009
rect 8043 1989 8063 2009
rect 8165 1989 8185 2009
rect 8261 1989 8281 2009
rect 324 1812 344 1832
rect 420 1812 440 1832
rect 542 1812 562 1832
rect 638 1812 658 1832
rect 748 1812 768 1832
rect 844 1812 864 1832
rect 2480 1750 2500 1770
rect 2576 1750 2596 1770
rect 2686 1750 2706 1770
rect 2782 1750 2802 1770
rect 2904 1750 2924 1770
rect 4688 1825 4708 1845
rect 3000 1750 3020 1770
rect 4784 1825 4804 1845
rect 4906 1825 4926 1845
rect 5002 1825 5022 1845
rect 5112 1825 5132 1845
rect 5208 1825 5228 1845
rect 6844 1763 6864 1783
rect 6940 1763 6960 1783
rect 7050 1763 7070 1783
rect 7146 1763 7166 1783
rect 7268 1763 7288 1783
rect 7364 1763 7384 1783
rect 1203 1432 1223 1452
rect 1299 1432 1319 1452
rect 1421 1432 1441 1452
rect 1517 1432 1537 1452
rect 1627 1432 1647 1452
rect 1723 1432 1743 1452
rect 3359 1370 3379 1390
rect 3455 1370 3475 1390
rect 3565 1370 3585 1390
rect 3661 1370 3681 1390
rect 3783 1370 3803 1390
rect 5567 1445 5587 1465
rect 3879 1370 3899 1390
rect 5663 1445 5683 1465
rect 5785 1445 5805 1465
rect 5881 1445 5901 1465
rect 5991 1445 6011 1465
rect 6087 1445 6107 1465
rect 7723 1383 7743 1403
rect 7819 1383 7839 1403
rect 7929 1383 7949 1403
rect 8025 1383 8045 1403
rect 8147 1383 8167 1403
rect 8243 1383 8263 1403
rect 306 1206 326 1226
rect 402 1206 422 1226
rect 524 1206 544 1226
rect 620 1206 640 1226
rect 730 1206 750 1226
rect 826 1206 846 1226
rect 4670 1219 4690 1239
rect 2562 1142 2582 1162
rect 2658 1142 2678 1162
rect 2768 1142 2788 1162
rect 2864 1142 2884 1162
rect 2986 1142 3006 1162
rect 4766 1219 4786 1239
rect 4888 1219 4908 1239
rect 4984 1219 5004 1239
rect 5094 1219 5114 1239
rect 5190 1219 5210 1239
rect 3082 1142 3102 1162
rect 1104 1022 1124 1042
rect 1200 1022 1220 1042
rect 1322 1022 1342 1042
rect 1418 1022 1438 1042
rect 1528 1022 1548 1042
rect 1624 1022 1644 1042
rect 6926 1155 6946 1175
rect 7022 1155 7042 1175
rect 7132 1155 7152 1175
rect 7228 1155 7248 1175
rect 7350 1155 7370 1175
rect 7446 1155 7466 1175
rect 5468 1035 5488 1055
rect 3360 958 3380 978
rect 3456 958 3476 978
rect 3566 958 3586 978
rect 3662 958 3682 978
rect 3784 958 3804 978
rect 5564 1035 5584 1055
rect 5686 1035 5706 1055
rect 5782 1035 5802 1055
rect 5892 1035 5912 1055
rect 5988 1035 6008 1055
rect 3880 958 3900 978
rect 7724 971 7744 991
rect 7820 971 7840 991
rect 7930 971 7950 991
rect 8026 971 8046 991
rect 8148 971 8168 991
rect 8244 971 8264 991
rect 307 794 327 814
rect 403 794 423 814
rect 525 794 545 814
rect 621 794 641 814
rect 731 794 751 814
rect 827 794 847 814
rect 4671 807 4691 827
rect 4767 807 4787 827
rect 4889 807 4909 827
rect 4985 807 5005 827
rect 5095 807 5115 827
rect 5191 807 5211 827
rect 1520 218 1540 238
rect 1616 218 1636 238
rect 1738 218 1758 238
rect 1834 218 1854 238
rect 1944 218 1964 238
rect 2040 218 2060 238
rect 5884 231 5904 251
rect 4009 144 4029 164
rect 4105 144 4125 164
rect 4227 144 4247 164
rect 4323 144 4343 164
rect 4433 144 4453 164
rect 5980 231 6000 251
rect 6102 231 6122 251
rect 6198 231 6218 251
rect 6308 231 6328 251
rect 6404 231 6424 251
rect 4529 144 4549 164
<< poly >>
rect 3518 8677 3568 8693
rect 3726 8677 3776 8693
rect 3944 8677 3994 8693
rect 7882 8690 7932 8706
rect 8090 8690 8140 8706
rect 8308 8690 8358 8706
rect 3518 8605 3568 8635
rect 3518 8585 3525 8605
rect 3545 8585 3568 8605
rect 3518 8558 3568 8585
rect 3726 8603 3776 8635
rect 3726 8583 3743 8603
rect 3763 8583 3776 8603
rect 3726 8558 3776 8583
rect 3944 8606 3994 8635
rect 3944 8586 3961 8606
rect 3981 8586 3994 8606
rect 3944 8558 3994 8586
rect 7882 8618 7932 8648
rect 7882 8598 7889 8618
rect 7909 8598 7932 8618
rect 2721 8449 2771 8465
rect 2929 8449 2979 8465
rect 3147 8449 3197 8465
rect 7882 8571 7932 8598
rect 8090 8616 8140 8648
rect 8090 8596 8107 8616
rect 8127 8596 8140 8616
rect 8090 8571 8140 8596
rect 8308 8619 8358 8648
rect 8308 8599 8325 8619
rect 8345 8599 8358 8619
rect 8308 8571 8358 8599
rect 3518 8445 3568 8458
rect 3726 8445 3776 8458
rect 3944 8445 3994 8458
rect 7085 8462 7135 8478
rect 7293 8462 7343 8478
rect 7511 8462 7561 8478
rect 7882 8458 7932 8471
rect 8090 8458 8140 8471
rect 8308 8458 8358 8471
rect 465 8390 515 8403
rect 683 8390 733 8403
rect 891 8390 941 8403
rect 2721 8377 2771 8407
rect 2721 8357 2728 8377
rect 2748 8357 2771 8377
rect 2721 8330 2771 8357
rect 2929 8375 2979 8407
rect 2929 8355 2946 8375
rect 2966 8355 2979 8375
rect 2929 8330 2979 8355
rect 3147 8378 3197 8407
rect 3147 8358 3164 8378
rect 3184 8358 3197 8378
rect 4829 8403 4879 8416
rect 5047 8403 5097 8416
rect 5255 8403 5305 8416
rect 3147 8330 3197 8358
rect 465 8262 515 8290
rect 465 8242 478 8262
rect 498 8242 515 8262
rect 465 8213 515 8242
rect 683 8265 733 8290
rect 683 8245 696 8265
rect 716 8245 733 8265
rect 683 8213 733 8245
rect 891 8263 941 8290
rect 891 8243 914 8263
rect 934 8243 941 8263
rect 891 8213 941 8243
rect 7085 8390 7135 8420
rect 7085 8370 7092 8390
rect 7112 8370 7135 8390
rect 7085 8343 7135 8370
rect 7293 8388 7343 8420
rect 7293 8368 7310 8388
rect 7330 8368 7343 8388
rect 7293 8343 7343 8368
rect 7511 8391 7561 8420
rect 7511 8371 7528 8391
rect 7548 8371 7561 8391
rect 7511 8343 7561 8371
rect 3519 8265 3569 8281
rect 3727 8265 3777 8281
rect 3945 8265 3995 8281
rect 1263 8206 1313 8219
rect 1481 8206 1531 8219
rect 1689 8206 1739 8219
rect 2721 8217 2771 8230
rect 2929 8217 2979 8230
rect 3147 8217 3197 8230
rect 4829 8275 4879 8303
rect 465 8155 515 8171
rect 683 8155 733 8171
rect 891 8155 941 8171
rect 3519 8193 3569 8223
rect 3519 8173 3526 8193
rect 3546 8173 3569 8193
rect 3519 8146 3569 8173
rect 3727 8191 3777 8223
rect 3727 8171 3744 8191
rect 3764 8171 3777 8191
rect 3727 8146 3777 8171
rect 3945 8194 3995 8223
rect 3945 8174 3962 8194
rect 3982 8174 3995 8194
rect 4829 8255 4842 8275
rect 4862 8255 4879 8275
rect 4829 8226 4879 8255
rect 5047 8278 5097 8303
rect 5047 8258 5060 8278
rect 5080 8258 5097 8278
rect 5047 8226 5097 8258
rect 5255 8276 5305 8303
rect 5255 8256 5278 8276
rect 5298 8256 5305 8276
rect 5255 8226 5305 8256
rect 7883 8278 7933 8294
rect 8091 8278 8141 8294
rect 8309 8278 8359 8294
rect 3945 8146 3995 8174
rect 5627 8219 5677 8232
rect 5845 8219 5895 8232
rect 6053 8219 6103 8232
rect 7085 8230 7135 8243
rect 7293 8230 7343 8243
rect 7511 8230 7561 8243
rect 4829 8168 4879 8184
rect 5047 8168 5097 8184
rect 5255 8168 5305 8184
rect 1263 8078 1313 8106
rect 1263 8058 1276 8078
rect 1296 8058 1313 8078
rect 1263 8029 1313 8058
rect 1481 8081 1531 8106
rect 1481 8061 1494 8081
rect 1514 8061 1531 8081
rect 1481 8029 1531 8061
rect 1689 8079 1739 8106
rect 1689 8059 1712 8079
rect 1732 8059 1739 8079
rect 1689 8029 1739 8059
rect 2622 8039 2672 8055
rect 2830 8039 2880 8055
rect 3048 8039 3098 8055
rect 7883 8206 7933 8236
rect 7883 8186 7890 8206
rect 7910 8186 7933 8206
rect 7883 8159 7933 8186
rect 8091 8204 8141 8236
rect 8091 8184 8108 8204
rect 8128 8184 8141 8204
rect 8091 8159 8141 8184
rect 8309 8207 8359 8236
rect 8309 8187 8326 8207
rect 8346 8187 8359 8207
rect 8309 8159 8359 8187
rect 5627 8091 5677 8119
rect 466 7978 516 7991
rect 684 7978 734 7991
rect 892 7978 942 7991
rect 3519 8033 3569 8046
rect 3727 8033 3777 8046
rect 3945 8033 3995 8046
rect 5627 8071 5640 8091
rect 5660 8071 5677 8091
rect 5627 8042 5677 8071
rect 5845 8094 5895 8119
rect 5845 8074 5858 8094
rect 5878 8074 5895 8094
rect 5845 8042 5895 8074
rect 6053 8092 6103 8119
rect 6053 8072 6076 8092
rect 6096 8072 6103 8092
rect 6053 8042 6103 8072
rect 6986 8052 7036 8068
rect 7194 8052 7244 8068
rect 7412 8052 7462 8068
rect 1263 7971 1313 7987
rect 1481 7971 1531 7987
rect 1689 7971 1739 7987
rect 2622 7967 2672 7997
rect 2622 7947 2629 7967
rect 2649 7947 2672 7967
rect 2622 7920 2672 7947
rect 2830 7965 2880 7997
rect 2830 7945 2847 7965
rect 2867 7945 2880 7965
rect 2830 7920 2880 7945
rect 3048 7968 3098 7997
rect 4830 7991 4880 8004
rect 5048 7991 5098 8004
rect 5256 7991 5306 8004
rect 7883 8046 7933 8059
rect 8091 8046 8141 8059
rect 8309 8046 8359 8059
rect 3048 7948 3065 7968
rect 3085 7948 3098 7968
rect 3048 7920 3098 7948
rect 466 7850 516 7878
rect 466 7830 479 7850
rect 499 7830 516 7850
rect 466 7801 516 7830
rect 684 7853 734 7878
rect 684 7833 697 7853
rect 717 7833 734 7853
rect 684 7801 734 7833
rect 892 7851 942 7878
rect 892 7831 915 7851
rect 935 7831 942 7851
rect 892 7801 942 7831
rect 5627 7984 5677 8000
rect 5845 7984 5895 8000
rect 6053 7984 6103 8000
rect 6986 7980 7036 8010
rect 6986 7960 6993 7980
rect 7013 7960 7036 7980
rect 6986 7933 7036 7960
rect 7194 7978 7244 8010
rect 7194 7958 7211 7978
rect 7231 7958 7244 7978
rect 7194 7933 7244 7958
rect 7412 7981 7462 8010
rect 7412 7961 7429 7981
rect 7449 7961 7462 7981
rect 7412 7933 7462 7961
rect 4830 7863 4880 7891
rect 2622 7807 2672 7820
rect 2830 7807 2880 7820
rect 3048 7807 3098 7820
rect 4830 7843 4843 7863
rect 4863 7843 4880 7863
rect 4830 7814 4880 7843
rect 5048 7866 5098 7891
rect 5048 7846 5061 7866
rect 5081 7846 5098 7866
rect 5048 7814 5098 7846
rect 5256 7864 5306 7891
rect 5256 7844 5279 7864
rect 5299 7844 5306 7864
rect 5256 7814 5306 7844
rect 6986 7820 7036 7833
rect 7194 7820 7244 7833
rect 7412 7820 7462 7833
rect 466 7743 516 7759
rect 684 7743 734 7759
rect 892 7743 942 7759
rect 4830 7756 4880 7772
rect 5048 7756 5098 7772
rect 5256 7756 5306 7772
rect 3501 7659 3551 7675
rect 3709 7659 3759 7675
rect 3927 7659 3977 7675
rect 7865 7672 7915 7688
rect 8073 7672 8123 7688
rect 8291 7672 8341 7688
rect 1345 7598 1395 7611
rect 1563 7598 1613 7611
rect 1771 7598 1821 7611
rect 3501 7587 3551 7617
rect 3501 7567 3508 7587
rect 3528 7567 3551 7587
rect 3501 7540 3551 7567
rect 3709 7585 3759 7617
rect 3709 7565 3726 7585
rect 3746 7565 3759 7585
rect 3709 7540 3759 7565
rect 3927 7588 3977 7617
rect 3927 7568 3944 7588
rect 3964 7568 3977 7588
rect 5709 7611 5759 7624
rect 5927 7611 5977 7624
rect 6135 7611 6185 7624
rect 3927 7540 3977 7568
rect 1345 7470 1395 7498
rect 1345 7450 1358 7470
rect 1378 7450 1395 7470
rect 1345 7421 1395 7450
rect 1563 7473 1613 7498
rect 1563 7453 1576 7473
rect 1596 7453 1613 7473
rect 1563 7421 1613 7453
rect 1771 7471 1821 7498
rect 1771 7451 1794 7471
rect 1814 7451 1821 7471
rect 1771 7421 1821 7451
rect 2704 7431 2754 7447
rect 2912 7431 2962 7447
rect 3130 7431 3180 7447
rect 7865 7600 7915 7630
rect 7865 7580 7872 7600
rect 7892 7580 7915 7600
rect 7865 7553 7915 7580
rect 8073 7598 8123 7630
rect 8073 7578 8090 7598
rect 8110 7578 8123 7598
rect 8073 7553 8123 7578
rect 8291 7601 8341 7630
rect 8291 7581 8308 7601
rect 8328 7581 8341 7601
rect 8291 7553 8341 7581
rect 5709 7483 5759 7511
rect 5709 7463 5722 7483
rect 5742 7463 5759 7483
rect 448 7372 498 7385
rect 666 7372 716 7385
rect 874 7372 924 7385
rect 3501 7427 3551 7440
rect 3709 7427 3759 7440
rect 3927 7427 3977 7440
rect 5709 7434 5759 7463
rect 5927 7486 5977 7511
rect 5927 7466 5940 7486
rect 5960 7466 5977 7486
rect 5927 7434 5977 7466
rect 6135 7484 6185 7511
rect 6135 7464 6158 7484
rect 6178 7464 6185 7484
rect 6135 7434 6185 7464
rect 7068 7444 7118 7460
rect 7276 7444 7326 7460
rect 7494 7444 7544 7460
rect 1345 7363 1395 7379
rect 1563 7363 1613 7379
rect 1771 7363 1821 7379
rect 2704 7359 2754 7389
rect 2704 7339 2711 7359
rect 2731 7339 2754 7359
rect 2704 7312 2754 7339
rect 2912 7357 2962 7389
rect 2912 7337 2929 7357
rect 2949 7337 2962 7357
rect 2912 7312 2962 7337
rect 3130 7360 3180 7389
rect 3130 7340 3147 7360
rect 3167 7340 3180 7360
rect 4812 7385 4862 7398
rect 5030 7385 5080 7398
rect 5238 7385 5288 7398
rect 7865 7440 7915 7453
rect 8073 7440 8123 7453
rect 8291 7440 8341 7453
rect 3130 7312 3180 7340
rect 448 7244 498 7272
rect 448 7224 461 7244
rect 481 7224 498 7244
rect 448 7195 498 7224
rect 666 7247 716 7272
rect 666 7227 679 7247
rect 699 7227 716 7247
rect 666 7195 716 7227
rect 874 7245 924 7272
rect 874 7225 897 7245
rect 917 7225 924 7245
rect 874 7195 924 7225
rect 5709 7376 5759 7392
rect 5927 7376 5977 7392
rect 6135 7376 6185 7392
rect 7068 7372 7118 7402
rect 7068 7352 7075 7372
rect 7095 7352 7118 7372
rect 7068 7325 7118 7352
rect 7276 7370 7326 7402
rect 7276 7350 7293 7370
rect 7313 7350 7326 7370
rect 7276 7325 7326 7350
rect 7494 7373 7544 7402
rect 7494 7353 7511 7373
rect 7531 7353 7544 7373
rect 7494 7325 7544 7353
rect 3502 7247 3552 7263
rect 3710 7247 3760 7263
rect 3928 7247 3978 7263
rect 1246 7188 1296 7201
rect 1464 7188 1514 7201
rect 1672 7188 1722 7201
rect 2704 7199 2754 7212
rect 2912 7199 2962 7212
rect 3130 7199 3180 7212
rect 4812 7257 4862 7285
rect 448 7137 498 7153
rect 666 7137 716 7153
rect 874 7137 924 7153
rect 3502 7175 3552 7205
rect 3502 7155 3509 7175
rect 3529 7155 3552 7175
rect 3502 7128 3552 7155
rect 3710 7173 3760 7205
rect 3710 7153 3727 7173
rect 3747 7153 3760 7173
rect 3710 7128 3760 7153
rect 3928 7176 3978 7205
rect 3928 7156 3945 7176
rect 3965 7156 3978 7176
rect 4812 7237 4825 7257
rect 4845 7237 4862 7257
rect 4812 7208 4862 7237
rect 5030 7260 5080 7285
rect 5030 7240 5043 7260
rect 5063 7240 5080 7260
rect 5030 7208 5080 7240
rect 5238 7258 5288 7285
rect 5238 7238 5261 7258
rect 5281 7238 5288 7258
rect 5238 7208 5288 7238
rect 7866 7260 7916 7276
rect 8074 7260 8124 7276
rect 8292 7260 8342 7276
rect 3928 7128 3978 7156
rect 5610 7201 5660 7214
rect 5828 7201 5878 7214
rect 6036 7201 6086 7214
rect 7068 7212 7118 7225
rect 7276 7212 7326 7225
rect 7494 7212 7544 7225
rect 4812 7150 4862 7166
rect 5030 7150 5080 7166
rect 5238 7150 5288 7166
rect 1246 7060 1296 7088
rect 1246 7040 1259 7060
rect 1279 7040 1296 7060
rect 1246 7011 1296 7040
rect 1464 7063 1514 7088
rect 1464 7043 1477 7063
rect 1497 7043 1514 7063
rect 1464 7011 1514 7043
rect 1672 7061 1722 7088
rect 1672 7041 1695 7061
rect 1715 7041 1722 7061
rect 1672 7011 1722 7041
rect 2539 7023 2589 7039
rect 2747 7023 2797 7039
rect 2965 7023 3015 7039
rect 7866 7188 7916 7218
rect 7866 7168 7873 7188
rect 7893 7168 7916 7188
rect 7866 7141 7916 7168
rect 8074 7186 8124 7218
rect 8074 7166 8091 7186
rect 8111 7166 8124 7186
rect 8074 7141 8124 7166
rect 8292 7189 8342 7218
rect 8292 7169 8309 7189
rect 8329 7169 8342 7189
rect 8292 7141 8342 7169
rect 5610 7073 5660 7101
rect 449 6960 499 6973
rect 667 6960 717 6973
rect 875 6960 925 6973
rect 3502 7015 3552 7028
rect 3710 7015 3760 7028
rect 3928 7015 3978 7028
rect 5610 7053 5623 7073
rect 5643 7053 5660 7073
rect 5610 7024 5660 7053
rect 5828 7076 5878 7101
rect 5828 7056 5841 7076
rect 5861 7056 5878 7076
rect 5828 7024 5878 7056
rect 6036 7074 6086 7101
rect 6036 7054 6059 7074
rect 6079 7054 6086 7074
rect 6036 7024 6086 7054
rect 6903 7036 6953 7052
rect 7111 7036 7161 7052
rect 7329 7036 7379 7052
rect 1246 6953 1296 6969
rect 1464 6953 1514 6969
rect 1672 6953 1722 6969
rect 2539 6951 2589 6981
rect 2539 6931 2546 6951
rect 2566 6931 2589 6951
rect 2539 6904 2589 6931
rect 2747 6949 2797 6981
rect 2747 6929 2764 6949
rect 2784 6929 2797 6949
rect 2747 6904 2797 6929
rect 2965 6952 3015 6981
rect 4813 6973 4863 6986
rect 5031 6973 5081 6986
rect 5239 6973 5289 6986
rect 7866 7028 7916 7041
rect 8074 7028 8124 7041
rect 8292 7028 8342 7041
rect 2965 6932 2982 6952
rect 3002 6932 3015 6952
rect 2965 6904 3015 6932
rect 449 6832 499 6860
rect 449 6812 462 6832
rect 482 6812 499 6832
rect 449 6783 499 6812
rect 667 6835 717 6860
rect 667 6815 680 6835
rect 700 6815 717 6835
rect 667 6783 717 6815
rect 875 6833 925 6860
rect 875 6813 898 6833
rect 918 6813 925 6833
rect 875 6783 925 6813
rect 5610 6966 5660 6982
rect 5828 6966 5878 6982
rect 6036 6966 6086 6982
rect 6903 6964 6953 6994
rect 6903 6944 6910 6964
rect 6930 6944 6953 6964
rect 6903 6917 6953 6944
rect 7111 6962 7161 6994
rect 7111 6942 7128 6962
rect 7148 6942 7161 6962
rect 7111 6917 7161 6942
rect 7329 6965 7379 6994
rect 7329 6945 7346 6965
rect 7366 6945 7379 6965
rect 7329 6917 7379 6945
rect 4813 6845 4863 6873
rect 2539 6791 2589 6804
rect 2747 6791 2797 6804
rect 2965 6791 3015 6804
rect 4813 6825 4826 6845
rect 4846 6825 4863 6845
rect 4813 6796 4863 6825
rect 5031 6848 5081 6873
rect 5031 6828 5044 6848
rect 5064 6828 5081 6848
rect 5031 6796 5081 6828
rect 5239 6846 5289 6873
rect 5239 6826 5262 6846
rect 5282 6826 5289 6846
rect 5239 6796 5289 6826
rect 6903 6804 6953 6817
rect 7111 6804 7161 6817
rect 7329 6804 7379 6817
rect 449 6725 499 6741
rect 667 6725 717 6741
rect 875 6725 925 6741
rect 4813 6738 4863 6754
rect 5031 6738 5081 6754
rect 5239 6738 5289 6754
rect 3481 6641 3531 6657
rect 3689 6641 3739 6657
rect 3907 6641 3957 6657
rect 7845 6654 7895 6670
rect 8053 6654 8103 6670
rect 8271 6654 8321 6670
rect 1391 6578 1441 6591
rect 1609 6578 1659 6591
rect 1817 6578 1867 6591
rect 3481 6569 3531 6599
rect 3481 6549 3488 6569
rect 3508 6549 3531 6569
rect 3481 6522 3531 6549
rect 3689 6567 3739 6599
rect 3689 6547 3706 6567
rect 3726 6547 3739 6567
rect 3689 6522 3739 6547
rect 3907 6570 3957 6599
rect 3907 6550 3924 6570
rect 3944 6550 3957 6570
rect 5755 6591 5805 6604
rect 5973 6591 6023 6604
rect 6181 6591 6231 6604
rect 3907 6522 3957 6550
rect 1391 6450 1441 6478
rect 1391 6430 1404 6450
rect 1424 6430 1441 6450
rect 1391 6401 1441 6430
rect 1609 6453 1659 6478
rect 1609 6433 1622 6453
rect 1642 6433 1659 6453
rect 1609 6401 1659 6433
rect 1817 6451 1867 6478
rect 1817 6431 1840 6451
rect 1860 6431 1867 6451
rect 1817 6401 1867 6431
rect 2684 6413 2734 6429
rect 2892 6413 2942 6429
rect 3110 6413 3160 6429
rect 7845 6582 7895 6612
rect 7845 6562 7852 6582
rect 7872 6562 7895 6582
rect 7845 6535 7895 6562
rect 8053 6580 8103 6612
rect 8053 6560 8070 6580
rect 8090 6560 8103 6580
rect 8053 6535 8103 6560
rect 8271 6583 8321 6612
rect 8271 6563 8288 6583
rect 8308 6563 8321 6583
rect 8271 6535 8321 6563
rect 5755 6463 5805 6491
rect 5755 6443 5768 6463
rect 5788 6443 5805 6463
rect 428 6354 478 6367
rect 646 6354 696 6367
rect 854 6354 904 6367
rect 3481 6409 3531 6422
rect 3689 6409 3739 6422
rect 3907 6409 3957 6422
rect 5755 6414 5805 6443
rect 5973 6466 6023 6491
rect 5973 6446 5986 6466
rect 6006 6446 6023 6466
rect 5973 6414 6023 6446
rect 6181 6464 6231 6491
rect 6181 6444 6204 6464
rect 6224 6444 6231 6464
rect 6181 6414 6231 6444
rect 7048 6426 7098 6442
rect 7256 6426 7306 6442
rect 7474 6426 7524 6442
rect 1391 6343 1441 6359
rect 1609 6343 1659 6359
rect 1817 6343 1867 6359
rect 2684 6341 2734 6371
rect 2684 6321 2691 6341
rect 2711 6321 2734 6341
rect 2684 6294 2734 6321
rect 2892 6339 2942 6371
rect 2892 6319 2909 6339
rect 2929 6319 2942 6339
rect 2892 6294 2942 6319
rect 3110 6342 3160 6371
rect 3110 6322 3127 6342
rect 3147 6322 3160 6342
rect 4792 6367 4842 6380
rect 5010 6367 5060 6380
rect 5218 6367 5268 6380
rect 7845 6422 7895 6435
rect 8053 6422 8103 6435
rect 8271 6422 8321 6435
rect 3110 6294 3160 6322
rect 428 6226 478 6254
rect 428 6206 441 6226
rect 461 6206 478 6226
rect 428 6177 478 6206
rect 646 6229 696 6254
rect 646 6209 659 6229
rect 679 6209 696 6229
rect 646 6177 696 6209
rect 854 6227 904 6254
rect 854 6207 877 6227
rect 897 6207 904 6227
rect 854 6177 904 6207
rect 5755 6356 5805 6372
rect 5973 6356 6023 6372
rect 6181 6356 6231 6372
rect 7048 6354 7098 6384
rect 7048 6334 7055 6354
rect 7075 6334 7098 6354
rect 7048 6307 7098 6334
rect 7256 6352 7306 6384
rect 7256 6332 7273 6352
rect 7293 6332 7306 6352
rect 7256 6307 7306 6332
rect 7474 6355 7524 6384
rect 7474 6335 7491 6355
rect 7511 6335 7524 6355
rect 7474 6307 7524 6335
rect 3482 6229 3532 6245
rect 3690 6229 3740 6245
rect 3908 6229 3958 6245
rect 1226 6170 1276 6183
rect 1444 6170 1494 6183
rect 1652 6170 1702 6183
rect 2684 6181 2734 6194
rect 2892 6181 2942 6194
rect 3110 6181 3160 6194
rect 4792 6239 4842 6267
rect 428 6119 478 6135
rect 646 6119 696 6135
rect 854 6119 904 6135
rect 3482 6157 3532 6187
rect 3482 6137 3489 6157
rect 3509 6137 3532 6157
rect 3482 6110 3532 6137
rect 3690 6155 3740 6187
rect 3690 6135 3707 6155
rect 3727 6135 3740 6155
rect 3690 6110 3740 6135
rect 3908 6158 3958 6187
rect 3908 6138 3925 6158
rect 3945 6138 3958 6158
rect 4792 6219 4805 6239
rect 4825 6219 4842 6239
rect 4792 6190 4842 6219
rect 5010 6242 5060 6267
rect 5010 6222 5023 6242
rect 5043 6222 5060 6242
rect 5010 6190 5060 6222
rect 5218 6240 5268 6267
rect 5218 6220 5241 6240
rect 5261 6220 5268 6240
rect 5218 6190 5268 6220
rect 7846 6242 7896 6258
rect 8054 6242 8104 6258
rect 8272 6242 8322 6258
rect 3908 6110 3958 6138
rect 5590 6183 5640 6196
rect 5808 6183 5858 6196
rect 6016 6183 6066 6196
rect 7048 6194 7098 6207
rect 7256 6194 7306 6207
rect 7474 6194 7524 6207
rect 4792 6132 4842 6148
rect 5010 6132 5060 6148
rect 5218 6132 5268 6148
rect 1226 6042 1276 6070
rect 1226 6022 1239 6042
rect 1259 6022 1276 6042
rect 1226 5993 1276 6022
rect 1444 6045 1494 6070
rect 1444 6025 1457 6045
rect 1477 6025 1494 6045
rect 1444 5993 1494 6025
rect 1652 6043 1702 6070
rect 1652 6023 1675 6043
rect 1695 6023 1702 6043
rect 1652 5993 1702 6023
rect 2585 6003 2635 6019
rect 2793 6003 2843 6019
rect 3011 6003 3061 6019
rect 7846 6170 7896 6200
rect 7846 6150 7853 6170
rect 7873 6150 7896 6170
rect 7846 6123 7896 6150
rect 8054 6168 8104 6200
rect 8054 6148 8071 6168
rect 8091 6148 8104 6168
rect 8054 6123 8104 6148
rect 8272 6171 8322 6200
rect 8272 6151 8289 6171
rect 8309 6151 8322 6171
rect 8272 6123 8322 6151
rect 5590 6055 5640 6083
rect 429 5942 479 5955
rect 647 5942 697 5955
rect 855 5942 905 5955
rect 3482 5997 3532 6010
rect 3690 5997 3740 6010
rect 3908 5997 3958 6010
rect 5590 6035 5603 6055
rect 5623 6035 5640 6055
rect 5590 6006 5640 6035
rect 5808 6058 5858 6083
rect 5808 6038 5821 6058
rect 5841 6038 5858 6058
rect 5808 6006 5858 6038
rect 6016 6056 6066 6083
rect 6016 6036 6039 6056
rect 6059 6036 6066 6056
rect 6016 6006 6066 6036
rect 6949 6016 6999 6032
rect 7157 6016 7207 6032
rect 7375 6016 7425 6032
rect 1226 5935 1276 5951
rect 1444 5935 1494 5951
rect 1652 5935 1702 5951
rect 2585 5931 2635 5961
rect 2585 5911 2592 5931
rect 2612 5911 2635 5931
rect 2585 5884 2635 5911
rect 2793 5929 2843 5961
rect 2793 5909 2810 5929
rect 2830 5909 2843 5929
rect 2793 5884 2843 5909
rect 3011 5932 3061 5961
rect 4793 5955 4843 5968
rect 5011 5955 5061 5968
rect 5219 5955 5269 5968
rect 7846 6010 7896 6023
rect 8054 6010 8104 6023
rect 8272 6010 8322 6023
rect 3011 5912 3028 5932
rect 3048 5912 3061 5932
rect 3011 5884 3061 5912
rect 429 5814 479 5842
rect 429 5794 442 5814
rect 462 5794 479 5814
rect 429 5765 479 5794
rect 647 5817 697 5842
rect 647 5797 660 5817
rect 680 5797 697 5817
rect 647 5765 697 5797
rect 855 5815 905 5842
rect 855 5795 878 5815
rect 898 5795 905 5815
rect 855 5765 905 5795
rect 5590 5948 5640 5964
rect 5808 5948 5858 5964
rect 6016 5948 6066 5964
rect 6949 5944 6999 5974
rect 6949 5924 6956 5944
rect 6976 5924 6999 5944
rect 6949 5897 6999 5924
rect 7157 5942 7207 5974
rect 7157 5922 7174 5942
rect 7194 5922 7207 5942
rect 7157 5897 7207 5922
rect 7375 5945 7425 5974
rect 7375 5925 7392 5945
rect 7412 5925 7425 5945
rect 7375 5897 7425 5925
rect 4793 5827 4843 5855
rect 2585 5771 2635 5784
rect 2793 5771 2843 5784
rect 3011 5771 3061 5784
rect 4793 5807 4806 5827
rect 4826 5807 4843 5827
rect 4793 5778 4843 5807
rect 5011 5830 5061 5855
rect 5011 5810 5024 5830
rect 5044 5810 5061 5830
rect 5011 5778 5061 5810
rect 5219 5828 5269 5855
rect 5219 5808 5242 5828
rect 5262 5808 5269 5828
rect 5219 5778 5269 5808
rect 6949 5784 6999 5797
rect 7157 5784 7207 5797
rect 7375 5784 7425 5797
rect 429 5707 479 5723
rect 647 5707 697 5723
rect 855 5707 905 5723
rect 4793 5720 4843 5736
rect 5011 5720 5061 5736
rect 5219 5720 5269 5736
rect 3464 5623 3514 5639
rect 3672 5623 3722 5639
rect 3890 5623 3940 5639
rect 7828 5636 7878 5652
rect 8036 5636 8086 5652
rect 8254 5636 8304 5652
rect 1308 5562 1358 5575
rect 1526 5562 1576 5575
rect 1734 5562 1784 5575
rect 3464 5551 3514 5581
rect 3464 5531 3471 5551
rect 3491 5531 3514 5551
rect 3464 5504 3514 5531
rect 3672 5549 3722 5581
rect 3672 5529 3689 5549
rect 3709 5529 3722 5549
rect 3672 5504 3722 5529
rect 3890 5552 3940 5581
rect 3890 5532 3907 5552
rect 3927 5532 3940 5552
rect 5672 5575 5722 5588
rect 5890 5575 5940 5588
rect 6098 5575 6148 5588
rect 3890 5504 3940 5532
rect 1308 5434 1358 5462
rect 1308 5414 1321 5434
rect 1341 5414 1358 5434
rect 1308 5385 1358 5414
rect 1526 5437 1576 5462
rect 1526 5417 1539 5437
rect 1559 5417 1576 5437
rect 1526 5385 1576 5417
rect 1734 5435 1784 5462
rect 1734 5415 1757 5435
rect 1777 5415 1784 5435
rect 1734 5385 1784 5415
rect 2667 5395 2717 5411
rect 2875 5395 2925 5411
rect 3093 5395 3143 5411
rect 7828 5564 7878 5594
rect 7828 5544 7835 5564
rect 7855 5544 7878 5564
rect 7828 5517 7878 5544
rect 8036 5562 8086 5594
rect 8036 5542 8053 5562
rect 8073 5542 8086 5562
rect 8036 5517 8086 5542
rect 8254 5565 8304 5594
rect 8254 5545 8271 5565
rect 8291 5545 8304 5565
rect 8254 5517 8304 5545
rect 5672 5447 5722 5475
rect 5672 5427 5685 5447
rect 5705 5427 5722 5447
rect 411 5336 461 5349
rect 629 5336 679 5349
rect 837 5336 887 5349
rect 3464 5391 3514 5404
rect 3672 5391 3722 5404
rect 3890 5391 3940 5404
rect 5672 5398 5722 5427
rect 5890 5450 5940 5475
rect 5890 5430 5903 5450
rect 5923 5430 5940 5450
rect 5890 5398 5940 5430
rect 6098 5448 6148 5475
rect 6098 5428 6121 5448
rect 6141 5428 6148 5448
rect 6098 5398 6148 5428
rect 7031 5408 7081 5424
rect 7239 5408 7289 5424
rect 7457 5408 7507 5424
rect 1308 5327 1358 5343
rect 1526 5327 1576 5343
rect 1734 5327 1784 5343
rect 2667 5323 2717 5353
rect 2667 5303 2674 5323
rect 2694 5303 2717 5323
rect 2667 5276 2717 5303
rect 2875 5321 2925 5353
rect 2875 5301 2892 5321
rect 2912 5301 2925 5321
rect 2875 5276 2925 5301
rect 3093 5324 3143 5353
rect 3093 5304 3110 5324
rect 3130 5304 3143 5324
rect 4775 5349 4825 5362
rect 4993 5349 5043 5362
rect 5201 5349 5251 5362
rect 7828 5404 7878 5417
rect 8036 5404 8086 5417
rect 8254 5404 8304 5417
rect 3093 5276 3143 5304
rect 411 5208 461 5236
rect 411 5188 424 5208
rect 444 5188 461 5208
rect 411 5159 461 5188
rect 629 5211 679 5236
rect 629 5191 642 5211
rect 662 5191 679 5211
rect 629 5159 679 5191
rect 837 5209 887 5236
rect 837 5189 860 5209
rect 880 5189 887 5209
rect 837 5159 887 5189
rect 5672 5340 5722 5356
rect 5890 5340 5940 5356
rect 6098 5340 6148 5356
rect 7031 5336 7081 5366
rect 7031 5316 7038 5336
rect 7058 5316 7081 5336
rect 7031 5289 7081 5316
rect 7239 5334 7289 5366
rect 7239 5314 7256 5334
rect 7276 5314 7289 5334
rect 7239 5289 7289 5314
rect 7457 5337 7507 5366
rect 7457 5317 7474 5337
rect 7494 5317 7507 5337
rect 7457 5289 7507 5317
rect 3465 5211 3515 5227
rect 3673 5211 3723 5227
rect 3891 5211 3941 5227
rect 1209 5152 1259 5165
rect 1427 5152 1477 5165
rect 1635 5152 1685 5165
rect 2667 5163 2717 5176
rect 2875 5163 2925 5176
rect 3093 5163 3143 5176
rect 4775 5221 4825 5249
rect 411 5101 461 5117
rect 629 5101 679 5117
rect 837 5101 887 5117
rect 3465 5139 3515 5169
rect 3465 5119 3472 5139
rect 3492 5119 3515 5139
rect 3465 5092 3515 5119
rect 3673 5137 3723 5169
rect 3673 5117 3690 5137
rect 3710 5117 3723 5137
rect 3673 5092 3723 5117
rect 3891 5140 3941 5169
rect 3891 5120 3908 5140
rect 3928 5120 3941 5140
rect 4775 5201 4788 5221
rect 4808 5201 4825 5221
rect 4775 5172 4825 5201
rect 4993 5224 5043 5249
rect 4993 5204 5006 5224
rect 5026 5204 5043 5224
rect 4993 5172 5043 5204
rect 5201 5222 5251 5249
rect 5201 5202 5224 5222
rect 5244 5202 5251 5222
rect 5201 5172 5251 5202
rect 7829 5224 7879 5240
rect 8037 5224 8087 5240
rect 8255 5224 8305 5240
rect 3891 5092 3941 5120
rect 5573 5165 5623 5178
rect 5791 5165 5841 5178
rect 5999 5165 6049 5178
rect 7031 5176 7081 5189
rect 7239 5176 7289 5189
rect 7457 5176 7507 5189
rect 4775 5114 4825 5130
rect 4993 5114 5043 5130
rect 5201 5114 5251 5130
rect 1209 5024 1259 5052
rect 1209 5004 1222 5024
rect 1242 5004 1259 5024
rect 1209 4975 1259 5004
rect 1427 5027 1477 5052
rect 1427 5007 1440 5027
rect 1460 5007 1477 5027
rect 1427 4975 1477 5007
rect 1635 5025 1685 5052
rect 1635 5005 1658 5025
rect 1678 5005 1685 5025
rect 1635 4975 1685 5005
rect 2363 4989 2413 5005
rect 2571 4989 2621 5005
rect 2789 4989 2839 5005
rect 7829 5152 7879 5182
rect 7829 5132 7836 5152
rect 7856 5132 7879 5152
rect 7829 5105 7879 5132
rect 8037 5150 8087 5182
rect 8037 5130 8054 5150
rect 8074 5130 8087 5150
rect 8037 5105 8087 5130
rect 8255 5153 8305 5182
rect 8255 5133 8272 5153
rect 8292 5133 8305 5153
rect 8255 5105 8305 5133
rect 5573 5037 5623 5065
rect 412 4924 462 4937
rect 630 4924 680 4937
rect 838 4924 888 4937
rect 3465 4979 3515 4992
rect 3673 4979 3723 4992
rect 3891 4979 3941 4992
rect 5573 5017 5586 5037
rect 5606 5017 5623 5037
rect 5573 4988 5623 5017
rect 5791 5040 5841 5065
rect 5791 5020 5804 5040
rect 5824 5020 5841 5040
rect 5791 4988 5841 5020
rect 5999 5038 6049 5065
rect 5999 5018 6022 5038
rect 6042 5018 6049 5038
rect 5999 4988 6049 5018
rect 6727 5002 6777 5018
rect 6935 5002 6985 5018
rect 7153 5002 7203 5018
rect 1209 4917 1259 4933
rect 1427 4917 1477 4933
rect 1635 4917 1685 4933
rect 2363 4917 2413 4947
rect 2363 4897 2370 4917
rect 2390 4897 2413 4917
rect 2363 4870 2413 4897
rect 2571 4915 2621 4947
rect 2571 4895 2588 4915
rect 2608 4895 2621 4915
rect 2571 4870 2621 4895
rect 2789 4918 2839 4947
rect 4776 4937 4826 4950
rect 4994 4937 5044 4950
rect 5202 4937 5252 4950
rect 7829 4992 7879 5005
rect 8037 4992 8087 5005
rect 8255 4992 8305 5005
rect 2789 4898 2806 4918
rect 2826 4898 2839 4918
rect 2789 4870 2839 4898
rect 412 4796 462 4824
rect 412 4776 425 4796
rect 445 4776 462 4796
rect 412 4747 462 4776
rect 630 4799 680 4824
rect 630 4779 643 4799
rect 663 4779 680 4799
rect 630 4747 680 4779
rect 838 4797 888 4824
rect 838 4777 861 4797
rect 881 4777 888 4797
rect 838 4747 888 4777
rect 5573 4930 5623 4946
rect 5791 4930 5841 4946
rect 5999 4930 6049 4946
rect 6727 4930 6777 4960
rect 6727 4910 6734 4930
rect 6754 4910 6777 4930
rect 6727 4883 6777 4910
rect 6935 4928 6985 4960
rect 6935 4908 6952 4928
rect 6972 4908 6985 4928
rect 6935 4883 6985 4908
rect 7153 4931 7203 4960
rect 7153 4911 7170 4931
rect 7190 4911 7203 4931
rect 7153 4883 7203 4911
rect 4776 4809 4826 4837
rect 2363 4757 2413 4770
rect 2571 4757 2621 4770
rect 2789 4757 2839 4770
rect 4776 4789 4789 4809
rect 4809 4789 4826 4809
rect 4776 4760 4826 4789
rect 4994 4812 5044 4837
rect 4994 4792 5007 4812
rect 5027 4792 5044 4812
rect 4994 4760 5044 4792
rect 5202 4810 5252 4837
rect 5202 4790 5225 4810
rect 5245 4790 5252 4810
rect 5202 4760 5252 4790
rect 6727 4770 6777 4783
rect 6935 4770 6985 4783
rect 7153 4770 7203 4783
rect 412 4689 462 4705
rect 630 4689 680 4705
rect 838 4689 888 4705
rect 4776 4702 4826 4718
rect 4994 4702 5044 4718
rect 5202 4702 5252 4718
rect 3445 4605 3495 4621
rect 3653 4605 3703 4621
rect 3871 4605 3921 4621
rect 7809 4618 7859 4634
rect 8017 4618 8067 4634
rect 8235 4618 8285 4634
rect 1494 4540 1544 4553
rect 1712 4540 1762 4553
rect 1920 4540 1970 4553
rect 3445 4533 3495 4563
rect 3445 4513 3452 4533
rect 3472 4513 3495 4533
rect 3445 4486 3495 4513
rect 3653 4531 3703 4563
rect 3653 4511 3670 4531
rect 3690 4511 3703 4531
rect 3653 4486 3703 4511
rect 3871 4534 3921 4563
rect 3871 4514 3888 4534
rect 3908 4514 3921 4534
rect 5858 4553 5908 4566
rect 6076 4553 6126 4566
rect 6284 4553 6334 4566
rect 3871 4486 3921 4514
rect 1494 4412 1544 4440
rect 1494 4392 1507 4412
rect 1527 4392 1544 4412
rect 1494 4363 1544 4392
rect 1712 4415 1762 4440
rect 1712 4395 1725 4415
rect 1745 4395 1762 4415
rect 1712 4363 1762 4395
rect 1920 4413 1970 4440
rect 1920 4393 1943 4413
rect 1963 4393 1970 4413
rect 1920 4363 1970 4393
rect 2648 4377 2698 4393
rect 2856 4377 2906 4393
rect 3074 4377 3124 4393
rect 7809 4546 7859 4576
rect 7809 4526 7816 4546
rect 7836 4526 7859 4546
rect 7809 4499 7859 4526
rect 8017 4544 8067 4576
rect 8017 4524 8034 4544
rect 8054 4524 8067 4544
rect 8017 4499 8067 4524
rect 8235 4547 8285 4576
rect 8235 4527 8252 4547
rect 8272 4527 8285 4547
rect 8235 4499 8285 4527
rect 5858 4425 5908 4453
rect 5858 4405 5871 4425
rect 5891 4405 5908 4425
rect 392 4318 442 4331
rect 610 4318 660 4331
rect 818 4318 868 4331
rect 3445 4373 3495 4386
rect 3653 4373 3703 4386
rect 3871 4373 3921 4386
rect 5858 4376 5908 4405
rect 6076 4428 6126 4453
rect 6076 4408 6089 4428
rect 6109 4408 6126 4428
rect 6076 4376 6126 4408
rect 6284 4426 6334 4453
rect 6284 4406 6307 4426
rect 6327 4406 6334 4426
rect 6284 4376 6334 4406
rect 7012 4390 7062 4406
rect 7220 4390 7270 4406
rect 7438 4390 7488 4406
rect 1494 4305 1544 4321
rect 1712 4305 1762 4321
rect 1920 4305 1970 4321
rect 2648 4305 2698 4335
rect 2648 4285 2655 4305
rect 2675 4285 2698 4305
rect 2648 4258 2698 4285
rect 2856 4303 2906 4335
rect 2856 4283 2873 4303
rect 2893 4283 2906 4303
rect 2856 4258 2906 4283
rect 3074 4306 3124 4335
rect 3074 4286 3091 4306
rect 3111 4286 3124 4306
rect 4756 4331 4806 4344
rect 4974 4331 5024 4344
rect 5182 4331 5232 4344
rect 7809 4386 7859 4399
rect 8017 4386 8067 4399
rect 8235 4386 8285 4399
rect 3074 4258 3124 4286
rect 392 4190 442 4218
rect 392 4170 405 4190
rect 425 4170 442 4190
rect 392 4141 442 4170
rect 610 4193 660 4218
rect 610 4173 623 4193
rect 643 4173 660 4193
rect 610 4141 660 4173
rect 818 4191 868 4218
rect 818 4171 841 4191
rect 861 4171 868 4191
rect 818 4141 868 4171
rect 5858 4318 5908 4334
rect 6076 4318 6126 4334
rect 6284 4318 6334 4334
rect 7012 4318 7062 4348
rect 7012 4298 7019 4318
rect 7039 4298 7062 4318
rect 7012 4271 7062 4298
rect 7220 4316 7270 4348
rect 7220 4296 7237 4316
rect 7257 4296 7270 4316
rect 7220 4271 7270 4296
rect 7438 4319 7488 4348
rect 7438 4299 7455 4319
rect 7475 4299 7488 4319
rect 7438 4271 7488 4299
rect 3446 4193 3496 4209
rect 3654 4193 3704 4209
rect 3872 4193 3922 4209
rect 1190 4134 1240 4147
rect 1408 4134 1458 4147
rect 1616 4134 1666 4147
rect 2648 4145 2698 4158
rect 2856 4145 2906 4158
rect 3074 4145 3124 4158
rect 4756 4203 4806 4231
rect 392 4083 442 4099
rect 610 4083 660 4099
rect 818 4083 868 4099
rect 3446 4121 3496 4151
rect 3446 4101 3453 4121
rect 3473 4101 3496 4121
rect 3446 4074 3496 4101
rect 3654 4119 3704 4151
rect 3654 4099 3671 4119
rect 3691 4099 3704 4119
rect 3654 4074 3704 4099
rect 3872 4122 3922 4151
rect 3872 4102 3889 4122
rect 3909 4102 3922 4122
rect 4756 4183 4769 4203
rect 4789 4183 4806 4203
rect 4756 4154 4806 4183
rect 4974 4206 5024 4231
rect 4974 4186 4987 4206
rect 5007 4186 5024 4206
rect 4974 4154 5024 4186
rect 5182 4204 5232 4231
rect 5182 4184 5205 4204
rect 5225 4184 5232 4204
rect 5182 4154 5232 4184
rect 7810 4206 7860 4222
rect 8018 4206 8068 4222
rect 8236 4206 8286 4222
rect 3872 4074 3922 4102
rect 5554 4147 5604 4160
rect 5772 4147 5822 4160
rect 5980 4147 6030 4160
rect 7012 4158 7062 4171
rect 7220 4158 7270 4171
rect 7438 4158 7488 4171
rect 4756 4096 4806 4112
rect 4974 4096 5024 4112
rect 5182 4096 5232 4112
rect 1190 4006 1240 4034
rect 1190 3986 1203 4006
rect 1223 3986 1240 4006
rect 1190 3957 1240 3986
rect 1408 4009 1458 4034
rect 1408 3989 1421 4009
rect 1441 3989 1458 4009
rect 1408 3957 1458 3989
rect 1616 4007 1666 4034
rect 1616 3987 1639 4007
rect 1659 3987 1666 4007
rect 1616 3957 1666 3987
rect 2549 3967 2599 3983
rect 2757 3967 2807 3983
rect 2975 3967 3025 3983
rect 7810 4134 7860 4164
rect 7810 4114 7817 4134
rect 7837 4114 7860 4134
rect 7810 4087 7860 4114
rect 8018 4132 8068 4164
rect 8018 4112 8035 4132
rect 8055 4112 8068 4132
rect 8018 4087 8068 4112
rect 8236 4135 8286 4164
rect 8236 4115 8253 4135
rect 8273 4115 8286 4135
rect 8236 4087 8286 4115
rect 5554 4019 5604 4047
rect 393 3906 443 3919
rect 611 3906 661 3919
rect 819 3906 869 3919
rect 3446 3961 3496 3974
rect 3654 3961 3704 3974
rect 3872 3961 3922 3974
rect 5554 3999 5567 4019
rect 5587 3999 5604 4019
rect 5554 3970 5604 3999
rect 5772 4022 5822 4047
rect 5772 4002 5785 4022
rect 5805 4002 5822 4022
rect 5772 3970 5822 4002
rect 5980 4020 6030 4047
rect 5980 4000 6003 4020
rect 6023 4000 6030 4020
rect 5980 3970 6030 4000
rect 6913 3980 6963 3996
rect 7121 3980 7171 3996
rect 7339 3980 7389 3996
rect 1190 3899 1240 3915
rect 1408 3899 1458 3915
rect 1616 3899 1666 3915
rect 2549 3895 2599 3925
rect 2549 3875 2556 3895
rect 2576 3875 2599 3895
rect 2549 3848 2599 3875
rect 2757 3893 2807 3925
rect 2757 3873 2774 3893
rect 2794 3873 2807 3893
rect 2757 3848 2807 3873
rect 2975 3896 3025 3925
rect 4757 3919 4807 3932
rect 4975 3919 5025 3932
rect 5183 3919 5233 3932
rect 7810 3974 7860 3987
rect 8018 3974 8068 3987
rect 8236 3974 8286 3987
rect 2975 3876 2992 3896
rect 3012 3876 3025 3896
rect 2975 3848 3025 3876
rect 393 3778 443 3806
rect 393 3758 406 3778
rect 426 3758 443 3778
rect 393 3729 443 3758
rect 611 3781 661 3806
rect 611 3761 624 3781
rect 644 3761 661 3781
rect 611 3729 661 3761
rect 819 3779 869 3806
rect 819 3759 842 3779
rect 862 3759 869 3779
rect 819 3729 869 3759
rect 5554 3912 5604 3928
rect 5772 3912 5822 3928
rect 5980 3912 6030 3928
rect 6913 3908 6963 3938
rect 6913 3888 6920 3908
rect 6940 3888 6963 3908
rect 6913 3861 6963 3888
rect 7121 3906 7171 3938
rect 7121 3886 7138 3906
rect 7158 3886 7171 3906
rect 7121 3861 7171 3886
rect 7339 3909 7389 3938
rect 7339 3889 7356 3909
rect 7376 3889 7389 3909
rect 7339 3861 7389 3889
rect 4757 3791 4807 3819
rect 2549 3735 2599 3748
rect 2757 3735 2807 3748
rect 2975 3735 3025 3748
rect 4757 3771 4770 3791
rect 4790 3771 4807 3791
rect 4757 3742 4807 3771
rect 4975 3794 5025 3819
rect 4975 3774 4988 3794
rect 5008 3774 5025 3794
rect 4975 3742 5025 3774
rect 5183 3792 5233 3819
rect 5183 3772 5206 3792
rect 5226 3772 5233 3792
rect 5183 3742 5233 3772
rect 6913 3748 6963 3761
rect 7121 3748 7171 3761
rect 7339 3748 7389 3761
rect 393 3671 443 3687
rect 611 3671 661 3687
rect 819 3671 869 3687
rect 4757 3684 4807 3700
rect 4975 3684 5025 3700
rect 5183 3684 5233 3700
rect 3428 3587 3478 3603
rect 3636 3587 3686 3603
rect 3854 3587 3904 3603
rect 7792 3600 7842 3616
rect 8000 3600 8050 3616
rect 8218 3600 8268 3616
rect 1272 3526 1322 3539
rect 1490 3526 1540 3539
rect 1698 3526 1748 3539
rect 3428 3515 3478 3545
rect 3428 3495 3435 3515
rect 3455 3495 3478 3515
rect 3428 3468 3478 3495
rect 3636 3513 3686 3545
rect 3636 3493 3653 3513
rect 3673 3493 3686 3513
rect 3636 3468 3686 3493
rect 3854 3516 3904 3545
rect 3854 3496 3871 3516
rect 3891 3496 3904 3516
rect 5636 3539 5686 3552
rect 5854 3539 5904 3552
rect 6062 3539 6112 3552
rect 3854 3468 3904 3496
rect 1272 3398 1322 3426
rect 1272 3378 1285 3398
rect 1305 3378 1322 3398
rect 1272 3349 1322 3378
rect 1490 3401 1540 3426
rect 1490 3381 1503 3401
rect 1523 3381 1540 3401
rect 1490 3349 1540 3381
rect 1698 3399 1748 3426
rect 1698 3379 1721 3399
rect 1741 3379 1748 3399
rect 1698 3349 1748 3379
rect 2631 3359 2681 3375
rect 2839 3359 2889 3375
rect 3057 3359 3107 3375
rect 7792 3528 7842 3558
rect 7792 3508 7799 3528
rect 7819 3508 7842 3528
rect 7792 3481 7842 3508
rect 8000 3526 8050 3558
rect 8000 3506 8017 3526
rect 8037 3506 8050 3526
rect 8000 3481 8050 3506
rect 8218 3529 8268 3558
rect 8218 3509 8235 3529
rect 8255 3509 8268 3529
rect 8218 3481 8268 3509
rect 5636 3411 5686 3439
rect 5636 3391 5649 3411
rect 5669 3391 5686 3411
rect 375 3300 425 3313
rect 593 3300 643 3313
rect 801 3300 851 3313
rect 3428 3355 3478 3368
rect 3636 3355 3686 3368
rect 3854 3355 3904 3368
rect 5636 3362 5686 3391
rect 5854 3414 5904 3439
rect 5854 3394 5867 3414
rect 5887 3394 5904 3414
rect 5854 3362 5904 3394
rect 6062 3412 6112 3439
rect 6062 3392 6085 3412
rect 6105 3392 6112 3412
rect 6062 3362 6112 3392
rect 6995 3372 7045 3388
rect 7203 3372 7253 3388
rect 7421 3372 7471 3388
rect 1272 3291 1322 3307
rect 1490 3291 1540 3307
rect 1698 3291 1748 3307
rect 2631 3287 2681 3317
rect 2631 3267 2638 3287
rect 2658 3267 2681 3287
rect 2631 3240 2681 3267
rect 2839 3285 2889 3317
rect 2839 3265 2856 3285
rect 2876 3265 2889 3285
rect 2839 3240 2889 3265
rect 3057 3288 3107 3317
rect 3057 3268 3074 3288
rect 3094 3268 3107 3288
rect 4739 3313 4789 3326
rect 4957 3313 5007 3326
rect 5165 3313 5215 3326
rect 7792 3368 7842 3381
rect 8000 3368 8050 3381
rect 8218 3368 8268 3381
rect 3057 3240 3107 3268
rect 375 3172 425 3200
rect 375 3152 388 3172
rect 408 3152 425 3172
rect 375 3123 425 3152
rect 593 3175 643 3200
rect 593 3155 606 3175
rect 626 3155 643 3175
rect 593 3123 643 3155
rect 801 3173 851 3200
rect 801 3153 824 3173
rect 844 3153 851 3173
rect 801 3123 851 3153
rect 5636 3304 5686 3320
rect 5854 3304 5904 3320
rect 6062 3304 6112 3320
rect 6995 3300 7045 3330
rect 6995 3280 7002 3300
rect 7022 3280 7045 3300
rect 6995 3253 7045 3280
rect 7203 3298 7253 3330
rect 7203 3278 7220 3298
rect 7240 3278 7253 3298
rect 7203 3253 7253 3278
rect 7421 3301 7471 3330
rect 7421 3281 7438 3301
rect 7458 3281 7471 3301
rect 7421 3253 7471 3281
rect 3429 3175 3479 3191
rect 3637 3175 3687 3191
rect 3855 3175 3905 3191
rect 1173 3116 1223 3129
rect 1391 3116 1441 3129
rect 1599 3116 1649 3129
rect 2631 3127 2681 3140
rect 2839 3127 2889 3140
rect 3057 3127 3107 3140
rect 4739 3185 4789 3213
rect 375 3065 425 3081
rect 593 3065 643 3081
rect 801 3065 851 3081
rect 3429 3103 3479 3133
rect 3429 3083 3436 3103
rect 3456 3083 3479 3103
rect 3429 3056 3479 3083
rect 3637 3101 3687 3133
rect 3637 3081 3654 3101
rect 3674 3081 3687 3101
rect 3637 3056 3687 3081
rect 3855 3104 3905 3133
rect 3855 3084 3872 3104
rect 3892 3084 3905 3104
rect 4739 3165 4752 3185
rect 4772 3165 4789 3185
rect 4739 3136 4789 3165
rect 4957 3188 5007 3213
rect 4957 3168 4970 3188
rect 4990 3168 5007 3188
rect 4957 3136 5007 3168
rect 5165 3186 5215 3213
rect 5165 3166 5188 3186
rect 5208 3166 5215 3186
rect 5165 3136 5215 3166
rect 7793 3188 7843 3204
rect 8001 3188 8051 3204
rect 8219 3188 8269 3204
rect 3855 3056 3905 3084
rect 5537 3129 5587 3142
rect 5755 3129 5805 3142
rect 5963 3129 6013 3142
rect 6995 3140 7045 3153
rect 7203 3140 7253 3153
rect 7421 3140 7471 3153
rect 4739 3078 4789 3094
rect 4957 3078 5007 3094
rect 5165 3078 5215 3094
rect 1173 2988 1223 3016
rect 1173 2968 1186 2988
rect 1206 2968 1223 2988
rect 1173 2939 1223 2968
rect 1391 2991 1441 3016
rect 1391 2971 1404 2991
rect 1424 2971 1441 2991
rect 1391 2939 1441 2971
rect 1599 2989 1649 3016
rect 1599 2969 1622 2989
rect 1642 2969 1649 2989
rect 1599 2939 1649 2969
rect 2466 2951 2516 2967
rect 2674 2951 2724 2967
rect 2892 2951 2942 2967
rect 7793 3116 7843 3146
rect 7793 3096 7800 3116
rect 7820 3096 7843 3116
rect 7793 3069 7843 3096
rect 8001 3114 8051 3146
rect 8001 3094 8018 3114
rect 8038 3094 8051 3114
rect 8001 3069 8051 3094
rect 8219 3117 8269 3146
rect 8219 3097 8236 3117
rect 8256 3097 8269 3117
rect 8219 3069 8269 3097
rect 5537 3001 5587 3029
rect 376 2888 426 2901
rect 594 2888 644 2901
rect 802 2888 852 2901
rect 3429 2943 3479 2956
rect 3637 2943 3687 2956
rect 3855 2943 3905 2956
rect 5537 2981 5550 3001
rect 5570 2981 5587 3001
rect 5537 2952 5587 2981
rect 5755 3004 5805 3029
rect 5755 2984 5768 3004
rect 5788 2984 5805 3004
rect 5755 2952 5805 2984
rect 5963 3002 6013 3029
rect 5963 2982 5986 3002
rect 6006 2982 6013 3002
rect 5963 2952 6013 2982
rect 6830 2964 6880 2980
rect 7038 2964 7088 2980
rect 7256 2964 7306 2980
rect 1173 2881 1223 2897
rect 1391 2881 1441 2897
rect 1599 2881 1649 2897
rect 2466 2879 2516 2909
rect 2466 2859 2473 2879
rect 2493 2859 2516 2879
rect 2466 2832 2516 2859
rect 2674 2877 2724 2909
rect 2674 2857 2691 2877
rect 2711 2857 2724 2877
rect 2674 2832 2724 2857
rect 2892 2880 2942 2909
rect 4740 2901 4790 2914
rect 4958 2901 5008 2914
rect 5166 2901 5216 2914
rect 7793 2956 7843 2969
rect 8001 2956 8051 2969
rect 8219 2956 8269 2969
rect 2892 2860 2909 2880
rect 2929 2860 2942 2880
rect 2892 2832 2942 2860
rect 376 2760 426 2788
rect 376 2740 389 2760
rect 409 2740 426 2760
rect 376 2711 426 2740
rect 594 2763 644 2788
rect 594 2743 607 2763
rect 627 2743 644 2763
rect 594 2711 644 2743
rect 802 2761 852 2788
rect 802 2741 825 2761
rect 845 2741 852 2761
rect 802 2711 852 2741
rect 5537 2894 5587 2910
rect 5755 2894 5805 2910
rect 5963 2894 6013 2910
rect 6830 2892 6880 2922
rect 6830 2872 6837 2892
rect 6857 2872 6880 2892
rect 6830 2845 6880 2872
rect 7038 2890 7088 2922
rect 7038 2870 7055 2890
rect 7075 2870 7088 2890
rect 7038 2845 7088 2870
rect 7256 2893 7306 2922
rect 7256 2873 7273 2893
rect 7293 2873 7306 2893
rect 7256 2845 7306 2873
rect 4740 2773 4790 2801
rect 2466 2719 2516 2732
rect 2674 2719 2724 2732
rect 2892 2719 2942 2732
rect 4740 2753 4753 2773
rect 4773 2753 4790 2773
rect 4740 2724 4790 2753
rect 4958 2776 5008 2801
rect 4958 2756 4971 2776
rect 4991 2756 5008 2776
rect 4958 2724 5008 2756
rect 5166 2774 5216 2801
rect 5166 2754 5189 2774
rect 5209 2754 5216 2774
rect 5166 2724 5216 2754
rect 6830 2732 6880 2745
rect 7038 2732 7088 2745
rect 7256 2732 7306 2745
rect 376 2653 426 2669
rect 594 2653 644 2669
rect 802 2653 852 2669
rect 4740 2666 4790 2682
rect 4958 2666 5008 2682
rect 5166 2666 5216 2682
rect 3408 2569 3458 2585
rect 3616 2569 3666 2585
rect 3834 2569 3884 2585
rect 7772 2582 7822 2598
rect 7980 2582 8030 2598
rect 8198 2582 8248 2598
rect 1318 2506 1368 2519
rect 1536 2506 1586 2519
rect 1744 2506 1794 2519
rect 3408 2497 3458 2527
rect 3408 2477 3415 2497
rect 3435 2477 3458 2497
rect 3408 2450 3458 2477
rect 3616 2495 3666 2527
rect 3616 2475 3633 2495
rect 3653 2475 3666 2495
rect 3616 2450 3666 2475
rect 3834 2498 3884 2527
rect 3834 2478 3851 2498
rect 3871 2478 3884 2498
rect 5682 2519 5732 2532
rect 5900 2519 5950 2532
rect 6108 2519 6158 2532
rect 3834 2450 3884 2478
rect 1318 2378 1368 2406
rect 1318 2358 1331 2378
rect 1351 2358 1368 2378
rect 1318 2329 1368 2358
rect 1536 2381 1586 2406
rect 1536 2361 1549 2381
rect 1569 2361 1586 2381
rect 1536 2329 1586 2361
rect 1744 2379 1794 2406
rect 1744 2359 1767 2379
rect 1787 2359 1794 2379
rect 1744 2329 1794 2359
rect 2611 2341 2661 2357
rect 2819 2341 2869 2357
rect 3037 2341 3087 2357
rect 7772 2510 7822 2540
rect 7772 2490 7779 2510
rect 7799 2490 7822 2510
rect 7772 2463 7822 2490
rect 7980 2508 8030 2540
rect 7980 2488 7997 2508
rect 8017 2488 8030 2508
rect 7980 2463 8030 2488
rect 8198 2511 8248 2540
rect 8198 2491 8215 2511
rect 8235 2491 8248 2511
rect 8198 2463 8248 2491
rect 5682 2391 5732 2419
rect 5682 2371 5695 2391
rect 5715 2371 5732 2391
rect 355 2282 405 2295
rect 573 2282 623 2295
rect 781 2282 831 2295
rect 3408 2337 3458 2350
rect 3616 2337 3666 2350
rect 3834 2337 3884 2350
rect 5682 2342 5732 2371
rect 5900 2394 5950 2419
rect 5900 2374 5913 2394
rect 5933 2374 5950 2394
rect 5900 2342 5950 2374
rect 6108 2392 6158 2419
rect 6108 2372 6131 2392
rect 6151 2372 6158 2392
rect 6108 2342 6158 2372
rect 6975 2354 7025 2370
rect 7183 2354 7233 2370
rect 7401 2354 7451 2370
rect 1318 2271 1368 2287
rect 1536 2271 1586 2287
rect 1744 2271 1794 2287
rect 2611 2269 2661 2299
rect 2611 2249 2618 2269
rect 2638 2249 2661 2269
rect 2611 2222 2661 2249
rect 2819 2267 2869 2299
rect 2819 2247 2836 2267
rect 2856 2247 2869 2267
rect 2819 2222 2869 2247
rect 3037 2270 3087 2299
rect 3037 2250 3054 2270
rect 3074 2250 3087 2270
rect 4719 2295 4769 2308
rect 4937 2295 4987 2308
rect 5145 2295 5195 2308
rect 7772 2350 7822 2363
rect 7980 2350 8030 2363
rect 8198 2350 8248 2363
rect 3037 2222 3087 2250
rect 355 2154 405 2182
rect 355 2134 368 2154
rect 388 2134 405 2154
rect 355 2105 405 2134
rect 573 2157 623 2182
rect 573 2137 586 2157
rect 606 2137 623 2157
rect 573 2105 623 2137
rect 781 2155 831 2182
rect 781 2135 804 2155
rect 824 2135 831 2155
rect 781 2105 831 2135
rect 5682 2284 5732 2300
rect 5900 2284 5950 2300
rect 6108 2284 6158 2300
rect 6975 2282 7025 2312
rect 6975 2262 6982 2282
rect 7002 2262 7025 2282
rect 6975 2235 7025 2262
rect 7183 2280 7233 2312
rect 7183 2260 7200 2280
rect 7220 2260 7233 2280
rect 7183 2235 7233 2260
rect 7401 2283 7451 2312
rect 7401 2263 7418 2283
rect 7438 2263 7451 2283
rect 7401 2235 7451 2263
rect 3409 2157 3459 2173
rect 3617 2157 3667 2173
rect 3835 2157 3885 2173
rect 1153 2098 1203 2111
rect 1371 2098 1421 2111
rect 1579 2098 1629 2111
rect 2611 2109 2661 2122
rect 2819 2109 2869 2122
rect 3037 2109 3087 2122
rect 4719 2167 4769 2195
rect 355 2047 405 2063
rect 573 2047 623 2063
rect 781 2047 831 2063
rect 3409 2085 3459 2115
rect 3409 2065 3416 2085
rect 3436 2065 3459 2085
rect 3409 2038 3459 2065
rect 3617 2083 3667 2115
rect 3617 2063 3634 2083
rect 3654 2063 3667 2083
rect 3617 2038 3667 2063
rect 3835 2086 3885 2115
rect 3835 2066 3852 2086
rect 3872 2066 3885 2086
rect 4719 2147 4732 2167
rect 4752 2147 4769 2167
rect 4719 2118 4769 2147
rect 4937 2170 4987 2195
rect 4937 2150 4950 2170
rect 4970 2150 4987 2170
rect 4937 2118 4987 2150
rect 5145 2168 5195 2195
rect 5145 2148 5168 2168
rect 5188 2148 5195 2168
rect 5145 2118 5195 2148
rect 7773 2170 7823 2186
rect 7981 2170 8031 2186
rect 8199 2170 8249 2186
rect 3835 2038 3885 2066
rect 5517 2111 5567 2124
rect 5735 2111 5785 2124
rect 5943 2111 5993 2124
rect 6975 2122 7025 2135
rect 7183 2122 7233 2135
rect 7401 2122 7451 2135
rect 4719 2060 4769 2076
rect 4937 2060 4987 2076
rect 5145 2060 5195 2076
rect 1153 1970 1203 1998
rect 1153 1950 1166 1970
rect 1186 1950 1203 1970
rect 1153 1921 1203 1950
rect 1371 1973 1421 1998
rect 1371 1953 1384 1973
rect 1404 1953 1421 1973
rect 1371 1921 1421 1953
rect 1579 1971 1629 1998
rect 1579 1951 1602 1971
rect 1622 1951 1629 1971
rect 1579 1921 1629 1951
rect 2512 1931 2562 1947
rect 2720 1931 2770 1947
rect 2938 1931 2988 1947
rect 7773 2098 7823 2128
rect 7773 2078 7780 2098
rect 7800 2078 7823 2098
rect 7773 2051 7823 2078
rect 7981 2096 8031 2128
rect 7981 2076 7998 2096
rect 8018 2076 8031 2096
rect 7981 2051 8031 2076
rect 8199 2099 8249 2128
rect 8199 2079 8216 2099
rect 8236 2079 8249 2099
rect 8199 2051 8249 2079
rect 5517 1983 5567 2011
rect 356 1870 406 1883
rect 574 1870 624 1883
rect 782 1870 832 1883
rect 3409 1925 3459 1938
rect 3617 1925 3667 1938
rect 3835 1925 3885 1938
rect 5517 1963 5530 1983
rect 5550 1963 5567 1983
rect 5517 1934 5567 1963
rect 5735 1986 5785 2011
rect 5735 1966 5748 1986
rect 5768 1966 5785 1986
rect 5735 1934 5785 1966
rect 5943 1984 5993 2011
rect 5943 1964 5966 1984
rect 5986 1964 5993 1984
rect 5943 1934 5993 1964
rect 6876 1944 6926 1960
rect 7084 1944 7134 1960
rect 7302 1944 7352 1960
rect 1153 1863 1203 1879
rect 1371 1863 1421 1879
rect 1579 1863 1629 1879
rect 2512 1859 2562 1889
rect 2512 1839 2519 1859
rect 2539 1839 2562 1859
rect 2512 1812 2562 1839
rect 2720 1857 2770 1889
rect 2720 1837 2737 1857
rect 2757 1837 2770 1857
rect 2720 1812 2770 1837
rect 2938 1860 2988 1889
rect 4720 1883 4770 1896
rect 4938 1883 4988 1896
rect 5146 1883 5196 1896
rect 7773 1938 7823 1951
rect 7981 1938 8031 1951
rect 8199 1938 8249 1951
rect 2938 1840 2955 1860
rect 2975 1840 2988 1860
rect 2938 1812 2988 1840
rect 356 1742 406 1770
rect 356 1722 369 1742
rect 389 1722 406 1742
rect 356 1693 406 1722
rect 574 1745 624 1770
rect 574 1725 587 1745
rect 607 1725 624 1745
rect 574 1693 624 1725
rect 782 1743 832 1770
rect 782 1723 805 1743
rect 825 1723 832 1743
rect 782 1693 832 1723
rect 5517 1876 5567 1892
rect 5735 1876 5785 1892
rect 5943 1876 5993 1892
rect 6876 1872 6926 1902
rect 6876 1852 6883 1872
rect 6903 1852 6926 1872
rect 6876 1825 6926 1852
rect 7084 1870 7134 1902
rect 7084 1850 7101 1870
rect 7121 1850 7134 1870
rect 7084 1825 7134 1850
rect 7302 1873 7352 1902
rect 7302 1853 7319 1873
rect 7339 1853 7352 1873
rect 7302 1825 7352 1853
rect 4720 1755 4770 1783
rect 2512 1699 2562 1712
rect 2720 1699 2770 1712
rect 2938 1699 2988 1712
rect 4720 1735 4733 1755
rect 4753 1735 4770 1755
rect 4720 1706 4770 1735
rect 4938 1758 4988 1783
rect 4938 1738 4951 1758
rect 4971 1738 4988 1758
rect 4938 1706 4988 1738
rect 5146 1756 5196 1783
rect 5146 1736 5169 1756
rect 5189 1736 5196 1756
rect 5146 1706 5196 1736
rect 6876 1712 6926 1725
rect 7084 1712 7134 1725
rect 7302 1712 7352 1725
rect 356 1635 406 1651
rect 574 1635 624 1651
rect 782 1635 832 1651
rect 4720 1648 4770 1664
rect 4938 1648 4988 1664
rect 5146 1648 5196 1664
rect 3391 1551 3441 1567
rect 3599 1551 3649 1567
rect 3817 1551 3867 1567
rect 7755 1564 7805 1580
rect 7963 1564 8013 1580
rect 8181 1564 8231 1580
rect 1235 1490 1285 1503
rect 1453 1490 1503 1503
rect 1661 1490 1711 1503
rect 3391 1479 3441 1509
rect 3391 1459 3398 1479
rect 3418 1459 3441 1479
rect 3391 1432 3441 1459
rect 3599 1477 3649 1509
rect 3599 1457 3616 1477
rect 3636 1457 3649 1477
rect 3599 1432 3649 1457
rect 3817 1480 3867 1509
rect 3817 1460 3834 1480
rect 3854 1460 3867 1480
rect 5599 1503 5649 1516
rect 5817 1503 5867 1516
rect 6025 1503 6075 1516
rect 3817 1432 3867 1460
rect 1235 1362 1285 1390
rect 1235 1342 1248 1362
rect 1268 1342 1285 1362
rect 1235 1313 1285 1342
rect 1453 1365 1503 1390
rect 1453 1345 1466 1365
rect 1486 1345 1503 1365
rect 1453 1313 1503 1345
rect 1661 1363 1711 1390
rect 1661 1343 1684 1363
rect 1704 1343 1711 1363
rect 1661 1313 1711 1343
rect 2594 1323 2644 1339
rect 2802 1323 2852 1339
rect 3020 1323 3070 1339
rect 7755 1492 7805 1522
rect 7755 1472 7762 1492
rect 7782 1472 7805 1492
rect 7755 1445 7805 1472
rect 7963 1490 8013 1522
rect 7963 1470 7980 1490
rect 8000 1470 8013 1490
rect 7963 1445 8013 1470
rect 8181 1493 8231 1522
rect 8181 1473 8198 1493
rect 8218 1473 8231 1493
rect 8181 1445 8231 1473
rect 5599 1375 5649 1403
rect 5599 1355 5612 1375
rect 5632 1355 5649 1375
rect 338 1264 388 1277
rect 556 1264 606 1277
rect 764 1264 814 1277
rect 3391 1319 3441 1332
rect 3599 1319 3649 1332
rect 3817 1319 3867 1332
rect 5599 1326 5649 1355
rect 5817 1378 5867 1403
rect 5817 1358 5830 1378
rect 5850 1358 5867 1378
rect 5817 1326 5867 1358
rect 6025 1376 6075 1403
rect 6025 1356 6048 1376
rect 6068 1356 6075 1376
rect 6025 1326 6075 1356
rect 6958 1336 7008 1352
rect 7166 1336 7216 1352
rect 7384 1336 7434 1352
rect 1235 1255 1285 1271
rect 1453 1255 1503 1271
rect 1661 1255 1711 1271
rect 2594 1251 2644 1281
rect 2594 1231 2601 1251
rect 2621 1231 2644 1251
rect 2594 1204 2644 1231
rect 2802 1249 2852 1281
rect 2802 1229 2819 1249
rect 2839 1229 2852 1249
rect 2802 1204 2852 1229
rect 3020 1252 3070 1281
rect 3020 1232 3037 1252
rect 3057 1232 3070 1252
rect 4702 1277 4752 1290
rect 4920 1277 4970 1290
rect 5128 1277 5178 1290
rect 7755 1332 7805 1345
rect 7963 1332 8013 1345
rect 8181 1332 8231 1345
rect 3020 1204 3070 1232
rect 338 1136 388 1164
rect 338 1116 351 1136
rect 371 1116 388 1136
rect 338 1087 388 1116
rect 556 1139 606 1164
rect 556 1119 569 1139
rect 589 1119 606 1139
rect 556 1087 606 1119
rect 764 1137 814 1164
rect 764 1117 787 1137
rect 807 1117 814 1137
rect 764 1087 814 1117
rect 5599 1268 5649 1284
rect 5817 1268 5867 1284
rect 6025 1268 6075 1284
rect 6958 1264 7008 1294
rect 6958 1244 6965 1264
rect 6985 1244 7008 1264
rect 6958 1217 7008 1244
rect 7166 1262 7216 1294
rect 7166 1242 7183 1262
rect 7203 1242 7216 1262
rect 7166 1217 7216 1242
rect 7384 1265 7434 1294
rect 7384 1245 7401 1265
rect 7421 1245 7434 1265
rect 7384 1217 7434 1245
rect 3392 1139 3442 1155
rect 3600 1139 3650 1155
rect 3818 1139 3868 1155
rect 1136 1080 1186 1093
rect 1354 1080 1404 1093
rect 1562 1080 1612 1093
rect 2594 1091 2644 1104
rect 2802 1091 2852 1104
rect 3020 1091 3070 1104
rect 4702 1149 4752 1177
rect 338 1029 388 1045
rect 556 1029 606 1045
rect 764 1029 814 1045
rect 3392 1067 3442 1097
rect 3392 1047 3399 1067
rect 3419 1047 3442 1067
rect 3392 1020 3442 1047
rect 3600 1065 3650 1097
rect 3600 1045 3617 1065
rect 3637 1045 3650 1065
rect 3600 1020 3650 1045
rect 3818 1068 3868 1097
rect 3818 1048 3835 1068
rect 3855 1048 3868 1068
rect 4702 1129 4715 1149
rect 4735 1129 4752 1149
rect 4702 1100 4752 1129
rect 4920 1152 4970 1177
rect 4920 1132 4933 1152
rect 4953 1132 4970 1152
rect 4920 1100 4970 1132
rect 5128 1150 5178 1177
rect 5128 1130 5151 1150
rect 5171 1130 5178 1150
rect 5128 1100 5178 1130
rect 7756 1152 7806 1168
rect 7964 1152 8014 1168
rect 8182 1152 8232 1168
rect 3818 1020 3868 1048
rect 5500 1093 5550 1106
rect 5718 1093 5768 1106
rect 5926 1093 5976 1106
rect 6958 1104 7008 1117
rect 7166 1104 7216 1117
rect 7384 1104 7434 1117
rect 4702 1042 4752 1058
rect 4920 1042 4970 1058
rect 5128 1042 5178 1058
rect 1136 952 1186 980
rect 1136 932 1149 952
rect 1169 932 1186 952
rect 1136 903 1186 932
rect 1354 955 1404 980
rect 1354 935 1367 955
rect 1387 935 1404 955
rect 1354 903 1404 935
rect 1562 953 1612 980
rect 1562 933 1585 953
rect 1605 933 1612 953
rect 1562 903 1612 933
rect 7756 1080 7806 1110
rect 7756 1060 7763 1080
rect 7783 1060 7806 1080
rect 7756 1033 7806 1060
rect 7964 1078 8014 1110
rect 7964 1058 7981 1078
rect 8001 1058 8014 1078
rect 7964 1033 8014 1058
rect 8182 1081 8232 1110
rect 8182 1061 8199 1081
rect 8219 1061 8232 1081
rect 8182 1033 8232 1061
rect 5500 965 5550 993
rect 3392 907 3442 920
rect 3600 907 3650 920
rect 3818 907 3868 920
rect 5500 945 5513 965
rect 5533 945 5550 965
rect 5500 916 5550 945
rect 5718 968 5768 993
rect 5718 948 5731 968
rect 5751 948 5768 968
rect 5718 916 5768 948
rect 5926 966 5976 993
rect 5926 946 5949 966
rect 5969 946 5976 966
rect 5926 916 5976 946
rect 7756 920 7806 933
rect 7964 920 8014 933
rect 8182 920 8232 933
rect 339 852 389 865
rect 557 852 607 865
rect 765 852 815 865
rect 1136 845 1186 861
rect 1354 845 1404 861
rect 1562 845 1612 861
rect 4703 865 4753 878
rect 4921 865 4971 878
rect 5129 865 5179 878
rect 339 724 389 752
rect 339 704 352 724
rect 372 704 389 724
rect 339 675 389 704
rect 557 727 607 752
rect 557 707 570 727
rect 590 707 607 727
rect 557 675 607 707
rect 765 725 815 752
rect 5500 858 5550 874
rect 5718 858 5768 874
rect 5926 858 5976 874
rect 765 705 788 725
rect 808 705 815 725
rect 765 675 815 705
rect 4703 737 4753 765
rect 4703 717 4716 737
rect 4736 717 4753 737
rect 4703 688 4753 717
rect 4921 740 4971 765
rect 4921 720 4934 740
rect 4954 720 4971 740
rect 4921 688 4971 720
rect 5129 738 5179 765
rect 5129 718 5152 738
rect 5172 718 5179 738
rect 5129 688 5179 718
rect 339 617 389 633
rect 557 617 607 633
rect 765 617 815 633
rect 4703 630 4753 646
rect 4921 630 4971 646
rect 5129 630 5179 646
rect 5916 289 5966 302
rect 6134 289 6184 302
rect 6342 289 6392 302
rect 1552 276 1602 289
rect 1770 276 1820 289
rect 1978 276 2028 289
rect 4041 202 4091 215
rect 4259 202 4309 215
rect 4467 202 4517 215
rect 1552 148 1602 176
rect 1552 128 1565 148
rect 1585 128 1602 148
rect 1552 99 1602 128
rect 1770 151 1820 176
rect 1770 131 1783 151
rect 1803 131 1820 151
rect 1770 99 1820 131
rect 1978 149 2028 176
rect 1978 129 2001 149
rect 2021 129 2028 149
rect 1978 99 2028 129
rect 5916 161 5966 189
rect 5916 141 5929 161
rect 5949 141 5966 161
rect 5916 112 5966 141
rect 6134 164 6184 189
rect 6134 144 6147 164
rect 6167 144 6184 164
rect 6134 112 6184 144
rect 6342 162 6392 189
rect 6342 142 6365 162
rect 6385 142 6392 162
rect 6342 112 6392 142
rect 4041 74 4091 102
rect 1552 41 1602 57
rect 1770 41 1820 57
rect 1978 41 2028 57
rect 4041 54 4054 74
rect 4074 54 4091 74
rect 4041 25 4091 54
rect 4259 77 4309 102
rect 4259 57 4272 77
rect 4292 57 4309 77
rect 4259 25 4309 57
rect 4467 75 4517 102
rect 4467 55 4490 75
rect 4510 55 4517 75
rect 4467 25 4517 55
rect 5916 54 5966 70
rect 6134 54 6184 70
rect 6342 54 6392 70
rect 4041 -33 4091 -17
rect 4259 -33 4309 -17
rect 4467 -33 4517 -17
<< polycont >>
rect 3525 8585 3545 8605
rect 3743 8583 3763 8603
rect 3961 8586 3981 8606
rect 7889 8598 7909 8618
rect 8107 8596 8127 8616
rect 8325 8599 8345 8619
rect 2728 8357 2748 8377
rect 2946 8355 2966 8375
rect 3164 8358 3184 8378
rect 478 8242 498 8262
rect 696 8245 716 8265
rect 914 8243 934 8263
rect 7092 8370 7112 8390
rect 7310 8368 7330 8388
rect 7528 8371 7548 8391
rect 3526 8173 3546 8193
rect 3744 8171 3764 8191
rect 3962 8174 3982 8194
rect 4842 8255 4862 8275
rect 5060 8258 5080 8278
rect 5278 8256 5298 8276
rect 1276 8058 1296 8078
rect 1494 8061 1514 8081
rect 1712 8059 1732 8079
rect 7890 8186 7910 8206
rect 8108 8184 8128 8204
rect 8326 8187 8346 8207
rect 5640 8071 5660 8091
rect 5858 8074 5878 8094
rect 6076 8072 6096 8092
rect 2629 7947 2649 7967
rect 2847 7945 2867 7965
rect 3065 7948 3085 7968
rect 479 7830 499 7850
rect 697 7833 717 7853
rect 915 7831 935 7851
rect 6993 7960 7013 7980
rect 7211 7958 7231 7978
rect 7429 7961 7449 7981
rect 4843 7843 4863 7863
rect 5061 7846 5081 7866
rect 5279 7844 5299 7864
rect 3508 7567 3528 7587
rect 3726 7565 3746 7585
rect 3944 7568 3964 7588
rect 1358 7450 1378 7470
rect 1576 7453 1596 7473
rect 1794 7451 1814 7471
rect 7872 7580 7892 7600
rect 8090 7578 8110 7598
rect 8308 7581 8328 7601
rect 5722 7463 5742 7483
rect 5940 7466 5960 7486
rect 6158 7464 6178 7484
rect 2711 7339 2731 7359
rect 2929 7337 2949 7357
rect 3147 7340 3167 7360
rect 461 7224 481 7244
rect 679 7227 699 7247
rect 897 7225 917 7245
rect 7075 7352 7095 7372
rect 7293 7350 7313 7370
rect 7511 7353 7531 7373
rect 3509 7155 3529 7175
rect 3727 7153 3747 7173
rect 3945 7156 3965 7176
rect 4825 7237 4845 7257
rect 5043 7240 5063 7260
rect 5261 7238 5281 7258
rect 1259 7040 1279 7060
rect 1477 7043 1497 7063
rect 1695 7041 1715 7061
rect 7873 7168 7893 7188
rect 8091 7166 8111 7186
rect 8309 7169 8329 7189
rect 5623 7053 5643 7073
rect 5841 7056 5861 7076
rect 6059 7054 6079 7074
rect 2546 6931 2566 6951
rect 2764 6929 2784 6949
rect 2982 6932 3002 6952
rect 462 6812 482 6832
rect 680 6815 700 6835
rect 898 6813 918 6833
rect 6910 6944 6930 6964
rect 7128 6942 7148 6962
rect 7346 6945 7366 6965
rect 4826 6825 4846 6845
rect 5044 6828 5064 6848
rect 5262 6826 5282 6846
rect 3488 6549 3508 6569
rect 3706 6547 3726 6567
rect 3924 6550 3944 6570
rect 1404 6430 1424 6450
rect 1622 6433 1642 6453
rect 1840 6431 1860 6451
rect 7852 6562 7872 6582
rect 8070 6560 8090 6580
rect 8288 6563 8308 6583
rect 5768 6443 5788 6463
rect 5986 6446 6006 6466
rect 6204 6444 6224 6464
rect 2691 6321 2711 6341
rect 2909 6319 2929 6339
rect 3127 6322 3147 6342
rect 441 6206 461 6226
rect 659 6209 679 6229
rect 877 6207 897 6227
rect 7055 6334 7075 6354
rect 7273 6332 7293 6352
rect 7491 6335 7511 6355
rect 3489 6137 3509 6157
rect 3707 6135 3727 6155
rect 3925 6138 3945 6158
rect 4805 6219 4825 6239
rect 5023 6222 5043 6242
rect 5241 6220 5261 6240
rect 1239 6022 1259 6042
rect 1457 6025 1477 6045
rect 1675 6023 1695 6043
rect 7853 6150 7873 6170
rect 8071 6148 8091 6168
rect 8289 6151 8309 6171
rect 5603 6035 5623 6055
rect 5821 6038 5841 6058
rect 6039 6036 6059 6056
rect 2592 5911 2612 5931
rect 2810 5909 2830 5929
rect 3028 5912 3048 5932
rect 442 5794 462 5814
rect 660 5797 680 5817
rect 878 5795 898 5815
rect 6956 5924 6976 5944
rect 7174 5922 7194 5942
rect 7392 5925 7412 5945
rect 4806 5807 4826 5827
rect 5024 5810 5044 5830
rect 5242 5808 5262 5828
rect 3471 5531 3491 5551
rect 3689 5529 3709 5549
rect 3907 5532 3927 5552
rect 1321 5414 1341 5434
rect 1539 5417 1559 5437
rect 1757 5415 1777 5435
rect 7835 5544 7855 5564
rect 8053 5542 8073 5562
rect 8271 5545 8291 5565
rect 5685 5427 5705 5447
rect 5903 5430 5923 5450
rect 6121 5428 6141 5448
rect 2674 5303 2694 5323
rect 2892 5301 2912 5321
rect 3110 5304 3130 5324
rect 424 5188 444 5208
rect 642 5191 662 5211
rect 860 5189 880 5209
rect 7038 5316 7058 5336
rect 7256 5314 7276 5334
rect 7474 5317 7494 5337
rect 3472 5119 3492 5139
rect 3690 5117 3710 5137
rect 3908 5120 3928 5140
rect 4788 5201 4808 5221
rect 5006 5204 5026 5224
rect 5224 5202 5244 5222
rect 1222 5004 1242 5024
rect 1440 5007 1460 5027
rect 1658 5005 1678 5025
rect 7836 5132 7856 5152
rect 8054 5130 8074 5150
rect 8272 5133 8292 5153
rect 5586 5017 5606 5037
rect 5804 5020 5824 5040
rect 6022 5018 6042 5038
rect 2370 4897 2390 4917
rect 2588 4895 2608 4915
rect 2806 4898 2826 4918
rect 425 4776 445 4796
rect 643 4779 663 4799
rect 861 4777 881 4797
rect 6734 4910 6754 4930
rect 6952 4908 6972 4928
rect 7170 4911 7190 4931
rect 4789 4789 4809 4809
rect 5007 4792 5027 4812
rect 5225 4790 5245 4810
rect 3452 4513 3472 4533
rect 3670 4511 3690 4531
rect 3888 4514 3908 4534
rect 1507 4392 1527 4412
rect 1725 4395 1745 4415
rect 1943 4393 1963 4413
rect 7816 4526 7836 4546
rect 8034 4524 8054 4544
rect 8252 4527 8272 4547
rect 5871 4405 5891 4425
rect 6089 4408 6109 4428
rect 6307 4406 6327 4426
rect 2655 4285 2675 4305
rect 2873 4283 2893 4303
rect 3091 4286 3111 4306
rect 405 4170 425 4190
rect 623 4173 643 4193
rect 841 4171 861 4191
rect 7019 4298 7039 4318
rect 7237 4296 7257 4316
rect 7455 4299 7475 4319
rect 3453 4101 3473 4121
rect 3671 4099 3691 4119
rect 3889 4102 3909 4122
rect 4769 4183 4789 4203
rect 4987 4186 5007 4206
rect 5205 4184 5225 4204
rect 1203 3986 1223 4006
rect 1421 3989 1441 4009
rect 1639 3987 1659 4007
rect 7817 4114 7837 4134
rect 8035 4112 8055 4132
rect 8253 4115 8273 4135
rect 5567 3999 5587 4019
rect 5785 4002 5805 4022
rect 6003 4000 6023 4020
rect 2556 3875 2576 3895
rect 2774 3873 2794 3893
rect 2992 3876 3012 3896
rect 406 3758 426 3778
rect 624 3761 644 3781
rect 842 3759 862 3779
rect 6920 3888 6940 3908
rect 7138 3886 7158 3906
rect 7356 3889 7376 3909
rect 4770 3771 4790 3791
rect 4988 3774 5008 3794
rect 5206 3772 5226 3792
rect 3435 3495 3455 3515
rect 3653 3493 3673 3513
rect 3871 3496 3891 3516
rect 1285 3378 1305 3398
rect 1503 3381 1523 3401
rect 1721 3379 1741 3399
rect 7799 3508 7819 3528
rect 8017 3506 8037 3526
rect 8235 3509 8255 3529
rect 5649 3391 5669 3411
rect 5867 3394 5887 3414
rect 6085 3392 6105 3412
rect 2638 3267 2658 3287
rect 2856 3265 2876 3285
rect 3074 3268 3094 3288
rect 388 3152 408 3172
rect 606 3155 626 3175
rect 824 3153 844 3173
rect 7002 3280 7022 3300
rect 7220 3278 7240 3298
rect 7438 3281 7458 3301
rect 3436 3083 3456 3103
rect 3654 3081 3674 3101
rect 3872 3084 3892 3104
rect 4752 3165 4772 3185
rect 4970 3168 4990 3188
rect 5188 3166 5208 3186
rect 1186 2968 1206 2988
rect 1404 2971 1424 2991
rect 1622 2969 1642 2989
rect 7800 3096 7820 3116
rect 8018 3094 8038 3114
rect 8236 3097 8256 3117
rect 5550 2981 5570 3001
rect 5768 2984 5788 3004
rect 5986 2982 6006 3002
rect 2473 2859 2493 2879
rect 2691 2857 2711 2877
rect 2909 2860 2929 2880
rect 389 2740 409 2760
rect 607 2743 627 2763
rect 825 2741 845 2761
rect 6837 2872 6857 2892
rect 7055 2870 7075 2890
rect 7273 2873 7293 2893
rect 4753 2753 4773 2773
rect 4971 2756 4991 2776
rect 5189 2754 5209 2774
rect 3415 2477 3435 2497
rect 3633 2475 3653 2495
rect 3851 2478 3871 2498
rect 1331 2358 1351 2378
rect 1549 2361 1569 2381
rect 1767 2359 1787 2379
rect 7779 2490 7799 2510
rect 7997 2488 8017 2508
rect 8215 2491 8235 2511
rect 5695 2371 5715 2391
rect 5913 2374 5933 2394
rect 6131 2372 6151 2392
rect 2618 2249 2638 2269
rect 2836 2247 2856 2267
rect 3054 2250 3074 2270
rect 368 2134 388 2154
rect 586 2137 606 2157
rect 804 2135 824 2155
rect 6982 2262 7002 2282
rect 7200 2260 7220 2280
rect 7418 2263 7438 2283
rect 3416 2065 3436 2085
rect 3634 2063 3654 2083
rect 3852 2066 3872 2086
rect 4732 2147 4752 2167
rect 4950 2150 4970 2170
rect 5168 2148 5188 2168
rect 1166 1950 1186 1970
rect 1384 1953 1404 1973
rect 1602 1951 1622 1971
rect 7780 2078 7800 2098
rect 7998 2076 8018 2096
rect 8216 2079 8236 2099
rect 5530 1963 5550 1983
rect 5748 1966 5768 1986
rect 5966 1964 5986 1984
rect 2519 1839 2539 1859
rect 2737 1837 2757 1857
rect 2955 1840 2975 1860
rect 369 1722 389 1742
rect 587 1725 607 1745
rect 805 1723 825 1743
rect 6883 1852 6903 1872
rect 7101 1850 7121 1870
rect 7319 1853 7339 1873
rect 4733 1735 4753 1755
rect 4951 1738 4971 1758
rect 5169 1736 5189 1756
rect 3398 1459 3418 1479
rect 3616 1457 3636 1477
rect 3834 1460 3854 1480
rect 1248 1342 1268 1362
rect 1466 1345 1486 1365
rect 1684 1343 1704 1363
rect 7762 1472 7782 1492
rect 7980 1470 8000 1490
rect 8198 1473 8218 1493
rect 5612 1355 5632 1375
rect 5830 1358 5850 1378
rect 6048 1356 6068 1376
rect 2601 1231 2621 1251
rect 2819 1229 2839 1249
rect 3037 1232 3057 1252
rect 351 1116 371 1136
rect 569 1119 589 1139
rect 787 1117 807 1137
rect 6965 1244 6985 1264
rect 7183 1242 7203 1262
rect 7401 1245 7421 1265
rect 3399 1047 3419 1067
rect 3617 1045 3637 1065
rect 3835 1048 3855 1068
rect 4715 1129 4735 1149
rect 4933 1132 4953 1152
rect 5151 1130 5171 1150
rect 1149 932 1169 952
rect 1367 935 1387 955
rect 1585 933 1605 953
rect 7763 1060 7783 1080
rect 7981 1058 8001 1078
rect 8199 1061 8219 1081
rect 5513 945 5533 965
rect 5731 948 5751 968
rect 5949 946 5969 966
rect 352 704 372 724
rect 570 707 590 727
rect 788 705 808 725
rect 4716 717 4736 737
rect 4934 720 4954 740
rect 5152 718 5172 738
rect 1565 128 1585 148
rect 1783 131 1803 151
rect 2001 129 2021 149
rect 5929 141 5949 161
rect 6147 144 6167 164
rect 6365 142 6385 162
rect 4054 54 4074 74
rect 4272 57 4292 77
rect 4490 55 4510 75
<< ndiffres >>
rect 4181 8670 4238 8689
rect 4181 8652 4199 8670
rect 4217 8667 4238 8670
rect 4217 8652 4332 8667
rect 240 8612 301 8628
rect 145 8608 301 8612
rect 145 8590 263 8608
rect 281 8590 301 8608
rect 145 8569 301 8590
rect 145 8568 245 8569
rect 146 8532 188 8568
rect 4181 8629 4332 8652
rect 8545 8683 8602 8702
rect 8545 8665 8563 8683
rect 8581 8680 8602 8683
rect 8581 8665 8696 8680
rect 4290 8593 4332 8629
rect 4604 8625 4665 8641
rect 4509 8621 4665 8625
rect 4509 8603 4627 8621
rect 4645 8603 4665 8621
rect 4233 8592 4333 8593
rect 4177 8571 4333 8592
rect 4509 8582 4665 8603
rect 4509 8581 4609 8582
rect 146 8509 297 8532
rect 146 8494 261 8509
rect 240 8491 261 8494
rect 279 8491 297 8509
rect 240 8472 297 8491
rect 4177 8553 4197 8571
rect 4215 8553 4333 8571
rect 4177 8549 4333 8553
rect 4177 8533 4238 8549
rect 4510 8545 4552 8581
rect 8545 8642 8696 8665
rect 8654 8606 8696 8642
rect 8597 8605 8697 8606
rect 8541 8584 8697 8605
rect 4510 8522 4661 8545
rect 4510 8507 4625 8522
rect 4604 8504 4625 8507
rect 4643 8504 4661 8522
rect 4604 8485 4661 8504
rect 4174 8452 4231 8471
rect 8541 8566 8561 8584
rect 8579 8566 8697 8584
rect 8541 8562 8697 8566
rect 8541 8546 8602 8562
rect 4174 8434 4192 8452
rect 4210 8449 4231 8452
rect 4210 8434 4325 8449
rect 4174 8411 4325 8434
rect 8538 8465 8595 8484
rect 8538 8447 8556 8465
rect 8574 8462 8595 8465
rect 8574 8447 8689 8462
rect 8538 8424 8689 8447
rect 235 8288 296 8304
rect 4283 8375 4325 8411
rect 4226 8374 4326 8375
rect 4170 8353 4326 8374
rect 4170 8335 4190 8353
rect 4208 8335 4326 8353
rect 4170 8331 4326 8335
rect 140 8284 296 8288
rect 140 8266 258 8284
rect 276 8266 296 8284
rect 140 8245 296 8266
rect 140 8244 240 8245
rect 141 8208 183 8244
rect 4170 8315 4231 8331
rect 4599 8301 4660 8317
rect 8647 8388 8689 8424
rect 8590 8387 8690 8388
rect 8534 8366 8690 8387
rect 8534 8348 8554 8366
rect 8572 8348 8690 8366
rect 8534 8344 8690 8348
rect 4504 8297 4660 8301
rect 4168 8269 4225 8288
rect 141 8185 292 8208
rect 141 8170 256 8185
rect 235 8167 256 8170
rect 274 8167 292 8185
rect 4168 8251 4186 8269
rect 4204 8266 4225 8269
rect 4504 8279 4622 8297
rect 4640 8279 4660 8297
rect 4204 8251 4319 8266
rect 4504 8258 4660 8279
rect 4504 8257 4604 8258
rect 4168 8228 4319 8251
rect 235 8148 292 8167
rect 229 8105 290 8121
rect 4277 8192 4319 8228
rect 4505 8221 4547 8257
rect 8534 8328 8595 8344
rect 8532 8282 8589 8301
rect 4505 8198 4656 8221
rect 4220 8191 4320 8192
rect 4164 8170 4320 8191
rect 4505 8183 4620 8198
rect 4164 8152 4184 8170
rect 4202 8152 4320 8170
rect 4599 8180 4620 8183
rect 4638 8180 4656 8198
rect 8532 8264 8550 8282
rect 8568 8279 8589 8282
rect 8568 8264 8683 8279
rect 8532 8241 8683 8264
rect 4599 8161 4656 8180
rect 4164 8148 4320 8152
rect 134 8101 290 8105
rect 134 8083 252 8101
rect 270 8083 290 8101
rect 134 8062 290 8083
rect 134 8061 234 8062
rect 135 8025 177 8061
rect 4164 8132 4225 8148
rect 4593 8118 4654 8134
rect 8641 8205 8683 8241
rect 8584 8204 8684 8205
rect 8528 8183 8684 8204
rect 8528 8165 8548 8183
rect 8566 8165 8684 8183
rect 8528 8161 8684 8165
rect 4498 8114 4654 8118
rect 4498 8096 4616 8114
rect 4634 8096 4654 8114
rect 4498 8075 4654 8096
rect 4498 8074 4598 8075
rect 135 8002 286 8025
rect 135 7987 250 8002
rect 229 7984 250 7987
rect 268 7984 286 8002
rect 229 7965 286 7984
rect 4499 8038 4541 8074
rect 8528 8145 8589 8161
rect 4499 8015 4650 8038
rect 4499 8000 4614 8015
rect 4593 7997 4614 8000
rect 4632 7997 4650 8015
rect 222 7887 283 7903
rect 127 7883 283 7887
rect 127 7865 245 7883
rect 263 7865 283 7883
rect 4593 7978 4650 7997
rect 4163 7945 4220 7964
rect 4163 7927 4181 7945
rect 4199 7942 4220 7945
rect 4199 7927 4314 7942
rect 127 7844 283 7865
rect 127 7843 227 7844
rect 128 7807 170 7843
rect 128 7784 279 7807
rect 4163 7904 4314 7927
rect 4272 7868 4314 7904
rect 4586 7900 4647 7916
rect 4491 7896 4647 7900
rect 4491 7878 4609 7896
rect 4627 7878 4647 7896
rect 8527 7958 8584 7977
rect 8527 7940 8545 7958
rect 8563 7955 8584 7958
rect 8563 7940 8678 7955
rect 4215 7867 4315 7868
rect 4159 7846 4315 7867
rect 4491 7857 4647 7878
rect 4491 7856 4591 7857
rect 4159 7828 4179 7846
rect 4197 7828 4315 7846
rect 4159 7824 4315 7828
rect 4159 7808 4220 7824
rect 4492 7820 4534 7856
rect 128 7769 243 7784
rect 222 7766 243 7769
rect 261 7766 279 7784
rect 222 7747 279 7766
rect 4492 7797 4643 7820
rect 8527 7917 8678 7940
rect 8636 7881 8678 7917
rect 8579 7880 8679 7881
rect 8523 7859 8679 7880
rect 8523 7841 8543 7859
rect 8561 7841 8679 7859
rect 8523 7837 8679 7841
rect 8523 7821 8584 7837
rect 4492 7782 4607 7797
rect 4586 7779 4607 7782
rect 4625 7779 4643 7797
rect 4586 7760 4643 7779
rect 4164 7652 4221 7671
rect 4164 7634 4182 7652
rect 4200 7649 4221 7652
rect 4200 7634 4315 7649
rect 223 7594 284 7610
rect 128 7590 284 7594
rect 128 7572 246 7590
rect 264 7572 284 7590
rect 128 7551 284 7572
rect 128 7550 228 7551
rect 129 7514 171 7550
rect 129 7491 280 7514
rect 4164 7611 4315 7634
rect 8528 7665 8585 7684
rect 8528 7647 8546 7665
rect 8564 7662 8585 7665
rect 8564 7647 8679 7662
rect 4273 7575 4315 7611
rect 4587 7607 4648 7623
rect 4492 7603 4648 7607
rect 4492 7585 4610 7603
rect 4628 7585 4648 7603
rect 4216 7574 4316 7575
rect 4160 7553 4316 7574
rect 4492 7564 4648 7585
rect 4492 7563 4592 7564
rect 129 7476 244 7491
rect 223 7473 244 7476
rect 262 7473 280 7491
rect 223 7454 280 7473
rect 4160 7535 4180 7553
rect 4198 7535 4316 7553
rect 4160 7531 4316 7535
rect 4160 7515 4221 7531
rect 4493 7527 4535 7563
rect 4493 7504 4644 7527
rect 8528 7624 8679 7647
rect 8637 7588 8679 7624
rect 8580 7587 8680 7588
rect 8524 7566 8680 7587
rect 4493 7489 4608 7504
rect 4587 7486 4608 7489
rect 4626 7486 4644 7504
rect 4587 7467 4644 7486
rect 4157 7434 4214 7453
rect 8524 7548 8544 7566
rect 8562 7548 8680 7566
rect 8524 7544 8680 7548
rect 8524 7528 8585 7544
rect 4157 7416 4175 7434
rect 4193 7431 4214 7434
rect 4193 7416 4308 7431
rect 4157 7393 4308 7416
rect 218 7270 279 7286
rect 4266 7357 4308 7393
rect 8521 7447 8578 7466
rect 8521 7429 8539 7447
rect 8557 7444 8578 7447
rect 8557 7429 8672 7444
rect 8521 7406 8672 7429
rect 4209 7356 4309 7357
rect 4153 7335 4309 7356
rect 4153 7317 4173 7335
rect 4191 7317 4309 7335
rect 4153 7313 4309 7317
rect 123 7266 279 7270
rect 123 7248 241 7266
rect 259 7248 279 7266
rect 123 7227 279 7248
rect 123 7226 223 7227
rect 124 7190 166 7226
rect 4153 7297 4214 7313
rect 4582 7283 4643 7299
rect 8630 7370 8672 7406
rect 8573 7369 8673 7370
rect 8517 7348 8673 7369
rect 8517 7330 8537 7348
rect 8555 7330 8673 7348
rect 8517 7326 8673 7330
rect 4487 7279 4643 7283
rect 4151 7251 4208 7270
rect 124 7167 275 7190
rect 124 7152 239 7167
rect 218 7149 239 7152
rect 257 7149 275 7167
rect 4151 7233 4169 7251
rect 4187 7248 4208 7251
rect 4487 7261 4605 7279
rect 4623 7261 4643 7279
rect 4187 7233 4302 7248
rect 4487 7240 4643 7261
rect 4487 7239 4587 7240
rect 4151 7210 4302 7233
rect 218 7130 275 7149
rect 212 7087 273 7103
rect 4260 7174 4302 7210
rect 4488 7203 4530 7239
rect 8517 7310 8578 7326
rect 8515 7264 8572 7283
rect 4488 7180 4639 7203
rect 4203 7173 4303 7174
rect 4147 7152 4303 7173
rect 4488 7165 4603 7180
rect 4147 7134 4167 7152
rect 4185 7134 4303 7152
rect 4582 7162 4603 7165
rect 4621 7162 4639 7180
rect 8515 7246 8533 7264
rect 8551 7261 8572 7264
rect 8551 7246 8666 7261
rect 8515 7223 8666 7246
rect 4582 7143 4639 7162
rect 4147 7130 4303 7134
rect 117 7083 273 7087
rect 117 7065 235 7083
rect 253 7065 273 7083
rect 117 7044 273 7065
rect 117 7043 217 7044
rect 118 7007 160 7043
rect 4147 7114 4208 7130
rect 4576 7100 4637 7116
rect 8624 7187 8666 7223
rect 8567 7186 8667 7187
rect 8511 7165 8667 7186
rect 8511 7147 8531 7165
rect 8549 7147 8667 7165
rect 8511 7143 8667 7147
rect 4481 7096 4637 7100
rect 4481 7078 4599 7096
rect 4617 7078 4637 7096
rect 4481 7057 4637 7078
rect 4481 7056 4581 7057
rect 118 6984 269 7007
rect 118 6969 233 6984
rect 212 6966 233 6969
rect 251 6966 269 6984
rect 212 6947 269 6966
rect 4482 7020 4524 7056
rect 8511 7127 8572 7143
rect 4482 6997 4633 7020
rect 4482 6982 4597 6997
rect 205 6869 266 6885
rect 110 6865 266 6869
rect 110 6847 228 6865
rect 246 6847 266 6865
rect 4576 6979 4597 6982
rect 4615 6979 4633 6997
rect 4576 6960 4633 6979
rect 4146 6927 4203 6946
rect 4146 6909 4164 6927
rect 4182 6924 4203 6927
rect 4182 6909 4297 6924
rect 110 6826 266 6847
rect 110 6825 210 6826
rect 111 6789 153 6825
rect 111 6766 262 6789
rect 4146 6886 4297 6909
rect 4255 6850 4297 6886
rect 4569 6882 4630 6898
rect 4474 6878 4630 6882
rect 4474 6860 4592 6878
rect 4610 6860 4630 6878
rect 8510 6940 8567 6959
rect 8510 6922 8528 6940
rect 8546 6937 8567 6940
rect 8546 6922 8661 6937
rect 4198 6849 4298 6850
rect 4142 6828 4298 6849
rect 4474 6839 4630 6860
rect 4474 6838 4574 6839
rect 4142 6810 4162 6828
rect 4180 6810 4298 6828
rect 4142 6806 4298 6810
rect 4142 6790 4203 6806
rect 4475 6802 4517 6838
rect 111 6751 226 6766
rect 205 6748 226 6751
rect 244 6748 262 6766
rect 205 6729 262 6748
rect 4475 6779 4626 6802
rect 8510 6899 8661 6922
rect 8619 6863 8661 6899
rect 8562 6862 8662 6863
rect 8506 6841 8662 6862
rect 8506 6823 8526 6841
rect 8544 6823 8662 6841
rect 8506 6819 8662 6823
rect 8506 6803 8567 6819
rect 4475 6764 4590 6779
rect 4569 6761 4590 6764
rect 4608 6761 4626 6779
rect 4569 6742 4626 6761
rect 4144 6634 4201 6653
rect 4144 6616 4162 6634
rect 4180 6631 4201 6634
rect 4180 6616 4295 6631
rect 203 6576 264 6592
rect 108 6572 264 6576
rect 108 6554 226 6572
rect 244 6554 264 6572
rect 108 6533 264 6554
rect 108 6532 208 6533
rect 109 6496 151 6532
rect 109 6473 260 6496
rect 4144 6593 4295 6616
rect 8508 6647 8565 6666
rect 8508 6629 8526 6647
rect 8544 6644 8565 6647
rect 8544 6629 8659 6644
rect 4253 6557 4295 6593
rect 4567 6589 4628 6605
rect 4472 6585 4628 6589
rect 4472 6567 4590 6585
rect 4608 6567 4628 6585
rect 4196 6556 4296 6557
rect 4140 6535 4296 6556
rect 4472 6546 4628 6567
rect 4472 6545 4572 6546
rect 109 6458 224 6473
rect 203 6455 224 6458
rect 242 6455 260 6473
rect 203 6436 260 6455
rect 4140 6517 4160 6535
rect 4178 6517 4296 6535
rect 4140 6513 4296 6517
rect 4140 6497 4201 6513
rect 4473 6509 4515 6545
rect 4473 6486 4624 6509
rect 8508 6606 8659 6629
rect 8617 6570 8659 6606
rect 8560 6569 8660 6570
rect 8504 6548 8660 6569
rect 4473 6471 4588 6486
rect 4567 6468 4588 6471
rect 4606 6468 4624 6486
rect 4567 6449 4624 6468
rect 4137 6416 4194 6435
rect 4137 6398 4155 6416
rect 4173 6413 4194 6416
rect 8504 6530 8524 6548
rect 8542 6530 8660 6548
rect 8504 6526 8660 6530
rect 8504 6510 8565 6526
rect 4173 6398 4288 6413
rect 4137 6375 4288 6398
rect 198 6252 259 6268
rect 4246 6339 4288 6375
rect 8501 6429 8558 6448
rect 8501 6411 8519 6429
rect 8537 6426 8558 6429
rect 8537 6411 8652 6426
rect 8501 6388 8652 6411
rect 4189 6338 4289 6339
rect 4133 6317 4289 6338
rect 4133 6299 4153 6317
rect 4171 6299 4289 6317
rect 4133 6295 4289 6299
rect 103 6248 259 6252
rect 103 6230 221 6248
rect 239 6230 259 6248
rect 103 6209 259 6230
rect 103 6208 203 6209
rect 104 6172 146 6208
rect 4133 6279 4194 6295
rect 4562 6265 4623 6281
rect 8610 6352 8652 6388
rect 8553 6351 8653 6352
rect 8497 6330 8653 6351
rect 8497 6312 8517 6330
rect 8535 6312 8653 6330
rect 8497 6308 8653 6312
rect 4467 6261 4623 6265
rect 4131 6233 4188 6252
rect 104 6149 255 6172
rect 104 6134 219 6149
rect 198 6131 219 6134
rect 237 6131 255 6149
rect 4131 6215 4149 6233
rect 4167 6230 4188 6233
rect 4467 6243 4585 6261
rect 4603 6243 4623 6261
rect 4167 6215 4282 6230
rect 4467 6222 4623 6243
rect 4467 6221 4567 6222
rect 4131 6192 4282 6215
rect 198 6112 255 6131
rect 192 6069 253 6085
rect 4240 6156 4282 6192
rect 4468 6185 4510 6221
rect 8497 6292 8558 6308
rect 8495 6246 8552 6265
rect 4468 6162 4619 6185
rect 4183 6155 4283 6156
rect 4127 6134 4283 6155
rect 4468 6147 4583 6162
rect 4127 6116 4147 6134
rect 4165 6116 4283 6134
rect 4562 6144 4583 6147
rect 4601 6144 4619 6162
rect 8495 6228 8513 6246
rect 8531 6243 8552 6246
rect 8531 6228 8646 6243
rect 8495 6205 8646 6228
rect 4562 6125 4619 6144
rect 4127 6112 4283 6116
rect 97 6065 253 6069
rect 97 6047 215 6065
rect 233 6047 253 6065
rect 97 6026 253 6047
rect 97 6025 197 6026
rect 98 5989 140 6025
rect 4127 6096 4188 6112
rect 4556 6082 4617 6098
rect 8604 6169 8646 6205
rect 8547 6168 8647 6169
rect 8491 6147 8647 6168
rect 8491 6129 8511 6147
rect 8529 6129 8647 6147
rect 8491 6125 8647 6129
rect 4461 6078 4617 6082
rect 4461 6060 4579 6078
rect 4597 6060 4617 6078
rect 4461 6039 4617 6060
rect 4461 6038 4561 6039
rect 98 5966 249 5989
rect 98 5951 213 5966
rect 192 5948 213 5951
rect 231 5948 249 5966
rect 192 5929 249 5948
rect 4462 6002 4504 6038
rect 8491 6109 8552 6125
rect 4462 5979 4613 6002
rect 4462 5964 4577 5979
rect 4556 5961 4577 5964
rect 4595 5961 4613 5979
rect 185 5851 246 5867
rect 90 5847 246 5851
rect 90 5829 208 5847
rect 226 5829 246 5847
rect 4556 5942 4613 5961
rect 4126 5909 4183 5928
rect 4126 5891 4144 5909
rect 4162 5906 4183 5909
rect 4162 5891 4277 5906
rect 90 5808 246 5829
rect 90 5807 190 5808
rect 91 5771 133 5807
rect 91 5748 242 5771
rect 4126 5868 4277 5891
rect 4235 5832 4277 5868
rect 4549 5864 4610 5880
rect 4454 5860 4610 5864
rect 4454 5842 4572 5860
rect 4590 5842 4610 5860
rect 8490 5922 8547 5941
rect 8490 5904 8508 5922
rect 8526 5919 8547 5922
rect 8526 5904 8641 5919
rect 4178 5831 4278 5832
rect 4122 5810 4278 5831
rect 4454 5821 4610 5842
rect 4454 5820 4554 5821
rect 4122 5792 4142 5810
rect 4160 5792 4278 5810
rect 4122 5788 4278 5792
rect 4122 5772 4183 5788
rect 4455 5784 4497 5820
rect 91 5733 206 5748
rect 185 5730 206 5733
rect 224 5730 242 5748
rect 185 5711 242 5730
rect 4455 5761 4606 5784
rect 8490 5881 8641 5904
rect 8599 5845 8641 5881
rect 8542 5844 8642 5845
rect 8486 5823 8642 5844
rect 8486 5805 8506 5823
rect 8524 5805 8642 5823
rect 8486 5801 8642 5805
rect 8486 5785 8547 5801
rect 4455 5746 4570 5761
rect 4549 5743 4570 5746
rect 4588 5743 4606 5761
rect 4549 5724 4606 5743
rect 4127 5616 4184 5635
rect 4127 5598 4145 5616
rect 4163 5613 4184 5616
rect 4163 5598 4278 5613
rect 186 5558 247 5574
rect 91 5554 247 5558
rect 91 5536 209 5554
rect 227 5536 247 5554
rect 91 5515 247 5536
rect 91 5514 191 5515
rect 92 5478 134 5514
rect 92 5455 243 5478
rect 4127 5575 4278 5598
rect 8491 5629 8548 5648
rect 8491 5611 8509 5629
rect 8527 5626 8548 5629
rect 8527 5611 8642 5626
rect 4236 5539 4278 5575
rect 4550 5571 4611 5587
rect 4455 5567 4611 5571
rect 4455 5549 4573 5567
rect 4591 5549 4611 5567
rect 4179 5538 4279 5539
rect 4123 5517 4279 5538
rect 4455 5528 4611 5549
rect 4455 5527 4555 5528
rect 92 5440 207 5455
rect 186 5437 207 5440
rect 225 5437 243 5455
rect 186 5418 243 5437
rect 4123 5499 4143 5517
rect 4161 5499 4279 5517
rect 4123 5495 4279 5499
rect 4123 5479 4184 5495
rect 4456 5491 4498 5527
rect 4456 5468 4607 5491
rect 8491 5588 8642 5611
rect 8600 5552 8642 5588
rect 8543 5551 8643 5552
rect 8487 5530 8643 5551
rect 4456 5453 4571 5468
rect 4550 5450 4571 5453
rect 4589 5450 4607 5468
rect 4550 5431 4607 5450
rect 4120 5398 4177 5417
rect 8487 5512 8507 5530
rect 8525 5512 8643 5530
rect 8487 5508 8643 5512
rect 8487 5492 8548 5508
rect 4120 5380 4138 5398
rect 4156 5395 4177 5398
rect 4156 5380 4271 5395
rect 4120 5357 4271 5380
rect 181 5234 242 5250
rect 4229 5321 4271 5357
rect 8484 5411 8541 5430
rect 8484 5393 8502 5411
rect 8520 5408 8541 5411
rect 8520 5393 8635 5408
rect 8484 5370 8635 5393
rect 4172 5320 4272 5321
rect 4116 5299 4272 5320
rect 4116 5281 4136 5299
rect 4154 5281 4272 5299
rect 4116 5277 4272 5281
rect 86 5230 242 5234
rect 86 5212 204 5230
rect 222 5212 242 5230
rect 86 5191 242 5212
rect 86 5190 186 5191
rect 87 5154 129 5190
rect 4116 5261 4177 5277
rect 4545 5247 4606 5263
rect 8593 5334 8635 5370
rect 8536 5333 8636 5334
rect 8480 5312 8636 5333
rect 8480 5294 8500 5312
rect 8518 5294 8636 5312
rect 8480 5290 8636 5294
rect 4450 5243 4606 5247
rect 4114 5215 4171 5234
rect 87 5131 238 5154
rect 87 5116 202 5131
rect 181 5113 202 5116
rect 220 5113 238 5131
rect 4114 5197 4132 5215
rect 4150 5212 4171 5215
rect 4450 5225 4568 5243
rect 4586 5225 4606 5243
rect 4150 5197 4265 5212
rect 4450 5204 4606 5225
rect 4450 5203 4550 5204
rect 4114 5174 4265 5197
rect 181 5094 238 5113
rect 175 5051 236 5067
rect 4223 5138 4265 5174
rect 4451 5167 4493 5203
rect 8480 5274 8541 5290
rect 8478 5228 8535 5247
rect 4451 5144 4602 5167
rect 4166 5137 4266 5138
rect 4110 5116 4266 5137
rect 4451 5129 4566 5144
rect 4110 5098 4130 5116
rect 4148 5098 4266 5116
rect 4545 5126 4566 5129
rect 4584 5126 4602 5144
rect 8478 5210 8496 5228
rect 8514 5225 8535 5228
rect 8514 5210 8629 5225
rect 8478 5187 8629 5210
rect 4545 5107 4602 5126
rect 4110 5094 4266 5098
rect 80 5047 236 5051
rect 80 5029 198 5047
rect 216 5029 236 5047
rect 80 5008 236 5029
rect 80 5007 180 5008
rect 81 4971 123 5007
rect 4110 5078 4171 5094
rect 4539 5064 4600 5080
rect 8587 5151 8629 5187
rect 8530 5150 8630 5151
rect 8474 5129 8630 5150
rect 8474 5111 8494 5129
rect 8512 5111 8630 5129
rect 8474 5107 8630 5111
rect 4444 5060 4600 5064
rect 4444 5042 4562 5060
rect 4580 5042 4600 5060
rect 4444 5021 4600 5042
rect 4444 5020 4544 5021
rect 81 4948 232 4971
rect 81 4933 196 4948
rect 175 4930 196 4933
rect 214 4930 232 4948
rect 175 4911 232 4930
rect 4445 4984 4487 5020
rect 8474 5091 8535 5107
rect 4445 4961 4596 4984
rect 168 4833 229 4849
rect 73 4829 229 4833
rect 73 4811 191 4829
rect 209 4811 229 4829
rect 4445 4946 4560 4961
rect 4539 4943 4560 4946
rect 4578 4943 4596 4961
rect 4539 4924 4596 4943
rect 4109 4891 4166 4910
rect 4109 4873 4127 4891
rect 4145 4888 4166 4891
rect 4145 4873 4260 4888
rect 73 4790 229 4811
rect 73 4789 173 4790
rect 74 4753 116 4789
rect 74 4730 225 4753
rect 4109 4850 4260 4873
rect 4218 4814 4260 4850
rect 4532 4846 4593 4862
rect 4437 4842 4593 4846
rect 4437 4824 4555 4842
rect 4573 4824 4593 4842
rect 8473 4904 8530 4923
rect 8473 4886 8491 4904
rect 8509 4901 8530 4904
rect 8509 4886 8624 4901
rect 4161 4813 4261 4814
rect 4105 4792 4261 4813
rect 4437 4803 4593 4824
rect 4437 4802 4537 4803
rect 4105 4774 4125 4792
rect 4143 4774 4261 4792
rect 4105 4770 4261 4774
rect 4105 4754 4166 4770
rect 4438 4766 4480 4802
rect 74 4715 189 4730
rect 168 4712 189 4715
rect 207 4712 225 4730
rect 168 4693 225 4712
rect 4438 4743 4589 4766
rect 8473 4863 8624 4886
rect 8582 4827 8624 4863
rect 8525 4826 8625 4827
rect 8469 4805 8625 4826
rect 8469 4787 8489 4805
rect 8507 4787 8625 4805
rect 8469 4783 8625 4787
rect 8469 4767 8530 4783
rect 4438 4728 4553 4743
rect 4532 4725 4553 4728
rect 4571 4725 4589 4743
rect 4532 4706 4589 4725
rect 4108 4598 4165 4617
rect 4108 4580 4126 4598
rect 4144 4595 4165 4598
rect 4144 4580 4259 4595
rect 167 4540 228 4556
rect 72 4536 228 4540
rect 72 4518 190 4536
rect 208 4518 228 4536
rect 72 4497 228 4518
rect 72 4496 172 4497
rect 73 4460 115 4496
rect 73 4437 224 4460
rect 4108 4557 4259 4580
rect 8472 4611 8529 4630
rect 8472 4593 8490 4611
rect 8508 4608 8529 4611
rect 8508 4593 8623 4608
rect 4217 4521 4259 4557
rect 4531 4553 4592 4569
rect 4436 4549 4592 4553
rect 4436 4531 4554 4549
rect 4572 4531 4592 4549
rect 4160 4520 4260 4521
rect 4104 4499 4260 4520
rect 4436 4510 4592 4531
rect 4436 4509 4536 4510
rect 73 4422 188 4437
rect 167 4419 188 4422
rect 206 4419 224 4437
rect 167 4400 224 4419
rect 4104 4481 4124 4499
rect 4142 4481 4260 4499
rect 4104 4477 4260 4481
rect 4104 4461 4165 4477
rect 4437 4473 4479 4509
rect 4437 4450 4588 4473
rect 8472 4570 8623 4593
rect 8581 4534 8623 4570
rect 8524 4533 8624 4534
rect 8468 4512 8624 4533
rect 4437 4435 4552 4450
rect 4531 4432 4552 4435
rect 4570 4432 4588 4450
rect 4531 4413 4588 4432
rect 4101 4380 4158 4399
rect 4101 4362 4119 4380
rect 4137 4377 4158 4380
rect 4137 4362 4252 4377
rect 8468 4494 8488 4512
rect 8506 4494 8624 4512
rect 8468 4490 8624 4494
rect 8468 4474 8529 4490
rect 4101 4339 4252 4362
rect 162 4216 223 4232
rect 4210 4303 4252 4339
rect 8465 4393 8522 4412
rect 8465 4375 8483 4393
rect 8501 4390 8522 4393
rect 8501 4375 8616 4390
rect 8465 4352 8616 4375
rect 4153 4302 4253 4303
rect 4097 4281 4253 4302
rect 4097 4263 4117 4281
rect 4135 4263 4253 4281
rect 4097 4259 4253 4263
rect 67 4212 223 4216
rect 67 4194 185 4212
rect 203 4194 223 4212
rect 67 4173 223 4194
rect 67 4172 167 4173
rect 68 4136 110 4172
rect 4097 4243 4158 4259
rect 4526 4229 4587 4245
rect 8574 4316 8616 4352
rect 8517 4315 8617 4316
rect 8461 4294 8617 4315
rect 8461 4276 8481 4294
rect 8499 4276 8617 4294
rect 8461 4272 8617 4276
rect 4431 4225 4587 4229
rect 4095 4197 4152 4216
rect 68 4113 219 4136
rect 68 4098 183 4113
rect 162 4095 183 4098
rect 201 4095 219 4113
rect 4095 4179 4113 4197
rect 4131 4194 4152 4197
rect 4431 4207 4549 4225
rect 4567 4207 4587 4225
rect 4131 4179 4246 4194
rect 4431 4186 4587 4207
rect 4431 4185 4531 4186
rect 4095 4156 4246 4179
rect 162 4076 219 4095
rect 156 4033 217 4049
rect 4204 4120 4246 4156
rect 4432 4149 4474 4185
rect 8461 4256 8522 4272
rect 8459 4210 8516 4229
rect 4432 4126 4583 4149
rect 4147 4119 4247 4120
rect 4091 4098 4247 4119
rect 4432 4111 4547 4126
rect 4091 4080 4111 4098
rect 4129 4080 4247 4098
rect 4526 4108 4547 4111
rect 4565 4108 4583 4126
rect 8459 4192 8477 4210
rect 8495 4207 8516 4210
rect 8495 4192 8610 4207
rect 8459 4169 8610 4192
rect 4526 4089 4583 4108
rect 4091 4076 4247 4080
rect 61 4029 217 4033
rect 61 4011 179 4029
rect 197 4011 217 4029
rect 61 3990 217 4011
rect 61 3989 161 3990
rect 62 3953 104 3989
rect 4091 4060 4152 4076
rect 4520 4046 4581 4062
rect 8568 4133 8610 4169
rect 8511 4132 8611 4133
rect 8455 4111 8611 4132
rect 8455 4093 8475 4111
rect 8493 4093 8611 4111
rect 8455 4089 8611 4093
rect 4425 4042 4581 4046
rect 4425 4024 4543 4042
rect 4561 4024 4581 4042
rect 4425 4003 4581 4024
rect 4425 4002 4525 4003
rect 62 3930 213 3953
rect 62 3915 177 3930
rect 156 3912 177 3915
rect 195 3912 213 3930
rect 156 3893 213 3912
rect 4426 3966 4468 4002
rect 8455 4073 8516 4089
rect 4426 3943 4577 3966
rect 4426 3928 4541 3943
rect 4520 3925 4541 3928
rect 4559 3925 4577 3943
rect 149 3815 210 3831
rect 54 3811 210 3815
rect 54 3793 172 3811
rect 190 3793 210 3811
rect 4520 3906 4577 3925
rect 4090 3873 4147 3892
rect 4090 3855 4108 3873
rect 4126 3870 4147 3873
rect 4126 3855 4241 3870
rect 54 3772 210 3793
rect 54 3771 154 3772
rect 55 3735 97 3771
rect 55 3712 206 3735
rect 4090 3832 4241 3855
rect 4199 3796 4241 3832
rect 4513 3828 4574 3844
rect 4418 3824 4574 3828
rect 4418 3806 4536 3824
rect 4554 3806 4574 3824
rect 8454 3886 8511 3905
rect 8454 3868 8472 3886
rect 8490 3883 8511 3886
rect 8490 3868 8605 3883
rect 4142 3795 4242 3796
rect 4086 3774 4242 3795
rect 4418 3785 4574 3806
rect 4418 3784 4518 3785
rect 4086 3756 4106 3774
rect 4124 3756 4242 3774
rect 4086 3752 4242 3756
rect 4086 3736 4147 3752
rect 4419 3748 4461 3784
rect 55 3697 170 3712
rect 149 3694 170 3697
rect 188 3694 206 3712
rect 149 3675 206 3694
rect 4419 3725 4570 3748
rect 8454 3845 8605 3868
rect 8563 3809 8605 3845
rect 8506 3808 8606 3809
rect 8450 3787 8606 3808
rect 8450 3769 8470 3787
rect 8488 3769 8606 3787
rect 8450 3765 8606 3769
rect 8450 3749 8511 3765
rect 4419 3710 4534 3725
rect 4513 3707 4534 3710
rect 4552 3707 4570 3725
rect 4513 3688 4570 3707
rect 4091 3580 4148 3599
rect 4091 3562 4109 3580
rect 4127 3577 4148 3580
rect 4127 3562 4242 3577
rect 150 3522 211 3538
rect 55 3518 211 3522
rect 55 3500 173 3518
rect 191 3500 211 3518
rect 55 3479 211 3500
rect 55 3478 155 3479
rect 56 3442 98 3478
rect 56 3419 207 3442
rect 4091 3539 4242 3562
rect 8455 3593 8512 3612
rect 8455 3575 8473 3593
rect 8491 3590 8512 3593
rect 8491 3575 8606 3590
rect 4200 3503 4242 3539
rect 4514 3535 4575 3551
rect 4419 3531 4575 3535
rect 4419 3513 4537 3531
rect 4555 3513 4575 3531
rect 4143 3502 4243 3503
rect 4087 3481 4243 3502
rect 4419 3492 4575 3513
rect 4419 3491 4519 3492
rect 56 3404 171 3419
rect 150 3401 171 3404
rect 189 3401 207 3419
rect 150 3382 207 3401
rect 4087 3463 4107 3481
rect 4125 3463 4243 3481
rect 4087 3459 4243 3463
rect 4087 3443 4148 3459
rect 4420 3455 4462 3491
rect 4420 3432 4571 3455
rect 8455 3552 8606 3575
rect 8564 3516 8606 3552
rect 8507 3515 8607 3516
rect 8451 3494 8607 3515
rect 4420 3417 4535 3432
rect 4514 3414 4535 3417
rect 4553 3414 4571 3432
rect 4514 3395 4571 3414
rect 4084 3362 4141 3381
rect 8451 3476 8471 3494
rect 8489 3476 8607 3494
rect 8451 3472 8607 3476
rect 8451 3456 8512 3472
rect 4084 3344 4102 3362
rect 4120 3359 4141 3362
rect 4120 3344 4235 3359
rect 4084 3321 4235 3344
rect 145 3198 206 3214
rect 4193 3285 4235 3321
rect 8448 3375 8505 3394
rect 8448 3357 8466 3375
rect 8484 3372 8505 3375
rect 8484 3357 8599 3372
rect 8448 3334 8599 3357
rect 4136 3284 4236 3285
rect 4080 3263 4236 3284
rect 4080 3245 4100 3263
rect 4118 3245 4236 3263
rect 4080 3241 4236 3245
rect 50 3194 206 3198
rect 50 3176 168 3194
rect 186 3176 206 3194
rect 50 3155 206 3176
rect 50 3154 150 3155
rect 51 3118 93 3154
rect 4080 3225 4141 3241
rect 4509 3211 4570 3227
rect 8557 3298 8599 3334
rect 8500 3297 8600 3298
rect 8444 3276 8600 3297
rect 8444 3258 8464 3276
rect 8482 3258 8600 3276
rect 8444 3254 8600 3258
rect 4414 3207 4570 3211
rect 4078 3179 4135 3198
rect 51 3095 202 3118
rect 51 3080 166 3095
rect 145 3077 166 3080
rect 184 3077 202 3095
rect 4078 3161 4096 3179
rect 4114 3176 4135 3179
rect 4414 3189 4532 3207
rect 4550 3189 4570 3207
rect 4114 3161 4229 3176
rect 4414 3168 4570 3189
rect 4414 3167 4514 3168
rect 4078 3138 4229 3161
rect 145 3058 202 3077
rect 139 3015 200 3031
rect 4187 3102 4229 3138
rect 4415 3131 4457 3167
rect 8444 3238 8505 3254
rect 8442 3192 8499 3211
rect 4415 3108 4566 3131
rect 4130 3101 4230 3102
rect 4074 3080 4230 3101
rect 4415 3093 4530 3108
rect 4074 3062 4094 3080
rect 4112 3062 4230 3080
rect 4509 3090 4530 3093
rect 4548 3090 4566 3108
rect 8442 3174 8460 3192
rect 8478 3189 8499 3192
rect 8478 3174 8593 3189
rect 8442 3151 8593 3174
rect 4509 3071 4566 3090
rect 4074 3058 4230 3062
rect 44 3011 200 3015
rect 44 2993 162 3011
rect 180 2993 200 3011
rect 44 2972 200 2993
rect 44 2971 144 2972
rect 45 2935 87 2971
rect 4074 3042 4135 3058
rect 4503 3028 4564 3044
rect 8551 3115 8593 3151
rect 8494 3114 8594 3115
rect 8438 3093 8594 3114
rect 8438 3075 8458 3093
rect 8476 3075 8594 3093
rect 8438 3071 8594 3075
rect 4408 3024 4564 3028
rect 4408 3006 4526 3024
rect 4544 3006 4564 3024
rect 4408 2985 4564 3006
rect 4408 2984 4508 2985
rect 45 2912 196 2935
rect 45 2897 160 2912
rect 139 2894 160 2897
rect 178 2894 196 2912
rect 139 2875 196 2894
rect 4409 2948 4451 2984
rect 8438 3055 8499 3071
rect 4409 2925 4560 2948
rect 4409 2910 4524 2925
rect 132 2797 193 2813
rect 37 2793 193 2797
rect 37 2775 155 2793
rect 173 2775 193 2793
rect 4503 2907 4524 2910
rect 4542 2907 4560 2925
rect 4503 2888 4560 2907
rect 4073 2855 4130 2874
rect 4073 2837 4091 2855
rect 4109 2852 4130 2855
rect 4109 2837 4224 2852
rect 37 2754 193 2775
rect 37 2753 137 2754
rect 38 2717 80 2753
rect 38 2694 189 2717
rect 4073 2814 4224 2837
rect 4182 2778 4224 2814
rect 4496 2810 4557 2826
rect 4401 2806 4557 2810
rect 4401 2788 4519 2806
rect 4537 2788 4557 2806
rect 8437 2868 8494 2887
rect 8437 2850 8455 2868
rect 8473 2865 8494 2868
rect 8473 2850 8588 2865
rect 4125 2777 4225 2778
rect 4069 2756 4225 2777
rect 4401 2767 4557 2788
rect 4401 2766 4501 2767
rect 4069 2738 4089 2756
rect 4107 2738 4225 2756
rect 4069 2734 4225 2738
rect 4069 2718 4130 2734
rect 4402 2730 4444 2766
rect 38 2679 153 2694
rect 132 2676 153 2679
rect 171 2676 189 2694
rect 132 2657 189 2676
rect 4402 2707 4553 2730
rect 8437 2827 8588 2850
rect 8546 2791 8588 2827
rect 8489 2790 8589 2791
rect 8433 2769 8589 2790
rect 8433 2751 8453 2769
rect 8471 2751 8589 2769
rect 8433 2747 8589 2751
rect 8433 2731 8494 2747
rect 4402 2692 4517 2707
rect 4496 2689 4517 2692
rect 4535 2689 4553 2707
rect 4496 2670 4553 2689
rect 4071 2562 4128 2581
rect 4071 2544 4089 2562
rect 4107 2559 4128 2562
rect 4107 2544 4222 2559
rect 130 2504 191 2520
rect 35 2500 191 2504
rect 35 2482 153 2500
rect 171 2482 191 2500
rect 35 2461 191 2482
rect 35 2460 135 2461
rect 36 2424 78 2460
rect 36 2401 187 2424
rect 4071 2521 4222 2544
rect 8435 2575 8492 2594
rect 8435 2557 8453 2575
rect 8471 2572 8492 2575
rect 8471 2557 8586 2572
rect 4180 2485 4222 2521
rect 4494 2517 4555 2533
rect 4399 2513 4555 2517
rect 4399 2495 4517 2513
rect 4535 2495 4555 2513
rect 4123 2484 4223 2485
rect 4067 2463 4223 2484
rect 4399 2474 4555 2495
rect 4399 2473 4499 2474
rect 36 2386 151 2401
rect 130 2383 151 2386
rect 169 2383 187 2401
rect 130 2364 187 2383
rect 4067 2445 4087 2463
rect 4105 2445 4223 2463
rect 4067 2441 4223 2445
rect 4067 2425 4128 2441
rect 4400 2437 4442 2473
rect 4400 2414 4551 2437
rect 8435 2534 8586 2557
rect 8544 2498 8586 2534
rect 8487 2497 8587 2498
rect 8431 2476 8587 2497
rect 4400 2399 4515 2414
rect 4494 2396 4515 2399
rect 4533 2396 4551 2414
rect 4494 2377 4551 2396
rect 4064 2344 4121 2363
rect 4064 2326 4082 2344
rect 4100 2341 4121 2344
rect 8431 2458 8451 2476
rect 8469 2458 8587 2476
rect 8431 2454 8587 2458
rect 8431 2438 8492 2454
rect 4100 2326 4215 2341
rect 4064 2303 4215 2326
rect 125 2180 186 2196
rect 4173 2267 4215 2303
rect 8428 2357 8485 2376
rect 8428 2339 8446 2357
rect 8464 2354 8485 2357
rect 8464 2339 8579 2354
rect 8428 2316 8579 2339
rect 4116 2266 4216 2267
rect 4060 2245 4216 2266
rect 4060 2227 4080 2245
rect 4098 2227 4216 2245
rect 4060 2223 4216 2227
rect 30 2176 186 2180
rect 30 2158 148 2176
rect 166 2158 186 2176
rect 30 2137 186 2158
rect 30 2136 130 2137
rect 31 2100 73 2136
rect 4060 2207 4121 2223
rect 4489 2193 4550 2209
rect 8537 2280 8579 2316
rect 8480 2279 8580 2280
rect 8424 2258 8580 2279
rect 8424 2240 8444 2258
rect 8462 2240 8580 2258
rect 8424 2236 8580 2240
rect 4394 2189 4550 2193
rect 4058 2161 4115 2180
rect 31 2077 182 2100
rect 31 2062 146 2077
rect 125 2059 146 2062
rect 164 2059 182 2077
rect 4058 2143 4076 2161
rect 4094 2158 4115 2161
rect 4394 2171 4512 2189
rect 4530 2171 4550 2189
rect 4094 2143 4209 2158
rect 4394 2150 4550 2171
rect 4394 2149 4494 2150
rect 4058 2120 4209 2143
rect 125 2040 182 2059
rect 119 1997 180 2013
rect 4167 2084 4209 2120
rect 4395 2113 4437 2149
rect 8424 2220 8485 2236
rect 8422 2174 8479 2193
rect 4395 2090 4546 2113
rect 4110 2083 4210 2084
rect 4054 2062 4210 2083
rect 4395 2075 4510 2090
rect 4054 2044 4074 2062
rect 4092 2044 4210 2062
rect 4489 2072 4510 2075
rect 4528 2072 4546 2090
rect 8422 2156 8440 2174
rect 8458 2171 8479 2174
rect 8458 2156 8573 2171
rect 8422 2133 8573 2156
rect 4489 2053 4546 2072
rect 4054 2040 4210 2044
rect 24 1993 180 1997
rect 24 1975 142 1993
rect 160 1975 180 1993
rect 24 1954 180 1975
rect 24 1953 124 1954
rect 25 1917 67 1953
rect 4054 2024 4115 2040
rect 4483 2010 4544 2026
rect 8531 2097 8573 2133
rect 8474 2096 8574 2097
rect 8418 2075 8574 2096
rect 8418 2057 8438 2075
rect 8456 2057 8574 2075
rect 8418 2053 8574 2057
rect 4388 2006 4544 2010
rect 4388 1988 4506 2006
rect 4524 1988 4544 2006
rect 4388 1967 4544 1988
rect 4388 1966 4488 1967
rect 25 1894 176 1917
rect 25 1879 140 1894
rect 119 1876 140 1879
rect 158 1876 176 1894
rect 119 1857 176 1876
rect 4389 1930 4431 1966
rect 8418 2037 8479 2053
rect 4389 1907 4540 1930
rect 4389 1892 4504 1907
rect 4483 1889 4504 1892
rect 4522 1889 4540 1907
rect 112 1779 173 1795
rect 17 1775 173 1779
rect 17 1757 135 1775
rect 153 1757 173 1775
rect 4483 1870 4540 1889
rect 4053 1837 4110 1856
rect 4053 1819 4071 1837
rect 4089 1834 4110 1837
rect 4089 1819 4204 1834
rect 17 1736 173 1757
rect 17 1735 117 1736
rect 18 1699 60 1735
rect 18 1676 169 1699
rect 4053 1796 4204 1819
rect 4162 1760 4204 1796
rect 4476 1792 4537 1808
rect 4381 1788 4537 1792
rect 4381 1770 4499 1788
rect 4517 1770 4537 1788
rect 8417 1850 8474 1869
rect 8417 1832 8435 1850
rect 8453 1847 8474 1850
rect 8453 1832 8568 1847
rect 4105 1759 4205 1760
rect 4049 1738 4205 1759
rect 4381 1749 4537 1770
rect 4381 1748 4481 1749
rect 4049 1720 4069 1738
rect 4087 1720 4205 1738
rect 4049 1716 4205 1720
rect 4049 1700 4110 1716
rect 4382 1712 4424 1748
rect 18 1661 133 1676
rect 112 1658 133 1661
rect 151 1658 169 1676
rect 112 1639 169 1658
rect 4382 1689 4533 1712
rect 8417 1809 8568 1832
rect 8526 1773 8568 1809
rect 8469 1772 8569 1773
rect 8413 1751 8569 1772
rect 8413 1733 8433 1751
rect 8451 1733 8569 1751
rect 8413 1729 8569 1733
rect 8413 1713 8474 1729
rect 4382 1674 4497 1689
rect 4476 1671 4497 1674
rect 4515 1671 4533 1689
rect 4476 1652 4533 1671
rect 4054 1544 4111 1563
rect 4054 1526 4072 1544
rect 4090 1541 4111 1544
rect 4090 1526 4205 1541
rect 113 1486 174 1502
rect 18 1482 174 1486
rect 18 1464 136 1482
rect 154 1464 174 1482
rect 18 1443 174 1464
rect 18 1442 118 1443
rect 19 1406 61 1442
rect 19 1383 170 1406
rect 4054 1503 4205 1526
rect 8418 1557 8475 1576
rect 8418 1539 8436 1557
rect 8454 1554 8475 1557
rect 8454 1539 8569 1554
rect 4163 1467 4205 1503
rect 4477 1499 4538 1515
rect 4382 1495 4538 1499
rect 4382 1477 4500 1495
rect 4518 1477 4538 1495
rect 4106 1466 4206 1467
rect 4050 1445 4206 1466
rect 4382 1456 4538 1477
rect 4382 1455 4482 1456
rect 19 1368 134 1383
rect 113 1365 134 1368
rect 152 1365 170 1383
rect 113 1346 170 1365
rect 4050 1427 4070 1445
rect 4088 1427 4206 1445
rect 4050 1423 4206 1427
rect 4050 1407 4111 1423
rect 4383 1419 4425 1455
rect 4383 1396 4534 1419
rect 8418 1516 8569 1539
rect 8527 1480 8569 1516
rect 8470 1479 8570 1480
rect 8414 1458 8570 1479
rect 4383 1381 4498 1396
rect 4477 1378 4498 1381
rect 4516 1378 4534 1396
rect 4477 1359 4534 1378
rect 4047 1326 4104 1345
rect 8414 1440 8434 1458
rect 8452 1440 8570 1458
rect 8414 1436 8570 1440
rect 8414 1420 8475 1436
rect 4047 1308 4065 1326
rect 4083 1323 4104 1326
rect 4083 1308 4198 1323
rect 4047 1285 4198 1308
rect 108 1162 169 1178
rect 4156 1249 4198 1285
rect 8411 1339 8468 1358
rect 8411 1321 8429 1339
rect 8447 1336 8468 1339
rect 8447 1321 8562 1336
rect 8411 1298 8562 1321
rect 4099 1248 4199 1249
rect 4043 1227 4199 1248
rect 4043 1209 4063 1227
rect 4081 1209 4199 1227
rect 4043 1205 4199 1209
rect 13 1158 169 1162
rect 13 1140 131 1158
rect 149 1140 169 1158
rect 13 1119 169 1140
rect 13 1118 113 1119
rect 14 1082 56 1118
rect 4043 1189 4104 1205
rect 4472 1175 4533 1191
rect 8520 1262 8562 1298
rect 8463 1261 8563 1262
rect 8407 1240 8563 1261
rect 8407 1222 8427 1240
rect 8445 1222 8563 1240
rect 8407 1218 8563 1222
rect 4377 1171 4533 1175
rect 4041 1143 4098 1162
rect 14 1059 165 1082
rect 14 1044 129 1059
rect 108 1041 129 1044
rect 147 1041 165 1059
rect 4041 1125 4059 1143
rect 4077 1140 4098 1143
rect 4377 1153 4495 1171
rect 4513 1153 4533 1171
rect 4077 1125 4192 1140
rect 4377 1132 4533 1153
rect 4377 1131 4477 1132
rect 4041 1102 4192 1125
rect 108 1022 165 1041
rect 102 979 163 995
rect 4150 1066 4192 1102
rect 4378 1095 4420 1131
rect 8407 1202 8468 1218
rect 8405 1156 8462 1175
rect 4378 1072 4529 1095
rect 4093 1065 4193 1066
rect 4037 1044 4193 1065
rect 4378 1057 4493 1072
rect 4037 1026 4057 1044
rect 4075 1026 4193 1044
rect 4472 1054 4493 1057
rect 4511 1054 4529 1072
rect 8405 1138 8423 1156
rect 8441 1153 8462 1156
rect 8441 1138 8556 1153
rect 8405 1115 8556 1138
rect 4472 1035 4529 1054
rect 4037 1022 4193 1026
rect 7 975 163 979
rect 7 957 125 975
rect 143 957 163 975
rect 7 936 163 957
rect 7 935 107 936
rect 8 899 50 935
rect 4037 1006 4098 1022
rect 4466 992 4527 1008
rect 8514 1079 8556 1115
rect 8457 1078 8557 1079
rect 8401 1057 8557 1078
rect 8401 1039 8421 1057
rect 8439 1039 8557 1057
rect 8401 1035 8557 1039
rect 4371 988 4527 992
rect 4371 970 4489 988
rect 4507 970 4527 988
rect 4371 949 4527 970
rect 4371 948 4471 949
rect 4372 912 4414 948
rect 8401 1019 8462 1035
rect 8 876 159 899
rect 8 861 123 876
rect 102 858 123 861
rect 141 858 159 876
rect 102 839 159 858
rect 4372 889 4523 912
rect 4372 874 4487 889
rect 4466 871 4487 874
rect 4505 871 4523 889
rect 95 761 156 777
rect 0 757 156 761
rect 0 739 118 757
rect 136 739 156 757
rect 4466 852 4523 871
rect 4036 819 4093 838
rect 4036 801 4054 819
rect 4072 816 4093 819
rect 4072 801 4187 816
rect 4036 778 4187 801
rect 0 718 156 739
rect 0 717 100 718
rect 1 681 43 717
rect 1 658 152 681
rect 4145 742 4187 778
rect 4459 774 4520 790
rect 4364 770 4520 774
rect 4364 752 4482 770
rect 4500 752 4520 770
rect 8400 832 8457 851
rect 8400 814 8418 832
rect 8436 829 8457 832
rect 8436 814 8551 829
rect 8400 791 8551 814
rect 4088 741 4188 742
rect 4032 720 4188 741
rect 4364 731 4520 752
rect 4364 730 4464 731
rect 4032 702 4052 720
rect 4070 702 4188 720
rect 4032 698 4188 702
rect 4032 682 4093 698
rect 4365 694 4407 730
rect 1 643 116 658
rect 95 640 116 643
rect 134 640 152 658
rect 95 621 152 640
rect 4365 671 4516 694
rect 8509 755 8551 791
rect 8452 754 8552 755
rect 8396 733 8552 754
rect 8396 715 8416 733
rect 8434 715 8552 733
rect 8396 711 8552 715
rect 8396 695 8457 711
rect 4365 656 4480 671
rect 4459 653 4480 656
rect 4498 653 4516 671
rect 4459 634 4516 653
<< locali >>
rect 2875 8749 2915 8757
rect 2875 8727 2883 8749
rect 2907 8727 2915 8749
rect 3779 8752 4235 8787
rect 7239 8762 7279 8770
rect 253 8608 300 8724
rect 253 8590 263 8608
rect 281 8590 300 8608
rect 253 8586 300 8590
rect 254 8581 291 8586
rect 242 8519 294 8521
rect 240 8515 673 8519
rect 240 8509 679 8515
rect 240 8491 261 8509
rect 279 8491 679 8509
rect 240 8473 679 8491
rect 242 8284 294 8473
rect 640 8448 679 8473
rect 2480 8498 2517 8504
rect 2480 8479 2488 8498
rect 2509 8479 2517 8498
rect 2480 8471 2517 8479
rect 424 8423 611 8447
rect 640 8428 1035 8448
rect 1055 8428 1058 8448
rect 640 8423 1058 8428
rect 424 8352 461 8423
rect 640 8422 983 8423
rect 640 8419 679 8422
rect 945 8421 982 8422
rect 576 8362 607 8363
rect 424 8332 433 8352
rect 453 8332 461 8352
rect 424 8322 461 8332
rect 520 8352 607 8362
rect 520 8332 529 8352
rect 549 8332 607 8352
rect 520 8323 607 8332
rect 520 8322 557 8323
rect 242 8266 258 8284
rect 276 8266 294 8284
rect 576 8272 607 8323
rect 642 8352 679 8419
rect 794 8362 830 8363
rect 642 8332 651 8352
rect 671 8332 679 8352
rect 642 8322 679 8332
rect 738 8352 886 8362
rect 986 8359 1082 8361
rect 738 8332 747 8352
rect 767 8332 857 8352
rect 877 8332 886 8352
rect 738 8323 886 8332
rect 944 8352 1082 8359
rect 944 8332 953 8352
rect 973 8332 1082 8352
rect 944 8323 1082 8332
rect 738 8322 775 8323
rect 468 8269 509 8270
rect 242 8248 294 8266
rect 360 8262 509 8269
rect 360 8242 419 8262
rect 439 8242 478 8262
rect 498 8242 509 8262
rect 360 8234 509 8242
rect 576 8265 733 8272
rect 576 8245 696 8265
rect 716 8245 733 8265
rect 576 8235 733 8245
rect 576 8234 611 8235
rect 576 8213 607 8234
rect 794 8213 830 8323
rect 849 8322 886 8323
rect 945 8322 982 8323
rect 905 8263 995 8269
rect 905 8243 914 8263
rect 934 8261 995 8263
rect 934 8243 959 8261
rect 905 8241 959 8243
rect 979 8241 995 8261
rect 905 8235 995 8241
rect 419 8212 456 8213
rect 418 8203 456 8212
rect 246 8185 286 8195
rect 246 8167 256 8185
rect 274 8167 286 8185
rect 418 8183 427 8203
rect 447 8183 456 8203
rect 418 8175 456 8183
rect 522 8207 607 8213
rect 637 8212 674 8213
rect 522 8187 530 8207
rect 550 8187 607 8207
rect 522 8179 607 8187
rect 636 8203 674 8212
rect 636 8183 645 8203
rect 665 8183 674 8203
rect 522 8178 558 8179
rect 636 8175 674 8183
rect 740 8207 884 8213
rect 740 8187 748 8207
rect 768 8187 801 8207
rect 821 8187 856 8207
rect 876 8187 884 8207
rect 740 8179 884 8187
rect 740 8178 776 8179
rect 848 8178 884 8179
rect 950 8212 987 8213
rect 950 8211 988 8212
rect 950 8203 1014 8211
rect 950 8183 959 8203
rect 979 8189 1014 8203
rect 1034 8189 1037 8209
rect 979 8184 1037 8189
rect 979 8183 1014 8184
rect 246 8111 286 8167
rect 419 8146 456 8175
rect 420 8144 456 8146
rect 420 8122 611 8144
rect 637 8143 674 8175
rect 950 8171 1014 8183
rect 1054 8145 1081 8323
rect 913 8143 1081 8145
rect 637 8133 1081 8143
rect 1222 8239 1409 8263
rect 1440 8244 1833 8264
rect 1853 8244 1856 8264
rect 1440 8239 1856 8244
rect 1222 8168 1259 8239
rect 1440 8238 1781 8239
rect 1374 8178 1405 8179
rect 1222 8148 1231 8168
rect 1251 8148 1259 8168
rect 1222 8138 1259 8148
rect 1318 8168 1405 8178
rect 1318 8148 1327 8168
rect 1347 8148 1405 8168
rect 1318 8139 1405 8148
rect 1318 8138 1355 8139
rect 243 8106 286 8111
rect 634 8117 1081 8133
rect 634 8111 662 8117
rect 913 8116 1081 8117
rect 243 8103 393 8106
rect 634 8103 661 8111
rect 243 8101 661 8103
rect 243 8083 252 8101
rect 270 8083 661 8101
rect 1374 8088 1405 8139
rect 1440 8168 1477 8238
rect 1743 8237 1780 8238
rect 1592 8178 1628 8179
rect 1440 8148 1449 8168
rect 1469 8148 1477 8168
rect 1440 8138 1477 8148
rect 1536 8168 1684 8178
rect 1784 8175 1880 8177
rect 1536 8148 1545 8168
rect 1565 8148 1655 8168
rect 1675 8148 1684 8168
rect 1536 8139 1684 8148
rect 1742 8168 1880 8175
rect 1742 8148 1751 8168
rect 1771 8148 1880 8168
rect 1742 8139 1880 8148
rect 1536 8138 1573 8139
rect 1266 8085 1307 8086
rect 243 8080 661 8083
rect 243 8074 286 8080
rect 246 8071 286 8074
rect 1158 8078 1307 8085
rect 643 8062 683 8063
rect 354 8045 683 8062
rect 1158 8058 1217 8078
rect 1237 8058 1276 8078
rect 1296 8058 1307 8078
rect 1158 8050 1307 8058
rect 1374 8081 1531 8088
rect 1374 8061 1494 8081
rect 1514 8061 1531 8081
rect 1374 8051 1531 8061
rect 1374 8050 1409 8051
rect 238 8002 281 8013
rect 238 7984 250 8002
rect 268 7984 281 8002
rect 238 7958 281 7984
rect 354 7958 381 8045
rect 643 8036 683 8045
rect 238 7937 381 7958
rect 425 8010 459 8026
rect 643 8016 1036 8036
rect 1056 8016 1059 8036
rect 1374 8029 1405 8050
rect 1592 8029 1628 8139
rect 1647 8138 1684 8139
rect 1743 8138 1780 8139
rect 1703 8079 1793 8085
rect 1703 8059 1712 8079
rect 1732 8077 1793 8079
rect 1732 8059 1757 8077
rect 1703 8057 1757 8059
rect 1777 8057 1793 8077
rect 1703 8051 1793 8057
rect 1217 8028 1254 8029
rect 643 8011 1059 8016
rect 1216 8019 1254 8028
rect 643 8010 984 8011
rect 425 7940 462 8010
rect 577 7950 608 7951
rect 238 7935 375 7937
rect 238 7893 281 7935
rect 425 7920 434 7940
rect 454 7920 462 7940
rect 425 7910 462 7920
rect 521 7940 608 7950
rect 521 7920 530 7940
rect 550 7920 608 7940
rect 521 7911 608 7920
rect 521 7910 558 7911
rect 236 7883 281 7893
rect 236 7865 245 7883
rect 263 7865 281 7883
rect 236 7859 281 7865
rect 577 7860 608 7911
rect 643 7940 680 8010
rect 946 8009 983 8010
rect 1216 7999 1225 8019
rect 1245 7999 1254 8019
rect 1216 7991 1254 7999
rect 1320 8023 1405 8029
rect 1435 8028 1472 8029
rect 1320 8003 1328 8023
rect 1348 8003 1405 8023
rect 1320 7995 1405 8003
rect 1434 8019 1472 8028
rect 1434 7999 1443 8019
rect 1463 7999 1472 8019
rect 1320 7994 1356 7995
rect 1434 7991 1472 7999
rect 1538 8023 1682 8029
rect 1538 8003 1546 8023
rect 1566 8004 1598 8023
rect 1619 8004 1654 8023
rect 1566 8003 1654 8004
rect 1674 8003 1682 8023
rect 1538 7995 1682 8003
rect 1538 7994 1574 7995
rect 1646 7994 1682 7995
rect 1748 8028 1785 8029
rect 1748 8027 1786 8028
rect 1748 8019 1812 8027
rect 1748 7999 1757 8019
rect 1777 8005 1812 8019
rect 1832 8005 1835 8025
rect 1777 8000 1835 8005
rect 1777 7999 1812 8000
rect 1217 7962 1254 7991
rect 1218 7960 1254 7962
rect 795 7950 831 7951
rect 643 7920 652 7940
rect 672 7920 680 7940
rect 643 7910 680 7920
rect 739 7940 887 7950
rect 987 7947 1083 7949
rect 739 7920 748 7940
rect 768 7920 858 7940
rect 878 7920 887 7940
rect 739 7911 887 7920
rect 945 7940 1083 7947
rect 945 7920 954 7940
rect 974 7920 1083 7940
rect 1218 7938 1409 7960
rect 1435 7959 1472 7991
rect 1748 7987 1812 7999
rect 1852 7961 1879 8139
rect 2484 8138 2517 8471
rect 2581 8503 2749 8504
rect 2875 8503 2915 8727
rect 3378 8731 3546 8732
rect 3779 8731 3824 8752
rect 3378 8705 3824 8731
rect 3378 8703 3546 8705
rect 3742 8704 3824 8705
rect 3959 8704 4040 8730
rect 4184 8717 4665 8752
rect 7239 8740 7247 8762
rect 7271 8740 7279 8762
rect 3378 8525 3405 8703
rect 3445 8665 3509 8677
rect 3785 8673 3822 8704
rect 4003 8673 4040 8704
rect 4187 8698 4226 8717
rect 4185 8679 4226 8698
rect 3445 8664 3480 8665
rect 3422 8659 3480 8664
rect 3422 8639 3425 8659
rect 3445 8645 3480 8659
rect 3500 8645 3509 8665
rect 3445 8637 3509 8645
rect 3471 8636 3509 8637
rect 3472 8635 3509 8636
rect 3575 8669 3611 8670
rect 3683 8669 3719 8670
rect 3575 8661 3719 8669
rect 3575 8641 3583 8661
rect 3603 8657 3691 8661
rect 3603 8641 3647 8657
rect 3575 8637 3647 8641
rect 3667 8641 3691 8657
rect 3711 8641 3719 8661
rect 3667 8637 3719 8641
rect 3575 8635 3719 8637
rect 3785 8665 3823 8673
rect 3901 8669 3937 8670
rect 3785 8645 3794 8665
rect 3814 8645 3823 8665
rect 3785 8636 3823 8645
rect 3852 8661 3937 8669
rect 3852 8641 3909 8661
rect 3929 8641 3937 8661
rect 3785 8635 3822 8636
rect 3852 8635 3937 8641
rect 4003 8665 4041 8673
rect 4003 8645 4012 8665
rect 4032 8645 4041 8665
rect 4003 8636 4041 8645
rect 4185 8670 4227 8679
rect 4185 8652 4199 8670
rect 4217 8652 4227 8670
rect 4185 8644 4227 8652
rect 4190 8642 4227 8644
rect 4003 8635 4040 8636
rect 3464 8607 3554 8613
rect 3464 8587 3480 8607
rect 3500 8605 3554 8607
rect 3500 8587 3525 8605
rect 3464 8585 3525 8587
rect 3545 8585 3554 8605
rect 3464 8579 3554 8585
rect 3477 8525 3514 8526
rect 3573 8525 3610 8526
rect 3629 8525 3665 8635
rect 3852 8614 3883 8635
rect 4617 8621 4664 8717
rect 3848 8613 3883 8614
rect 3726 8603 3883 8613
rect 3726 8583 3743 8603
rect 3763 8583 3883 8603
rect 3726 8576 3883 8583
rect 3950 8606 4099 8614
rect 3950 8586 3961 8606
rect 3981 8586 4020 8606
rect 4040 8586 4099 8606
rect 4617 8603 4627 8621
rect 4645 8603 4664 8621
rect 4617 8599 4664 8603
rect 4618 8594 4655 8599
rect 3950 8579 4099 8586
rect 3950 8578 3991 8579
rect 4187 8577 4224 8580
rect 3684 8525 3721 8526
rect 3377 8516 3515 8525
rect 2581 8477 3025 8503
rect 2581 8475 2749 8477
rect 2581 8297 2608 8475
rect 2648 8437 2712 8449
rect 2988 8445 3025 8477
rect 3051 8476 3242 8498
rect 3377 8496 3486 8516
rect 3506 8496 3515 8516
rect 3377 8489 3515 8496
rect 3573 8516 3721 8525
rect 3573 8496 3582 8516
rect 3602 8496 3692 8516
rect 3712 8496 3721 8516
rect 3377 8487 3473 8489
rect 3573 8486 3721 8496
rect 3780 8516 3817 8526
rect 3780 8496 3788 8516
rect 3808 8496 3817 8516
rect 3629 8485 3665 8486
rect 3206 8474 3242 8476
rect 3206 8445 3243 8474
rect 2648 8436 2683 8437
rect 2625 8431 2683 8436
rect 2625 8411 2628 8431
rect 2648 8417 2683 8431
rect 2703 8417 2712 8437
rect 2648 8411 2712 8417
rect 2625 8409 2712 8411
rect 2625 8405 2652 8409
rect 2674 8408 2712 8409
rect 2675 8407 2712 8408
rect 2778 8441 2814 8442
rect 2886 8441 2922 8442
rect 2778 8434 2922 8441
rect 2778 8433 2840 8434
rect 2778 8413 2786 8433
rect 2806 8416 2840 8433
rect 2859 8433 2922 8434
rect 2859 8416 2894 8433
rect 2806 8413 2894 8416
rect 2914 8413 2922 8433
rect 2778 8407 2922 8413
rect 2988 8437 3026 8445
rect 3104 8441 3140 8442
rect 2988 8417 2997 8437
rect 3017 8417 3026 8437
rect 2988 8408 3026 8417
rect 3055 8433 3140 8441
rect 3055 8413 3112 8433
rect 3132 8413 3140 8433
rect 2988 8407 3025 8408
rect 3055 8407 3140 8413
rect 3206 8437 3244 8445
rect 3206 8417 3215 8437
rect 3235 8417 3244 8437
rect 3477 8426 3514 8427
rect 3780 8426 3817 8496
rect 3852 8525 3883 8576
rect 4179 8571 4224 8577
rect 4179 8553 4197 8571
rect 4215 8553 4224 8571
rect 4179 8543 4224 8553
rect 3902 8525 3939 8526
rect 3852 8516 3939 8525
rect 3852 8496 3910 8516
rect 3930 8496 3939 8516
rect 3852 8486 3939 8496
rect 3998 8516 4035 8526
rect 3998 8496 4006 8516
rect 4026 8496 4035 8516
rect 4179 8501 4222 8543
rect 4606 8532 4658 8534
rect 4085 8499 4222 8501
rect 3852 8485 3883 8486
rect 3998 8426 4035 8496
rect 3476 8425 3817 8426
rect 3206 8408 3244 8417
rect 3401 8420 3817 8425
rect 3206 8407 3243 8408
rect 2667 8379 2757 8385
rect 2667 8359 2683 8379
rect 2703 8377 2757 8379
rect 2703 8359 2728 8377
rect 2667 8357 2728 8359
rect 2748 8357 2757 8377
rect 2667 8351 2757 8357
rect 2680 8297 2717 8298
rect 2776 8297 2813 8298
rect 2832 8297 2868 8407
rect 3055 8386 3086 8407
rect 3401 8400 3404 8420
rect 3424 8400 3817 8420
rect 4001 8410 4035 8426
rect 4079 8478 4222 8499
rect 4604 8528 5037 8532
rect 4604 8522 5043 8528
rect 4604 8504 4625 8522
rect 4643 8504 5043 8522
rect 4604 8486 5043 8504
rect 3777 8391 3817 8400
rect 4079 8391 4106 8478
rect 4179 8452 4222 8478
rect 4179 8434 4192 8452
rect 4210 8434 4222 8452
rect 4179 8423 4222 8434
rect 3051 8385 3086 8386
rect 2929 8375 3086 8385
rect 2929 8355 2946 8375
rect 2966 8355 3086 8375
rect 2929 8348 3086 8355
rect 3153 8378 3299 8386
rect 3153 8358 3164 8378
rect 3184 8358 3223 8378
rect 3243 8358 3299 8378
rect 3777 8374 4106 8391
rect 3777 8373 3817 8374
rect 3153 8351 3299 8358
rect 4174 8362 4214 8365
rect 4174 8356 4217 8362
rect 3799 8353 4217 8356
rect 3153 8350 3194 8351
rect 2887 8297 2924 8298
rect 2580 8288 2718 8297
rect 2580 8268 2689 8288
rect 2709 8268 2718 8288
rect 2580 8261 2718 8268
rect 2776 8288 2924 8297
rect 2776 8268 2785 8288
rect 2805 8268 2895 8288
rect 2915 8268 2924 8288
rect 2580 8259 2676 8261
rect 2776 8258 2924 8268
rect 2983 8288 3020 8298
rect 2983 8268 2991 8288
rect 3011 8268 3020 8288
rect 2832 8257 2868 8258
rect 2680 8198 2717 8199
rect 2983 8198 3020 8268
rect 3055 8297 3086 8348
rect 3799 8335 4190 8353
rect 4208 8335 4217 8353
rect 3799 8333 4217 8335
rect 3799 8325 3826 8333
rect 4067 8330 4217 8333
rect 3379 8319 3547 8320
rect 3798 8319 3826 8325
rect 3379 8303 3826 8319
rect 4174 8325 4217 8330
rect 3105 8297 3142 8298
rect 3055 8288 3142 8297
rect 3055 8268 3113 8288
rect 3133 8268 3142 8288
rect 3055 8258 3142 8268
rect 3201 8288 3238 8298
rect 3201 8268 3209 8288
rect 3229 8268 3238 8288
rect 3055 8257 3086 8258
rect 2679 8197 3020 8198
rect 3201 8197 3238 8268
rect 2604 8192 3020 8197
rect 2604 8172 2607 8192
rect 2627 8172 3020 8192
rect 3051 8173 3238 8197
rect 3379 8293 3823 8303
rect 3379 8291 3547 8293
rect 2479 8093 2521 8138
rect 3379 8113 3406 8291
rect 3446 8253 3510 8265
rect 3786 8261 3823 8293
rect 3849 8292 4040 8314
rect 4004 8290 4040 8292
rect 4004 8261 4041 8290
rect 4174 8269 4214 8325
rect 3446 8252 3481 8253
rect 3423 8247 3481 8252
rect 3423 8227 3426 8247
rect 3446 8233 3481 8247
rect 3501 8233 3510 8253
rect 3446 8225 3510 8233
rect 3472 8224 3510 8225
rect 3473 8223 3510 8224
rect 3576 8257 3612 8258
rect 3684 8257 3720 8258
rect 3576 8249 3720 8257
rect 3576 8229 3584 8249
rect 3604 8229 3639 8249
rect 3659 8229 3692 8249
rect 3712 8229 3720 8249
rect 3576 8223 3720 8229
rect 3786 8253 3824 8261
rect 3902 8257 3938 8258
rect 3786 8233 3795 8253
rect 3815 8233 3824 8253
rect 3786 8224 3824 8233
rect 3853 8249 3938 8257
rect 3853 8229 3910 8249
rect 3930 8229 3938 8249
rect 3786 8223 3823 8224
rect 3853 8223 3938 8229
rect 4004 8253 4042 8261
rect 4004 8233 4013 8253
rect 4033 8233 4042 8253
rect 4174 8251 4186 8269
rect 4204 8251 4214 8269
rect 4606 8297 4658 8486
rect 5004 8461 5043 8486
rect 6844 8511 6881 8517
rect 6844 8492 6852 8511
rect 6873 8492 6881 8511
rect 6844 8484 6881 8492
rect 4788 8436 4975 8460
rect 5004 8441 5399 8461
rect 5419 8441 5422 8461
rect 5004 8436 5422 8441
rect 4788 8365 4825 8436
rect 5004 8435 5347 8436
rect 5004 8432 5043 8435
rect 5309 8434 5346 8435
rect 4940 8375 4971 8376
rect 4788 8345 4797 8365
rect 4817 8345 4825 8365
rect 4788 8335 4825 8345
rect 4884 8365 4971 8375
rect 4884 8345 4893 8365
rect 4913 8345 4971 8365
rect 4884 8336 4971 8345
rect 4884 8335 4921 8336
rect 4606 8279 4622 8297
rect 4640 8279 4658 8297
rect 4940 8285 4971 8336
rect 5006 8365 5043 8432
rect 5158 8375 5194 8376
rect 5006 8345 5015 8365
rect 5035 8345 5043 8365
rect 5006 8335 5043 8345
rect 5102 8365 5250 8375
rect 5350 8372 5446 8374
rect 5102 8345 5111 8365
rect 5131 8345 5221 8365
rect 5241 8345 5250 8365
rect 5102 8336 5250 8345
rect 5308 8365 5446 8372
rect 5308 8345 5317 8365
rect 5337 8345 5446 8365
rect 5308 8336 5446 8345
rect 5102 8335 5139 8336
rect 4832 8282 4873 8283
rect 4606 8261 4658 8279
rect 4724 8275 4873 8282
rect 4174 8241 4214 8251
rect 4724 8255 4783 8275
rect 4803 8255 4842 8275
rect 4862 8255 4873 8275
rect 4724 8247 4873 8255
rect 4940 8278 5097 8285
rect 4940 8258 5060 8278
rect 5080 8258 5097 8278
rect 4940 8248 5097 8258
rect 4940 8247 4975 8248
rect 4004 8224 4042 8233
rect 4940 8226 4971 8247
rect 5158 8226 5194 8336
rect 5213 8335 5250 8336
rect 5309 8335 5346 8336
rect 5269 8276 5359 8282
rect 5269 8256 5278 8276
rect 5298 8274 5359 8276
rect 5298 8256 5323 8274
rect 5269 8254 5323 8256
rect 5343 8254 5359 8274
rect 5269 8248 5359 8254
rect 4783 8225 4820 8226
rect 4004 8223 4041 8224
rect 3465 8195 3555 8201
rect 3465 8175 3481 8195
rect 3501 8193 3555 8195
rect 3501 8175 3526 8193
rect 3465 8173 3526 8175
rect 3546 8173 3555 8193
rect 3465 8167 3555 8173
rect 3478 8113 3515 8114
rect 3574 8113 3611 8114
rect 3630 8113 3666 8223
rect 3853 8202 3884 8223
rect 4782 8216 4820 8225
rect 3849 8201 3884 8202
rect 3727 8191 3884 8201
rect 3727 8171 3744 8191
rect 3764 8171 3884 8191
rect 3727 8164 3884 8171
rect 3951 8194 4100 8202
rect 3951 8174 3962 8194
rect 3982 8174 4021 8194
rect 4041 8174 4100 8194
rect 4610 8198 4650 8208
rect 3951 8167 4100 8174
rect 4166 8170 4218 8188
rect 3951 8166 3992 8167
rect 3685 8113 3722 8114
rect 3378 8104 3516 8113
rect 2850 8093 2883 8095
rect 2479 8081 2926 8093
rect 1711 7959 1879 7961
rect 1435 7933 1879 7959
rect 945 7911 1083 7920
rect 739 7910 776 7911
rect 236 7856 273 7859
rect 469 7857 510 7858
rect 361 7850 510 7857
rect 361 7830 420 7850
rect 440 7830 479 7850
rect 499 7830 510 7850
rect 361 7822 510 7830
rect 577 7853 734 7860
rect 577 7833 697 7853
rect 717 7833 734 7853
rect 577 7823 734 7833
rect 577 7822 612 7823
rect 577 7801 608 7822
rect 795 7801 831 7911
rect 850 7910 887 7911
rect 946 7910 983 7911
rect 906 7851 996 7857
rect 906 7831 915 7851
rect 935 7849 996 7851
rect 935 7831 960 7849
rect 906 7829 960 7831
rect 980 7829 996 7849
rect 906 7823 996 7829
rect 420 7800 457 7801
rect 233 7792 270 7794
rect 233 7784 275 7792
rect 233 7766 243 7784
rect 261 7766 275 7784
rect 233 7757 275 7766
rect 419 7791 457 7800
rect 419 7771 428 7791
rect 448 7771 457 7791
rect 419 7763 457 7771
rect 523 7795 608 7801
rect 638 7800 675 7801
rect 523 7775 531 7795
rect 551 7775 608 7795
rect 523 7767 608 7775
rect 637 7791 675 7800
rect 637 7771 646 7791
rect 666 7771 675 7791
rect 523 7766 559 7767
rect 637 7763 675 7771
rect 741 7799 885 7801
rect 741 7795 793 7799
rect 741 7775 749 7795
rect 769 7779 793 7795
rect 813 7795 885 7799
rect 813 7779 857 7795
rect 769 7775 857 7779
rect 877 7775 885 7795
rect 741 7767 885 7775
rect 741 7766 777 7767
rect 849 7766 885 7767
rect 951 7800 988 7801
rect 951 7799 989 7800
rect 951 7791 1015 7799
rect 951 7771 960 7791
rect 980 7777 1015 7791
rect 1035 7777 1038 7797
rect 980 7772 1038 7777
rect 980 7771 1015 7772
rect 234 7732 275 7757
rect 420 7732 457 7763
rect 638 7732 675 7763
rect 951 7759 1015 7771
rect 1055 7733 1082 7911
rect 234 7705 283 7732
rect 419 7706 468 7732
rect 637 7731 718 7732
rect 914 7731 1082 7733
rect 637 7706 1082 7731
rect 638 7705 1082 7706
rect 236 7672 283 7705
rect 639 7672 679 7705
rect 914 7704 1082 7705
rect 1545 7709 1585 7933
rect 1711 7932 1879 7933
rect 2482 8067 2926 8081
rect 2482 8065 2650 8067
rect 2482 7887 2509 8065
rect 2549 8027 2613 8039
rect 2889 8035 2926 8067
rect 2952 8066 3143 8088
rect 3378 8084 3487 8104
rect 3507 8084 3516 8104
rect 3378 8077 3516 8084
rect 3574 8104 3722 8113
rect 3574 8084 3583 8104
rect 3603 8084 3693 8104
rect 3713 8084 3722 8104
rect 3378 8075 3474 8077
rect 3574 8074 3722 8084
rect 3781 8104 3818 8114
rect 3781 8084 3789 8104
rect 3809 8084 3818 8104
rect 3630 8073 3666 8074
rect 3107 8064 3143 8066
rect 3107 8035 3144 8064
rect 2549 8026 2584 8027
rect 2526 8021 2584 8026
rect 2526 8001 2529 8021
rect 2549 8007 2584 8021
rect 2604 8007 2613 8027
rect 2549 7999 2613 8007
rect 2575 7998 2613 7999
rect 2576 7997 2613 7998
rect 2679 8031 2715 8032
rect 2787 8031 2823 8032
rect 2679 8025 2823 8031
rect 2679 8023 2740 8025
rect 2679 8003 2687 8023
rect 2707 8008 2740 8023
rect 2759 8023 2823 8025
rect 2759 8008 2795 8023
rect 2707 8003 2795 8008
rect 2815 8003 2823 8023
rect 2679 7997 2823 8003
rect 2889 8027 2927 8035
rect 3005 8031 3041 8032
rect 2889 8007 2898 8027
rect 2918 8007 2927 8027
rect 2889 7998 2927 8007
rect 2956 8023 3041 8031
rect 2956 8003 3013 8023
rect 3033 8003 3041 8023
rect 2889 7997 2926 7998
rect 2956 7997 3041 8003
rect 3107 8027 3145 8035
rect 3107 8007 3116 8027
rect 3136 8007 3145 8027
rect 3781 8017 3818 8084
rect 3853 8113 3884 8164
rect 4166 8152 4184 8170
rect 4202 8152 4218 8170
rect 3903 8113 3940 8114
rect 3853 8104 3940 8113
rect 3853 8084 3911 8104
rect 3931 8084 3940 8104
rect 3853 8074 3940 8084
rect 3999 8104 4036 8114
rect 3999 8084 4007 8104
rect 4027 8084 4036 8104
rect 3853 8073 3884 8074
rect 3478 8014 3515 8015
rect 3781 8014 3820 8017
rect 3477 8013 3820 8014
rect 3999 8013 4036 8084
rect 3107 7998 3145 8007
rect 3402 8008 3820 8013
rect 3107 7997 3144 7998
rect 2568 7969 2658 7975
rect 2568 7949 2584 7969
rect 2604 7967 2658 7969
rect 2604 7949 2629 7967
rect 2568 7947 2629 7949
rect 2649 7947 2658 7967
rect 2568 7941 2658 7947
rect 2581 7887 2618 7888
rect 2677 7887 2714 7888
rect 2733 7887 2769 7997
rect 2956 7976 2987 7997
rect 3402 7988 3405 8008
rect 3425 7988 3820 8008
rect 3849 7989 4036 8013
rect 2952 7975 2987 7976
rect 2830 7965 2987 7975
rect 2830 7945 2847 7965
rect 2867 7945 2987 7965
rect 2830 7938 2987 7945
rect 3054 7968 3203 7976
rect 3054 7948 3065 7968
rect 3085 7948 3124 7968
rect 3144 7948 3203 7968
rect 3054 7941 3203 7948
rect 3781 7963 3820 7988
rect 4166 7963 4218 8152
rect 4610 8180 4620 8198
rect 4638 8180 4650 8198
rect 4782 8196 4791 8216
rect 4811 8196 4820 8216
rect 4782 8188 4820 8196
rect 4886 8220 4971 8226
rect 5001 8225 5038 8226
rect 4886 8200 4894 8220
rect 4914 8200 4971 8220
rect 4886 8192 4971 8200
rect 5000 8216 5038 8225
rect 5000 8196 5009 8216
rect 5029 8196 5038 8216
rect 4886 8191 4922 8192
rect 5000 8188 5038 8196
rect 5104 8220 5248 8226
rect 5104 8200 5112 8220
rect 5132 8200 5165 8220
rect 5185 8200 5220 8220
rect 5240 8200 5248 8220
rect 5104 8192 5248 8200
rect 5104 8191 5140 8192
rect 5212 8191 5248 8192
rect 5314 8225 5351 8226
rect 5314 8224 5352 8225
rect 5314 8216 5378 8224
rect 5314 8196 5323 8216
rect 5343 8202 5378 8216
rect 5398 8202 5401 8222
rect 5343 8197 5401 8202
rect 5343 8196 5378 8197
rect 4610 8124 4650 8180
rect 4783 8159 4820 8188
rect 4784 8157 4820 8159
rect 4784 8135 4975 8157
rect 5001 8156 5038 8188
rect 5314 8184 5378 8196
rect 5418 8158 5445 8336
rect 5277 8156 5445 8158
rect 5001 8146 5445 8156
rect 5586 8252 5773 8276
rect 5804 8257 6197 8277
rect 6217 8257 6220 8277
rect 5804 8252 6220 8257
rect 5586 8181 5623 8252
rect 5804 8251 6145 8252
rect 5738 8191 5769 8192
rect 5586 8161 5595 8181
rect 5615 8161 5623 8181
rect 5586 8151 5623 8161
rect 5682 8181 5769 8191
rect 5682 8161 5691 8181
rect 5711 8161 5769 8181
rect 5682 8152 5769 8161
rect 5682 8151 5719 8152
rect 4607 8119 4650 8124
rect 4998 8130 5445 8146
rect 4998 8124 5026 8130
rect 5277 8129 5445 8130
rect 4607 8116 4757 8119
rect 4998 8116 5025 8124
rect 4607 8114 5025 8116
rect 4607 8096 4616 8114
rect 4634 8096 5025 8114
rect 5738 8101 5769 8152
rect 5804 8181 5841 8251
rect 6107 8250 6144 8251
rect 5956 8191 5992 8192
rect 5804 8161 5813 8181
rect 5833 8161 5841 8181
rect 5804 8151 5841 8161
rect 5900 8181 6048 8191
rect 6148 8188 6244 8190
rect 5900 8161 5909 8181
rect 5929 8161 6019 8181
rect 6039 8161 6048 8181
rect 5900 8152 6048 8161
rect 6106 8181 6244 8188
rect 6106 8161 6115 8181
rect 6135 8161 6244 8181
rect 6106 8152 6244 8161
rect 5900 8151 5937 8152
rect 5630 8098 5671 8099
rect 4607 8093 5025 8096
rect 4607 8087 4650 8093
rect 4610 8084 4650 8087
rect 5522 8091 5671 8098
rect 5007 8075 5047 8076
rect 4718 8058 5047 8075
rect 5522 8071 5581 8091
rect 5601 8071 5640 8091
rect 5660 8071 5671 8091
rect 5522 8063 5671 8071
rect 5738 8094 5895 8101
rect 5738 8074 5858 8094
rect 5878 8074 5895 8094
rect 5738 8064 5895 8074
rect 5738 8063 5773 8064
rect 4602 8015 4645 8026
rect 4602 7997 4614 8015
rect 4632 7997 4645 8015
rect 4602 7971 4645 7997
rect 4718 7971 4745 8058
rect 5007 8049 5047 8058
rect 3781 7945 4220 7963
rect 3054 7940 3095 7941
rect 2788 7887 2825 7888
rect 2481 7878 2619 7887
rect 2481 7858 2590 7878
rect 2610 7858 2619 7878
rect 2481 7851 2619 7858
rect 2677 7878 2825 7887
rect 2677 7858 2686 7878
rect 2706 7858 2796 7878
rect 2816 7858 2825 7878
rect 2481 7849 2577 7851
rect 2677 7848 2825 7858
rect 2884 7878 2921 7888
rect 2884 7858 2892 7878
rect 2912 7858 2921 7878
rect 2733 7847 2769 7848
rect 2581 7788 2618 7789
rect 2884 7788 2921 7858
rect 2956 7887 2987 7938
rect 3781 7927 4181 7945
rect 4199 7927 4220 7945
rect 3781 7921 4220 7927
rect 3787 7917 4220 7921
rect 4602 7950 4745 7971
rect 4789 8023 4823 8039
rect 5007 8029 5400 8049
rect 5420 8029 5423 8049
rect 5738 8042 5769 8063
rect 5956 8042 5992 8152
rect 6011 8151 6048 8152
rect 6107 8151 6144 8152
rect 6067 8092 6157 8098
rect 6067 8072 6076 8092
rect 6096 8090 6157 8092
rect 6096 8072 6121 8090
rect 6067 8070 6121 8072
rect 6141 8070 6157 8090
rect 6067 8064 6157 8070
rect 5581 8041 5618 8042
rect 5007 8024 5423 8029
rect 5580 8032 5618 8041
rect 5007 8023 5348 8024
rect 4789 7953 4826 8023
rect 4941 7963 4972 7964
rect 4602 7948 4739 7950
rect 4166 7915 4218 7917
rect 4602 7906 4645 7948
rect 4789 7933 4798 7953
rect 4818 7933 4826 7953
rect 4789 7923 4826 7933
rect 4885 7953 4972 7963
rect 4885 7933 4894 7953
rect 4914 7933 4972 7953
rect 4885 7924 4972 7933
rect 4885 7923 4922 7924
rect 4600 7896 4645 7906
rect 3006 7887 3043 7888
rect 2956 7878 3043 7887
rect 2956 7858 3014 7878
rect 3034 7858 3043 7878
rect 2956 7848 3043 7858
rect 3102 7878 3139 7888
rect 3102 7858 3110 7878
rect 3130 7858 3139 7878
rect 4600 7878 4609 7896
rect 4627 7878 4645 7896
rect 4600 7872 4645 7878
rect 4941 7873 4972 7924
rect 5007 7953 5044 8023
rect 5310 8022 5347 8023
rect 5580 8012 5589 8032
rect 5609 8012 5618 8032
rect 5580 8004 5618 8012
rect 5684 8036 5769 8042
rect 5799 8041 5836 8042
rect 5684 8016 5692 8036
rect 5712 8016 5769 8036
rect 5684 8008 5769 8016
rect 5798 8032 5836 8041
rect 5798 8012 5807 8032
rect 5827 8012 5836 8032
rect 5684 8007 5720 8008
rect 5798 8004 5836 8012
rect 5902 8036 6046 8042
rect 5902 8016 5910 8036
rect 5930 8017 5962 8036
rect 5983 8017 6018 8036
rect 5930 8016 6018 8017
rect 6038 8016 6046 8036
rect 5902 8008 6046 8016
rect 5902 8007 5938 8008
rect 6010 8007 6046 8008
rect 6112 8041 6149 8042
rect 6112 8040 6150 8041
rect 6112 8032 6176 8040
rect 6112 8012 6121 8032
rect 6141 8018 6176 8032
rect 6196 8018 6199 8038
rect 6141 8013 6199 8018
rect 6141 8012 6176 8013
rect 5581 7975 5618 8004
rect 5582 7973 5618 7975
rect 5159 7963 5195 7964
rect 5007 7933 5016 7953
rect 5036 7933 5044 7953
rect 5007 7923 5044 7933
rect 5103 7953 5251 7963
rect 5351 7960 5447 7962
rect 5103 7933 5112 7953
rect 5132 7933 5222 7953
rect 5242 7933 5251 7953
rect 5103 7924 5251 7933
rect 5309 7953 5447 7960
rect 5309 7933 5318 7953
rect 5338 7933 5447 7953
rect 5582 7951 5773 7973
rect 5799 7972 5836 8004
rect 6112 8000 6176 8012
rect 6216 7974 6243 8152
rect 6848 8151 6881 8484
rect 6945 8516 7113 8517
rect 7239 8516 7279 8740
rect 7742 8744 7910 8745
rect 7742 8743 8186 8744
rect 8549 8743 8590 8744
rect 7742 8718 8590 8743
rect 7742 8716 7910 8718
rect 8106 8717 8590 8718
rect 7742 8538 7769 8716
rect 7809 8678 7873 8690
rect 8149 8686 8186 8717
rect 8367 8686 8404 8717
rect 8549 8692 8590 8717
rect 7809 8677 7844 8678
rect 7786 8672 7844 8677
rect 7786 8652 7789 8672
rect 7809 8658 7844 8672
rect 7864 8658 7873 8678
rect 7809 8650 7873 8658
rect 7835 8649 7873 8650
rect 7836 8648 7873 8649
rect 7939 8682 7975 8683
rect 8047 8682 8083 8683
rect 7939 8674 8083 8682
rect 7939 8654 7947 8674
rect 7967 8670 8055 8674
rect 7967 8654 8011 8670
rect 7939 8650 8011 8654
rect 8031 8654 8055 8670
rect 8075 8654 8083 8674
rect 8031 8650 8083 8654
rect 7939 8648 8083 8650
rect 8149 8678 8187 8686
rect 8265 8682 8301 8683
rect 8149 8658 8158 8678
rect 8178 8658 8187 8678
rect 8149 8649 8187 8658
rect 8216 8674 8301 8682
rect 8216 8654 8273 8674
rect 8293 8654 8301 8674
rect 8149 8648 8186 8649
rect 8216 8648 8301 8654
rect 8367 8678 8405 8686
rect 8367 8658 8376 8678
rect 8396 8658 8405 8678
rect 8367 8649 8405 8658
rect 8549 8683 8591 8692
rect 8549 8665 8563 8683
rect 8581 8665 8591 8683
rect 8549 8657 8591 8665
rect 8554 8655 8591 8657
rect 8367 8648 8404 8649
rect 7828 8620 7918 8626
rect 7828 8600 7844 8620
rect 7864 8618 7918 8620
rect 7864 8600 7889 8618
rect 7828 8598 7889 8600
rect 7909 8598 7918 8618
rect 7828 8592 7918 8598
rect 7841 8538 7878 8539
rect 7937 8538 7974 8539
rect 7993 8538 8029 8648
rect 8216 8627 8247 8648
rect 8212 8626 8247 8627
rect 8090 8616 8247 8626
rect 8090 8596 8107 8616
rect 8127 8596 8247 8616
rect 8090 8589 8247 8596
rect 8314 8619 8463 8627
rect 8314 8599 8325 8619
rect 8345 8599 8384 8619
rect 8404 8599 8463 8619
rect 8314 8592 8463 8599
rect 8314 8591 8355 8592
rect 8551 8590 8588 8593
rect 8048 8538 8085 8539
rect 7741 8529 7879 8538
rect 6945 8490 7389 8516
rect 6945 8488 7113 8490
rect 6945 8310 6972 8488
rect 7012 8450 7076 8462
rect 7352 8458 7389 8490
rect 7415 8489 7606 8511
rect 7741 8509 7850 8529
rect 7870 8509 7879 8529
rect 7741 8502 7879 8509
rect 7937 8529 8085 8538
rect 7937 8509 7946 8529
rect 7966 8509 8056 8529
rect 8076 8509 8085 8529
rect 7741 8500 7837 8502
rect 7937 8499 8085 8509
rect 8144 8529 8181 8539
rect 8144 8509 8152 8529
rect 8172 8509 8181 8529
rect 7993 8498 8029 8499
rect 7570 8487 7606 8489
rect 7570 8458 7607 8487
rect 7012 8449 7047 8450
rect 6989 8444 7047 8449
rect 6989 8424 6992 8444
rect 7012 8430 7047 8444
rect 7067 8430 7076 8450
rect 7012 8424 7076 8430
rect 6989 8422 7076 8424
rect 6989 8418 7016 8422
rect 7038 8421 7076 8422
rect 7039 8420 7076 8421
rect 7142 8454 7178 8455
rect 7250 8454 7286 8455
rect 7142 8447 7286 8454
rect 7142 8446 7204 8447
rect 7142 8426 7150 8446
rect 7170 8429 7204 8446
rect 7223 8446 7286 8447
rect 7223 8429 7258 8446
rect 7170 8426 7258 8429
rect 7278 8426 7286 8446
rect 7142 8420 7286 8426
rect 7352 8450 7390 8458
rect 7468 8454 7504 8455
rect 7352 8430 7361 8450
rect 7381 8430 7390 8450
rect 7352 8421 7390 8430
rect 7419 8446 7504 8454
rect 7419 8426 7476 8446
rect 7496 8426 7504 8446
rect 7352 8420 7389 8421
rect 7419 8420 7504 8426
rect 7570 8450 7608 8458
rect 7570 8430 7579 8450
rect 7599 8430 7608 8450
rect 7841 8439 7878 8440
rect 8144 8439 8181 8509
rect 8216 8538 8247 8589
rect 8543 8584 8588 8590
rect 8543 8566 8561 8584
rect 8579 8566 8588 8584
rect 8543 8556 8588 8566
rect 8266 8538 8303 8539
rect 8216 8529 8303 8538
rect 8216 8509 8274 8529
rect 8294 8509 8303 8529
rect 8216 8499 8303 8509
rect 8362 8529 8399 8539
rect 8362 8509 8370 8529
rect 8390 8509 8399 8529
rect 8543 8514 8586 8556
rect 8449 8512 8586 8514
rect 8216 8498 8247 8499
rect 8362 8439 8399 8509
rect 7840 8438 8181 8439
rect 7570 8421 7608 8430
rect 7765 8433 8181 8438
rect 7570 8420 7607 8421
rect 7031 8392 7121 8398
rect 7031 8372 7047 8392
rect 7067 8390 7121 8392
rect 7067 8372 7092 8390
rect 7031 8370 7092 8372
rect 7112 8370 7121 8390
rect 7031 8364 7121 8370
rect 7044 8310 7081 8311
rect 7140 8310 7177 8311
rect 7196 8310 7232 8420
rect 7419 8399 7450 8420
rect 7765 8413 7768 8433
rect 7788 8413 8181 8433
rect 8365 8423 8399 8439
rect 8443 8491 8586 8512
rect 8141 8404 8181 8413
rect 8443 8404 8470 8491
rect 8543 8465 8586 8491
rect 8543 8447 8556 8465
rect 8574 8447 8586 8465
rect 8543 8436 8586 8447
rect 7415 8398 7450 8399
rect 7293 8388 7450 8398
rect 7293 8368 7310 8388
rect 7330 8368 7450 8388
rect 7293 8361 7450 8368
rect 7517 8391 7663 8399
rect 7517 8371 7528 8391
rect 7548 8371 7587 8391
rect 7607 8371 7663 8391
rect 8141 8387 8470 8404
rect 8141 8386 8181 8387
rect 7517 8364 7663 8371
rect 8538 8375 8578 8378
rect 8538 8369 8581 8375
rect 8163 8366 8581 8369
rect 7517 8363 7558 8364
rect 7251 8310 7288 8311
rect 6944 8301 7082 8310
rect 6944 8281 7053 8301
rect 7073 8281 7082 8301
rect 6944 8274 7082 8281
rect 7140 8301 7288 8310
rect 7140 8281 7149 8301
rect 7169 8281 7259 8301
rect 7279 8281 7288 8301
rect 6944 8272 7040 8274
rect 7140 8271 7288 8281
rect 7347 8301 7384 8311
rect 7347 8281 7355 8301
rect 7375 8281 7384 8301
rect 7196 8270 7232 8271
rect 7044 8211 7081 8212
rect 7347 8211 7384 8281
rect 7419 8310 7450 8361
rect 8163 8348 8554 8366
rect 8572 8348 8581 8366
rect 8163 8346 8581 8348
rect 8163 8338 8190 8346
rect 8431 8343 8581 8346
rect 7743 8332 7911 8333
rect 8162 8332 8190 8338
rect 7743 8316 8190 8332
rect 8538 8338 8581 8343
rect 7469 8310 7506 8311
rect 7419 8301 7506 8310
rect 7419 8281 7477 8301
rect 7497 8281 7506 8301
rect 7419 8271 7506 8281
rect 7565 8301 7602 8311
rect 7565 8281 7573 8301
rect 7593 8281 7602 8301
rect 7419 8270 7450 8271
rect 7043 8210 7384 8211
rect 7565 8210 7602 8281
rect 6968 8205 7384 8210
rect 6968 8185 6971 8205
rect 6991 8185 7384 8205
rect 7415 8186 7602 8210
rect 7743 8306 8187 8316
rect 7743 8304 7911 8306
rect 6843 8106 6885 8151
rect 7743 8126 7770 8304
rect 7810 8266 7874 8278
rect 8150 8274 8187 8306
rect 8213 8305 8404 8327
rect 8368 8303 8404 8305
rect 8368 8274 8405 8303
rect 8538 8282 8578 8338
rect 7810 8265 7845 8266
rect 7787 8260 7845 8265
rect 7787 8240 7790 8260
rect 7810 8246 7845 8260
rect 7865 8246 7874 8266
rect 7810 8238 7874 8246
rect 7836 8237 7874 8238
rect 7837 8236 7874 8237
rect 7940 8270 7976 8271
rect 8048 8270 8084 8271
rect 7940 8262 8084 8270
rect 7940 8242 7948 8262
rect 7968 8242 8003 8262
rect 8023 8242 8056 8262
rect 8076 8242 8084 8262
rect 7940 8236 8084 8242
rect 8150 8266 8188 8274
rect 8266 8270 8302 8271
rect 8150 8246 8159 8266
rect 8179 8246 8188 8266
rect 8150 8237 8188 8246
rect 8217 8262 8302 8270
rect 8217 8242 8274 8262
rect 8294 8242 8302 8262
rect 8150 8236 8187 8237
rect 8217 8236 8302 8242
rect 8368 8266 8406 8274
rect 8368 8246 8377 8266
rect 8397 8246 8406 8266
rect 8538 8264 8550 8282
rect 8568 8264 8578 8282
rect 8538 8254 8578 8264
rect 8368 8237 8406 8246
rect 8368 8236 8405 8237
rect 7829 8208 7919 8214
rect 7829 8188 7845 8208
rect 7865 8206 7919 8208
rect 7865 8188 7890 8206
rect 7829 8186 7890 8188
rect 7910 8186 7919 8206
rect 7829 8180 7919 8186
rect 7842 8126 7879 8127
rect 7938 8126 7975 8127
rect 7994 8126 8030 8236
rect 8217 8215 8248 8236
rect 8213 8214 8248 8215
rect 8091 8204 8248 8214
rect 8091 8184 8108 8204
rect 8128 8184 8248 8204
rect 8091 8177 8248 8184
rect 8315 8207 8464 8215
rect 8315 8187 8326 8207
rect 8346 8187 8385 8207
rect 8405 8187 8464 8207
rect 8315 8180 8464 8187
rect 8530 8183 8582 8201
rect 8315 8179 8356 8180
rect 8049 8126 8086 8127
rect 7742 8117 7880 8126
rect 7214 8106 7247 8108
rect 6843 8094 7290 8106
rect 6075 7972 6243 7974
rect 5799 7946 6243 7972
rect 5309 7924 5447 7933
rect 5103 7923 5140 7924
rect 4600 7869 4637 7872
rect 4833 7870 4874 7871
rect 2956 7847 2987 7848
rect 2580 7787 2921 7788
rect 3102 7787 3139 7858
rect 4725 7863 4874 7870
rect 4169 7850 4206 7855
rect 4160 7846 4207 7850
rect 4160 7828 4179 7846
rect 4197 7828 4207 7846
rect 4725 7843 4784 7863
rect 4804 7843 4843 7863
rect 4863 7843 4874 7863
rect 4725 7835 4874 7843
rect 4941 7866 5098 7873
rect 4941 7846 5061 7866
rect 5081 7846 5098 7866
rect 4941 7836 5098 7846
rect 4941 7835 4976 7836
rect 2505 7782 2921 7787
rect 2505 7762 2508 7782
rect 2528 7762 2921 7782
rect 2952 7763 3139 7787
rect 3764 7785 3804 7790
rect 4160 7785 4207 7828
rect 4941 7814 4972 7835
rect 5159 7814 5195 7924
rect 5214 7923 5251 7924
rect 5310 7923 5347 7924
rect 5270 7864 5360 7870
rect 5270 7844 5279 7864
rect 5299 7862 5360 7864
rect 5299 7844 5324 7862
rect 5270 7842 5324 7844
rect 5344 7842 5360 7862
rect 5270 7836 5360 7842
rect 4784 7813 4821 7814
rect 3764 7746 4207 7785
rect 4597 7805 4634 7807
rect 4597 7797 4639 7805
rect 4597 7779 4607 7797
rect 4625 7779 4639 7797
rect 4597 7770 4639 7779
rect 4783 7804 4821 7813
rect 4783 7784 4792 7804
rect 4812 7784 4821 7804
rect 4783 7776 4821 7784
rect 4887 7808 4972 7814
rect 5002 7813 5039 7814
rect 4887 7788 4895 7808
rect 4915 7788 4972 7808
rect 4887 7780 4972 7788
rect 5001 7804 5039 7813
rect 5001 7784 5010 7804
rect 5030 7784 5039 7804
rect 4887 7779 4923 7780
rect 5001 7776 5039 7784
rect 5105 7812 5249 7814
rect 5105 7808 5157 7812
rect 5105 7788 5113 7808
rect 5133 7792 5157 7808
rect 5177 7808 5249 7812
rect 5177 7792 5221 7808
rect 5133 7788 5221 7792
rect 5241 7788 5249 7808
rect 5105 7780 5249 7788
rect 5105 7779 5141 7780
rect 5213 7779 5249 7780
rect 5315 7813 5352 7814
rect 5315 7812 5353 7813
rect 5315 7804 5379 7812
rect 5315 7784 5324 7804
rect 5344 7790 5379 7804
rect 5399 7790 5402 7810
rect 5344 7785 5402 7790
rect 5344 7784 5379 7785
rect 1545 7687 1553 7709
rect 1577 7687 1585 7709
rect 1545 7679 1585 7687
rect 2858 7731 2898 7739
rect 2858 7709 2866 7731
rect 2890 7709 2898 7731
rect 236 7633 679 7672
rect 236 7590 283 7633
rect 639 7628 679 7633
rect 1304 7631 1491 7655
rect 1522 7636 1915 7656
rect 1935 7636 1938 7656
rect 1522 7631 1938 7636
rect 236 7572 246 7590
rect 264 7572 283 7590
rect 236 7568 283 7572
rect 237 7563 274 7568
rect 1304 7560 1341 7631
rect 1522 7630 1863 7631
rect 1456 7570 1487 7571
rect 1304 7540 1313 7560
rect 1333 7540 1341 7560
rect 1304 7530 1341 7540
rect 1400 7560 1487 7570
rect 1400 7540 1409 7560
rect 1429 7540 1487 7560
rect 1400 7531 1487 7540
rect 1400 7530 1437 7531
rect 225 7501 277 7503
rect 223 7497 656 7501
rect 223 7491 662 7497
rect 223 7473 244 7491
rect 262 7473 662 7491
rect 1456 7480 1487 7531
rect 1522 7560 1559 7630
rect 1825 7629 1862 7630
rect 1674 7570 1710 7571
rect 1522 7540 1531 7560
rect 1551 7540 1559 7560
rect 1522 7530 1559 7540
rect 1618 7560 1766 7570
rect 1866 7567 1962 7569
rect 1618 7540 1627 7560
rect 1647 7540 1737 7560
rect 1757 7540 1766 7560
rect 1618 7531 1766 7540
rect 1824 7560 1962 7567
rect 1824 7540 1833 7560
rect 1853 7540 1962 7560
rect 1824 7531 1962 7540
rect 1618 7530 1655 7531
rect 1348 7477 1389 7478
rect 223 7455 662 7473
rect 225 7266 277 7455
rect 623 7430 662 7455
rect 1240 7470 1389 7477
rect 1240 7450 1299 7470
rect 1319 7450 1358 7470
rect 1378 7450 1389 7470
rect 1240 7442 1389 7450
rect 1456 7473 1613 7480
rect 1456 7453 1576 7473
rect 1596 7453 1613 7473
rect 1456 7443 1613 7453
rect 1456 7442 1491 7443
rect 407 7405 594 7429
rect 623 7410 1018 7430
rect 1038 7410 1041 7430
rect 1456 7421 1487 7442
rect 1674 7421 1710 7531
rect 1729 7530 1766 7531
rect 1825 7530 1862 7531
rect 1785 7471 1875 7477
rect 1785 7451 1794 7471
rect 1814 7469 1875 7471
rect 1814 7451 1839 7469
rect 1785 7449 1839 7451
rect 1859 7449 1875 7469
rect 1785 7443 1875 7449
rect 1299 7420 1336 7421
rect 623 7405 1041 7410
rect 1298 7411 1336 7420
rect 407 7334 444 7405
rect 623 7404 966 7405
rect 623 7401 662 7404
rect 928 7403 965 7404
rect 559 7344 590 7345
rect 407 7314 416 7334
rect 436 7314 444 7334
rect 407 7304 444 7314
rect 503 7334 590 7344
rect 503 7314 512 7334
rect 532 7314 590 7334
rect 503 7305 590 7314
rect 503 7304 540 7305
rect 225 7248 241 7266
rect 259 7248 277 7266
rect 559 7254 590 7305
rect 625 7334 662 7401
rect 1298 7391 1307 7411
rect 1327 7391 1336 7411
rect 1298 7383 1336 7391
rect 1402 7415 1487 7421
rect 1517 7420 1554 7421
rect 1402 7395 1410 7415
rect 1430 7395 1487 7415
rect 1402 7387 1487 7395
rect 1516 7411 1554 7420
rect 1516 7391 1525 7411
rect 1545 7391 1554 7411
rect 1402 7386 1438 7387
rect 1516 7383 1554 7391
rect 1620 7416 1764 7421
rect 1620 7415 1682 7416
rect 1620 7395 1628 7415
rect 1648 7397 1682 7415
rect 1703 7415 1764 7416
rect 1703 7397 1736 7415
rect 1648 7395 1736 7397
rect 1756 7395 1764 7415
rect 1620 7387 1764 7395
rect 1620 7386 1656 7387
rect 1728 7386 1764 7387
rect 1830 7420 1867 7421
rect 1830 7419 1868 7420
rect 1830 7411 1894 7419
rect 1830 7391 1839 7411
rect 1859 7397 1894 7411
rect 1914 7397 1917 7417
rect 1859 7392 1917 7397
rect 1859 7391 1894 7392
rect 1299 7354 1336 7383
rect 1300 7352 1336 7354
rect 777 7344 813 7345
rect 625 7314 634 7334
rect 654 7314 662 7334
rect 625 7304 662 7314
rect 721 7334 869 7344
rect 969 7341 1065 7343
rect 721 7314 730 7334
rect 750 7314 840 7334
rect 860 7314 869 7334
rect 721 7305 869 7314
rect 927 7334 1065 7341
rect 927 7314 936 7334
rect 956 7314 1065 7334
rect 1300 7330 1491 7352
rect 1517 7351 1554 7383
rect 1830 7379 1894 7391
rect 1934 7353 1961 7531
rect 1793 7351 1961 7353
rect 1517 7337 1961 7351
rect 2564 7485 2732 7486
rect 2858 7485 2898 7709
rect 3361 7713 3529 7714
rect 3764 7713 3804 7746
rect 4160 7713 4207 7746
rect 4598 7745 4639 7770
rect 4784 7745 4821 7776
rect 5002 7745 5039 7776
rect 5315 7772 5379 7784
rect 5419 7746 5446 7924
rect 4598 7718 4647 7745
rect 4783 7719 4832 7745
rect 5001 7744 5082 7745
rect 5278 7744 5446 7746
rect 5001 7719 5446 7744
rect 5002 7718 5446 7719
rect 3361 7712 3805 7713
rect 3361 7687 3806 7712
rect 3361 7685 3529 7687
rect 3725 7686 3806 7687
rect 3975 7686 4024 7712
rect 4160 7686 4209 7713
rect 3361 7507 3388 7685
rect 3428 7647 3492 7659
rect 3768 7655 3805 7686
rect 3986 7655 4023 7686
rect 4168 7661 4209 7686
rect 4600 7685 4647 7718
rect 5003 7685 5043 7718
rect 5278 7717 5446 7718
rect 5909 7722 5949 7946
rect 6075 7945 6243 7946
rect 6846 8080 7290 8094
rect 6846 8078 7014 8080
rect 6846 7900 6873 8078
rect 6913 8040 6977 8052
rect 7253 8048 7290 8080
rect 7316 8079 7507 8101
rect 7742 8097 7851 8117
rect 7871 8097 7880 8117
rect 7742 8090 7880 8097
rect 7938 8117 8086 8126
rect 7938 8097 7947 8117
rect 7967 8097 8057 8117
rect 8077 8097 8086 8117
rect 7742 8088 7838 8090
rect 7938 8087 8086 8097
rect 8145 8117 8182 8127
rect 8145 8097 8153 8117
rect 8173 8097 8182 8117
rect 7994 8086 8030 8087
rect 7471 8077 7507 8079
rect 7471 8048 7508 8077
rect 6913 8039 6948 8040
rect 6890 8034 6948 8039
rect 6890 8014 6893 8034
rect 6913 8020 6948 8034
rect 6968 8020 6977 8040
rect 6913 8012 6977 8020
rect 6939 8011 6977 8012
rect 6940 8010 6977 8011
rect 7043 8044 7079 8045
rect 7151 8044 7187 8045
rect 7043 8038 7187 8044
rect 7043 8036 7104 8038
rect 7043 8016 7051 8036
rect 7071 8021 7104 8036
rect 7123 8036 7187 8038
rect 7123 8021 7159 8036
rect 7071 8016 7159 8021
rect 7179 8016 7187 8036
rect 7043 8010 7187 8016
rect 7253 8040 7291 8048
rect 7369 8044 7405 8045
rect 7253 8020 7262 8040
rect 7282 8020 7291 8040
rect 7253 8011 7291 8020
rect 7320 8036 7405 8044
rect 7320 8016 7377 8036
rect 7397 8016 7405 8036
rect 7253 8010 7290 8011
rect 7320 8010 7405 8016
rect 7471 8040 7509 8048
rect 7471 8020 7480 8040
rect 7500 8020 7509 8040
rect 8145 8030 8182 8097
rect 8217 8126 8248 8177
rect 8530 8165 8548 8183
rect 8566 8165 8582 8183
rect 8267 8126 8304 8127
rect 8217 8117 8304 8126
rect 8217 8097 8275 8117
rect 8295 8097 8304 8117
rect 8217 8087 8304 8097
rect 8363 8117 8400 8127
rect 8363 8097 8371 8117
rect 8391 8097 8400 8117
rect 8217 8086 8248 8087
rect 7842 8027 7879 8028
rect 8145 8027 8184 8030
rect 7841 8026 8184 8027
rect 8363 8026 8400 8097
rect 7471 8011 7509 8020
rect 7766 8021 8184 8026
rect 7471 8010 7508 8011
rect 6932 7982 7022 7988
rect 6932 7962 6948 7982
rect 6968 7980 7022 7982
rect 6968 7962 6993 7980
rect 6932 7960 6993 7962
rect 7013 7960 7022 7980
rect 6932 7954 7022 7960
rect 6945 7900 6982 7901
rect 7041 7900 7078 7901
rect 7097 7900 7133 8010
rect 7320 7989 7351 8010
rect 7766 8001 7769 8021
rect 7789 8001 8184 8021
rect 8213 8002 8400 8026
rect 7316 7988 7351 7989
rect 7194 7978 7351 7988
rect 7194 7958 7211 7978
rect 7231 7958 7351 7978
rect 7194 7951 7351 7958
rect 7418 7981 7567 7989
rect 7418 7961 7429 7981
rect 7449 7961 7488 7981
rect 7508 7961 7567 7981
rect 7418 7954 7567 7961
rect 8145 7976 8184 8001
rect 8530 7976 8582 8165
rect 8145 7958 8584 7976
rect 7418 7953 7459 7954
rect 7152 7900 7189 7901
rect 6845 7891 6983 7900
rect 6845 7871 6954 7891
rect 6974 7871 6983 7891
rect 6845 7864 6983 7871
rect 7041 7891 7189 7900
rect 7041 7871 7050 7891
rect 7070 7871 7160 7891
rect 7180 7871 7189 7891
rect 6845 7862 6941 7864
rect 7041 7861 7189 7871
rect 7248 7891 7285 7901
rect 7248 7871 7256 7891
rect 7276 7871 7285 7891
rect 7097 7860 7133 7861
rect 6945 7801 6982 7802
rect 7248 7801 7285 7871
rect 7320 7900 7351 7951
rect 8145 7940 8545 7958
rect 8563 7940 8584 7958
rect 8145 7934 8584 7940
rect 8151 7930 8584 7934
rect 8530 7928 8582 7930
rect 7370 7900 7407 7901
rect 7320 7891 7407 7900
rect 7320 7871 7378 7891
rect 7398 7871 7407 7891
rect 7320 7861 7407 7871
rect 7466 7891 7503 7901
rect 7466 7871 7474 7891
rect 7494 7871 7503 7891
rect 7320 7860 7351 7861
rect 6944 7800 7285 7801
rect 7466 7800 7503 7871
rect 8533 7863 8570 7868
rect 8524 7859 8571 7863
rect 8524 7841 8543 7859
rect 8561 7841 8571 7859
rect 6869 7795 7285 7800
rect 6869 7775 6872 7795
rect 6892 7775 7285 7795
rect 7316 7776 7503 7800
rect 8128 7798 8168 7803
rect 8524 7798 8571 7841
rect 8128 7759 8571 7798
rect 5909 7700 5917 7722
rect 5941 7700 5949 7722
rect 5909 7692 5949 7700
rect 7222 7744 7262 7752
rect 7222 7722 7230 7744
rect 7254 7722 7262 7744
rect 3428 7646 3463 7647
rect 3405 7641 3463 7646
rect 3405 7621 3408 7641
rect 3428 7627 3463 7641
rect 3483 7627 3492 7647
rect 3428 7619 3492 7627
rect 3454 7618 3492 7619
rect 3455 7617 3492 7618
rect 3558 7651 3594 7652
rect 3666 7651 3702 7652
rect 3558 7643 3702 7651
rect 3558 7623 3566 7643
rect 3586 7639 3674 7643
rect 3586 7623 3630 7639
rect 3558 7619 3630 7623
rect 3650 7623 3674 7639
rect 3694 7623 3702 7643
rect 3650 7619 3702 7623
rect 3558 7617 3702 7619
rect 3768 7647 3806 7655
rect 3884 7651 3920 7652
rect 3768 7627 3777 7647
rect 3797 7627 3806 7647
rect 3768 7618 3806 7627
rect 3835 7643 3920 7651
rect 3835 7623 3892 7643
rect 3912 7623 3920 7643
rect 3768 7617 3805 7618
rect 3835 7617 3920 7623
rect 3986 7647 4024 7655
rect 3986 7627 3995 7647
rect 4015 7627 4024 7647
rect 3986 7618 4024 7627
rect 4168 7652 4210 7661
rect 4168 7634 4182 7652
rect 4200 7634 4210 7652
rect 4168 7626 4210 7634
rect 4173 7624 4210 7626
rect 4600 7646 5043 7685
rect 3986 7617 4023 7618
rect 3447 7589 3537 7595
rect 3447 7569 3463 7589
rect 3483 7587 3537 7589
rect 3483 7569 3508 7587
rect 3447 7567 3508 7569
rect 3528 7567 3537 7587
rect 3447 7561 3537 7567
rect 3460 7507 3497 7508
rect 3556 7507 3593 7508
rect 3612 7507 3648 7617
rect 3835 7596 3866 7617
rect 4600 7603 4647 7646
rect 5003 7641 5043 7646
rect 5668 7644 5855 7668
rect 5886 7649 6279 7669
rect 6299 7649 6302 7669
rect 5886 7644 6302 7649
rect 3831 7595 3866 7596
rect 3709 7585 3866 7595
rect 3709 7565 3726 7585
rect 3746 7565 3866 7585
rect 3709 7558 3866 7565
rect 3933 7588 4082 7596
rect 3933 7568 3944 7588
rect 3964 7568 4003 7588
rect 4023 7568 4082 7588
rect 4600 7585 4610 7603
rect 4628 7585 4647 7603
rect 4600 7581 4647 7585
rect 4601 7576 4638 7581
rect 3933 7561 4082 7568
rect 5668 7573 5705 7644
rect 5886 7643 6227 7644
rect 5820 7583 5851 7584
rect 3933 7560 3974 7561
rect 4170 7559 4207 7562
rect 3667 7507 3704 7508
rect 3360 7498 3498 7507
rect 2564 7459 3008 7485
rect 2564 7457 2732 7459
rect 1517 7325 1964 7337
rect 1560 7323 1593 7325
rect 927 7305 1065 7314
rect 721 7304 758 7305
rect 451 7251 492 7252
rect 225 7230 277 7248
rect 343 7244 492 7251
rect 343 7224 402 7244
rect 422 7224 461 7244
rect 481 7224 492 7244
rect 343 7216 492 7224
rect 559 7247 716 7254
rect 559 7227 679 7247
rect 699 7227 716 7247
rect 559 7217 716 7227
rect 559 7216 594 7217
rect 559 7195 590 7216
rect 777 7195 813 7305
rect 832 7304 869 7305
rect 928 7304 965 7305
rect 888 7245 978 7251
rect 888 7225 897 7245
rect 917 7243 978 7245
rect 917 7225 942 7243
rect 888 7223 942 7225
rect 962 7223 978 7243
rect 888 7217 978 7223
rect 402 7194 439 7195
rect 401 7185 439 7194
rect 229 7167 269 7177
rect 229 7149 239 7167
rect 257 7149 269 7167
rect 401 7165 410 7185
rect 430 7165 439 7185
rect 401 7157 439 7165
rect 505 7189 590 7195
rect 620 7194 657 7195
rect 505 7169 513 7189
rect 533 7169 590 7189
rect 505 7161 590 7169
rect 619 7185 657 7194
rect 619 7165 628 7185
rect 648 7165 657 7185
rect 505 7160 541 7161
rect 619 7157 657 7165
rect 723 7189 867 7195
rect 723 7169 731 7189
rect 751 7169 784 7189
rect 804 7169 839 7189
rect 859 7169 867 7189
rect 723 7161 867 7169
rect 723 7160 759 7161
rect 831 7160 867 7161
rect 933 7194 970 7195
rect 933 7193 971 7194
rect 933 7185 997 7193
rect 933 7165 942 7185
rect 962 7171 997 7185
rect 1017 7171 1020 7191
rect 962 7166 1020 7171
rect 962 7165 997 7166
rect 229 7093 269 7149
rect 402 7128 439 7157
rect 403 7126 439 7128
rect 403 7104 594 7126
rect 620 7125 657 7157
rect 933 7153 997 7165
rect 1037 7127 1064 7305
rect 1922 7280 1964 7325
rect 896 7125 1064 7127
rect 620 7115 1064 7125
rect 1205 7221 1392 7245
rect 1423 7226 1816 7246
rect 1836 7226 1839 7246
rect 1423 7221 1839 7226
rect 1205 7150 1242 7221
rect 1423 7220 1764 7221
rect 1357 7160 1388 7161
rect 1205 7130 1214 7150
rect 1234 7130 1242 7150
rect 1205 7120 1242 7130
rect 1301 7150 1388 7160
rect 1301 7130 1310 7150
rect 1330 7130 1388 7150
rect 1301 7121 1388 7130
rect 1301 7120 1338 7121
rect 226 7088 269 7093
rect 617 7099 1064 7115
rect 617 7093 645 7099
rect 896 7098 1064 7099
rect 226 7085 376 7088
rect 617 7085 644 7093
rect 226 7083 644 7085
rect 226 7065 235 7083
rect 253 7065 644 7083
rect 1357 7070 1388 7121
rect 1423 7150 1460 7220
rect 1726 7219 1763 7220
rect 1575 7160 1611 7161
rect 1423 7130 1432 7150
rect 1452 7130 1460 7150
rect 1423 7120 1460 7130
rect 1519 7150 1667 7160
rect 1767 7157 1863 7159
rect 1519 7130 1528 7150
rect 1548 7130 1638 7150
rect 1658 7130 1667 7150
rect 1519 7121 1667 7130
rect 1725 7150 1863 7157
rect 1725 7130 1734 7150
rect 1754 7130 1863 7150
rect 1725 7121 1863 7130
rect 1519 7120 1556 7121
rect 1249 7067 1290 7068
rect 226 7062 644 7065
rect 226 7056 269 7062
rect 229 7053 269 7056
rect 1144 7060 1290 7067
rect 626 7044 666 7045
rect 337 7027 666 7044
rect 1144 7040 1200 7060
rect 1220 7040 1259 7060
rect 1279 7040 1290 7060
rect 1144 7032 1290 7040
rect 1357 7063 1514 7070
rect 1357 7043 1477 7063
rect 1497 7043 1514 7063
rect 1357 7033 1514 7043
rect 1357 7032 1392 7033
rect 221 6984 264 6995
rect 221 6966 233 6984
rect 251 6966 264 6984
rect 221 6940 264 6966
rect 337 6940 364 7027
rect 626 7018 666 7027
rect 221 6919 364 6940
rect 408 6992 442 7008
rect 626 6998 1019 7018
rect 1039 6998 1042 7018
rect 1357 7011 1388 7032
rect 1575 7011 1611 7121
rect 1630 7120 1667 7121
rect 1726 7120 1763 7121
rect 1686 7061 1776 7067
rect 1686 7041 1695 7061
rect 1715 7059 1776 7061
rect 1715 7041 1740 7059
rect 1686 7039 1740 7041
rect 1760 7039 1776 7059
rect 1686 7033 1776 7039
rect 1200 7010 1237 7011
rect 626 6993 1042 6998
rect 1199 7001 1237 7010
rect 626 6992 967 6993
rect 408 6922 445 6992
rect 560 6932 591 6933
rect 221 6917 358 6919
rect 221 6875 264 6917
rect 408 6902 417 6922
rect 437 6902 445 6922
rect 408 6892 445 6902
rect 504 6922 591 6932
rect 504 6902 513 6922
rect 533 6902 591 6922
rect 504 6893 591 6902
rect 504 6892 541 6893
rect 219 6865 264 6875
rect 219 6847 228 6865
rect 246 6847 264 6865
rect 219 6841 264 6847
rect 560 6842 591 6893
rect 626 6922 663 6992
rect 929 6991 966 6992
rect 1199 6981 1208 7001
rect 1228 6981 1237 7001
rect 1199 6973 1237 6981
rect 1303 7005 1388 7011
rect 1418 7010 1455 7011
rect 1303 6985 1311 7005
rect 1331 6985 1388 7005
rect 1303 6977 1388 6985
rect 1417 7001 1455 7010
rect 1417 6981 1426 7001
rect 1446 6981 1455 7001
rect 1303 6976 1339 6977
rect 1417 6973 1455 6981
rect 1521 7005 1665 7011
rect 1521 6985 1529 7005
rect 1549 7002 1637 7005
rect 1549 6985 1584 7002
rect 1521 6984 1584 6985
rect 1603 6985 1637 7002
rect 1657 6985 1665 7005
rect 1603 6984 1665 6985
rect 1521 6977 1665 6984
rect 1521 6976 1557 6977
rect 1629 6976 1665 6977
rect 1731 7010 1768 7011
rect 1731 7009 1769 7010
rect 1791 7009 1818 7013
rect 1731 7007 1818 7009
rect 1731 7001 1795 7007
rect 1731 6981 1740 7001
rect 1760 6987 1795 7001
rect 1815 6987 1818 7007
rect 1760 6982 1818 6987
rect 1760 6981 1795 6982
rect 1200 6944 1237 6973
rect 1201 6942 1237 6944
rect 778 6932 814 6933
rect 626 6902 635 6922
rect 655 6902 663 6922
rect 626 6892 663 6902
rect 722 6922 870 6932
rect 970 6929 1066 6931
rect 722 6902 731 6922
rect 751 6902 841 6922
rect 861 6902 870 6922
rect 722 6893 870 6902
rect 928 6922 1066 6929
rect 928 6902 937 6922
rect 957 6902 1066 6922
rect 1201 6920 1392 6942
rect 1418 6941 1455 6973
rect 1731 6969 1795 6981
rect 1835 6943 1862 7121
rect 1694 6941 1862 6943
rect 1418 6915 1862 6941
rect 928 6893 1066 6902
rect 722 6892 759 6893
rect 219 6838 256 6841
rect 452 6839 493 6840
rect 344 6832 493 6839
rect 344 6812 403 6832
rect 423 6812 462 6832
rect 482 6812 493 6832
rect 344 6804 493 6812
rect 560 6835 717 6842
rect 560 6815 680 6835
rect 700 6815 717 6835
rect 560 6805 717 6815
rect 560 6804 595 6805
rect 560 6783 591 6804
rect 778 6783 814 6893
rect 833 6892 870 6893
rect 929 6892 966 6893
rect 889 6833 979 6839
rect 889 6813 898 6833
rect 918 6831 979 6833
rect 918 6813 943 6831
rect 889 6811 943 6813
rect 963 6811 979 6831
rect 889 6805 979 6811
rect 403 6782 440 6783
rect 215 6774 253 6776
rect 215 6766 258 6774
rect 215 6748 226 6766
rect 244 6748 258 6766
rect 215 6721 258 6748
rect 402 6773 440 6782
rect 402 6753 411 6773
rect 431 6753 440 6773
rect 402 6745 440 6753
rect 506 6777 591 6783
rect 621 6782 658 6783
rect 506 6757 514 6777
rect 534 6757 591 6777
rect 506 6749 591 6757
rect 620 6773 658 6782
rect 620 6753 629 6773
rect 649 6753 658 6773
rect 506 6748 542 6749
rect 620 6745 658 6753
rect 724 6781 868 6783
rect 724 6777 776 6781
rect 724 6757 732 6777
rect 752 6761 776 6777
rect 796 6777 868 6781
rect 796 6761 840 6777
rect 752 6757 840 6761
rect 860 6757 868 6777
rect 724 6749 868 6757
rect 724 6748 760 6749
rect 832 6748 868 6749
rect 934 6782 971 6783
rect 934 6781 972 6782
rect 934 6773 998 6781
rect 934 6753 943 6773
rect 963 6759 998 6773
rect 1018 6759 1021 6779
rect 963 6754 1021 6759
rect 963 6753 998 6754
rect 216 6714 258 6721
rect 403 6714 440 6745
rect 621 6714 658 6745
rect 934 6741 998 6753
rect 1038 6715 1065 6893
rect 216 6674 261 6714
rect 403 6689 548 6714
rect 621 6713 701 6714
rect 897 6713 1065 6715
rect 621 6697 1065 6713
rect 405 6688 548 6689
rect 620 6687 1065 6697
rect 216 6653 263 6674
rect 620 6653 661 6687
rect 897 6686 1065 6687
rect 1528 6691 1568 6915
rect 1694 6914 1862 6915
rect 1926 6947 1959 7280
rect 2564 7279 2591 7457
rect 2631 7419 2695 7431
rect 2971 7427 3008 7459
rect 3034 7458 3225 7480
rect 3360 7478 3469 7498
rect 3489 7478 3498 7498
rect 3360 7471 3498 7478
rect 3556 7498 3704 7507
rect 3556 7478 3565 7498
rect 3585 7478 3675 7498
rect 3695 7478 3704 7498
rect 3360 7469 3456 7471
rect 3556 7468 3704 7478
rect 3763 7498 3800 7508
rect 3763 7478 3771 7498
rect 3791 7478 3800 7498
rect 3612 7467 3648 7468
rect 3189 7456 3225 7458
rect 3189 7427 3226 7456
rect 2631 7418 2666 7419
rect 2608 7413 2666 7418
rect 2608 7393 2611 7413
rect 2631 7399 2666 7413
rect 2686 7399 2695 7419
rect 2631 7391 2695 7399
rect 2657 7390 2695 7391
rect 2658 7389 2695 7390
rect 2761 7423 2797 7424
rect 2869 7423 2905 7424
rect 2761 7415 2905 7423
rect 2761 7395 2769 7415
rect 2789 7414 2877 7415
rect 2789 7395 2824 7414
rect 2845 7395 2877 7414
rect 2897 7395 2905 7415
rect 2761 7389 2905 7395
rect 2971 7419 3009 7427
rect 3087 7423 3123 7424
rect 2971 7399 2980 7419
rect 3000 7399 3009 7419
rect 2971 7390 3009 7399
rect 3038 7415 3123 7423
rect 3038 7395 3095 7415
rect 3115 7395 3123 7415
rect 2971 7389 3008 7390
rect 3038 7389 3123 7395
rect 3189 7419 3227 7427
rect 3189 7399 3198 7419
rect 3218 7399 3227 7419
rect 3460 7408 3497 7409
rect 3763 7408 3800 7478
rect 3835 7507 3866 7558
rect 4162 7553 4207 7559
rect 4162 7535 4180 7553
rect 4198 7535 4207 7553
rect 5668 7553 5677 7573
rect 5697 7553 5705 7573
rect 5668 7543 5705 7553
rect 5764 7573 5851 7583
rect 5764 7553 5773 7573
rect 5793 7553 5851 7573
rect 5764 7544 5851 7553
rect 5764 7543 5801 7544
rect 4162 7525 4207 7535
rect 3885 7507 3922 7508
rect 3835 7498 3922 7507
rect 3835 7478 3893 7498
rect 3913 7478 3922 7498
rect 3835 7468 3922 7478
rect 3981 7498 4018 7508
rect 3981 7478 3989 7498
rect 4009 7478 4018 7498
rect 4162 7483 4205 7525
rect 4589 7514 4641 7516
rect 4068 7481 4205 7483
rect 3835 7467 3866 7468
rect 3981 7408 4018 7478
rect 3459 7407 3800 7408
rect 3189 7390 3227 7399
rect 3384 7402 3800 7407
rect 3189 7389 3226 7390
rect 2650 7361 2740 7367
rect 2650 7341 2666 7361
rect 2686 7359 2740 7361
rect 2686 7341 2711 7359
rect 2650 7339 2711 7341
rect 2731 7339 2740 7359
rect 2650 7333 2740 7339
rect 2663 7279 2700 7280
rect 2759 7279 2796 7280
rect 2815 7279 2851 7389
rect 3038 7368 3069 7389
rect 3384 7382 3387 7402
rect 3407 7382 3800 7402
rect 3984 7392 4018 7408
rect 4062 7460 4205 7481
rect 4587 7510 5020 7514
rect 4587 7504 5026 7510
rect 4587 7486 4608 7504
rect 4626 7486 5026 7504
rect 5820 7493 5851 7544
rect 5886 7573 5923 7643
rect 6189 7642 6226 7643
rect 6038 7583 6074 7584
rect 5886 7553 5895 7573
rect 5915 7553 5923 7573
rect 5886 7543 5923 7553
rect 5982 7573 6130 7583
rect 6230 7580 6326 7582
rect 5982 7553 5991 7573
rect 6011 7553 6101 7573
rect 6121 7553 6130 7573
rect 5982 7544 6130 7553
rect 6188 7573 6326 7580
rect 6188 7553 6197 7573
rect 6217 7553 6326 7573
rect 6188 7544 6326 7553
rect 5982 7543 6019 7544
rect 5712 7490 5753 7491
rect 4587 7468 5026 7486
rect 3760 7373 3800 7382
rect 4062 7373 4089 7460
rect 4162 7434 4205 7460
rect 4162 7416 4175 7434
rect 4193 7416 4205 7434
rect 4162 7405 4205 7416
rect 3034 7367 3069 7368
rect 2912 7357 3069 7367
rect 2912 7337 2929 7357
rect 2949 7337 3069 7357
rect 2912 7330 3069 7337
rect 3136 7360 3285 7368
rect 3136 7340 3147 7360
rect 3167 7340 3206 7360
rect 3226 7340 3285 7360
rect 3760 7356 4089 7373
rect 3760 7355 3800 7356
rect 3136 7333 3285 7340
rect 4157 7344 4197 7347
rect 4157 7338 4200 7344
rect 3782 7335 4200 7338
rect 3136 7332 3177 7333
rect 2870 7279 2907 7280
rect 2563 7270 2701 7279
rect 2426 7260 2462 7266
rect 2426 7242 2431 7260
rect 2453 7242 2462 7260
rect 2426 7238 2462 7242
rect 2563 7250 2672 7270
rect 2692 7250 2701 7270
rect 2563 7243 2701 7250
rect 2759 7270 2907 7279
rect 2759 7250 2768 7270
rect 2788 7250 2878 7270
rect 2898 7250 2907 7270
rect 2563 7241 2659 7243
rect 2759 7240 2907 7250
rect 2966 7270 3003 7280
rect 2966 7250 2974 7270
rect 2994 7250 3003 7270
rect 2815 7239 2851 7240
rect 2429 7079 2462 7238
rect 2663 7180 2700 7181
rect 2966 7180 3003 7250
rect 3038 7279 3069 7330
rect 3782 7317 4173 7335
rect 4191 7317 4200 7335
rect 3782 7315 4200 7317
rect 3782 7307 3809 7315
rect 4050 7312 4200 7315
rect 3362 7301 3530 7302
rect 3781 7301 3809 7307
rect 3362 7285 3809 7301
rect 4157 7307 4200 7312
rect 3088 7279 3125 7280
rect 3038 7270 3125 7279
rect 3038 7250 3096 7270
rect 3116 7250 3125 7270
rect 3038 7240 3125 7250
rect 3184 7270 3221 7280
rect 3184 7250 3192 7270
rect 3212 7250 3221 7270
rect 3038 7239 3069 7240
rect 2662 7179 3003 7180
rect 3184 7179 3221 7250
rect 2587 7174 3003 7179
rect 2587 7154 2590 7174
rect 2610 7154 3003 7174
rect 3034 7155 3221 7179
rect 3362 7275 3806 7285
rect 3362 7273 3530 7275
rect 3362 7095 3389 7273
rect 3429 7235 3493 7247
rect 3769 7243 3806 7275
rect 3832 7274 4023 7296
rect 3987 7272 4023 7274
rect 3987 7243 4024 7272
rect 4157 7251 4197 7307
rect 3429 7234 3464 7235
rect 3406 7229 3464 7234
rect 3406 7209 3409 7229
rect 3429 7215 3464 7229
rect 3484 7215 3493 7235
rect 3429 7207 3493 7215
rect 3455 7206 3493 7207
rect 3456 7205 3493 7206
rect 3559 7239 3595 7240
rect 3667 7239 3703 7240
rect 3559 7231 3703 7239
rect 3559 7211 3567 7231
rect 3587 7211 3622 7231
rect 3642 7211 3675 7231
rect 3695 7211 3703 7231
rect 3559 7205 3703 7211
rect 3769 7235 3807 7243
rect 3885 7239 3921 7240
rect 3769 7215 3778 7235
rect 3798 7215 3807 7235
rect 3769 7206 3807 7215
rect 3836 7231 3921 7239
rect 3836 7211 3893 7231
rect 3913 7211 3921 7231
rect 3769 7205 3806 7206
rect 3836 7205 3921 7211
rect 3987 7235 4025 7243
rect 3987 7215 3996 7235
rect 4016 7215 4025 7235
rect 4157 7233 4169 7251
rect 4187 7233 4197 7251
rect 4589 7279 4641 7468
rect 4987 7443 5026 7468
rect 5604 7483 5753 7490
rect 5604 7463 5663 7483
rect 5683 7463 5722 7483
rect 5742 7463 5753 7483
rect 5604 7455 5753 7463
rect 5820 7486 5977 7493
rect 5820 7466 5940 7486
rect 5960 7466 5977 7486
rect 5820 7456 5977 7466
rect 5820 7455 5855 7456
rect 4771 7418 4958 7442
rect 4987 7423 5382 7443
rect 5402 7423 5405 7443
rect 5820 7434 5851 7455
rect 6038 7434 6074 7544
rect 6093 7543 6130 7544
rect 6189 7543 6226 7544
rect 6149 7484 6239 7490
rect 6149 7464 6158 7484
rect 6178 7482 6239 7484
rect 6178 7464 6203 7482
rect 6149 7462 6203 7464
rect 6223 7462 6239 7482
rect 6149 7456 6239 7462
rect 5663 7433 5700 7434
rect 4987 7418 5405 7423
rect 5662 7424 5700 7433
rect 4771 7347 4808 7418
rect 4987 7417 5330 7418
rect 4987 7414 5026 7417
rect 5292 7416 5329 7417
rect 4923 7357 4954 7358
rect 4771 7327 4780 7347
rect 4800 7327 4808 7347
rect 4771 7317 4808 7327
rect 4867 7347 4954 7357
rect 4867 7327 4876 7347
rect 4896 7327 4954 7347
rect 4867 7318 4954 7327
rect 4867 7317 4904 7318
rect 4589 7261 4605 7279
rect 4623 7261 4641 7279
rect 4923 7267 4954 7318
rect 4989 7347 5026 7414
rect 5662 7404 5671 7424
rect 5691 7404 5700 7424
rect 5662 7396 5700 7404
rect 5766 7428 5851 7434
rect 5881 7433 5918 7434
rect 5766 7408 5774 7428
rect 5794 7408 5851 7428
rect 5766 7400 5851 7408
rect 5880 7424 5918 7433
rect 5880 7404 5889 7424
rect 5909 7404 5918 7424
rect 5766 7399 5802 7400
rect 5880 7396 5918 7404
rect 5984 7429 6128 7434
rect 5984 7428 6046 7429
rect 5984 7408 5992 7428
rect 6012 7410 6046 7428
rect 6067 7428 6128 7429
rect 6067 7410 6100 7428
rect 6012 7408 6100 7410
rect 6120 7408 6128 7428
rect 5984 7400 6128 7408
rect 5984 7399 6020 7400
rect 6092 7399 6128 7400
rect 6194 7433 6231 7434
rect 6194 7432 6232 7433
rect 6194 7424 6258 7432
rect 6194 7404 6203 7424
rect 6223 7410 6258 7424
rect 6278 7410 6281 7430
rect 6223 7405 6281 7410
rect 6223 7404 6258 7405
rect 5663 7367 5700 7396
rect 5664 7365 5700 7367
rect 5141 7357 5177 7358
rect 4989 7327 4998 7347
rect 5018 7327 5026 7347
rect 4989 7317 5026 7327
rect 5085 7347 5233 7357
rect 5333 7354 5429 7356
rect 5085 7327 5094 7347
rect 5114 7327 5204 7347
rect 5224 7327 5233 7347
rect 5085 7318 5233 7327
rect 5291 7347 5429 7354
rect 5291 7327 5300 7347
rect 5320 7327 5429 7347
rect 5664 7343 5855 7365
rect 5881 7364 5918 7396
rect 6194 7392 6258 7404
rect 6298 7366 6325 7544
rect 6157 7364 6325 7366
rect 5881 7350 6325 7364
rect 6928 7498 7096 7499
rect 7222 7498 7262 7722
rect 7725 7726 7893 7727
rect 8128 7726 8168 7759
rect 8524 7726 8571 7759
rect 7725 7725 8169 7726
rect 7725 7700 8170 7725
rect 7725 7698 7893 7700
rect 8089 7699 8170 7700
rect 8339 7699 8388 7725
rect 8524 7699 8573 7726
rect 7725 7520 7752 7698
rect 7792 7660 7856 7672
rect 8132 7668 8169 7699
rect 8350 7668 8387 7699
rect 8532 7674 8573 7699
rect 7792 7659 7827 7660
rect 7769 7654 7827 7659
rect 7769 7634 7772 7654
rect 7792 7640 7827 7654
rect 7847 7640 7856 7660
rect 7792 7632 7856 7640
rect 7818 7631 7856 7632
rect 7819 7630 7856 7631
rect 7922 7664 7958 7665
rect 8030 7664 8066 7665
rect 7922 7656 8066 7664
rect 7922 7636 7930 7656
rect 7950 7652 8038 7656
rect 7950 7636 7994 7652
rect 7922 7632 7994 7636
rect 8014 7636 8038 7652
rect 8058 7636 8066 7656
rect 8014 7632 8066 7636
rect 7922 7630 8066 7632
rect 8132 7660 8170 7668
rect 8248 7664 8284 7665
rect 8132 7640 8141 7660
rect 8161 7640 8170 7660
rect 8132 7631 8170 7640
rect 8199 7656 8284 7664
rect 8199 7636 8256 7656
rect 8276 7636 8284 7656
rect 8132 7630 8169 7631
rect 8199 7630 8284 7636
rect 8350 7660 8388 7668
rect 8350 7640 8359 7660
rect 8379 7640 8388 7660
rect 8350 7631 8388 7640
rect 8532 7665 8574 7674
rect 8532 7647 8546 7665
rect 8564 7647 8574 7665
rect 8532 7639 8574 7647
rect 8537 7637 8574 7639
rect 8350 7630 8387 7631
rect 7811 7602 7901 7608
rect 7811 7582 7827 7602
rect 7847 7600 7901 7602
rect 7847 7582 7872 7600
rect 7811 7580 7872 7582
rect 7892 7580 7901 7600
rect 7811 7574 7901 7580
rect 7824 7520 7861 7521
rect 7920 7520 7957 7521
rect 7976 7520 8012 7630
rect 8199 7609 8230 7630
rect 8195 7608 8230 7609
rect 8073 7598 8230 7608
rect 8073 7578 8090 7598
rect 8110 7578 8230 7598
rect 8073 7571 8230 7578
rect 8297 7601 8446 7609
rect 8297 7581 8308 7601
rect 8328 7581 8367 7601
rect 8387 7581 8446 7601
rect 8297 7574 8446 7581
rect 8297 7573 8338 7574
rect 8534 7572 8571 7575
rect 8031 7520 8068 7521
rect 7724 7511 7862 7520
rect 6928 7472 7372 7498
rect 6928 7470 7096 7472
rect 5881 7338 6328 7350
rect 5924 7336 5957 7338
rect 5291 7318 5429 7327
rect 5085 7317 5122 7318
rect 4815 7264 4856 7265
rect 4589 7243 4641 7261
rect 4707 7257 4856 7264
rect 4157 7223 4197 7233
rect 4707 7237 4766 7257
rect 4786 7237 4825 7257
rect 4845 7237 4856 7257
rect 4707 7229 4856 7237
rect 4923 7260 5080 7267
rect 4923 7240 5043 7260
rect 5063 7240 5080 7260
rect 4923 7230 5080 7240
rect 4923 7229 4958 7230
rect 3987 7206 4025 7215
rect 4923 7208 4954 7229
rect 5141 7208 5177 7318
rect 5196 7317 5233 7318
rect 5292 7317 5329 7318
rect 5252 7258 5342 7264
rect 5252 7238 5261 7258
rect 5281 7256 5342 7258
rect 5281 7238 5306 7256
rect 5252 7236 5306 7238
rect 5326 7236 5342 7256
rect 5252 7230 5342 7236
rect 4766 7207 4803 7208
rect 3987 7205 4024 7206
rect 3448 7177 3538 7183
rect 3448 7157 3464 7177
rect 3484 7175 3538 7177
rect 3484 7157 3509 7175
rect 3448 7155 3509 7157
rect 3529 7155 3538 7175
rect 3448 7149 3538 7155
rect 3461 7095 3498 7096
rect 3557 7095 3594 7096
rect 3613 7095 3649 7205
rect 3836 7184 3867 7205
rect 4765 7198 4803 7207
rect 3832 7183 3867 7184
rect 3710 7173 3867 7183
rect 3710 7153 3727 7173
rect 3747 7153 3867 7173
rect 3710 7146 3867 7153
rect 3934 7176 4083 7184
rect 3934 7156 3945 7176
rect 3965 7156 4004 7176
rect 4024 7156 4083 7176
rect 4593 7180 4633 7190
rect 3934 7149 4083 7156
rect 4149 7152 4201 7170
rect 3934 7148 3975 7149
rect 3668 7095 3705 7096
rect 3361 7086 3499 7095
rect 2428 7078 2465 7079
rect 2399 7077 2567 7078
rect 2693 7077 2733 7079
rect 2224 7068 2263 7074
rect 2224 7046 2232 7068
rect 2256 7046 2263 7068
rect 1926 6939 1963 6947
rect 1926 6920 1934 6939
rect 1955 6920 1963 6939
rect 1926 6914 1963 6920
rect 1528 6669 1536 6691
rect 1560 6669 1568 6691
rect 1528 6661 1568 6669
rect 216 6623 661 6653
rect 1699 6636 1764 6637
rect 216 6620 639 6623
rect 216 6572 263 6620
rect 216 6554 226 6572
rect 244 6554 263 6572
rect 216 6550 263 6554
rect 1350 6611 1537 6635
rect 1568 6616 1961 6636
rect 1981 6616 1984 6636
rect 1568 6611 1984 6616
rect 217 6545 254 6550
rect 1350 6540 1387 6611
rect 1568 6610 1909 6611
rect 1502 6550 1533 6551
rect 1350 6520 1359 6540
rect 1379 6520 1387 6540
rect 1350 6510 1387 6520
rect 1446 6540 1533 6550
rect 1446 6520 1455 6540
rect 1475 6520 1533 6540
rect 1446 6511 1533 6520
rect 1446 6510 1483 6511
rect 205 6483 257 6485
rect 203 6479 636 6483
rect 203 6473 642 6479
rect 203 6455 224 6473
rect 242 6455 642 6473
rect 1502 6460 1533 6511
rect 1568 6540 1605 6610
rect 1871 6609 1908 6610
rect 1720 6550 1756 6551
rect 1568 6520 1577 6540
rect 1597 6520 1605 6540
rect 1568 6510 1605 6520
rect 1664 6540 1812 6550
rect 1912 6547 2008 6549
rect 1664 6520 1673 6540
rect 1693 6520 1783 6540
rect 1803 6520 1812 6540
rect 1664 6511 1812 6520
rect 1870 6540 2008 6547
rect 1870 6520 1879 6540
rect 1899 6520 2008 6540
rect 1870 6511 2008 6520
rect 1664 6510 1701 6511
rect 1394 6457 1435 6458
rect 203 6437 642 6455
rect 205 6248 257 6437
rect 603 6412 642 6437
rect 1286 6450 1435 6457
rect 1286 6430 1345 6450
rect 1365 6430 1404 6450
rect 1424 6430 1435 6450
rect 1286 6422 1435 6430
rect 1502 6453 1659 6460
rect 1502 6433 1622 6453
rect 1642 6433 1659 6453
rect 1502 6423 1659 6433
rect 1502 6422 1537 6423
rect 387 6387 574 6411
rect 603 6392 998 6412
rect 1018 6392 1021 6412
rect 1502 6401 1533 6422
rect 1720 6401 1756 6511
rect 1775 6510 1812 6511
rect 1871 6510 1908 6511
rect 1831 6451 1921 6457
rect 1831 6431 1840 6451
rect 1860 6449 1921 6451
rect 1860 6431 1885 6449
rect 1831 6429 1885 6431
rect 1905 6429 1921 6449
rect 1831 6423 1921 6429
rect 1345 6400 1382 6401
rect 603 6387 1021 6392
rect 1344 6391 1382 6400
rect 387 6316 424 6387
rect 603 6386 946 6387
rect 603 6383 642 6386
rect 908 6385 945 6386
rect 539 6326 570 6327
rect 387 6296 396 6316
rect 416 6296 424 6316
rect 387 6286 424 6296
rect 483 6316 570 6326
rect 483 6296 492 6316
rect 512 6296 570 6316
rect 483 6287 570 6296
rect 483 6286 520 6287
rect 205 6230 221 6248
rect 239 6230 257 6248
rect 539 6236 570 6287
rect 605 6316 642 6383
rect 1344 6371 1353 6391
rect 1373 6371 1382 6391
rect 1344 6363 1382 6371
rect 1448 6395 1533 6401
rect 1563 6400 1600 6401
rect 1448 6375 1456 6395
rect 1476 6375 1533 6395
rect 1448 6367 1533 6375
rect 1562 6391 1600 6400
rect 1562 6371 1571 6391
rect 1591 6371 1600 6391
rect 1448 6366 1484 6367
rect 1562 6363 1600 6371
rect 1666 6395 1810 6401
rect 1666 6375 1674 6395
rect 1694 6394 1782 6395
rect 1694 6376 1729 6394
rect 1747 6376 1782 6394
rect 1694 6375 1782 6376
rect 1802 6375 1810 6395
rect 1666 6367 1810 6375
rect 1666 6366 1702 6367
rect 1774 6366 1810 6367
rect 1876 6400 1913 6401
rect 1876 6399 1914 6400
rect 1876 6391 1940 6399
rect 1876 6371 1885 6391
rect 1905 6377 1940 6391
rect 1960 6377 1963 6397
rect 1905 6372 1963 6377
rect 1905 6371 1940 6372
rect 1345 6334 1382 6363
rect 1346 6332 1382 6334
rect 757 6326 793 6327
rect 605 6296 614 6316
rect 634 6296 642 6316
rect 605 6286 642 6296
rect 701 6316 849 6326
rect 949 6323 1045 6325
rect 701 6296 710 6316
rect 730 6296 820 6316
rect 840 6296 849 6316
rect 701 6287 849 6296
rect 907 6316 1045 6323
rect 907 6296 916 6316
rect 936 6296 1045 6316
rect 1346 6310 1537 6332
rect 1563 6331 1600 6363
rect 1876 6359 1940 6371
rect 1980 6335 2007 6511
rect 1926 6333 2007 6335
rect 1839 6331 2007 6333
rect 1563 6305 2007 6331
rect 1673 6303 1713 6305
rect 1839 6304 2007 6305
rect 907 6287 1045 6296
rect 1948 6302 2007 6304
rect 701 6286 738 6287
rect 431 6233 472 6234
rect 205 6212 257 6230
rect 323 6226 472 6233
rect 323 6206 382 6226
rect 402 6206 441 6226
rect 461 6206 472 6226
rect 323 6198 472 6206
rect 539 6229 696 6236
rect 539 6209 659 6229
rect 679 6209 696 6229
rect 539 6199 696 6209
rect 539 6198 574 6199
rect 539 6177 570 6198
rect 757 6177 793 6287
rect 812 6286 849 6287
rect 908 6286 945 6287
rect 868 6227 958 6233
rect 868 6207 877 6227
rect 897 6225 958 6227
rect 897 6207 922 6225
rect 868 6205 922 6207
rect 942 6205 958 6225
rect 868 6199 958 6205
rect 382 6176 419 6177
rect 381 6167 419 6176
rect 209 6149 249 6159
rect 209 6131 219 6149
rect 237 6131 249 6149
rect 381 6147 390 6167
rect 410 6147 419 6167
rect 381 6139 419 6147
rect 485 6171 570 6177
rect 600 6176 637 6177
rect 485 6151 493 6171
rect 513 6151 570 6171
rect 485 6143 570 6151
rect 599 6167 637 6176
rect 599 6147 608 6167
rect 628 6147 637 6167
rect 485 6142 521 6143
rect 599 6139 637 6147
rect 703 6171 847 6177
rect 703 6151 711 6171
rect 731 6151 764 6171
rect 784 6151 819 6171
rect 839 6151 847 6171
rect 703 6143 847 6151
rect 703 6142 739 6143
rect 811 6142 847 6143
rect 913 6176 950 6177
rect 913 6175 951 6176
rect 913 6167 977 6175
rect 913 6147 922 6167
rect 942 6153 977 6167
rect 997 6153 1000 6173
rect 942 6148 1000 6153
rect 942 6147 977 6148
rect 209 6075 249 6131
rect 382 6110 419 6139
rect 383 6108 419 6110
rect 383 6086 574 6108
rect 600 6107 637 6139
rect 913 6135 977 6147
rect 1017 6109 1044 6287
rect 1948 6284 1977 6302
rect 876 6107 1044 6109
rect 600 6097 1044 6107
rect 1185 6203 1372 6227
rect 1403 6208 1796 6228
rect 1816 6208 1819 6228
rect 1403 6203 1819 6208
rect 1185 6132 1222 6203
rect 1403 6202 1744 6203
rect 1337 6142 1368 6143
rect 1185 6112 1194 6132
rect 1214 6112 1222 6132
rect 1185 6102 1222 6112
rect 1281 6132 1368 6142
rect 1281 6112 1290 6132
rect 1310 6112 1368 6132
rect 1281 6103 1368 6112
rect 1281 6102 1318 6103
rect 206 6070 249 6075
rect 597 6081 1044 6097
rect 597 6075 625 6081
rect 876 6080 1044 6081
rect 206 6067 356 6070
rect 597 6067 624 6075
rect 206 6065 624 6067
rect 206 6047 215 6065
rect 233 6047 624 6065
rect 1337 6052 1368 6103
rect 1403 6132 1440 6202
rect 1706 6201 1743 6202
rect 1555 6142 1591 6143
rect 1403 6112 1412 6132
rect 1432 6112 1440 6132
rect 1403 6102 1440 6112
rect 1499 6132 1647 6142
rect 1747 6139 1843 6141
rect 1499 6112 1508 6132
rect 1528 6112 1618 6132
rect 1638 6112 1647 6132
rect 1499 6103 1647 6112
rect 1705 6132 1843 6139
rect 1705 6112 1714 6132
rect 1734 6112 1843 6132
rect 1705 6103 1843 6112
rect 1499 6102 1536 6103
rect 1229 6049 1270 6050
rect 206 6044 624 6047
rect 206 6038 249 6044
rect 209 6035 249 6038
rect 1121 6042 1270 6049
rect 606 6026 646 6027
rect 317 6009 646 6026
rect 1121 6022 1180 6042
rect 1200 6022 1239 6042
rect 1259 6022 1270 6042
rect 1121 6014 1270 6022
rect 1337 6045 1494 6052
rect 1337 6025 1457 6045
rect 1477 6025 1494 6045
rect 1337 6015 1494 6025
rect 1337 6014 1372 6015
rect 201 5966 244 5977
rect 201 5948 213 5966
rect 231 5948 244 5966
rect 201 5922 244 5948
rect 317 5922 344 6009
rect 606 6000 646 6009
rect 201 5901 344 5922
rect 388 5974 422 5990
rect 606 5980 999 6000
rect 1019 5980 1022 6000
rect 1337 5993 1368 6014
rect 1555 5993 1591 6103
rect 1610 6102 1647 6103
rect 1706 6102 1743 6103
rect 1666 6043 1756 6049
rect 1666 6023 1675 6043
rect 1695 6041 1756 6043
rect 1695 6023 1720 6041
rect 1666 6021 1720 6023
rect 1740 6021 1756 6041
rect 1666 6015 1756 6021
rect 1180 5992 1217 5993
rect 606 5975 1022 5980
rect 1179 5983 1217 5992
rect 606 5974 947 5975
rect 388 5904 425 5974
rect 540 5914 571 5915
rect 201 5899 338 5901
rect 201 5857 244 5899
rect 388 5884 397 5904
rect 417 5884 425 5904
rect 388 5874 425 5884
rect 484 5904 571 5914
rect 484 5884 493 5904
rect 513 5884 571 5904
rect 484 5875 571 5884
rect 484 5874 521 5875
rect 199 5847 244 5857
rect 199 5829 208 5847
rect 226 5829 244 5847
rect 199 5823 244 5829
rect 540 5824 571 5875
rect 606 5904 643 5974
rect 909 5973 946 5974
rect 1179 5963 1188 5983
rect 1208 5963 1217 5983
rect 1179 5955 1217 5963
rect 1283 5987 1368 5993
rect 1398 5992 1435 5993
rect 1283 5967 1291 5987
rect 1311 5967 1368 5987
rect 1283 5959 1368 5967
rect 1397 5983 1435 5992
rect 1397 5963 1406 5983
rect 1426 5963 1435 5983
rect 1283 5958 1319 5959
rect 1397 5955 1435 5963
rect 1501 5987 1645 5993
rect 1501 5967 1509 5987
rect 1529 5968 1561 5987
rect 1582 5968 1617 5987
rect 1529 5967 1617 5968
rect 1637 5967 1645 5987
rect 1501 5959 1645 5967
rect 1501 5958 1537 5959
rect 1609 5958 1645 5959
rect 1711 5992 1748 5993
rect 1711 5991 1749 5992
rect 1711 5983 1775 5991
rect 1711 5963 1720 5983
rect 1740 5969 1775 5983
rect 1795 5969 1798 5989
rect 1740 5964 1798 5969
rect 1740 5963 1775 5964
rect 1180 5926 1217 5955
rect 1181 5924 1217 5926
rect 758 5914 794 5915
rect 606 5884 615 5904
rect 635 5884 643 5904
rect 606 5874 643 5884
rect 702 5904 850 5914
rect 950 5911 1046 5913
rect 702 5884 711 5904
rect 731 5884 821 5904
rect 841 5884 850 5904
rect 702 5875 850 5884
rect 908 5904 1046 5911
rect 908 5884 917 5904
rect 937 5884 1046 5904
rect 1181 5902 1372 5924
rect 1398 5923 1435 5955
rect 1711 5951 1775 5963
rect 1815 5925 1842 6103
rect 1674 5923 1842 5925
rect 1398 5897 1842 5923
rect 908 5875 1046 5884
rect 702 5874 739 5875
rect 199 5820 236 5823
rect 432 5821 473 5822
rect 324 5814 473 5821
rect 324 5794 383 5814
rect 403 5794 442 5814
rect 462 5794 473 5814
rect 324 5786 473 5794
rect 540 5817 697 5824
rect 540 5797 660 5817
rect 680 5797 697 5817
rect 540 5787 697 5797
rect 540 5786 575 5787
rect 540 5765 571 5786
rect 758 5765 794 5875
rect 813 5874 850 5875
rect 909 5874 946 5875
rect 869 5815 959 5821
rect 869 5795 878 5815
rect 898 5813 959 5815
rect 898 5795 923 5813
rect 869 5793 923 5795
rect 943 5793 959 5813
rect 869 5787 959 5793
rect 383 5764 420 5765
rect 196 5756 233 5758
rect 196 5748 238 5756
rect 196 5730 206 5748
rect 224 5730 238 5748
rect 196 5721 238 5730
rect 382 5755 420 5764
rect 382 5735 391 5755
rect 411 5735 420 5755
rect 382 5727 420 5735
rect 486 5759 571 5765
rect 601 5764 638 5765
rect 486 5739 494 5759
rect 514 5739 571 5759
rect 486 5731 571 5739
rect 600 5755 638 5764
rect 600 5735 609 5755
rect 629 5735 638 5755
rect 486 5730 522 5731
rect 600 5727 638 5735
rect 704 5763 848 5765
rect 704 5759 756 5763
rect 704 5739 712 5759
rect 732 5743 756 5759
rect 776 5759 848 5763
rect 776 5743 820 5759
rect 732 5739 820 5743
rect 840 5739 848 5759
rect 704 5731 848 5739
rect 704 5730 740 5731
rect 812 5730 848 5731
rect 914 5764 951 5765
rect 914 5763 952 5764
rect 914 5755 978 5763
rect 914 5735 923 5755
rect 943 5741 978 5755
rect 998 5741 1001 5761
rect 943 5736 1001 5741
rect 943 5735 978 5736
rect 197 5696 238 5721
rect 383 5696 420 5727
rect 601 5696 638 5727
rect 914 5723 978 5735
rect 1018 5697 1045 5875
rect 197 5669 246 5696
rect 382 5670 431 5696
rect 600 5695 681 5696
rect 877 5695 1045 5697
rect 600 5670 1045 5695
rect 601 5669 1045 5670
rect 199 5636 246 5669
rect 602 5636 642 5669
rect 877 5668 1045 5669
rect 1508 5673 1548 5897
rect 1674 5896 1842 5897
rect 1508 5651 1516 5673
rect 1540 5651 1548 5673
rect 1508 5643 1548 5651
rect 199 5597 642 5636
rect 199 5554 246 5597
rect 602 5592 642 5597
rect 1267 5595 1454 5619
rect 1485 5600 1878 5620
rect 1898 5600 1901 5620
rect 1485 5595 1901 5600
rect 199 5536 209 5554
rect 227 5536 246 5554
rect 199 5532 246 5536
rect 200 5527 237 5532
rect 1267 5524 1304 5595
rect 1485 5594 1826 5595
rect 1419 5534 1450 5535
rect 1267 5504 1276 5524
rect 1296 5504 1304 5524
rect 1267 5494 1304 5504
rect 1363 5524 1450 5534
rect 1363 5504 1372 5524
rect 1392 5504 1450 5524
rect 1363 5495 1450 5504
rect 1363 5494 1400 5495
rect 188 5465 240 5467
rect 186 5461 619 5465
rect 186 5455 625 5461
rect 186 5437 207 5455
rect 225 5437 625 5455
rect 1419 5444 1450 5495
rect 1485 5524 1522 5594
rect 1788 5593 1825 5594
rect 1637 5534 1673 5535
rect 1485 5504 1494 5524
rect 1514 5504 1522 5524
rect 1485 5494 1522 5504
rect 1581 5524 1729 5534
rect 1829 5531 1925 5533
rect 1581 5504 1590 5524
rect 1610 5504 1700 5524
rect 1720 5504 1729 5524
rect 1581 5495 1729 5504
rect 1787 5524 1925 5531
rect 1787 5504 1796 5524
rect 1816 5504 1925 5524
rect 1787 5495 1925 5504
rect 1581 5494 1618 5495
rect 1311 5441 1352 5442
rect 186 5419 625 5437
rect 188 5230 240 5419
rect 586 5394 625 5419
rect 1203 5434 1352 5441
rect 1203 5414 1262 5434
rect 1282 5414 1321 5434
rect 1341 5414 1352 5434
rect 1203 5406 1352 5414
rect 1419 5437 1576 5444
rect 1419 5417 1539 5437
rect 1559 5417 1576 5437
rect 1419 5407 1576 5417
rect 1419 5406 1454 5407
rect 370 5369 557 5393
rect 586 5374 981 5394
rect 1001 5374 1004 5394
rect 1419 5385 1450 5406
rect 1637 5385 1673 5495
rect 1692 5494 1729 5495
rect 1788 5494 1825 5495
rect 1748 5435 1838 5441
rect 1748 5415 1757 5435
rect 1777 5433 1838 5435
rect 1777 5415 1802 5433
rect 1748 5413 1802 5415
rect 1822 5413 1838 5433
rect 1748 5407 1838 5413
rect 1262 5384 1299 5385
rect 586 5369 1004 5374
rect 1261 5375 1299 5384
rect 370 5298 407 5369
rect 586 5368 929 5369
rect 586 5365 625 5368
rect 891 5367 928 5368
rect 522 5308 553 5309
rect 370 5278 379 5298
rect 399 5278 407 5298
rect 370 5268 407 5278
rect 466 5298 553 5308
rect 466 5278 475 5298
rect 495 5278 553 5298
rect 466 5269 553 5278
rect 466 5268 503 5269
rect 188 5212 204 5230
rect 222 5212 240 5230
rect 522 5218 553 5269
rect 588 5298 625 5365
rect 1261 5355 1270 5375
rect 1290 5355 1299 5375
rect 1261 5347 1299 5355
rect 1365 5379 1450 5385
rect 1480 5384 1517 5385
rect 1365 5359 1373 5379
rect 1393 5359 1450 5379
rect 1365 5351 1450 5359
rect 1479 5375 1517 5384
rect 1479 5355 1488 5375
rect 1508 5355 1517 5375
rect 1365 5350 1401 5351
rect 1479 5347 1517 5355
rect 1583 5379 1727 5385
rect 1583 5359 1591 5379
rect 1611 5374 1699 5379
rect 1611 5359 1647 5374
rect 1583 5357 1647 5359
rect 1666 5359 1699 5374
rect 1719 5359 1727 5379
rect 1666 5357 1727 5359
rect 1583 5351 1727 5357
rect 1583 5350 1619 5351
rect 1691 5350 1727 5351
rect 1793 5384 1830 5385
rect 1793 5383 1831 5384
rect 1793 5375 1857 5383
rect 1793 5355 1802 5375
rect 1822 5361 1857 5375
rect 1877 5361 1880 5381
rect 1822 5356 1880 5361
rect 1822 5355 1857 5356
rect 1262 5318 1299 5347
rect 1263 5316 1299 5318
rect 740 5308 776 5309
rect 588 5278 597 5298
rect 617 5278 625 5298
rect 588 5268 625 5278
rect 684 5298 832 5308
rect 932 5305 1028 5307
rect 684 5278 693 5298
rect 713 5278 803 5298
rect 823 5278 832 5298
rect 684 5269 832 5278
rect 890 5298 1028 5305
rect 890 5278 899 5298
rect 919 5278 1028 5298
rect 1263 5294 1454 5316
rect 1480 5315 1517 5347
rect 1793 5343 1857 5355
rect 1897 5317 1924 5495
rect 1756 5315 1924 5317
rect 1480 5301 1924 5315
rect 1948 5338 1976 6284
rect 1948 5308 1993 5338
rect 1480 5289 1927 5301
rect 1523 5287 1556 5289
rect 890 5269 1028 5278
rect 684 5268 721 5269
rect 414 5215 455 5216
rect 188 5194 240 5212
rect 306 5208 455 5215
rect 306 5188 365 5208
rect 385 5188 424 5208
rect 444 5188 455 5208
rect 306 5180 455 5188
rect 522 5211 679 5218
rect 522 5191 642 5211
rect 662 5191 679 5211
rect 522 5181 679 5191
rect 522 5180 557 5181
rect 522 5159 553 5180
rect 740 5159 776 5269
rect 795 5268 832 5269
rect 891 5268 928 5269
rect 851 5209 941 5215
rect 851 5189 860 5209
rect 880 5207 941 5209
rect 880 5189 905 5207
rect 851 5187 905 5189
rect 925 5187 941 5207
rect 851 5181 941 5187
rect 365 5158 402 5159
rect 364 5149 402 5158
rect 192 5131 232 5141
rect 192 5113 202 5131
rect 220 5113 232 5131
rect 364 5129 373 5149
rect 393 5129 402 5149
rect 364 5121 402 5129
rect 468 5153 553 5159
rect 583 5158 620 5159
rect 468 5133 476 5153
rect 496 5133 553 5153
rect 468 5125 553 5133
rect 582 5149 620 5158
rect 582 5129 591 5149
rect 611 5129 620 5149
rect 468 5124 504 5125
rect 582 5121 620 5129
rect 686 5153 830 5159
rect 686 5133 694 5153
rect 714 5133 747 5153
rect 767 5133 802 5153
rect 822 5133 830 5153
rect 686 5125 830 5133
rect 686 5124 722 5125
rect 794 5124 830 5125
rect 896 5158 933 5159
rect 896 5157 934 5158
rect 896 5149 960 5157
rect 896 5129 905 5149
rect 925 5135 960 5149
rect 980 5135 983 5155
rect 925 5130 983 5135
rect 925 5129 960 5130
rect 192 5057 232 5113
rect 365 5092 402 5121
rect 366 5090 402 5092
rect 366 5068 557 5090
rect 583 5089 620 5121
rect 896 5117 960 5129
rect 1000 5091 1027 5269
rect 1885 5244 1927 5289
rect 1948 5290 1959 5308
rect 1981 5290 1993 5308
rect 1948 5284 1993 5290
rect 1949 5283 1993 5284
rect 859 5089 1027 5091
rect 583 5079 1027 5089
rect 1168 5185 1355 5209
rect 1386 5190 1779 5210
rect 1799 5190 1802 5210
rect 1386 5185 1802 5190
rect 1168 5114 1205 5185
rect 1386 5184 1727 5185
rect 1320 5124 1351 5125
rect 1168 5094 1177 5114
rect 1197 5094 1205 5114
rect 1168 5084 1205 5094
rect 1264 5114 1351 5124
rect 1264 5094 1273 5114
rect 1293 5094 1351 5114
rect 1264 5085 1351 5094
rect 1264 5084 1301 5085
rect 189 5052 232 5057
rect 580 5063 1027 5079
rect 580 5057 608 5063
rect 859 5062 1027 5063
rect 189 5049 339 5052
rect 580 5049 607 5057
rect 189 5047 607 5049
rect 189 5029 198 5047
rect 216 5029 607 5047
rect 1320 5034 1351 5085
rect 1386 5114 1423 5184
rect 1689 5183 1726 5184
rect 1538 5124 1574 5125
rect 1386 5094 1395 5114
rect 1415 5094 1423 5114
rect 1386 5084 1423 5094
rect 1482 5114 1630 5124
rect 1730 5121 1826 5123
rect 1482 5094 1491 5114
rect 1511 5094 1601 5114
rect 1621 5094 1630 5114
rect 1482 5085 1630 5094
rect 1688 5114 1826 5121
rect 1688 5094 1697 5114
rect 1717 5094 1826 5114
rect 1688 5085 1826 5094
rect 1482 5084 1519 5085
rect 1212 5031 1253 5032
rect 189 5026 607 5029
rect 189 5020 232 5026
rect 192 5017 232 5020
rect 1107 5024 1253 5031
rect 589 5008 629 5009
rect 300 4991 629 5008
rect 1107 5004 1163 5024
rect 1183 5004 1222 5024
rect 1242 5004 1253 5024
rect 1107 4996 1253 5004
rect 1320 5027 1477 5034
rect 1320 5007 1440 5027
rect 1460 5007 1477 5027
rect 1320 4997 1477 5007
rect 1320 4996 1355 4997
rect 184 4948 227 4959
rect 184 4930 196 4948
rect 214 4930 227 4948
rect 184 4904 227 4930
rect 300 4904 327 4991
rect 589 4982 629 4991
rect 184 4883 327 4904
rect 371 4956 405 4972
rect 589 4962 982 4982
rect 1002 4962 1005 4982
rect 1320 4975 1351 4996
rect 1538 4975 1574 5085
rect 1593 5084 1630 5085
rect 1689 5084 1726 5085
rect 1649 5025 1739 5031
rect 1649 5005 1658 5025
rect 1678 5023 1739 5025
rect 1678 5005 1703 5023
rect 1649 5003 1703 5005
rect 1723 5003 1739 5023
rect 1649 4997 1739 5003
rect 1163 4974 1200 4975
rect 589 4957 1005 4962
rect 1162 4965 1200 4974
rect 589 4956 930 4957
rect 371 4886 408 4956
rect 523 4896 554 4897
rect 184 4881 321 4883
rect 184 4839 227 4881
rect 371 4866 380 4886
rect 400 4866 408 4886
rect 371 4856 408 4866
rect 467 4886 554 4896
rect 467 4866 476 4886
rect 496 4866 554 4886
rect 467 4857 554 4866
rect 467 4856 504 4857
rect 182 4829 227 4839
rect 182 4811 191 4829
rect 209 4811 227 4829
rect 182 4805 227 4811
rect 523 4806 554 4857
rect 589 4886 626 4956
rect 892 4955 929 4956
rect 1162 4945 1171 4965
rect 1191 4945 1200 4965
rect 1162 4937 1200 4945
rect 1266 4969 1351 4975
rect 1381 4974 1418 4975
rect 1266 4949 1274 4969
rect 1294 4949 1351 4969
rect 1266 4941 1351 4949
rect 1380 4965 1418 4974
rect 1380 4945 1389 4965
rect 1409 4945 1418 4965
rect 1266 4940 1302 4941
rect 1380 4937 1418 4945
rect 1484 4969 1628 4975
rect 1484 4949 1492 4969
rect 1512 4966 1600 4969
rect 1512 4949 1547 4966
rect 1484 4948 1547 4949
rect 1566 4949 1600 4966
rect 1620 4949 1628 4969
rect 1566 4948 1628 4949
rect 1484 4941 1628 4948
rect 1484 4940 1520 4941
rect 1592 4940 1628 4941
rect 1694 4974 1731 4975
rect 1694 4973 1732 4974
rect 1754 4973 1781 4977
rect 1694 4971 1781 4973
rect 1694 4965 1758 4971
rect 1694 4945 1703 4965
rect 1723 4951 1758 4965
rect 1778 4951 1781 4971
rect 1723 4946 1781 4951
rect 1723 4945 1758 4946
rect 1163 4908 1200 4937
rect 1164 4906 1200 4908
rect 741 4896 777 4897
rect 589 4866 598 4886
rect 618 4866 626 4886
rect 589 4856 626 4866
rect 685 4886 833 4896
rect 933 4893 1029 4895
rect 685 4866 694 4886
rect 714 4866 804 4886
rect 824 4866 833 4886
rect 685 4857 833 4866
rect 891 4886 1029 4893
rect 891 4866 900 4886
rect 920 4866 1029 4886
rect 1164 4884 1355 4906
rect 1381 4905 1418 4937
rect 1694 4933 1758 4945
rect 1798 4907 1825 5085
rect 1657 4905 1825 4907
rect 1381 4879 1825 4905
rect 891 4857 1029 4866
rect 685 4856 722 4857
rect 182 4802 219 4805
rect 415 4803 456 4804
rect 307 4796 456 4803
rect 307 4776 366 4796
rect 386 4776 425 4796
rect 445 4776 456 4796
rect 307 4768 456 4776
rect 523 4799 680 4806
rect 523 4779 643 4799
rect 663 4779 680 4799
rect 523 4769 680 4779
rect 523 4768 558 4769
rect 523 4747 554 4768
rect 741 4747 777 4857
rect 796 4856 833 4857
rect 892 4856 929 4857
rect 852 4797 942 4803
rect 852 4777 861 4797
rect 881 4795 942 4797
rect 881 4777 906 4795
rect 852 4775 906 4777
rect 926 4775 942 4795
rect 852 4769 942 4775
rect 366 4746 403 4747
rect 179 4738 216 4740
rect 179 4730 221 4738
rect 179 4712 189 4730
rect 207 4712 221 4730
rect 179 4703 221 4712
rect 365 4737 403 4746
rect 365 4717 374 4737
rect 394 4717 403 4737
rect 365 4709 403 4717
rect 469 4741 554 4747
rect 584 4746 621 4747
rect 469 4721 477 4741
rect 497 4721 554 4741
rect 469 4713 554 4721
rect 583 4737 621 4746
rect 583 4717 592 4737
rect 612 4717 621 4737
rect 469 4712 505 4713
rect 583 4709 621 4717
rect 687 4745 831 4747
rect 687 4741 739 4745
rect 687 4721 695 4741
rect 715 4725 739 4741
rect 759 4741 831 4745
rect 759 4725 803 4741
rect 715 4721 803 4725
rect 823 4721 831 4741
rect 687 4713 831 4721
rect 687 4712 723 4713
rect 795 4712 831 4713
rect 897 4746 934 4747
rect 897 4745 935 4746
rect 897 4737 961 4745
rect 897 4717 906 4737
rect 926 4723 961 4737
rect 981 4723 984 4743
rect 926 4718 984 4723
rect 926 4717 961 4718
rect 180 4678 221 4703
rect 366 4678 403 4709
rect 584 4678 621 4709
rect 897 4705 961 4717
rect 1001 4679 1028 4857
rect 180 4644 223 4678
rect 362 4652 429 4678
rect 584 4677 664 4678
rect 860 4677 1028 4679
rect 584 4651 1028 4677
rect 180 4633 227 4644
rect 584 4634 619 4651
rect 860 4650 1028 4651
rect 1491 4655 1531 4879
rect 1657 4878 1825 4879
rect 1889 4911 1922 5244
rect 2224 5231 2263 7046
rect 2399 7052 2843 7077
rect 2399 6871 2426 7052
rect 2568 7051 2843 7052
rect 2466 7011 2530 7023
rect 2806 7019 2843 7051
rect 2869 7050 3060 7072
rect 3361 7066 3470 7086
rect 3490 7066 3499 7086
rect 3361 7059 3499 7066
rect 3557 7086 3705 7095
rect 3557 7066 3566 7086
rect 3586 7066 3676 7086
rect 3696 7066 3705 7086
rect 3361 7057 3457 7059
rect 3557 7056 3705 7066
rect 3764 7086 3801 7096
rect 3764 7066 3772 7086
rect 3792 7066 3801 7086
rect 3613 7055 3649 7056
rect 3024 7048 3060 7050
rect 3024 7019 3061 7048
rect 2466 7010 2501 7011
rect 2443 7005 2501 7010
rect 2443 6985 2446 7005
rect 2466 6991 2501 7005
rect 2521 6991 2530 7011
rect 2466 6983 2530 6991
rect 2492 6982 2530 6983
rect 2493 6981 2530 6982
rect 2596 7015 2632 7016
rect 2704 7015 2740 7016
rect 2596 7007 2740 7015
rect 2596 6987 2604 7007
rect 2624 7005 2712 7007
rect 2624 6987 2657 7005
rect 2596 6983 2657 6987
rect 2680 6987 2712 7005
rect 2732 6987 2740 7007
rect 2680 6983 2740 6987
rect 2596 6981 2740 6983
rect 2806 7011 2844 7019
rect 2922 7015 2958 7016
rect 2806 6991 2815 7011
rect 2835 6991 2844 7011
rect 2806 6982 2844 6991
rect 2873 7007 2958 7015
rect 2873 6987 2930 7007
rect 2950 6987 2958 7007
rect 2806 6981 2843 6982
rect 2873 6981 2958 6987
rect 3024 7011 3062 7019
rect 3024 6991 3033 7011
rect 3053 6991 3062 7011
rect 3764 6999 3801 7066
rect 3836 7095 3867 7146
rect 4149 7134 4167 7152
rect 4185 7134 4201 7152
rect 3886 7095 3923 7096
rect 3836 7086 3923 7095
rect 3836 7066 3894 7086
rect 3914 7066 3923 7086
rect 3836 7056 3923 7066
rect 3982 7086 4019 7096
rect 3982 7066 3990 7086
rect 4010 7066 4019 7086
rect 3836 7055 3867 7056
rect 3461 6996 3498 6997
rect 3764 6996 3803 6999
rect 3460 6995 3803 6996
rect 3982 6995 4019 7066
rect 3024 6982 3062 6991
rect 3385 6990 3803 6995
rect 3024 6981 3061 6982
rect 2485 6953 2575 6959
rect 2485 6933 2501 6953
rect 2521 6951 2575 6953
rect 2521 6933 2546 6951
rect 2485 6931 2546 6933
rect 2566 6931 2575 6951
rect 2485 6925 2575 6931
rect 2498 6871 2535 6872
rect 2594 6871 2631 6872
rect 2650 6871 2686 6981
rect 2873 6960 2904 6981
rect 3385 6970 3388 6990
rect 3408 6970 3803 6990
rect 3832 6971 4019 6995
rect 2869 6959 2904 6960
rect 2747 6949 2904 6959
rect 2747 6929 2764 6949
rect 2784 6929 2904 6949
rect 2747 6922 2904 6929
rect 2971 6952 3120 6960
rect 2971 6932 2982 6952
rect 3002 6932 3041 6952
rect 3061 6932 3120 6952
rect 2971 6925 3120 6932
rect 3764 6945 3803 6970
rect 4149 6945 4201 7134
rect 4593 7162 4603 7180
rect 4621 7162 4633 7180
rect 4765 7178 4774 7198
rect 4794 7178 4803 7198
rect 4765 7170 4803 7178
rect 4869 7202 4954 7208
rect 4984 7207 5021 7208
rect 4869 7182 4877 7202
rect 4897 7182 4954 7202
rect 4869 7174 4954 7182
rect 4983 7198 5021 7207
rect 4983 7178 4992 7198
rect 5012 7178 5021 7198
rect 4869 7173 4905 7174
rect 4983 7170 5021 7178
rect 5087 7202 5231 7208
rect 5087 7182 5095 7202
rect 5115 7182 5148 7202
rect 5168 7182 5203 7202
rect 5223 7182 5231 7202
rect 5087 7174 5231 7182
rect 5087 7173 5123 7174
rect 5195 7173 5231 7174
rect 5297 7207 5334 7208
rect 5297 7206 5335 7207
rect 5297 7198 5361 7206
rect 5297 7178 5306 7198
rect 5326 7184 5361 7198
rect 5381 7184 5384 7204
rect 5326 7179 5384 7184
rect 5326 7178 5361 7179
rect 4593 7106 4633 7162
rect 4766 7141 4803 7170
rect 4767 7139 4803 7141
rect 4767 7117 4958 7139
rect 4984 7138 5021 7170
rect 5297 7166 5361 7178
rect 5401 7140 5428 7318
rect 6286 7293 6328 7338
rect 5260 7138 5428 7140
rect 4984 7128 5428 7138
rect 5569 7234 5756 7258
rect 5787 7239 6180 7259
rect 6200 7239 6203 7259
rect 5787 7234 6203 7239
rect 5569 7163 5606 7234
rect 5787 7233 6128 7234
rect 5721 7173 5752 7174
rect 5569 7143 5578 7163
rect 5598 7143 5606 7163
rect 5569 7133 5606 7143
rect 5665 7163 5752 7173
rect 5665 7143 5674 7163
rect 5694 7143 5752 7163
rect 5665 7134 5752 7143
rect 5665 7133 5702 7134
rect 4590 7101 4633 7106
rect 4981 7112 5428 7128
rect 4981 7106 5009 7112
rect 5260 7111 5428 7112
rect 4590 7098 4740 7101
rect 4981 7098 5008 7106
rect 4590 7096 5008 7098
rect 4590 7078 4599 7096
rect 4617 7078 5008 7096
rect 5721 7083 5752 7134
rect 5787 7163 5824 7233
rect 6090 7232 6127 7233
rect 5939 7173 5975 7174
rect 5787 7143 5796 7163
rect 5816 7143 5824 7163
rect 5787 7133 5824 7143
rect 5883 7163 6031 7173
rect 6131 7170 6227 7172
rect 5883 7143 5892 7163
rect 5912 7143 6002 7163
rect 6022 7143 6031 7163
rect 5883 7134 6031 7143
rect 6089 7163 6227 7170
rect 6089 7143 6098 7163
rect 6118 7143 6227 7163
rect 6089 7134 6227 7143
rect 5883 7133 5920 7134
rect 5613 7080 5654 7081
rect 4590 7075 5008 7078
rect 4590 7069 4633 7075
rect 4593 7066 4633 7069
rect 5508 7073 5654 7080
rect 4990 7057 5030 7058
rect 4701 7040 5030 7057
rect 5508 7053 5564 7073
rect 5584 7053 5623 7073
rect 5643 7053 5654 7073
rect 5508 7045 5654 7053
rect 5721 7076 5878 7083
rect 5721 7056 5841 7076
rect 5861 7056 5878 7076
rect 5721 7046 5878 7056
rect 5721 7045 5756 7046
rect 4585 6997 4628 7008
rect 4585 6979 4597 6997
rect 4615 6979 4628 6997
rect 4585 6953 4628 6979
rect 4701 6953 4728 7040
rect 4990 7031 5030 7040
rect 3764 6927 4203 6945
rect 2971 6924 3012 6925
rect 2705 6871 2742 6872
rect 2398 6862 2536 6871
rect 2398 6842 2507 6862
rect 2527 6842 2536 6862
rect 2398 6835 2536 6842
rect 2594 6862 2742 6871
rect 2594 6842 2603 6862
rect 2623 6842 2713 6862
rect 2733 6842 2742 6862
rect 2398 6833 2494 6835
rect 2594 6832 2742 6842
rect 2801 6862 2838 6872
rect 2801 6842 2809 6862
rect 2829 6842 2838 6862
rect 2650 6831 2686 6832
rect 2498 6772 2535 6773
rect 2801 6772 2838 6842
rect 2873 6871 2904 6922
rect 3764 6909 4164 6927
rect 4182 6909 4203 6927
rect 3764 6903 4203 6909
rect 3770 6899 4203 6903
rect 4585 6932 4728 6953
rect 4772 7005 4806 7021
rect 4990 7011 5383 7031
rect 5403 7011 5406 7031
rect 5721 7024 5752 7045
rect 5939 7024 5975 7134
rect 5994 7133 6031 7134
rect 6090 7133 6127 7134
rect 6050 7074 6140 7080
rect 6050 7054 6059 7074
rect 6079 7072 6140 7074
rect 6079 7054 6104 7072
rect 6050 7052 6104 7054
rect 6124 7052 6140 7072
rect 6050 7046 6140 7052
rect 5564 7023 5601 7024
rect 4990 7006 5406 7011
rect 5563 7014 5601 7023
rect 4990 7005 5331 7006
rect 4772 6935 4809 7005
rect 4924 6945 4955 6946
rect 4585 6930 4722 6932
rect 4149 6897 4201 6899
rect 4585 6888 4628 6930
rect 4772 6915 4781 6935
rect 4801 6915 4809 6935
rect 4772 6905 4809 6915
rect 4868 6935 4955 6945
rect 4868 6915 4877 6935
rect 4897 6915 4955 6935
rect 4868 6906 4955 6915
rect 4868 6905 4905 6906
rect 4583 6878 4628 6888
rect 2923 6871 2960 6872
rect 2873 6862 2960 6871
rect 2873 6842 2931 6862
rect 2951 6842 2960 6862
rect 2873 6832 2960 6842
rect 3019 6862 3056 6872
rect 3019 6842 3027 6862
rect 3047 6842 3056 6862
rect 4583 6860 4592 6878
rect 4610 6860 4628 6878
rect 4583 6854 4628 6860
rect 4924 6855 4955 6906
rect 4990 6935 5027 7005
rect 5293 7004 5330 7005
rect 5563 6994 5572 7014
rect 5592 6994 5601 7014
rect 5563 6986 5601 6994
rect 5667 7018 5752 7024
rect 5782 7023 5819 7024
rect 5667 6998 5675 7018
rect 5695 6998 5752 7018
rect 5667 6990 5752 6998
rect 5781 7014 5819 7023
rect 5781 6994 5790 7014
rect 5810 6994 5819 7014
rect 5667 6989 5703 6990
rect 5781 6986 5819 6994
rect 5885 7018 6029 7024
rect 5885 6998 5893 7018
rect 5913 7015 6001 7018
rect 5913 6998 5948 7015
rect 5885 6997 5948 6998
rect 5967 6998 6001 7015
rect 6021 6998 6029 7018
rect 5967 6997 6029 6998
rect 5885 6990 6029 6997
rect 5885 6989 5921 6990
rect 5993 6989 6029 6990
rect 6095 7023 6132 7024
rect 6095 7022 6133 7023
rect 6155 7022 6182 7026
rect 6095 7020 6182 7022
rect 6095 7014 6159 7020
rect 6095 6994 6104 7014
rect 6124 7000 6159 7014
rect 6179 7000 6182 7020
rect 6124 6995 6182 7000
rect 6124 6994 6159 6995
rect 5564 6957 5601 6986
rect 5565 6955 5601 6957
rect 5142 6945 5178 6946
rect 4990 6915 4999 6935
rect 5019 6915 5027 6935
rect 4990 6905 5027 6915
rect 5086 6935 5234 6945
rect 5334 6942 5430 6944
rect 5086 6915 5095 6935
rect 5115 6915 5205 6935
rect 5225 6915 5234 6935
rect 5086 6906 5234 6915
rect 5292 6935 5430 6942
rect 5292 6915 5301 6935
rect 5321 6915 5430 6935
rect 5565 6933 5756 6955
rect 5782 6954 5819 6986
rect 6095 6982 6159 6994
rect 6199 6956 6226 7134
rect 6058 6954 6226 6956
rect 5782 6928 6226 6954
rect 5292 6906 5430 6915
rect 5086 6905 5123 6906
rect 4583 6851 4620 6854
rect 4816 6852 4857 6853
rect 2873 6831 2904 6832
rect 2497 6771 2838 6772
rect 3019 6771 3056 6842
rect 4708 6845 4857 6852
rect 4152 6832 4189 6837
rect 2422 6766 2838 6771
rect 2422 6746 2425 6766
rect 2445 6746 2838 6766
rect 2869 6747 3056 6771
rect 4143 6828 4190 6832
rect 4143 6810 4162 6828
rect 4180 6810 4190 6828
rect 4708 6825 4767 6845
rect 4787 6825 4826 6845
rect 4846 6825 4857 6845
rect 4708 6817 4857 6825
rect 4924 6848 5081 6855
rect 4924 6828 5044 6848
rect 5064 6828 5081 6848
rect 4924 6818 5081 6828
rect 4924 6817 4959 6818
rect 4143 6762 4190 6810
rect 4924 6796 4955 6817
rect 5142 6796 5178 6906
rect 5197 6905 5234 6906
rect 5293 6905 5330 6906
rect 5253 6846 5343 6852
rect 5253 6826 5262 6846
rect 5282 6844 5343 6846
rect 5282 6826 5307 6844
rect 5253 6824 5307 6826
rect 5327 6824 5343 6844
rect 5253 6818 5343 6824
rect 4767 6795 4804 6796
rect 3767 6759 4190 6762
rect 2642 6745 2707 6746
rect 3745 6729 4190 6759
rect 4579 6787 4617 6789
rect 4579 6779 4622 6787
rect 4579 6761 4590 6779
rect 4608 6761 4622 6779
rect 4579 6734 4622 6761
rect 4766 6786 4804 6795
rect 4766 6766 4775 6786
rect 4795 6766 4804 6786
rect 4766 6758 4804 6766
rect 4870 6790 4955 6796
rect 4985 6795 5022 6796
rect 4870 6770 4878 6790
rect 4898 6770 4955 6790
rect 4870 6762 4955 6770
rect 4984 6786 5022 6795
rect 4984 6766 4993 6786
rect 5013 6766 5022 6786
rect 4870 6761 4906 6762
rect 4984 6758 5022 6766
rect 5088 6794 5232 6796
rect 5088 6790 5140 6794
rect 5088 6770 5096 6790
rect 5116 6774 5140 6790
rect 5160 6790 5232 6794
rect 5160 6774 5204 6790
rect 5116 6770 5204 6774
rect 5224 6770 5232 6790
rect 5088 6762 5232 6770
rect 5088 6761 5124 6762
rect 5196 6761 5232 6762
rect 5298 6795 5335 6796
rect 5298 6794 5336 6795
rect 5298 6786 5362 6794
rect 5298 6766 5307 6786
rect 5327 6772 5362 6786
rect 5382 6772 5385 6792
rect 5327 6767 5385 6772
rect 5327 6766 5362 6767
rect 2838 6713 2878 6721
rect 2838 6691 2846 6713
rect 2870 6691 2878 6713
rect 2443 6462 2480 6468
rect 2443 6443 2451 6462
rect 2472 6443 2480 6462
rect 2443 6435 2480 6443
rect 2447 6102 2480 6435
rect 2544 6467 2712 6468
rect 2838 6467 2878 6691
rect 3341 6695 3509 6696
rect 3745 6695 3786 6729
rect 4143 6708 4190 6729
rect 3341 6685 3786 6695
rect 3858 6693 4001 6694
rect 3341 6669 3785 6685
rect 3341 6667 3509 6669
rect 3705 6668 3785 6669
rect 3858 6668 4003 6693
rect 4145 6668 4190 6708
rect 3341 6489 3368 6667
rect 3408 6629 3472 6641
rect 3748 6637 3785 6668
rect 3966 6637 4003 6668
rect 4148 6661 4190 6668
rect 4580 6727 4622 6734
rect 4767 6727 4804 6758
rect 4985 6727 5022 6758
rect 5298 6754 5362 6766
rect 5402 6728 5429 6906
rect 4580 6687 4625 6727
rect 4767 6702 4912 6727
rect 4985 6726 5065 6727
rect 5261 6726 5429 6728
rect 4985 6710 5429 6726
rect 4769 6701 4912 6702
rect 4984 6700 5429 6710
rect 4580 6666 4627 6687
rect 4984 6666 5025 6700
rect 5261 6699 5429 6700
rect 5892 6704 5932 6928
rect 6058 6927 6226 6928
rect 6290 6960 6323 7293
rect 6928 7292 6955 7470
rect 6995 7432 7059 7444
rect 7335 7440 7372 7472
rect 7398 7471 7589 7493
rect 7724 7491 7833 7511
rect 7853 7491 7862 7511
rect 7724 7484 7862 7491
rect 7920 7511 8068 7520
rect 7920 7491 7929 7511
rect 7949 7491 8039 7511
rect 8059 7491 8068 7511
rect 7724 7482 7820 7484
rect 7920 7481 8068 7491
rect 8127 7511 8164 7521
rect 8127 7491 8135 7511
rect 8155 7491 8164 7511
rect 7976 7480 8012 7481
rect 7553 7469 7589 7471
rect 7553 7440 7590 7469
rect 6995 7431 7030 7432
rect 6972 7426 7030 7431
rect 6972 7406 6975 7426
rect 6995 7412 7030 7426
rect 7050 7412 7059 7432
rect 6995 7404 7059 7412
rect 7021 7403 7059 7404
rect 7022 7402 7059 7403
rect 7125 7436 7161 7437
rect 7233 7436 7269 7437
rect 7125 7428 7269 7436
rect 7125 7408 7133 7428
rect 7153 7427 7241 7428
rect 7153 7408 7188 7427
rect 7209 7408 7241 7427
rect 7261 7408 7269 7428
rect 7125 7402 7269 7408
rect 7335 7432 7373 7440
rect 7451 7436 7487 7437
rect 7335 7412 7344 7432
rect 7364 7412 7373 7432
rect 7335 7403 7373 7412
rect 7402 7428 7487 7436
rect 7402 7408 7459 7428
rect 7479 7408 7487 7428
rect 7335 7402 7372 7403
rect 7402 7402 7487 7408
rect 7553 7432 7591 7440
rect 7553 7412 7562 7432
rect 7582 7412 7591 7432
rect 7824 7421 7861 7422
rect 8127 7421 8164 7491
rect 8199 7520 8230 7571
rect 8526 7566 8571 7572
rect 8526 7548 8544 7566
rect 8562 7548 8571 7566
rect 8526 7538 8571 7548
rect 8249 7520 8286 7521
rect 8199 7511 8286 7520
rect 8199 7491 8257 7511
rect 8277 7491 8286 7511
rect 8199 7481 8286 7491
rect 8345 7511 8382 7521
rect 8345 7491 8353 7511
rect 8373 7491 8382 7511
rect 8526 7496 8569 7538
rect 8432 7494 8569 7496
rect 8199 7480 8230 7481
rect 8345 7421 8382 7491
rect 7823 7420 8164 7421
rect 7553 7403 7591 7412
rect 7748 7415 8164 7420
rect 7553 7402 7590 7403
rect 7014 7374 7104 7380
rect 7014 7354 7030 7374
rect 7050 7372 7104 7374
rect 7050 7354 7075 7372
rect 7014 7352 7075 7354
rect 7095 7352 7104 7372
rect 7014 7346 7104 7352
rect 7027 7292 7064 7293
rect 7123 7292 7160 7293
rect 7179 7292 7215 7402
rect 7402 7381 7433 7402
rect 7748 7395 7751 7415
rect 7771 7395 8164 7415
rect 8348 7405 8382 7421
rect 8426 7473 8569 7494
rect 8124 7386 8164 7395
rect 8426 7386 8453 7473
rect 8526 7447 8569 7473
rect 8526 7429 8539 7447
rect 8557 7429 8569 7447
rect 8526 7418 8569 7429
rect 7398 7380 7433 7381
rect 7276 7370 7433 7380
rect 7276 7350 7293 7370
rect 7313 7350 7433 7370
rect 7276 7343 7433 7350
rect 7500 7373 7649 7381
rect 7500 7353 7511 7373
rect 7531 7353 7570 7373
rect 7590 7353 7649 7373
rect 8124 7369 8453 7386
rect 8124 7368 8164 7369
rect 7500 7346 7649 7353
rect 8521 7357 8561 7360
rect 8521 7351 8564 7357
rect 8146 7348 8564 7351
rect 7500 7345 7541 7346
rect 7234 7292 7271 7293
rect 6927 7283 7065 7292
rect 6790 7273 6826 7279
rect 6790 7255 6795 7273
rect 6817 7255 6826 7273
rect 6790 7251 6826 7255
rect 6927 7263 7036 7283
rect 7056 7263 7065 7283
rect 6927 7256 7065 7263
rect 7123 7283 7271 7292
rect 7123 7263 7132 7283
rect 7152 7263 7242 7283
rect 7262 7263 7271 7283
rect 6927 7254 7023 7256
rect 7123 7253 7271 7263
rect 7330 7283 7367 7293
rect 7330 7263 7338 7283
rect 7358 7263 7367 7283
rect 7179 7252 7215 7253
rect 6793 7092 6826 7251
rect 7027 7193 7064 7194
rect 7330 7193 7367 7263
rect 7402 7292 7433 7343
rect 8146 7330 8537 7348
rect 8555 7330 8564 7348
rect 8146 7328 8564 7330
rect 8146 7320 8173 7328
rect 8414 7325 8564 7328
rect 7726 7314 7894 7315
rect 8145 7314 8173 7320
rect 7726 7298 8173 7314
rect 8521 7320 8564 7325
rect 7452 7292 7489 7293
rect 7402 7283 7489 7292
rect 7402 7263 7460 7283
rect 7480 7263 7489 7283
rect 7402 7253 7489 7263
rect 7548 7283 7585 7293
rect 7548 7263 7556 7283
rect 7576 7263 7585 7283
rect 7402 7252 7433 7253
rect 7026 7192 7367 7193
rect 7548 7192 7585 7263
rect 6951 7187 7367 7192
rect 6951 7167 6954 7187
rect 6974 7167 7367 7187
rect 7398 7168 7585 7192
rect 7726 7288 8170 7298
rect 7726 7286 7894 7288
rect 7726 7108 7753 7286
rect 7793 7248 7857 7260
rect 8133 7256 8170 7288
rect 8196 7287 8387 7309
rect 8351 7285 8387 7287
rect 8351 7256 8388 7285
rect 8521 7264 8561 7320
rect 7793 7247 7828 7248
rect 7770 7242 7828 7247
rect 7770 7222 7773 7242
rect 7793 7228 7828 7242
rect 7848 7228 7857 7248
rect 7793 7220 7857 7228
rect 7819 7219 7857 7220
rect 7820 7218 7857 7219
rect 7923 7252 7959 7253
rect 8031 7252 8067 7253
rect 7923 7244 8067 7252
rect 7923 7224 7931 7244
rect 7951 7224 7986 7244
rect 8006 7224 8039 7244
rect 8059 7224 8067 7244
rect 7923 7218 8067 7224
rect 8133 7248 8171 7256
rect 8249 7252 8285 7253
rect 8133 7228 8142 7248
rect 8162 7228 8171 7248
rect 8133 7219 8171 7228
rect 8200 7244 8285 7252
rect 8200 7224 8257 7244
rect 8277 7224 8285 7244
rect 8133 7218 8170 7219
rect 8200 7218 8285 7224
rect 8351 7248 8389 7256
rect 8351 7228 8360 7248
rect 8380 7228 8389 7248
rect 8521 7246 8533 7264
rect 8551 7246 8561 7264
rect 8521 7236 8561 7246
rect 8351 7219 8389 7228
rect 8351 7218 8388 7219
rect 7812 7190 7902 7196
rect 7812 7170 7828 7190
rect 7848 7188 7902 7190
rect 7848 7170 7873 7188
rect 7812 7168 7873 7170
rect 7893 7168 7902 7188
rect 7812 7162 7902 7168
rect 7825 7108 7862 7109
rect 7921 7108 7958 7109
rect 7977 7108 8013 7218
rect 8200 7197 8231 7218
rect 8196 7196 8231 7197
rect 8074 7186 8231 7196
rect 8074 7166 8091 7186
rect 8111 7166 8231 7186
rect 8074 7159 8231 7166
rect 8298 7189 8447 7197
rect 8298 7169 8309 7189
rect 8329 7169 8368 7189
rect 8388 7169 8447 7189
rect 8298 7162 8447 7169
rect 8513 7165 8565 7183
rect 8298 7161 8339 7162
rect 8032 7108 8069 7109
rect 7725 7099 7863 7108
rect 6792 7091 6829 7092
rect 6763 7090 6931 7091
rect 7057 7090 7097 7092
rect 6588 7081 6627 7087
rect 6588 7059 6596 7081
rect 6620 7059 6627 7081
rect 6290 6952 6327 6960
rect 6290 6933 6298 6952
rect 6319 6933 6327 6952
rect 6290 6927 6327 6933
rect 5892 6682 5900 6704
rect 5924 6682 5932 6704
rect 5892 6674 5932 6682
rect 3408 6628 3443 6629
rect 3385 6623 3443 6628
rect 3385 6603 3388 6623
rect 3408 6609 3443 6623
rect 3463 6609 3472 6629
rect 3408 6601 3472 6609
rect 3434 6600 3472 6601
rect 3435 6599 3472 6600
rect 3538 6633 3574 6634
rect 3646 6633 3682 6634
rect 3538 6625 3682 6633
rect 3538 6605 3546 6625
rect 3566 6621 3654 6625
rect 3566 6605 3610 6621
rect 3538 6601 3610 6605
rect 3630 6605 3654 6621
rect 3674 6605 3682 6625
rect 3630 6601 3682 6605
rect 3538 6599 3682 6601
rect 3748 6629 3786 6637
rect 3864 6633 3900 6634
rect 3748 6609 3757 6629
rect 3777 6609 3786 6629
rect 3748 6600 3786 6609
rect 3815 6625 3900 6633
rect 3815 6605 3872 6625
rect 3892 6605 3900 6625
rect 3748 6599 3785 6600
rect 3815 6599 3900 6605
rect 3966 6629 4004 6637
rect 3966 6609 3975 6629
rect 3995 6609 4004 6629
rect 3966 6600 4004 6609
rect 4148 6634 4191 6661
rect 4148 6616 4162 6634
rect 4180 6616 4191 6634
rect 4148 6608 4191 6616
rect 4153 6606 4191 6608
rect 4580 6636 5025 6666
rect 6063 6649 6128 6650
rect 4580 6633 5003 6636
rect 3966 6599 4003 6600
rect 3427 6571 3517 6577
rect 3427 6551 3443 6571
rect 3463 6569 3517 6571
rect 3463 6551 3488 6569
rect 3427 6549 3488 6551
rect 3508 6549 3517 6569
rect 3427 6543 3517 6549
rect 3440 6489 3477 6490
rect 3536 6489 3573 6490
rect 3592 6489 3628 6599
rect 3815 6578 3846 6599
rect 4580 6585 4627 6633
rect 3811 6577 3846 6578
rect 3689 6567 3846 6577
rect 3689 6547 3706 6567
rect 3726 6547 3846 6567
rect 3689 6540 3846 6547
rect 3913 6570 4062 6578
rect 3913 6550 3924 6570
rect 3944 6550 3983 6570
rect 4003 6550 4062 6570
rect 4580 6567 4590 6585
rect 4608 6567 4627 6585
rect 4580 6563 4627 6567
rect 5714 6624 5901 6648
rect 5932 6629 6325 6649
rect 6345 6629 6348 6649
rect 5932 6624 6348 6629
rect 4581 6558 4618 6563
rect 3913 6543 4062 6550
rect 5714 6553 5751 6624
rect 5932 6623 6273 6624
rect 5866 6563 5897 6564
rect 3913 6542 3954 6543
rect 4150 6541 4187 6544
rect 3647 6489 3684 6490
rect 3340 6480 3478 6489
rect 2544 6441 2988 6467
rect 2544 6439 2712 6441
rect 2544 6261 2571 6439
rect 2611 6401 2675 6413
rect 2951 6409 2988 6441
rect 3014 6440 3205 6462
rect 3340 6460 3449 6480
rect 3469 6460 3478 6480
rect 3340 6453 3478 6460
rect 3536 6480 3684 6489
rect 3536 6460 3545 6480
rect 3565 6460 3655 6480
rect 3675 6460 3684 6480
rect 3340 6451 3436 6453
rect 3536 6450 3684 6460
rect 3743 6480 3780 6490
rect 3743 6460 3751 6480
rect 3771 6460 3780 6480
rect 3592 6449 3628 6450
rect 3169 6438 3205 6440
rect 3169 6409 3206 6438
rect 2611 6400 2646 6401
rect 2588 6395 2646 6400
rect 2588 6375 2591 6395
rect 2611 6381 2646 6395
rect 2666 6381 2675 6401
rect 2611 6375 2675 6381
rect 2588 6373 2675 6375
rect 2588 6369 2615 6373
rect 2637 6372 2675 6373
rect 2638 6371 2675 6372
rect 2741 6405 2777 6406
rect 2849 6405 2885 6406
rect 2741 6398 2885 6405
rect 2741 6397 2803 6398
rect 2741 6377 2749 6397
rect 2769 6380 2803 6397
rect 2822 6397 2885 6398
rect 2822 6380 2857 6397
rect 2769 6377 2857 6380
rect 2877 6377 2885 6397
rect 2741 6371 2885 6377
rect 2951 6401 2989 6409
rect 3067 6405 3103 6406
rect 2951 6381 2960 6401
rect 2980 6381 2989 6401
rect 2951 6372 2989 6381
rect 3018 6397 3103 6405
rect 3018 6377 3075 6397
rect 3095 6377 3103 6397
rect 2951 6371 2988 6372
rect 3018 6371 3103 6377
rect 3169 6401 3207 6409
rect 3169 6381 3178 6401
rect 3198 6381 3207 6401
rect 3440 6390 3477 6391
rect 3743 6390 3780 6460
rect 3815 6489 3846 6540
rect 4142 6535 4187 6541
rect 4142 6517 4160 6535
rect 4178 6517 4187 6535
rect 5714 6533 5723 6553
rect 5743 6533 5751 6553
rect 5714 6523 5751 6533
rect 5810 6553 5897 6563
rect 5810 6533 5819 6553
rect 5839 6533 5897 6553
rect 5810 6524 5897 6533
rect 5810 6523 5847 6524
rect 4142 6507 4187 6517
rect 3865 6489 3902 6490
rect 3815 6480 3902 6489
rect 3815 6460 3873 6480
rect 3893 6460 3902 6480
rect 3815 6450 3902 6460
rect 3961 6480 3998 6490
rect 3961 6460 3969 6480
rect 3989 6460 3998 6480
rect 4142 6465 4185 6507
rect 4569 6496 4621 6498
rect 4048 6463 4185 6465
rect 3815 6449 3846 6450
rect 3961 6390 3998 6460
rect 3439 6389 3780 6390
rect 3169 6372 3207 6381
rect 3364 6384 3780 6389
rect 3169 6371 3206 6372
rect 2630 6343 2720 6349
rect 2630 6323 2646 6343
rect 2666 6341 2720 6343
rect 2666 6323 2691 6341
rect 2630 6321 2691 6323
rect 2711 6321 2720 6341
rect 2630 6315 2720 6321
rect 2643 6261 2680 6262
rect 2739 6261 2776 6262
rect 2795 6261 2831 6371
rect 3018 6350 3049 6371
rect 3364 6364 3367 6384
rect 3387 6364 3780 6384
rect 3964 6374 3998 6390
rect 4042 6442 4185 6463
rect 4567 6492 5000 6496
rect 4567 6486 5006 6492
rect 4567 6468 4588 6486
rect 4606 6468 5006 6486
rect 5866 6473 5897 6524
rect 5932 6553 5969 6623
rect 6235 6622 6272 6623
rect 6084 6563 6120 6564
rect 5932 6533 5941 6553
rect 5961 6533 5969 6553
rect 5932 6523 5969 6533
rect 6028 6553 6176 6563
rect 6276 6560 6372 6562
rect 6028 6533 6037 6553
rect 6057 6533 6147 6553
rect 6167 6533 6176 6553
rect 6028 6524 6176 6533
rect 6234 6553 6372 6560
rect 6234 6533 6243 6553
rect 6263 6533 6372 6553
rect 6234 6524 6372 6533
rect 6028 6523 6065 6524
rect 5758 6470 5799 6471
rect 4567 6450 5006 6468
rect 3740 6355 3780 6364
rect 4042 6355 4069 6442
rect 4142 6416 4185 6442
rect 4142 6398 4155 6416
rect 4173 6398 4185 6416
rect 4142 6387 4185 6398
rect 3014 6349 3049 6350
rect 2892 6339 3049 6349
rect 2892 6319 2909 6339
rect 2929 6319 3049 6339
rect 2892 6312 3049 6319
rect 3116 6342 3262 6350
rect 3116 6322 3127 6342
rect 3147 6322 3186 6342
rect 3206 6322 3262 6342
rect 3740 6338 4069 6355
rect 3740 6337 3780 6338
rect 3116 6315 3262 6322
rect 4137 6326 4177 6329
rect 4137 6320 4180 6326
rect 3762 6317 4180 6320
rect 3116 6314 3157 6315
rect 2850 6261 2887 6262
rect 2543 6252 2681 6261
rect 2543 6232 2652 6252
rect 2672 6232 2681 6252
rect 2543 6225 2681 6232
rect 2739 6252 2887 6261
rect 2739 6232 2748 6252
rect 2768 6232 2858 6252
rect 2878 6232 2887 6252
rect 2543 6223 2639 6225
rect 2739 6222 2887 6232
rect 2946 6252 2983 6262
rect 2946 6232 2954 6252
rect 2974 6232 2983 6252
rect 2795 6221 2831 6222
rect 2643 6162 2680 6163
rect 2946 6162 2983 6232
rect 3018 6261 3049 6312
rect 3762 6299 4153 6317
rect 4171 6299 4180 6317
rect 3762 6297 4180 6299
rect 3762 6289 3789 6297
rect 4030 6294 4180 6297
rect 3342 6283 3510 6284
rect 3761 6283 3789 6289
rect 3342 6267 3789 6283
rect 4137 6289 4180 6294
rect 3068 6261 3105 6262
rect 3018 6252 3105 6261
rect 3018 6232 3076 6252
rect 3096 6232 3105 6252
rect 3018 6222 3105 6232
rect 3164 6252 3201 6262
rect 3164 6232 3172 6252
rect 3192 6232 3201 6252
rect 3018 6221 3049 6222
rect 2642 6161 2983 6162
rect 3164 6161 3201 6232
rect 2567 6156 2983 6161
rect 2567 6136 2570 6156
rect 2590 6136 2983 6156
rect 3014 6137 3201 6161
rect 3342 6257 3786 6267
rect 3342 6255 3510 6257
rect 2442 6057 2484 6102
rect 3342 6077 3369 6255
rect 3409 6217 3473 6229
rect 3749 6225 3786 6257
rect 3812 6256 4003 6278
rect 3967 6254 4003 6256
rect 3967 6225 4004 6254
rect 4137 6233 4177 6289
rect 3409 6216 3444 6217
rect 3386 6211 3444 6216
rect 3386 6191 3389 6211
rect 3409 6197 3444 6211
rect 3464 6197 3473 6217
rect 3409 6189 3473 6197
rect 3435 6188 3473 6189
rect 3436 6187 3473 6188
rect 3539 6221 3575 6222
rect 3647 6221 3683 6222
rect 3539 6213 3683 6221
rect 3539 6193 3547 6213
rect 3567 6193 3602 6213
rect 3622 6193 3655 6213
rect 3675 6193 3683 6213
rect 3539 6187 3683 6193
rect 3749 6217 3787 6225
rect 3865 6221 3901 6222
rect 3749 6197 3758 6217
rect 3778 6197 3787 6217
rect 3749 6188 3787 6197
rect 3816 6213 3901 6221
rect 3816 6193 3873 6213
rect 3893 6193 3901 6213
rect 3749 6187 3786 6188
rect 3816 6187 3901 6193
rect 3967 6217 4005 6225
rect 3967 6197 3976 6217
rect 3996 6197 4005 6217
rect 4137 6215 4149 6233
rect 4167 6215 4177 6233
rect 4569 6261 4621 6450
rect 4967 6425 5006 6450
rect 5650 6463 5799 6470
rect 5650 6443 5709 6463
rect 5729 6443 5768 6463
rect 5788 6443 5799 6463
rect 5650 6435 5799 6443
rect 5866 6466 6023 6473
rect 5866 6446 5986 6466
rect 6006 6446 6023 6466
rect 5866 6436 6023 6446
rect 5866 6435 5901 6436
rect 4751 6400 4938 6424
rect 4967 6405 5362 6425
rect 5382 6405 5385 6425
rect 5866 6414 5897 6435
rect 6084 6414 6120 6524
rect 6139 6523 6176 6524
rect 6235 6523 6272 6524
rect 6195 6464 6285 6470
rect 6195 6444 6204 6464
rect 6224 6462 6285 6464
rect 6224 6444 6249 6462
rect 6195 6442 6249 6444
rect 6269 6442 6285 6462
rect 6195 6436 6285 6442
rect 5709 6413 5746 6414
rect 4967 6400 5385 6405
rect 5708 6404 5746 6413
rect 4751 6329 4788 6400
rect 4967 6399 5310 6400
rect 4967 6396 5006 6399
rect 5272 6398 5309 6399
rect 4903 6339 4934 6340
rect 4751 6309 4760 6329
rect 4780 6309 4788 6329
rect 4751 6299 4788 6309
rect 4847 6329 4934 6339
rect 4847 6309 4856 6329
rect 4876 6309 4934 6329
rect 4847 6300 4934 6309
rect 4847 6299 4884 6300
rect 4569 6243 4585 6261
rect 4603 6243 4621 6261
rect 4903 6249 4934 6300
rect 4969 6329 5006 6396
rect 5708 6384 5717 6404
rect 5737 6384 5746 6404
rect 5708 6376 5746 6384
rect 5812 6408 5897 6414
rect 5927 6413 5964 6414
rect 5812 6388 5820 6408
rect 5840 6388 5897 6408
rect 5812 6380 5897 6388
rect 5926 6404 5964 6413
rect 5926 6384 5935 6404
rect 5955 6384 5964 6404
rect 5812 6379 5848 6380
rect 5926 6376 5964 6384
rect 6030 6408 6174 6414
rect 6030 6388 6038 6408
rect 6058 6407 6146 6408
rect 6058 6389 6093 6407
rect 6111 6389 6146 6407
rect 6058 6388 6146 6389
rect 6166 6388 6174 6408
rect 6030 6380 6174 6388
rect 6030 6379 6066 6380
rect 6138 6379 6174 6380
rect 6240 6413 6277 6414
rect 6240 6412 6278 6413
rect 6240 6404 6304 6412
rect 6240 6384 6249 6404
rect 6269 6390 6304 6404
rect 6324 6390 6327 6410
rect 6269 6385 6327 6390
rect 6269 6384 6304 6385
rect 5709 6347 5746 6376
rect 5710 6345 5746 6347
rect 5121 6339 5157 6340
rect 4969 6309 4978 6329
rect 4998 6309 5006 6329
rect 4969 6299 5006 6309
rect 5065 6329 5213 6339
rect 5313 6336 5409 6338
rect 5065 6309 5074 6329
rect 5094 6309 5184 6329
rect 5204 6309 5213 6329
rect 5065 6300 5213 6309
rect 5271 6329 5409 6336
rect 5271 6309 5280 6329
rect 5300 6309 5409 6329
rect 5710 6323 5901 6345
rect 5927 6344 5964 6376
rect 6240 6372 6304 6384
rect 6344 6348 6371 6524
rect 6290 6346 6371 6348
rect 6203 6344 6371 6346
rect 5927 6318 6371 6344
rect 6037 6316 6077 6318
rect 6203 6317 6371 6318
rect 5271 6300 5409 6309
rect 6312 6315 6371 6317
rect 5065 6299 5102 6300
rect 4795 6246 4836 6247
rect 4569 6225 4621 6243
rect 4687 6239 4836 6246
rect 4137 6205 4177 6215
rect 4687 6219 4746 6239
rect 4766 6219 4805 6239
rect 4825 6219 4836 6239
rect 4687 6211 4836 6219
rect 4903 6242 5060 6249
rect 4903 6222 5023 6242
rect 5043 6222 5060 6242
rect 4903 6212 5060 6222
rect 4903 6211 4938 6212
rect 3967 6188 4005 6197
rect 4903 6190 4934 6211
rect 5121 6190 5157 6300
rect 5176 6299 5213 6300
rect 5272 6299 5309 6300
rect 5232 6240 5322 6246
rect 5232 6220 5241 6240
rect 5261 6238 5322 6240
rect 5261 6220 5286 6238
rect 5232 6218 5286 6220
rect 5306 6218 5322 6238
rect 5232 6212 5322 6218
rect 4746 6189 4783 6190
rect 3967 6187 4004 6188
rect 3428 6159 3518 6165
rect 3428 6139 3444 6159
rect 3464 6157 3518 6159
rect 3464 6139 3489 6157
rect 3428 6137 3489 6139
rect 3509 6137 3518 6157
rect 3428 6131 3518 6137
rect 3441 6077 3478 6078
rect 3537 6077 3574 6078
rect 3593 6077 3629 6187
rect 3816 6166 3847 6187
rect 4745 6180 4783 6189
rect 3812 6165 3847 6166
rect 3690 6155 3847 6165
rect 3690 6135 3707 6155
rect 3727 6135 3847 6155
rect 3690 6128 3847 6135
rect 3914 6158 4063 6166
rect 3914 6138 3925 6158
rect 3945 6138 3984 6158
rect 4004 6138 4063 6158
rect 4573 6162 4613 6172
rect 3914 6131 4063 6138
rect 4129 6134 4181 6152
rect 3914 6130 3955 6131
rect 3648 6077 3685 6078
rect 3341 6068 3479 6077
rect 2813 6057 2846 6059
rect 2442 6045 2889 6057
rect 2445 6031 2889 6045
rect 2445 6029 2613 6031
rect 2445 5851 2472 6029
rect 2512 5991 2576 6003
rect 2852 5999 2889 6031
rect 2915 6030 3106 6052
rect 3341 6048 3450 6068
rect 3470 6048 3479 6068
rect 3341 6041 3479 6048
rect 3537 6068 3685 6077
rect 3537 6048 3546 6068
rect 3566 6048 3656 6068
rect 3676 6048 3685 6068
rect 3341 6039 3437 6041
rect 3537 6038 3685 6048
rect 3744 6068 3781 6078
rect 3744 6048 3752 6068
rect 3772 6048 3781 6068
rect 3593 6037 3629 6038
rect 3070 6028 3106 6030
rect 3070 5999 3107 6028
rect 2512 5990 2547 5991
rect 2489 5985 2547 5990
rect 2489 5965 2492 5985
rect 2512 5971 2547 5985
rect 2567 5971 2576 5991
rect 2512 5963 2576 5971
rect 2538 5962 2576 5963
rect 2539 5961 2576 5962
rect 2642 5995 2678 5996
rect 2750 5995 2786 5996
rect 2642 5987 2786 5995
rect 2642 5967 2650 5987
rect 2670 5985 2758 5987
rect 2670 5967 2703 5985
rect 2642 5966 2703 5967
rect 2724 5967 2758 5985
rect 2778 5967 2786 5987
rect 2724 5966 2786 5967
rect 2642 5961 2786 5966
rect 2852 5991 2890 5999
rect 2968 5995 3004 5996
rect 2852 5971 2861 5991
rect 2881 5971 2890 5991
rect 2852 5962 2890 5971
rect 2919 5987 3004 5995
rect 2919 5967 2976 5987
rect 2996 5967 3004 5987
rect 2852 5961 2889 5962
rect 2919 5961 3004 5967
rect 3070 5991 3108 5999
rect 3070 5971 3079 5991
rect 3099 5971 3108 5991
rect 3744 5981 3781 6048
rect 3816 6077 3847 6128
rect 4129 6116 4147 6134
rect 4165 6116 4181 6134
rect 3866 6077 3903 6078
rect 3816 6068 3903 6077
rect 3816 6048 3874 6068
rect 3894 6048 3903 6068
rect 3816 6038 3903 6048
rect 3962 6068 3999 6078
rect 3962 6048 3970 6068
rect 3990 6048 3999 6068
rect 3816 6037 3847 6038
rect 3441 5978 3478 5979
rect 3744 5978 3783 5981
rect 3440 5977 3783 5978
rect 3962 5977 3999 6048
rect 3070 5962 3108 5971
rect 3365 5972 3783 5977
rect 3070 5961 3107 5962
rect 2531 5933 2621 5939
rect 2531 5913 2547 5933
rect 2567 5931 2621 5933
rect 2567 5913 2592 5931
rect 2531 5911 2592 5913
rect 2612 5911 2621 5931
rect 2531 5905 2621 5911
rect 2544 5851 2581 5852
rect 2640 5851 2677 5852
rect 2696 5851 2732 5961
rect 2919 5940 2950 5961
rect 3365 5952 3368 5972
rect 3388 5952 3783 5972
rect 3812 5953 3999 5977
rect 2915 5939 2950 5940
rect 2793 5929 2950 5939
rect 2793 5909 2810 5929
rect 2830 5909 2950 5929
rect 2793 5902 2950 5909
rect 3017 5932 3166 5940
rect 3017 5912 3028 5932
rect 3048 5912 3087 5932
rect 3107 5912 3166 5932
rect 3017 5905 3166 5912
rect 3744 5927 3783 5952
rect 4129 5927 4181 6116
rect 4573 6144 4583 6162
rect 4601 6144 4613 6162
rect 4745 6160 4754 6180
rect 4774 6160 4783 6180
rect 4745 6152 4783 6160
rect 4849 6184 4934 6190
rect 4964 6189 5001 6190
rect 4849 6164 4857 6184
rect 4877 6164 4934 6184
rect 4849 6156 4934 6164
rect 4963 6180 5001 6189
rect 4963 6160 4972 6180
rect 4992 6160 5001 6180
rect 4849 6155 4885 6156
rect 4963 6152 5001 6160
rect 5067 6184 5211 6190
rect 5067 6164 5075 6184
rect 5095 6164 5128 6184
rect 5148 6164 5183 6184
rect 5203 6164 5211 6184
rect 5067 6156 5211 6164
rect 5067 6155 5103 6156
rect 5175 6155 5211 6156
rect 5277 6189 5314 6190
rect 5277 6188 5315 6189
rect 5277 6180 5341 6188
rect 5277 6160 5286 6180
rect 5306 6166 5341 6180
rect 5361 6166 5364 6186
rect 5306 6161 5364 6166
rect 5306 6160 5341 6161
rect 4573 6088 4613 6144
rect 4746 6123 4783 6152
rect 4747 6121 4783 6123
rect 4747 6099 4938 6121
rect 4964 6120 5001 6152
rect 5277 6148 5341 6160
rect 5381 6122 5408 6300
rect 6312 6297 6341 6315
rect 5240 6120 5408 6122
rect 4964 6110 5408 6120
rect 5549 6216 5736 6240
rect 5767 6221 6160 6241
rect 6180 6221 6183 6241
rect 5767 6216 6183 6221
rect 5549 6145 5586 6216
rect 5767 6215 6108 6216
rect 5701 6155 5732 6156
rect 5549 6125 5558 6145
rect 5578 6125 5586 6145
rect 5549 6115 5586 6125
rect 5645 6145 5732 6155
rect 5645 6125 5654 6145
rect 5674 6125 5732 6145
rect 5645 6116 5732 6125
rect 5645 6115 5682 6116
rect 4570 6083 4613 6088
rect 4961 6094 5408 6110
rect 4961 6088 4989 6094
rect 5240 6093 5408 6094
rect 4570 6080 4720 6083
rect 4961 6080 4988 6088
rect 4570 6078 4988 6080
rect 4570 6060 4579 6078
rect 4597 6060 4988 6078
rect 5701 6065 5732 6116
rect 5767 6145 5804 6215
rect 6070 6214 6107 6215
rect 5919 6155 5955 6156
rect 5767 6125 5776 6145
rect 5796 6125 5804 6145
rect 5767 6115 5804 6125
rect 5863 6145 6011 6155
rect 6111 6152 6207 6154
rect 5863 6125 5872 6145
rect 5892 6125 5982 6145
rect 6002 6125 6011 6145
rect 5863 6116 6011 6125
rect 6069 6145 6207 6152
rect 6069 6125 6078 6145
rect 6098 6125 6207 6145
rect 6069 6116 6207 6125
rect 5863 6115 5900 6116
rect 5593 6062 5634 6063
rect 4570 6057 4988 6060
rect 4570 6051 4613 6057
rect 4573 6048 4613 6051
rect 5485 6055 5634 6062
rect 4970 6039 5010 6040
rect 4681 6022 5010 6039
rect 5485 6035 5544 6055
rect 5564 6035 5603 6055
rect 5623 6035 5634 6055
rect 5485 6027 5634 6035
rect 5701 6058 5858 6065
rect 5701 6038 5821 6058
rect 5841 6038 5858 6058
rect 5701 6028 5858 6038
rect 5701 6027 5736 6028
rect 4565 5979 4608 5990
rect 4565 5961 4577 5979
rect 4595 5961 4608 5979
rect 4565 5935 4608 5961
rect 4681 5935 4708 6022
rect 4970 6013 5010 6022
rect 3744 5909 4183 5927
rect 3017 5904 3058 5905
rect 2751 5851 2788 5852
rect 2444 5842 2582 5851
rect 2444 5822 2553 5842
rect 2573 5822 2582 5842
rect 2444 5815 2582 5822
rect 2640 5842 2788 5851
rect 2640 5822 2649 5842
rect 2669 5822 2759 5842
rect 2779 5822 2788 5842
rect 2444 5813 2540 5815
rect 2640 5812 2788 5822
rect 2847 5842 2884 5852
rect 2847 5822 2855 5842
rect 2875 5822 2884 5842
rect 2696 5811 2732 5812
rect 2544 5752 2581 5753
rect 2847 5752 2884 5822
rect 2919 5851 2950 5902
rect 3744 5891 4144 5909
rect 4162 5891 4183 5909
rect 3744 5885 4183 5891
rect 3750 5881 4183 5885
rect 4565 5914 4708 5935
rect 4752 5987 4786 6003
rect 4970 5993 5363 6013
rect 5383 5993 5386 6013
rect 5701 6006 5732 6027
rect 5919 6006 5955 6116
rect 5974 6115 6011 6116
rect 6070 6115 6107 6116
rect 6030 6056 6120 6062
rect 6030 6036 6039 6056
rect 6059 6054 6120 6056
rect 6059 6036 6084 6054
rect 6030 6034 6084 6036
rect 6104 6034 6120 6054
rect 6030 6028 6120 6034
rect 5544 6005 5581 6006
rect 4970 5988 5386 5993
rect 5543 5996 5581 6005
rect 4970 5987 5311 5988
rect 4752 5917 4789 5987
rect 4904 5927 4935 5928
rect 4565 5912 4702 5914
rect 4129 5879 4181 5881
rect 4565 5870 4608 5912
rect 4752 5897 4761 5917
rect 4781 5897 4789 5917
rect 4752 5887 4789 5897
rect 4848 5917 4935 5927
rect 4848 5897 4857 5917
rect 4877 5897 4935 5917
rect 4848 5888 4935 5897
rect 4848 5887 4885 5888
rect 4563 5860 4608 5870
rect 2969 5851 3006 5852
rect 2919 5842 3006 5851
rect 2919 5822 2977 5842
rect 2997 5822 3006 5842
rect 2919 5812 3006 5822
rect 3065 5842 3102 5852
rect 3065 5822 3073 5842
rect 3093 5822 3102 5842
rect 4563 5842 4572 5860
rect 4590 5842 4608 5860
rect 4563 5836 4608 5842
rect 4904 5837 4935 5888
rect 4970 5917 5007 5987
rect 5273 5986 5310 5987
rect 5543 5976 5552 5996
rect 5572 5976 5581 5996
rect 5543 5968 5581 5976
rect 5647 6000 5732 6006
rect 5762 6005 5799 6006
rect 5647 5980 5655 6000
rect 5675 5980 5732 6000
rect 5647 5972 5732 5980
rect 5761 5996 5799 6005
rect 5761 5976 5770 5996
rect 5790 5976 5799 5996
rect 5647 5971 5683 5972
rect 5761 5968 5799 5976
rect 5865 6000 6009 6006
rect 5865 5980 5873 6000
rect 5893 5981 5925 6000
rect 5946 5981 5981 6000
rect 5893 5980 5981 5981
rect 6001 5980 6009 6000
rect 5865 5972 6009 5980
rect 5865 5971 5901 5972
rect 5973 5971 6009 5972
rect 6075 6005 6112 6006
rect 6075 6004 6113 6005
rect 6075 5996 6139 6004
rect 6075 5976 6084 5996
rect 6104 5982 6139 5996
rect 6159 5982 6162 6002
rect 6104 5977 6162 5982
rect 6104 5976 6139 5977
rect 5544 5939 5581 5968
rect 5545 5937 5581 5939
rect 5122 5927 5158 5928
rect 4970 5897 4979 5917
rect 4999 5897 5007 5917
rect 4970 5887 5007 5897
rect 5066 5917 5214 5927
rect 5314 5924 5410 5926
rect 5066 5897 5075 5917
rect 5095 5897 5185 5917
rect 5205 5897 5214 5917
rect 5066 5888 5214 5897
rect 5272 5917 5410 5924
rect 5272 5897 5281 5917
rect 5301 5897 5410 5917
rect 5545 5915 5736 5937
rect 5762 5936 5799 5968
rect 6075 5964 6139 5976
rect 6179 5938 6206 6116
rect 6038 5936 6206 5938
rect 5762 5910 6206 5936
rect 5272 5888 5410 5897
rect 5066 5887 5103 5888
rect 4563 5833 4600 5836
rect 4796 5834 4837 5835
rect 2919 5811 2950 5812
rect 2543 5751 2884 5752
rect 3065 5751 3102 5822
rect 4688 5827 4837 5834
rect 4132 5814 4169 5819
rect 4123 5810 4170 5814
rect 4123 5792 4142 5810
rect 4160 5792 4170 5810
rect 4688 5807 4747 5827
rect 4767 5807 4806 5827
rect 4826 5807 4837 5827
rect 4688 5799 4837 5807
rect 4904 5830 5061 5837
rect 4904 5810 5024 5830
rect 5044 5810 5061 5830
rect 4904 5800 5061 5810
rect 4904 5799 4939 5800
rect 2468 5746 2884 5751
rect 2468 5726 2471 5746
rect 2491 5726 2884 5746
rect 2915 5727 3102 5751
rect 3727 5749 3767 5754
rect 4123 5749 4170 5792
rect 4904 5778 4935 5799
rect 5122 5778 5158 5888
rect 5177 5887 5214 5888
rect 5273 5887 5310 5888
rect 5233 5828 5323 5834
rect 5233 5808 5242 5828
rect 5262 5826 5323 5828
rect 5262 5808 5287 5826
rect 5233 5806 5287 5808
rect 5307 5806 5323 5826
rect 5233 5800 5323 5806
rect 4747 5777 4784 5778
rect 3727 5710 4170 5749
rect 4560 5769 4597 5771
rect 4560 5761 4602 5769
rect 4560 5743 4570 5761
rect 4588 5743 4602 5761
rect 4560 5734 4602 5743
rect 4746 5768 4784 5777
rect 4746 5748 4755 5768
rect 4775 5748 4784 5768
rect 4746 5740 4784 5748
rect 4850 5772 4935 5778
rect 4965 5777 5002 5778
rect 4850 5752 4858 5772
rect 4878 5752 4935 5772
rect 4850 5744 4935 5752
rect 4964 5768 5002 5777
rect 4964 5748 4973 5768
rect 4993 5748 5002 5768
rect 4850 5743 4886 5744
rect 4964 5740 5002 5748
rect 5068 5776 5212 5778
rect 5068 5772 5120 5776
rect 5068 5752 5076 5772
rect 5096 5756 5120 5772
rect 5140 5772 5212 5776
rect 5140 5756 5184 5772
rect 5096 5752 5184 5756
rect 5204 5752 5212 5772
rect 5068 5744 5212 5752
rect 5068 5743 5104 5744
rect 5176 5743 5212 5744
rect 5278 5777 5315 5778
rect 5278 5776 5316 5777
rect 5278 5768 5342 5776
rect 5278 5748 5287 5768
rect 5307 5754 5342 5768
rect 5362 5754 5365 5774
rect 5307 5749 5365 5754
rect 5307 5748 5342 5749
rect 2821 5695 2861 5703
rect 2821 5673 2829 5695
rect 2853 5673 2861 5695
rect 2527 5449 2695 5450
rect 2821 5449 2861 5673
rect 3324 5677 3492 5678
rect 3727 5677 3767 5710
rect 4123 5677 4170 5710
rect 4561 5709 4602 5734
rect 4747 5709 4784 5740
rect 4965 5709 5002 5740
rect 5278 5736 5342 5748
rect 5382 5710 5409 5888
rect 4561 5682 4610 5709
rect 4746 5683 4795 5709
rect 4964 5708 5045 5709
rect 5241 5708 5409 5710
rect 4964 5683 5409 5708
rect 4965 5682 5409 5683
rect 3324 5676 3768 5677
rect 3324 5651 3769 5676
rect 3324 5649 3492 5651
rect 3688 5650 3769 5651
rect 3938 5650 3987 5676
rect 4123 5650 4172 5677
rect 3324 5471 3351 5649
rect 3391 5611 3455 5623
rect 3731 5619 3768 5650
rect 3949 5619 3986 5650
rect 4131 5625 4172 5650
rect 4563 5649 4610 5682
rect 4966 5649 5006 5682
rect 5241 5681 5409 5682
rect 5872 5686 5912 5910
rect 6038 5909 6206 5910
rect 5872 5664 5880 5686
rect 5904 5664 5912 5686
rect 5872 5656 5912 5664
rect 3391 5610 3426 5611
rect 3368 5605 3426 5610
rect 3368 5585 3371 5605
rect 3391 5591 3426 5605
rect 3446 5591 3455 5611
rect 3391 5583 3455 5591
rect 3417 5582 3455 5583
rect 3418 5581 3455 5582
rect 3521 5615 3557 5616
rect 3629 5615 3665 5616
rect 3521 5607 3665 5615
rect 3521 5587 3529 5607
rect 3549 5603 3637 5607
rect 3549 5587 3593 5603
rect 3521 5583 3593 5587
rect 3613 5587 3637 5603
rect 3657 5587 3665 5607
rect 3613 5583 3665 5587
rect 3521 5581 3665 5583
rect 3731 5611 3769 5619
rect 3847 5615 3883 5616
rect 3731 5591 3740 5611
rect 3760 5591 3769 5611
rect 3731 5582 3769 5591
rect 3798 5607 3883 5615
rect 3798 5587 3855 5607
rect 3875 5587 3883 5607
rect 3731 5581 3768 5582
rect 3798 5581 3883 5587
rect 3949 5611 3987 5619
rect 3949 5591 3958 5611
rect 3978 5591 3987 5611
rect 3949 5582 3987 5591
rect 4131 5616 4173 5625
rect 4131 5598 4145 5616
rect 4163 5598 4173 5616
rect 4131 5590 4173 5598
rect 4136 5588 4173 5590
rect 4563 5610 5006 5649
rect 3949 5581 3986 5582
rect 3410 5553 3500 5559
rect 3410 5533 3426 5553
rect 3446 5551 3500 5553
rect 3446 5533 3471 5551
rect 3410 5531 3471 5533
rect 3491 5531 3500 5551
rect 3410 5525 3500 5531
rect 3423 5471 3460 5472
rect 3519 5471 3556 5472
rect 3575 5471 3611 5581
rect 3798 5560 3829 5581
rect 4563 5567 4610 5610
rect 4966 5605 5006 5610
rect 5631 5608 5818 5632
rect 5849 5613 6242 5633
rect 6262 5613 6265 5633
rect 5849 5608 6265 5613
rect 3794 5559 3829 5560
rect 3672 5549 3829 5559
rect 3672 5529 3689 5549
rect 3709 5529 3829 5549
rect 3672 5522 3829 5529
rect 3896 5552 4045 5560
rect 3896 5532 3907 5552
rect 3927 5532 3966 5552
rect 3986 5532 4045 5552
rect 4563 5549 4573 5567
rect 4591 5549 4610 5567
rect 4563 5545 4610 5549
rect 4564 5540 4601 5545
rect 3896 5525 4045 5532
rect 5631 5537 5668 5608
rect 5849 5607 6190 5608
rect 5783 5547 5814 5548
rect 3896 5524 3937 5525
rect 4133 5523 4170 5526
rect 3630 5471 3667 5472
rect 3323 5462 3461 5471
rect 2527 5423 2971 5449
rect 2527 5421 2695 5423
rect 2527 5243 2554 5421
rect 2594 5383 2658 5395
rect 2934 5391 2971 5423
rect 2997 5422 3188 5444
rect 3323 5442 3432 5462
rect 3452 5442 3461 5462
rect 3323 5435 3461 5442
rect 3519 5462 3667 5471
rect 3519 5442 3528 5462
rect 3548 5442 3638 5462
rect 3658 5442 3667 5462
rect 3323 5433 3419 5435
rect 3519 5432 3667 5442
rect 3726 5462 3763 5472
rect 3726 5442 3734 5462
rect 3754 5442 3763 5462
rect 3575 5431 3611 5432
rect 3152 5420 3188 5422
rect 3152 5391 3189 5420
rect 2594 5382 2629 5383
rect 2571 5377 2629 5382
rect 2571 5357 2574 5377
rect 2594 5363 2629 5377
rect 2649 5363 2658 5383
rect 2594 5355 2658 5363
rect 2620 5354 2658 5355
rect 2621 5353 2658 5354
rect 2724 5387 2760 5388
rect 2832 5387 2868 5388
rect 2724 5379 2868 5387
rect 2724 5359 2732 5379
rect 2752 5378 2840 5379
rect 2752 5359 2787 5378
rect 2808 5359 2840 5378
rect 2860 5359 2868 5379
rect 2724 5353 2868 5359
rect 2934 5383 2972 5391
rect 3050 5387 3086 5388
rect 2934 5363 2943 5383
rect 2963 5363 2972 5383
rect 2934 5354 2972 5363
rect 3001 5379 3086 5387
rect 3001 5359 3058 5379
rect 3078 5359 3086 5379
rect 2934 5353 2971 5354
rect 3001 5353 3086 5359
rect 3152 5383 3190 5391
rect 3152 5363 3161 5383
rect 3181 5363 3190 5383
rect 3423 5372 3460 5373
rect 3726 5372 3763 5442
rect 3798 5471 3829 5522
rect 4125 5517 4170 5523
rect 4125 5499 4143 5517
rect 4161 5499 4170 5517
rect 5631 5517 5640 5537
rect 5660 5517 5668 5537
rect 5631 5507 5668 5517
rect 5727 5537 5814 5547
rect 5727 5517 5736 5537
rect 5756 5517 5814 5537
rect 5727 5508 5814 5517
rect 5727 5507 5764 5508
rect 4125 5489 4170 5499
rect 3848 5471 3885 5472
rect 3798 5462 3885 5471
rect 3798 5442 3856 5462
rect 3876 5442 3885 5462
rect 3798 5432 3885 5442
rect 3944 5462 3981 5472
rect 3944 5442 3952 5462
rect 3972 5442 3981 5462
rect 4125 5447 4168 5489
rect 4552 5478 4604 5480
rect 4031 5445 4168 5447
rect 3798 5431 3829 5432
rect 3944 5372 3981 5442
rect 3422 5371 3763 5372
rect 3152 5354 3190 5363
rect 3347 5366 3763 5371
rect 3152 5353 3189 5354
rect 2613 5325 2703 5331
rect 2613 5305 2629 5325
rect 2649 5323 2703 5325
rect 2649 5305 2674 5323
rect 2613 5303 2674 5305
rect 2694 5303 2703 5323
rect 2613 5297 2703 5303
rect 2626 5243 2663 5244
rect 2722 5243 2759 5244
rect 2778 5243 2814 5353
rect 3001 5332 3032 5353
rect 3347 5346 3350 5366
rect 3370 5346 3763 5366
rect 3947 5356 3981 5372
rect 4025 5424 4168 5445
rect 4550 5474 4983 5478
rect 4550 5468 4989 5474
rect 4550 5450 4571 5468
rect 4589 5450 4989 5468
rect 5783 5457 5814 5508
rect 5849 5537 5886 5607
rect 6152 5606 6189 5607
rect 6001 5547 6037 5548
rect 5849 5517 5858 5537
rect 5878 5517 5886 5537
rect 5849 5507 5886 5517
rect 5945 5537 6093 5547
rect 6193 5544 6289 5546
rect 5945 5517 5954 5537
rect 5974 5517 6064 5537
rect 6084 5517 6093 5537
rect 5945 5508 6093 5517
rect 6151 5537 6289 5544
rect 6151 5517 6160 5537
rect 6180 5517 6289 5537
rect 6151 5508 6289 5517
rect 5945 5507 5982 5508
rect 5675 5454 5716 5455
rect 4550 5432 4989 5450
rect 3723 5337 3763 5346
rect 4025 5337 4052 5424
rect 4125 5398 4168 5424
rect 4125 5380 4138 5398
rect 4156 5380 4168 5398
rect 4125 5369 4168 5380
rect 2997 5331 3032 5332
rect 2875 5321 3032 5331
rect 2875 5301 2892 5321
rect 2912 5301 3032 5321
rect 2875 5294 3032 5301
rect 3099 5324 3248 5332
rect 3099 5304 3110 5324
rect 3130 5304 3169 5324
rect 3189 5304 3248 5324
rect 3723 5320 4052 5337
rect 3723 5319 3763 5320
rect 3099 5297 3248 5304
rect 4120 5308 4160 5311
rect 4120 5302 4163 5308
rect 3745 5299 4163 5302
rect 3099 5296 3140 5297
rect 2833 5243 2870 5244
rect 2526 5234 2664 5243
rect 2224 5059 2264 5231
rect 2526 5214 2635 5234
rect 2655 5214 2664 5234
rect 2526 5207 2664 5214
rect 2722 5234 2870 5243
rect 2722 5214 2731 5234
rect 2751 5214 2841 5234
rect 2861 5214 2870 5234
rect 2526 5205 2622 5207
rect 2722 5204 2870 5214
rect 2929 5234 2966 5244
rect 2929 5214 2937 5234
rect 2957 5214 2966 5234
rect 2778 5203 2814 5204
rect 2626 5144 2663 5145
rect 2929 5144 2966 5214
rect 3001 5243 3032 5294
rect 3745 5281 4136 5299
rect 4154 5281 4163 5299
rect 3745 5279 4163 5281
rect 3745 5271 3772 5279
rect 4013 5276 4163 5279
rect 3325 5265 3493 5266
rect 3744 5265 3772 5271
rect 3325 5249 3772 5265
rect 4120 5271 4163 5276
rect 3051 5243 3088 5244
rect 3001 5234 3088 5243
rect 3001 5214 3059 5234
rect 3079 5214 3088 5234
rect 3001 5204 3088 5214
rect 3147 5234 3184 5244
rect 3147 5214 3155 5234
rect 3175 5214 3184 5234
rect 3001 5203 3032 5204
rect 2625 5143 2966 5144
rect 3147 5143 3184 5214
rect 2550 5138 2966 5143
rect 2550 5118 2553 5138
rect 2573 5118 2966 5138
rect 2997 5119 3184 5143
rect 3325 5239 3769 5249
rect 3325 5237 3493 5239
rect 3325 5059 3352 5237
rect 3392 5199 3456 5211
rect 3732 5207 3769 5239
rect 3795 5238 3986 5260
rect 3950 5236 3986 5238
rect 3950 5207 3987 5236
rect 4120 5215 4160 5271
rect 3392 5198 3427 5199
rect 3369 5193 3427 5198
rect 3369 5173 3372 5193
rect 3392 5179 3427 5193
rect 3447 5179 3456 5199
rect 3392 5171 3456 5179
rect 3418 5170 3456 5171
rect 3419 5169 3456 5170
rect 3522 5203 3558 5204
rect 3630 5203 3666 5204
rect 3522 5195 3666 5203
rect 3522 5175 3530 5195
rect 3550 5175 3585 5195
rect 3605 5175 3638 5195
rect 3658 5175 3666 5195
rect 3522 5169 3666 5175
rect 3732 5199 3770 5207
rect 3848 5203 3884 5204
rect 3732 5179 3741 5199
rect 3761 5179 3770 5199
rect 3732 5170 3770 5179
rect 3799 5195 3884 5203
rect 3799 5175 3856 5195
rect 3876 5175 3884 5195
rect 3732 5169 3769 5170
rect 3799 5169 3884 5175
rect 3950 5199 3988 5207
rect 3950 5179 3959 5199
rect 3979 5179 3988 5199
rect 4120 5197 4132 5215
rect 4150 5197 4160 5215
rect 4552 5243 4604 5432
rect 4950 5407 4989 5432
rect 5567 5447 5716 5454
rect 5567 5427 5626 5447
rect 5646 5427 5685 5447
rect 5705 5427 5716 5447
rect 5567 5419 5716 5427
rect 5783 5450 5940 5457
rect 5783 5430 5903 5450
rect 5923 5430 5940 5450
rect 5783 5420 5940 5430
rect 5783 5419 5818 5420
rect 4734 5382 4921 5406
rect 4950 5387 5345 5407
rect 5365 5387 5368 5407
rect 5783 5398 5814 5419
rect 6001 5398 6037 5508
rect 6056 5507 6093 5508
rect 6152 5507 6189 5508
rect 6112 5448 6202 5454
rect 6112 5428 6121 5448
rect 6141 5446 6202 5448
rect 6141 5428 6166 5446
rect 6112 5426 6166 5428
rect 6186 5426 6202 5446
rect 6112 5420 6202 5426
rect 5626 5397 5663 5398
rect 4950 5382 5368 5387
rect 5625 5388 5663 5397
rect 4734 5311 4771 5382
rect 4950 5381 5293 5382
rect 4950 5378 4989 5381
rect 5255 5380 5292 5381
rect 4886 5321 4917 5322
rect 4734 5291 4743 5311
rect 4763 5291 4771 5311
rect 4734 5281 4771 5291
rect 4830 5311 4917 5321
rect 4830 5291 4839 5311
rect 4859 5291 4917 5311
rect 4830 5282 4917 5291
rect 4830 5281 4867 5282
rect 4552 5225 4568 5243
rect 4586 5225 4604 5243
rect 4886 5231 4917 5282
rect 4952 5311 4989 5378
rect 5625 5368 5634 5388
rect 5654 5368 5663 5388
rect 5625 5360 5663 5368
rect 5729 5392 5814 5398
rect 5844 5397 5881 5398
rect 5729 5372 5737 5392
rect 5757 5372 5814 5392
rect 5729 5364 5814 5372
rect 5843 5388 5881 5397
rect 5843 5368 5852 5388
rect 5872 5368 5881 5388
rect 5729 5363 5765 5364
rect 5843 5360 5881 5368
rect 5947 5392 6091 5398
rect 5947 5372 5955 5392
rect 5975 5387 6063 5392
rect 5975 5372 6011 5387
rect 5947 5370 6011 5372
rect 6030 5372 6063 5387
rect 6083 5372 6091 5392
rect 6030 5370 6091 5372
rect 5947 5364 6091 5370
rect 5947 5363 5983 5364
rect 6055 5363 6091 5364
rect 6157 5397 6194 5398
rect 6157 5396 6195 5397
rect 6157 5388 6221 5396
rect 6157 5368 6166 5388
rect 6186 5374 6221 5388
rect 6241 5374 6244 5394
rect 6186 5369 6244 5374
rect 6186 5368 6221 5369
rect 5626 5331 5663 5360
rect 5627 5329 5663 5331
rect 5104 5321 5140 5322
rect 4952 5291 4961 5311
rect 4981 5291 4989 5311
rect 4952 5281 4989 5291
rect 5048 5311 5196 5321
rect 5296 5318 5392 5320
rect 5048 5291 5057 5311
rect 5077 5291 5167 5311
rect 5187 5291 5196 5311
rect 5048 5282 5196 5291
rect 5254 5311 5392 5318
rect 5254 5291 5263 5311
rect 5283 5291 5392 5311
rect 5627 5307 5818 5329
rect 5844 5328 5881 5360
rect 6157 5356 6221 5368
rect 6261 5330 6288 5508
rect 6120 5328 6288 5330
rect 5844 5314 6288 5328
rect 6312 5351 6340 6297
rect 6312 5321 6357 5351
rect 5844 5302 6291 5314
rect 5887 5300 5920 5302
rect 5254 5282 5392 5291
rect 5048 5281 5085 5282
rect 4778 5228 4819 5229
rect 4552 5207 4604 5225
rect 4670 5221 4819 5228
rect 4120 5187 4160 5197
rect 4670 5201 4729 5221
rect 4749 5201 4788 5221
rect 4808 5201 4819 5221
rect 4670 5193 4819 5201
rect 4886 5224 5043 5231
rect 4886 5204 5006 5224
rect 5026 5204 5043 5224
rect 4886 5194 5043 5204
rect 4886 5193 4921 5194
rect 3950 5170 3988 5179
rect 4886 5172 4917 5193
rect 5104 5172 5140 5282
rect 5159 5281 5196 5282
rect 5255 5281 5292 5282
rect 5215 5222 5305 5228
rect 5215 5202 5224 5222
rect 5244 5220 5305 5222
rect 5244 5202 5269 5220
rect 5215 5200 5269 5202
rect 5289 5200 5305 5220
rect 5215 5194 5305 5200
rect 4729 5171 4766 5172
rect 3950 5169 3987 5170
rect 3411 5141 3501 5147
rect 3411 5121 3427 5141
rect 3447 5139 3501 5141
rect 3447 5121 3472 5139
rect 3411 5119 3472 5121
rect 3492 5119 3501 5139
rect 3411 5113 3501 5119
rect 3424 5059 3461 5060
rect 3520 5059 3557 5060
rect 3576 5059 3612 5169
rect 3799 5148 3830 5169
rect 4728 5162 4766 5171
rect 3795 5147 3830 5148
rect 3673 5137 3830 5147
rect 3673 5117 3690 5137
rect 3710 5117 3830 5137
rect 3673 5110 3830 5117
rect 3897 5140 4046 5148
rect 3897 5120 3908 5140
rect 3928 5120 3967 5140
rect 3987 5120 4046 5140
rect 4556 5144 4596 5154
rect 3897 5113 4046 5120
rect 4112 5116 4164 5134
rect 3897 5112 3938 5113
rect 3631 5059 3668 5060
rect 2225 5044 2264 5059
rect 3324 5050 3462 5059
rect 2225 5043 2391 5044
rect 2517 5043 2557 5045
rect 2225 5017 2667 5043
rect 2225 5015 2391 5017
rect 1889 4903 1926 4911
rect 1889 4884 1897 4903
rect 1918 4884 1926 4903
rect 1889 4878 1926 4884
rect 2225 4837 2250 5015
rect 2290 4977 2354 4989
rect 2630 4985 2667 5017
rect 2693 5016 2884 5038
rect 3324 5030 3433 5050
rect 3453 5030 3462 5050
rect 3324 5023 3462 5030
rect 3520 5050 3668 5059
rect 3520 5030 3529 5050
rect 3549 5030 3639 5050
rect 3659 5030 3668 5050
rect 3324 5021 3420 5023
rect 3520 5020 3668 5030
rect 3727 5050 3764 5060
rect 3727 5030 3735 5050
rect 3755 5030 3764 5050
rect 3576 5019 3612 5020
rect 2848 5014 2884 5016
rect 2848 4985 2885 5014
rect 2290 4976 2325 4977
rect 2267 4971 2325 4976
rect 2267 4951 2270 4971
rect 2290 4957 2325 4971
rect 2345 4957 2354 4977
rect 2290 4949 2354 4957
rect 2316 4948 2354 4949
rect 2317 4947 2354 4948
rect 2420 4981 2456 4982
rect 2528 4981 2564 4982
rect 2420 4976 2564 4981
rect 2420 4973 2482 4976
rect 2420 4953 2428 4973
rect 2448 4953 2482 4973
rect 2420 4950 2482 4953
rect 2508 4973 2564 4976
rect 2508 4953 2536 4973
rect 2556 4953 2564 4973
rect 2508 4950 2564 4953
rect 2420 4947 2564 4950
rect 2630 4977 2668 4985
rect 2746 4981 2782 4982
rect 2630 4957 2639 4977
rect 2659 4957 2668 4977
rect 2630 4948 2668 4957
rect 2697 4973 2782 4981
rect 2697 4953 2754 4973
rect 2774 4953 2782 4973
rect 2630 4947 2667 4948
rect 2697 4947 2782 4953
rect 2848 4977 2886 4985
rect 2848 4957 2857 4977
rect 2877 4957 2886 4977
rect 3727 4963 3764 5030
rect 3799 5059 3830 5110
rect 4112 5098 4130 5116
rect 4148 5098 4164 5116
rect 3849 5059 3886 5060
rect 3799 5050 3886 5059
rect 3799 5030 3857 5050
rect 3877 5030 3886 5050
rect 3799 5020 3886 5030
rect 3945 5050 3982 5060
rect 3945 5030 3953 5050
rect 3973 5030 3982 5050
rect 3799 5019 3830 5020
rect 3424 4960 3461 4961
rect 3727 4960 3766 4963
rect 3423 4959 3766 4960
rect 3945 4959 3982 5030
rect 2848 4948 2886 4957
rect 3348 4954 3766 4959
rect 2848 4947 2885 4948
rect 2309 4919 2399 4925
rect 2309 4899 2325 4919
rect 2345 4917 2399 4919
rect 2345 4899 2370 4917
rect 2309 4897 2370 4899
rect 2390 4897 2399 4917
rect 2309 4891 2399 4897
rect 2322 4837 2359 4838
rect 2418 4837 2455 4838
rect 2474 4837 2510 4947
rect 2697 4926 2728 4947
rect 3348 4934 3351 4954
rect 3371 4934 3766 4954
rect 3795 4935 3982 4959
rect 2693 4925 2728 4926
rect 2571 4915 2728 4925
rect 2571 4895 2588 4915
rect 2608 4895 2728 4915
rect 2571 4888 2728 4895
rect 2795 4918 2944 4926
rect 2795 4898 2806 4918
rect 2826 4898 2865 4918
rect 2885 4898 2944 4918
rect 2795 4891 2944 4898
rect 3727 4909 3766 4934
rect 4112 4909 4164 5098
rect 4556 5126 4566 5144
rect 4584 5126 4596 5144
rect 4728 5142 4737 5162
rect 4757 5142 4766 5162
rect 4728 5134 4766 5142
rect 4832 5166 4917 5172
rect 4947 5171 4984 5172
rect 4832 5146 4840 5166
rect 4860 5146 4917 5166
rect 4832 5138 4917 5146
rect 4946 5162 4984 5171
rect 4946 5142 4955 5162
rect 4975 5142 4984 5162
rect 4832 5137 4868 5138
rect 4946 5134 4984 5142
rect 5050 5166 5194 5172
rect 5050 5146 5058 5166
rect 5078 5146 5111 5166
rect 5131 5146 5166 5166
rect 5186 5146 5194 5166
rect 5050 5138 5194 5146
rect 5050 5137 5086 5138
rect 5158 5137 5194 5138
rect 5260 5171 5297 5172
rect 5260 5170 5298 5171
rect 5260 5162 5324 5170
rect 5260 5142 5269 5162
rect 5289 5148 5324 5162
rect 5344 5148 5347 5168
rect 5289 5143 5347 5148
rect 5289 5142 5324 5143
rect 4556 5070 4596 5126
rect 4729 5105 4766 5134
rect 4730 5103 4766 5105
rect 4730 5081 4921 5103
rect 4947 5102 4984 5134
rect 5260 5130 5324 5142
rect 5364 5104 5391 5282
rect 6249 5257 6291 5302
rect 6312 5303 6323 5321
rect 6345 5303 6357 5321
rect 6312 5297 6357 5303
rect 6313 5296 6357 5297
rect 5223 5102 5391 5104
rect 4947 5092 5391 5102
rect 5532 5198 5719 5222
rect 5750 5203 6143 5223
rect 6163 5203 6166 5223
rect 5750 5198 6166 5203
rect 5532 5127 5569 5198
rect 5750 5197 6091 5198
rect 5684 5137 5715 5138
rect 5532 5107 5541 5127
rect 5561 5107 5569 5127
rect 5532 5097 5569 5107
rect 5628 5127 5715 5137
rect 5628 5107 5637 5127
rect 5657 5107 5715 5127
rect 5628 5098 5715 5107
rect 5628 5097 5665 5098
rect 4553 5065 4596 5070
rect 4944 5076 5391 5092
rect 4944 5070 4972 5076
rect 5223 5075 5391 5076
rect 4553 5062 4703 5065
rect 4944 5062 4971 5070
rect 4553 5060 4971 5062
rect 4553 5042 4562 5060
rect 4580 5042 4971 5060
rect 5684 5047 5715 5098
rect 5750 5127 5787 5197
rect 6053 5196 6090 5197
rect 5902 5137 5938 5138
rect 5750 5107 5759 5127
rect 5779 5107 5787 5127
rect 5750 5097 5787 5107
rect 5846 5127 5994 5137
rect 6094 5134 6190 5136
rect 5846 5107 5855 5127
rect 5875 5107 5965 5127
rect 5985 5107 5994 5127
rect 5846 5098 5994 5107
rect 6052 5127 6190 5134
rect 6052 5107 6061 5127
rect 6081 5107 6190 5127
rect 6052 5098 6190 5107
rect 5846 5097 5883 5098
rect 5576 5044 5617 5045
rect 4553 5039 4971 5042
rect 4553 5033 4596 5039
rect 4556 5030 4596 5033
rect 5471 5037 5617 5044
rect 4953 5021 4993 5022
rect 4664 5004 4993 5021
rect 5471 5017 5527 5037
rect 5547 5017 5586 5037
rect 5606 5017 5617 5037
rect 5471 5009 5617 5017
rect 5684 5040 5841 5047
rect 5684 5020 5804 5040
rect 5824 5020 5841 5040
rect 5684 5010 5841 5020
rect 5684 5009 5719 5010
rect 4548 4961 4591 4972
rect 4548 4943 4560 4961
rect 4578 4943 4591 4961
rect 4548 4917 4591 4943
rect 4664 4917 4691 5004
rect 4953 4995 4993 5004
rect 3727 4891 4166 4909
rect 2795 4890 2836 4891
rect 2529 4837 2566 4838
rect 2225 4828 2360 4837
rect 2225 4808 2331 4828
rect 2351 4808 2360 4828
rect 2225 4801 2360 4808
rect 2418 4828 2566 4837
rect 2418 4808 2427 4828
rect 2447 4808 2537 4828
rect 2557 4808 2566 4828
rect 2225 4799 2318 4801
rect 2418 4798 2566 4808
rect 2625 4828 2662 4838
rect 2625 4808 2633 4828
rect 2653 4808 2662 4828
rect 2474 4797 2510 4798
rect 2322 4738 2359 4739
rect 2625 4738 2662 4808
rect 2697 4837 2728 4888
rect 3727 4873 4127 4891
rect 4145 4873 4166 4891
rect 3727 4867 4166 4873
rect 3733 4863 4166 4867
rect 4548 4896 4691 4917
rect 4735 4969 4769 4985
rect 4953 4975 5346 4995
rect 5366 4975 5369 4995
rect 5684 4988 5715 5009
rect 5902 4988 5938 5098
rect 5957 5097 5994 5098
rect 6053 5097 6090 5098
rect 6013 5038 6103 5044
rect 6013 5018 6022 5038
rect 6042 5036 6103 5038
rect 6042 5018 6067 5036
rect 6013 5016 6067 5018
rect 6087 5016 6103 5036
rect 6013 5010 6103 5016
rect 5527 4987 5564 4988
rect 4953 4970 5369 4975
rect 5526 4978 5564 4987
rect 4953 4969 5294 4970
rect 4735 4899 4772 4969
rect 4887 4909 4918 4910
rect 4548 4894 4685 4896
rect 4112 4861 4164 4863
rect 4548 4852 4591 4894
rect 4735 4879 4744 4899
rect 4764 4879 4772 4899
rect 4735 4869 4772 4879
rect 4831 4899 4918 4909
rect 4831 4879 4840 4899
rect 4860 4879 4918 4899
rect 4831 4870 4918 4879
rect 4831 4869 4868 4870
rect 4546 4842 4591 4852
rect 2747 4837 2784 4838
rect 2697 4828 2784 4837
rect 2697 4808 2755 4828
rect 2775 4808 2784 4828
rect 2697 4798 2784 4808
rect 2843 4828 2880 4838
rect 2843 4808 2851 4828
rect 2871 4808 2880 4828
rect 4546 4824 4555 4842
rect 4573 4824 4591 4842
rect 4546 4818 4591 4824
rect 4887 4819 4918 4870
rect 4953 4899 4990 4969
rect 5256 4968 5293 4969
rect 5526 4958 5535 4978
rect 5555 4958 5564 4978
rect 5526 4950 5564 4958
rect 5630 4982 5715 4988
rect 5745 4987 5782 4988
rect 5630 4962 5638 4982
rect 5658 4962 5715 4982
rect 5630 4954 5715 4962
rect 5744 4978 5782 4987
rect 5744 4958 5753 4978
rect 5773 4958 5782 4978
rect 5630 4953 5666 4954
rect 5744 4950 5782 4958
rect 5848 4982 5992 4988
rect 5848 4962 5856 4982
rect 5876 4979 5964 4982
rect 5876 4962 5911 4979
rect 5848 4961 5911 4962
rect 5930 4962 5964 4979
rect 5984 4962 5992 4982
rect 5930 4961 5992 4962
rect 5848 4954 5992 4961
rect 5848 4953 5884 4954
rect 5956 4953 5992 4954
rect 6058 4987 6095 4988
rect 6058 4986 6096 4987
rect 6118 4986 6145 4990
rect 6058 4984 6145 4986
rect 6058 4978 6122 4984
rect 6058 4958 6067 4978
rect 6087 4964 6122 4978
rect 6142 4964 6145 4984
rect 6087 4959 6145 4964
rect 6087 4958 6122 4959
rect 5527 4921 5564 4950
rect 5528 4919 5564 4921
rect 5105 4909 5141 4910
rect 4953 4879 4962 4899
rect 4982 4879 4990 4899
rect 4953 4869 4990 4879
rect 5049 4899 5197 4909
rect 5297 4906 5393 4908
rect 5049 4879 5058 4899
rect 5078 4879 5168 4899
rect 5188 4879 5197 4899
rect 5049 4870 5197 4879
rect 5255 4899 5393 4906
rect 5255 4879 5264 4899
rect 5284 4879 5393 4899
rect 5528 4897 5719 4919
rect 5745 4918 5782 4950
rect 6058 4946 6122 4958
rect 6162 4920 6189 5098
rect 6021 4918 6189 4920
rect 5745 4892 6189 4918
rect 5255 4870 5393 4879
rect 5049 4869 5086 4870
rect 4546 4815 4583 4818
rect 4779 4816 4820 4817
rect 2697 4797 2728 4798
rect 2321 4737 2662 4738
rect 2843 4737 2880 4808
rect 4671 4809 4820 4816
rect 4115 4796 4152 4801
rect 2246 4732 2662 4737
rect 2246 4712 2249 4732
rect 2269 4712 2662 4732
rect 2693 4713 2880 4737
rect 4106 4792 4153 4796
rect 4106 4774 4125 4792
rect 4143 4774 4153 4792
rect 4671 4789 4730 4809
rect 4750 4789 4789 4809
rect 4809 4789 4820 4809
rect 4671 4781 4820 4789
rect 4887 4812 5044 4819
rect 4887 4792 5007 4812
rect 5027 4792 5044 4812
rect 4887 4782 5044 4792
rect 4887 4781 4922 4782
rect 3714 4715 3752 4716
rect 4106 4715 4153 4774
rect 4887 4760 4918 4781
rect 5105 4760 5141 4870
rect 5160 4869 5197 4870
rect 5256 4869 5293 4870
rect 5216 4810 5306 4816
rect 5216 4790 5225 4810
rect 5245 4808 5306 4810
rect 5245 4790 5270 4808
rect 5216 4788 5270 4790
rect 5290 4788 5306 4808
rect 5216 4782 5306 4788
rect 4730 4759 4767 4760
rect 4543 4751 4580 4753
rect 4543 4743 4585 4751
rect 4543 4725 4553 4743
rect 4571 4725 4585 4743
rect 4543 4716 4585 4725
rect 4729 4750 4767 4759
rect 4729 4730 4738 4750
rect 4758 4730 4767 4750
rect 4729 4722 4767 4730
rect 4833 4754 4918 4760
rect 4948 4759 4985 4760
rect 4833 4734 4841 4754
rect 4861 4734 4918 4754
rect 4833 4726 4918 4734
rect 4947 4750 4985 4759
rect 4947 4730 4956 4750
rect 4976 4730 4985 4750
rect 4833 4725 4869 4726
rect 4947 4722 4985 4730
rect 5051 4758 5195 4760
rect 5051 4754 5103 4758
rect 5051 4734 5059 4754
rect 5079 4738 5103 4754
rect 5123 4754 5195 4758
rect 5123 4738 5167 4754
rect 5079 4734 5167 4738
rect 5187 4734 5195 4754
rect 5051 4726 5195 4734
rect 5051 4725 5087 4726
rect 5159 4725 5195 4726
rect 5261 4759 5298 4760
rect 5261 4758 5299 4759
rect 5261 4750 5325 4758
rect 5261 4730 5270 4750
rect 5290 4736 5325 4750
rect 5345 4736 5348 4756
rect 5290 4731 5348 4736
rect 5290 4730 5325 4731
rect 2466 4711 2531 4712
rect 581 4633 619 4634
rect 180 4595 619 4633
rect 1491 4633 1499 4655
rect 1523 4633 1531 4655
rect 1491 4625 1531 4633
rect 2802 4677 2842 4685
rect 2802 4655 2810 4677
rect 2834 4655 2842 4677
rect 3714 4677 4153 4715
rect 3714 4676 3752 4677
rect 1802 4598 1867 4599
rect 180 4536 227 4595
rect 581 4594 619 4595
rect 180 4518 190 4536
rect 208 4518 227 4536
rect 180 4514 227 4518
rect 1453 4573 1640 4597
rect 1671 4578 2064 4598
rect 2084 4578 2087 4598
rect 1671 4573 2087 4578
rect 181 4509 218 4514
rect 1453 4502 1490 4573
rect 1671 4572 2012 4573
rect 1605 4512 1636 4513
rect 1453 4482 1462 4502
rect 1482 4482 1490 4502
rect 1453 4472 1490 4482
rect 1549 4502 1636 4512
rect 1549 4482 1558 4502
rect 1578 4482 1636 4502
rect 1549 4473 1636 4482
rect 1549 4472 1586 4473
rect 169 4447 221 4449
rect 167 4443 600 4447
rect 167 4437 606 4443
rect 167 4419 188 4437
rect 206 4419 606 4437
rect 1605 4422 1636 4473
rect 1671 4502 1708 4572
rect 1974 4571 2011 4572
rect 1823 4512 1859 4513
rect 1671 4482 1680 4502
rect 1700 4482 1708 4502
rect 1671 4472 1708 4482
rect 1767 4502 1915 4512
rect 2015 4509 2111 4511
rect 1767 4482 1776 4502
rect 1796 4482 1886 4502
rect 1906 4482 1915 4502
rect 1767 4473 1915 4482
rect 1973 4502 2111 4509
rect 1973 4482 1982 4502
rect 2002 4482 2111 4502
rect 1973 4473 2111 4482
rect 1767 4472 1804 4473
rect 1497 4419 1538 4420
rect 167 4401 606 4419
rect 169 4212 221 4401
rect 567 4376 606 4401
rect 1389 4412 1538 4419
rect 1389 4392 1448 4412
rect 1468 4392 1507 4412
rect 1527 4392 1538 4412
rect 1389 4384 1538 4392
rect 1605 4415 1762 4422
rect 1605 4395 1725 4415
rect 1745 4395 1762 4415
rect 1605 4385 1762 4395
rect 1605 4384 1640 4385
rect 351 4351 538 4375
rect 567 4356 962 4376
rect 982 4356 985 4376
rect 1605 4363 1636 4384
rect 1823 4363 1859 4473
rect 1878 4472 1915 4473
rect 1974 4472 2011 4473
rect 1934 4413 2024 4419
rect 1934 4393 1943 4413
rect 1963 4411 2024 4413
rect 1963 4393 1988 4411
rect 1934 4391 1988 4393
rect 2008 4391 2024 4411
rect 1934 4385 2024 4391
rect 1448 4362 1485 4363
rect 567 4351 985 4356
rect 1447 4353 1485 4362
rect 351 4280 388 4351
rect 567 4350 910 4351
rect 567 4347 606 4350
rect 872 4349 909 4350
rect 503 4290 534 4291
rect 351 4260 360 4280
rect 380 4260 388 4280
rect 351 4250 388 4260
rect 447 4280 534 4290
rect 447 4260 456 4280
rect 476 4260 534 4280
rect 447 4251 534 4260
rect 447 4250 484 4251
rect 169 4194 185 4212
rect 203 4194 221 4212
rect 503 4200 534 4251
rect 569 4280 606 4347
rect 1447 4333 1456 4353
rect 1476 4333 1485 4353
rect 1447 4325 1485 4333
rect 1551 4357 1636 4363
rect 1666 4362 1703 4363
rect 1551 4337 1559 4357
rect 1579 4337 1636 4357
rect 1551 4329 1636 4337
rect 1665 4353 1703 4362
rect 1665 4333 1674 4353
rect 1694 4333 1703 4353
rect 1551 4328 1587 4329
rect 1665 4325 1703 4333
rect 1769 4357 1913 4363
rect 1769 4337 1777 4357
rect 1797 4351 1885 4357
rect 1797 4337 1826 4351
rect 1769 4329 1826 4337
rect 1769 4328 1805 4329
rect 1849 4337 1885 4351
rect 1905 4337 1913 4357
rect 1849 4329 1913 4337
rect 1877 4328 1913 4329
rect 1979 4362 2016 4363
rect 1979 4361 2017 4362
rect 1979 4353 2043 4361
rect 1979 4333 1988 4353
rect 2008 4339 2043 4353
rect 2063 4339 2066 4359
rect 2008 4334 2066 4339
rect 2008 4333 2043 4334
rect 1448 4296 1485 4325
rect 1449 4294 1485 4296
rect 721 4290 757 4291
rect 569 4260 578 4280
rect 598 4260 606 4280
rect 569 4250 606 4260
rect 665 4280 813 4290
rect 913 4287 1009 4289
rect 665 4260 674 4280
rect 694 4260 784 4280
rect 804 4260 813 4280
rect 665 4251 813 4260
rect 871 4280 1009 4287
rect 871 4260 880 4280
rect 900 4260 1009 4280
rect 1449 4272 1640 4294
rect 1666 4293 1703 4325
rect 1979 4321 2043 4333
rect 2083 4295 2110 4473
rect 2407 4426 2444 4432
rect 2407 4407 2415 4426
rect 2436 4407 2444 4426
rect 2407 4399 2444 4407
rect 1942 4293 2110 4295
rect 1666 4267 2110 4293
rect 1776 4265 1816 4267
rect 1942 4266 2110 4267
rect 871 4251 1009 4260
rect 2069 4261 2110 4266
rect 665 4250 702 4251
rect 395 4197 436 4198
rect 169 4176 221 4194
rect 287 4190 436 4197
rect 287 4170 346 4190
rect 366 4170 405 4190
rect 425 4170 436 4190
rect 287 4162 436 4170
rect 503 4193 660 4200
rect 503 4173 623 4193
rect 643 4173 660 4193
rect 503 4163 660 4173
rect 503 4162 538 4163
rect 503 4141 534 4162
rect 721 4141 757 4251
rect 776 4250 813 4251
rect 872 4250 909 4251
rect 832 4191 922 4197
rect 832 4171 841 4191
rect 861 4189 922 4191
rect 861 4171 886 4189
rect 832 4169 886 4171
rect 906 4169 922 4189
rect 832 4163 922 4169
rect 346 4140 383 4141
rect 345 4131 383 4140
rect 173 4113 213 4123
rect 173 4095 183 4113
rect 201 4095 213 4113
rect 345 4111 354 4131
rect 374 4111 383 4131
rect 345 4103 383 4111
rect 449 4135 534 4141
rect 564 4140 601 4141
rect 449 4115 457 4135
rect 477 4115 534 4135
rect 449 4107 534 4115
rect 563 4131 601 4140
rect 563 4111 572 4131
rect 592 4111 601 4131
rect 449 4106 485 4107
rect 563 4103 601 4111
rect 667 4135 811 4141
rect 667 4115 675 4135
rect 695 4115 728 4135
rect 748 4115 783 4135
rect 803 4115 811 4135
rect 667 4107 811 4115
rect 667 4106 703 4107
rect 775 4106 811 4107
rect 877 4140 914 4141
rect 877 4139 915 4140
rect 877 4131 941 4139
rect 877 4111 886 4131
rect 906 4117 941 4131
rect 961 4117 964 4137
rect 906 4112 964 4117
rect 906 4111 941 4112
rect 173 4039 213 4095
rect 346 4074 383 4103
rect 347 4072 383 4074
rect 347 4050 538 4072
rect 564 4071 601 4103
rect 877 4099 941 4111
rect 981 4073 1008 4251
rect 840 4071 1008 4073
rect 564 4061 1008 4071
rect 1149 4167 1336 4191
rect 1367 4172 1760 4192
rect 1780 4172 1783 4192
rect 1367 4167 1783 4172
rect 1149 4096 1186 4167
rect 1367 4166 1708 4167
rect 1301 4106 1332 4107
rect 1149 4076 1158 4096
rect 1178 4076 1186 4096
rect 1149 4066 1186 4076
rect 1245 4096 1332 4106
rect 1245 4076 1254 4096
rect 1274 4076 1332 4096
rect 1245 4067 1332 4076
rect 1245 4066 1282 4067
rect 170 4034 213 4039
rect 561 4045 1008 4061
rect 561 4039 589 4045
rect 840 4044 1008 4045
rect 170 4031 320 4034
rect 561 4031 588 4039
rect 170 4029 588 4031
rect 170 4011 179 4029
rect 197 4011 588 4029
rect 1301 4016 1332 4067
rect 1367 4096 1404 4166
rect 1670 4165 1707 4166
rect 1519 4106 1555 4107
rect 1367 4076 1376 4096
rect 1396 4076 1404 4096
rect 1367 4066 1404 4076
rect 1463 4096 1611 4106
rect 1711 4103 1807 4105
rect 1463 4076 1472 4096
rect 1492 4076 1582 4096
rect 1602 4076 1611 4096
rect 1463 4067 1611 4076
rect 1669 4096 1807 4103
rect 1669 4076 1678 4096
rect 1698 4076 1807 4096
rect 2069 4079 2109 4261
rect 1669 4067 1807 4076
rect 1463 4066 1500 4067
rect 1193 4013 1234 4014
rect 170 4008 588 4011
rect 170 4002 213 4008
rect 173 3999 213 4002
rect 1085 4006 1234 4013
rect 570 3990 610 3991
rect 281 3973 610 3990
rect 1085 3986 1144 4006
rect 1164 3986 1203 4006
rect 1223 3986 1234 4006
rect 1085 3978 1234 3986
rect 1301 4009 1458 4016
rect 1301 3989 1421 4009
rect 1441 3989 1458 4009
rect 1301 3979 1458 3989
rect 1301 3978 1336 3979
rect 165 3930 208 3941
rect 165 3912 177 3930
rect 195 3912 208 3930
rect 165 3886 208 3912
rect 281 3886 308 3973
rect 570 3964 610 3973
rect 165 3865 308 3886
rect 352 3938 386 3954
rect 570 3944 963 3964
rect 983 3944 986 3964
rect 1301 3957 1332 3978
rect 1519 3957 1555 4067
rect 1574 4066 1611 4067
rect 1670 4066 1707 4067
rect 1630 4007 1720 4013
rect 1630 3987 1639 4007
rect 1659 4005 1720 4007
rect 1659 3987 1684 4005
rect 1630 3985 1684 3987
rect 1704 3985 1720 4005
rect 1630 3979 1720 3985
rect 1144 3956 1181 3957
rect 570 3939 986 3944
rect 1143 3947 1181 3956
rect 570 3938 911 3939
rect 352 3868 389 3938
rect 504 3878 535 3879
rect 165 3863 302 3865
rect 165 3821 208 3863
rect 352 3848 361 3868
rect 381 3848 389 3868
rect 352 3838 389 3848
rect 448 3868 535 3878
rect 448 3848 457 3868
rect 477 3848 535 3868
rect 448 3839 535 3848
rect 448 3838 485 3839
rect 163 3811 208 3821
rect 163 3793 172 3811
rect 190 3793 208 3811
rect 163 3787 208 3793
rect 504 3788 535 3839
rect 570 3868 607 3938
rect 873 3937 910 3938
rect 1143 3927 1152 3947
rect 1172 3927 1181 3947
rect 1143 3919 1181 3927
rect 1247 3951 1332 3957
rect 1362 3956 1399 3957
rect 1247 3931 1255 3951
rect 1275 3931 1332 3951
rect 1247 3923 1332 3931
rect 1361 3947 1399 3956
rect 1361 3927 1370 3947
rect 1390 3927 1399 3947
rect 1247 3922 1283 3923
rect 1361 3919 1399 3927
rect 1465 3951 1609 3957
rect 1465 3931 1473 3951
rect 1493 3932 1525 3951
rect 1546 3932 1581 3951
rect 1493 3931 1581 3932
rect 1601 3931 1609 3951
rect 1465 3923 1609 3931
rect 1465 3922 1501 3923
rect 1573 3922 1609 3923
rect 1675 3956 1712 3957
rect 1675 3955 1713 3956
rect 1675 3947 1739 3955
rect 1675 3927 1684 3947
rect 1704 3933 1739 3947
rect 1759 3933 1762 3953
rect 1704 3928 1762 3933
rect 1704 3927 1739 3928
rect 1144 3890 1181 3919
rect 1145 3888 1181 3890
rect 722 3878 758 3879
rect 570 3848 579 3868
rect 599 3848 607 3868
rect 570 3838 607 3848
rect 666 3868 814 3878
rect 914 3875 1010 3877
rect 666 3848 675 3868
rect 695 3848 785 3868
rect 805 3848 814 3868
rect 666 3839 814 3848
rect 872 3868 1010 3875
rect 872 3848 881 3868
rect 901 3848 1010 3868
rect 1145 3866 1336 3888
rect 1362 3887 1399 3919
rect 1675 3915 1739 3927
rect 1779 3889 1806 4067
rect 1638 3887 1806 3889
rect 1362 3861 1806 3887
rect 872 3839 1010 3848
rect 666 3838 703 3839
rect 163 3784 200 3787
rect 396 3785 437 3786
rect 288 3778 437 3785
rect 288 3758 347 3778
rect 367 3758 406 3778
rect 426 3758 437 3778
rect 288 3750 437 3758
rect 504 3781 661 3788
rect 504 3761 624 3781
rect 644 3761 661 3781
rect 504 3751 661 3761
rect 504 3750 539 3751
rect 504 3729 535 3750
rect 722 3729 758 3839
rect 777 3838 814 3839
rect 873 3838 910 3839
rect 833 3779 923 3785
rect 833 3759 842 3779
rect 862 3777 923 3779
rect 862 3759 887 3777
rect 833 3757 887 3759
rect 907 3757 923 3777
rect 833 3751 923 3757
rect 347 3728 384 3729
rect 160 3720 197 3722
rect 160 3712 202 3720
rect 160 3694 170 3712
rect 188 3694 202 3712
rect 160 3685 202 3694
rect 346 3719 384 3728
rect 346 3699 355 3719
rect 375 3699 384 3719
rect 346 3691 384 3699
rect 450 3723 535 3729
rect 565 3728 602 3729
rect 450 3703 458 3723
rect 478 3703 535 3723
rect 450 3695 535 3703
rect 564 3719 602 3728
rect 564 3699 573 3719
rect 593 3699 602 3719
rect 450 3694 486 3695
rect 564 3691 602 3699
rect 668 3727 812 3729
rect 668 3723 720 3727
rect 668 3703 676 3723
rect 696 3707 720 3723
rect 740 3723 812 3727
rect 740 3707 784 3723
rect 696 3703 784 3707
rect 804 3703 812 3723
rect 668 3695 812 3703
rect 668 3694 704 3695
rect 776 3694 812 3695
rect 878 3728 915 3729
rect 878 3727 916 3728
rect 878 3719 942 3727
rect 878 3699 887 3719
rect 907 3705 942 3719
rect 962 3705 965 3725
rect 907 3700 965 3705
rect 907 3699 942 3700
rect 161 3660 202 3685
rect 347 3660 384 3691
rect 565 3660 602 3691
rect 878 3687 942 3699
rect 982 3661 1009 3839
rect 161 3633 210 3660
rect 346 3634 395 3660
rect 564 3659 645 3660
rect 841 3659 1009 3661
rect 564 3634 1009 3659
rect 565 3633 1009 3634
rect 163 3600 210 3633
rect 566 3600 606 3633
rect 841 3632 1009 3633
rect 1472 3637 1512 3861
rect 1638 3860 1806 3861
rect 1472 3615 1480 3637
rect 1504 3615 1512 3637
rect 1472 3607 1512 3615
rect 163 3561 606 3600
rect 163 3518 210 3561
rect 566 3556 606 3561
rect 1231 3559 1418 3583
rect 1449 3564 1842 3584
rect 1862 3564 1865 3584
rect 1449 3559 1865 3564
rect 163 3500 173 3518
rect 191 3500 210 3518
rect 163 3496 210 3500
rect 164 3491 201 3496
rect 1231 3488 1268 3559
rect 1449 3558 1790 3559
rect 1383 3498 1414 3499
rect 1231 3468 1240 3488
rect 1260 3468 1268 3488
rect 1231 3458 1268 3468
rect 1327 3488 1414 3498
rect 1327 3468 1336 3488
rect 1356 3468 1414 3488
rect 1327 3459 1414 3468
rect 1327 3458 1364 3459
rect 152 3429 204 3431
rect 150 3425 583 3429
rect 150 3419 589 3425
rect 150 3401 171 3419
rect 189 3401 589 3419
rect 1383 3408 1414 3459
rect 1449 3488 1486 3558
rect 1752 3557 1789 3558
rect 1601 3498 1637 3499
rect 1449 3468 1458 3488
rect 1478 3468 1486 3488
rect 1449 3458 1486 3468
rect 1545 3488 1693 3498
rect 1793 3495 1889 3497
rect 1545 3468 1554 3488
rect 1574 3468 1664 3488
rect 1684 3468 1693 3488
rect 1545 3459 1693 3468
rect 1751 3488 1889 3495
rect 1751 3468 1760 3488
rect 1780 3468 1889 3488
rect 1751 3459 1889 3468
rect 1545 3458 1582 3459
rect 1275 3405 1316 3406
rect 150 3383 589 3401
rect 152 3194 204 3383
rect 550 3358 589 3383
rect 1167 3398 1316 3405
rect 1167 3378 1226 3398
rect 1246 3378 1285 3398
rect 1305 3378 1316 3398
rect 1167 3370 1316 3378
rect 1383 3401 1540 3408
rect 1383 3381 1503 3401
rect 1523 3381 1540 3401
rect 1383 3371 1540 3381
rect 1383 3370 1418 3371
rect 334 3333 521 3357
rect 550 3338 945 3358
rect 965 3338 968 3358
rect 1383 3349 1414 3370
rect 1601 3349 1637 3459
rect 1656 3458 1693 3459
rect 1752 3458 1789 3459
rect 1712 3399 1802 3405
rect 1712 3379 1721 3399
rect 1741 3397 1802 3399
rect 1741 3379 1766 3397
rect 1712 3377 1766 3379
rect 1786 3377 1802 3397
rect 1712 3371 1802 3377
rect 1226 3348 1263 3349
rect 550 3333 968 3338
rect 1225 3339 1263 3348
rect 334 3262 371 3333
rect 550 3332 893 3333
rect 550 3329 589 3332
rect 855 3331 892 3332
rect 486 3272 517 3273
rect 334 3242 343 3262
rect 363 3242 371 3262
rect 334 3232 371 3242
rect 430 3262 517 3272
rect 430 3242 439 3262
rect 459 3242 517 3262
rect 430 3233 517 3242
rect 430 3232 467 3233
rect 152 3176 168 3194
rect 186 3176 204 3194
rect 486 3182 517 3233
rect 552 3262 589 3329
rect 1225 3319 1234 3339
rect 1254 3319 1263 3339
rect 1225 3311 1263 3319
rect 1329 3343 1414 3349
rect 1444 3348 1481 3349
rect 1329 3323 1337 3343
rect 1357 3323 1414 3343
rect 1329 3315 1414 3323
rect 1443 3339 1481 3348
rect 1443 3319 1452 3339
rect 1472 3319 1481 3339
rect 1329 3314 1365 3315
rect 1443 3311 1481 3319
rect 1547 3344 1691 3349
rect 1547 3343 1609 3344
rect 1547 3323 1555 3343
rect 1575 3325 1609 3343
rect 1630 3343 1691 3344
rect 1630 3325 1663 3343
rect 1575 3323 1663 3325
rect 1683 3323 1691 3343
rect 1547 3315 1691 3323
rect 1547 3314 1583 3315
rect 1655 3314 1691 3315
rect 1757 3348 1794 3349
rect 1757 3347 1795 3348
rect 1757 3339 1821 3347
rect 1757 3319 1766 3339
rect 1786 3325 1821 3339
rect 1841 3325 1844 3345
rect 1786 3320 1844 3325
rect 1786 3319 1821 3320
rect 1226 3282 1263 3311
rect 1227 3280 1263 3282
rect 704 3272 740 3273
rect 552 3242 561 3262
rect 581 3242 589 3262
rect 552 3232 589 3242
rect 648 3262 796 3272
rect 896 3269 992 3271
rect 648 3242 657 3262
rect 677 3242 767 3262
rect 787 3242 796 3262
rect 648 3233 796 3242
rect 854 3262 992 3269
rect 854 3242 863 3262
rect 883 3242 992 3262
rect 1227 3258 1418 3280
rect 1444 3279 1481 3311
rect 1757 3307 1821 3319
rect 1861 3281 1888 3459
rect 1720 3279 1888 3281
rect 1444 3265 1888 3279
rect 1444 3253 1891 3265
rect 1487 3251 1520 3253
rect 854 3233 992 3242
rect 648 3232 685 3233
rect 378 3179 419 3180
rect 152 3158 204 3176
rect 270 3172 419 3179
rect 270 3152 329 3172
rect 349 3152 388 3172
rect 408 3152 419 3172
rect 270 3144 419 3152
rect 486 3175 643 3182
rect 486 3155 606 3175
rect 626 3155 643 3175
rect 486 3145 643 3155
rect 486 3144 521 3145
rect 486 3123 517 3144
rect 704 3123 740 3233
rect 759 3232 796 3233
rect 855 3232 892 3233
rect 815 3173 905 3179
rect 815 3153 824 3173
rect 844 3171 905 3173
rect 844 3153 869 3171
rect 815 3151 869 3153
rect 889 3151 905 3171
rect 815 3145 905 3151
rect 329 3122 366 3123
rect 328 3113 366 3122
rect 156 3095 196 3105
rect 156 3077 166 3095
rect 184 3077 196 3095
rect 328 3093 337 3113
rect 357 3093 366 3113
rect 328 3085 366 3093
rect 432 3117 517 3123
rect 547 3122 584 3123
rect 432 3097 440 3117
rect 460 3097 517 3117
rect 432 3089 517 3097
rect 546 3113 584 3122
rect 546 3093 555 3113
rect 575 3093 584 3113
rect 432 3088 468 3089
rect 546 3085 584 3093
rect 650 3117 794 3123
rect 650 3097 658 3117
rect 678 3097 711 3117
rect 731 3097 766 3117
rect 786 3097 794 3117
rect 650 3089 794 3097
rect 650 3088 686 3089
rect 758 3088 794 3089
rect 860 3122 897 3123
rect 860 3121 898 3122
rect 860 3113 924 3121
rect 860 3093 869 3113
rect 889 3099 924 3113
rect 944 3099 947 3119
rect 889 3094 947 3099
rect 889 3093 924 3094
rect 156 3021 196 3077
rect 329 3056 366 3085
rect 330 3054 366 3056
rect 330 3032 521 3054
rect 547 3053 584 3085
rect 860 3081 924 3093
rect 964 3055 991 3233
rect 1849 3208 1891 3253
rect 823 3053 991 3055
rect 547 3043 991 3053
rect 1132 3149 1319 3173
rect 1350 3154 1743 3174
rect 1763 3154 1766 3174
rect 1350 3149 1766 3154
rect 1132 3078 1169 3149
rect 1350 3148 1691 3149
rect 1284 3088 1315 3089
rect 1132 3058 1141 3078
rect 1161 3058 1169 3078
rect 1132 3048 1169 3058
rect 1228 3078 1315 3088
rect 1228 3058 1237 3078
rect 1257 3058 1315 3078
rect 1228 3049 1315 3058
rect 1228 3048 1265 3049
rect 153 3016 196 3021
rect 544 3027 991 3043
rect 544 3021 572 3027
rect 823 3026 991 3027
rect 153 3013 303 3016
rect 544 3013 571 3021
rect 153 3011 571 3013
rect 153 2993 162 3011
rect 180 2993 571 3011
rect 1284 2998 1315 3049
rect 1350 3078 1387 3148
rect 1653 3147 1690 3148
rect 1502 3088 1538 3089
rect 1350 3058 1359 3078
rect 1379 3058 1387 3078
rect 1350 3048 1387 3058
rect 1446 3078 1594 3088
rect 1694 3085 1790 3087
rect 1446 3058 1455 3078
rect 1475 3058 1565 3078
rect 1585 3058 1594 3078
rect 1446 3049 1594 3058
rect 1652 3078 1790 3085
rect 1652 3058 1661 3078
rect 1681 3058 1790 3078
rect 1652 3049 1790 3058
rect 1446 3048 1483 3049
rect 1176 2995 1217 2996
rect 153 2990 571 2993
rect 153 2984 196 2990
rect 156 2981 196 2984
rect 1071 2988 1217 2995
rect 553 2972 593 2973
rect 264 2955 593 2972
rect 1071 2968 1127 2988
rect 1147 2968 1186 2988
rect 1206 2968 1217 2988
rect 1071 2960 1217 2968
rect 1284 2991 1441 2998
rect 1284 2971 1404 2991
rect 1424 2971 1441 2991
rect 1284 2961 1441 2971
rect 1284 2960 1319 2961
rect 148 2912 191 2923
rect 148 2894 160 2912
rect 178 2894 191 2912
rect 148 2868 191 2894
rect 264 2868 291 2955
rect 553 2946 593 2955
rect 148 2847 291 2868
rect 335 2920 369 2936
rect 553 2926 946 2946
rect 966 2926 969 2946
rect 1284 2939 1315 2960
rect 1502 2939 1538 3049
rect 1557 3048 1594 3049
rect 1653 3048 1690 3049
rect 1613 2989 1703 2995
rect 1613 2969 1622 2989
rect 1642 2987 1703 2989
rect 1642 2969 1667 2987
rect 1613 2967 1667 2969
rect 1687 2967 1703 2987
rect 1613 2961 1703 2967
rect 1127 2938 1164 2939
rect 553 2921 969 2926
rect 1126 2929 1164 2938
rect 553 2920 894 2921
rect 335 2850 372 2920
rect 487 2860 518 2861
rect 148 2845 285 2847
rect 148 2803 191 2845
rect 335 2830 344 2850
rect 364 2830 372 2850
rect 335 2820 372 2830
rect 431 2850 518 2860
rect 431 2830 440 2850
rect 460 2830 518 2850
rect 431 2821 518 2830
rect 431 2820 468 2821
rect 146 2793 191 2803
rect 146 2775 155 2793
rect 173 2775 191 2793
rect 146 2769 191 2775
rect 487 2770 518 2821
rect 553 2850 590 2920
rect 856 2919 893 2920
rect 1126 2909 1135 2929
rect 1155 2909 1164 2929
rect 1126 2901 1164 2909
rect 1230 2933 1315 2939
rect 1345 2938 1382 2939
rect 1230 2913 1238 2933
rect 1258 2913 1315 2933
rect 1230 2905 1315 2913
rect 1344 2929 1382 2938
rect 1344 2909 1353 2929
rect 1373 2909 1382 2929
rect 1230 2904 1266 2905
rect 1344 2901 1382 2909
rect 1448 2933 1592 2939
rect 1448 2913 1456 2933
rect 1476 2930 1564 2933
rect 1476 2913 1511 2930
rect 1448 2912 1511 2913
rect 1530 2913 1564 2930
rect 1584 2913 1592 2933
rect 1530 2912 1592 2913
rect 1448 2905 1592 2912
rect 1448 2904 1484 2905
rect 1556 2904 1592 2905
rect 1658 2938 1695 2939
rect 1658 2937 1696 2938
rect 1718 2937 1745 2941
rect 1658 2935 1745 2937
rect 1658 2929 1722 2935
rect 1658 2909 1667 2929
rect 1687 2915 1722 2929
rect 1742 2915 1745 2935
rect 1687 2910 1745 2915
rect 1687 2909 1722 2910
rect 1127 2872 1164 2901
rect 1128 2870 1164 2872
rect 705 2860 741 2861
rect 553 2830 562 2850
rect 582 2830 590 2850
rect 553 2820 590 2830
rect 649 2850 797 2860
rect 897 2857 993 2859
rect 649 2830 658 2850
rect 678 2830 768 2850
rect 788 2830 797 2850
rect 649 2821 797 2830
rect 855 2850 993 2857
rect 855 2830 864 2850
rect 884 2830 993 2850
rect 1128 2848 1319 2870
rect 1345 2869 1382 2901
rect 1658 2897 1722 2909
rect 1762 2871 1789 3049
rect 1621 2869 1789 2871
rect 1345 2843 1789 2869
rect 855 2821 993 2830
rect 649 2820 686 2821
rect 146 2766 183 2769
rect 379 2767 420 2768
rect 271 2760 420 2767
rect 271 2740 330 2760
rect 350 2740 389 2760
rect 409 2740 420 2760
rect 271 2732 420 2740
rect 487 2763 644 2770
rect 487 2743 607 2763
rect 627 2743 644 2763
rect 487 2733 644 2743
rect 487 2732 522 2733
rect 487 2711 518 2732
rect 705 2711 741 2821
rect 760 2820 797 2821
rect 856 2820 893 2821
rect 816 2761 906 2767
rect 816 2741 825 2761
rect 845 2759 906 2761
rect 845 2741 870 2759
rect 816 2739 870 2741
rect 890 2739 906 2759
rect 816 2733 906 2739
rect 330 2710 367 2711
rect 142 2702 180 2704
rect 142 2694 185 2702
rect 142 2676 153 2694
rect 171 2676 185 2694
rect 142 2649 185 2676
rect 329 2701 367 2710
rect 329 2681 338 2701
rect 358 2681 367 2701
rect 329 2673 367 2681
rect 433 2705 518 2711
rect 548 2710 585 2711
rect 433 2685 441 2705
rect 461 2685 518 2705
rect 433 2677 518 2685
rect 547 2701 585 2710
rect 547 2681 556 2701
rect 576 2681 585 2701
rect 433 2676 469 2677
rect 547 2673 585 2681
rect 651 2709 795 2711
rect 651 2705 703 2709
rect 651 2685 659 2705
rect 679 2689 703 2705
rect 723 2705 795 2709
rect 723 2689 767 2705
rect 679 2685 767 2689
rect 787 2685 795 2705
rect 651 2677 795 2685
rect 651 2676 687 2677
rect 759 2676 795 2677
rect 861 2710 898 2711
rect 861 2709 899 2710
rect 861 2701 925 2709
rect 861 2681 870 2701
rect 890 2687 925 2701
rect 945 2687 948 2707
rect 890 2682 948 2687
rect 890 2681 925 2682
rect 143 2642 185 2649
rect 330 2642 367 2673
rect 548 2642 585 2673
rect 861 2669 925 2681
rect 965 2643 992 2821
rect 143 2602 188 2642
rect 330 2617 475 2642
rect 548 2641 628 2642
rect 824 2641 992 2643
rect 548 2625 992 2641
rect 332 2616 475 2617
rect 547 2615 992 2625
rect 143 2581 190 2602
rect 547 2581 588 2615
rect 824 2614 992 2615
rect 1455 2619 1495 2843
rect 1621 2842 1789 2843
rect 1853 2875 1886 3208
rect 1853 2867 1890 2875
rect 1853 2848 1861 2867
rect 1882 2848 1890 2867
rect 1853 2842 1890 2848
rect 1455 2597 1463 2619
rect 1487 2597 1495 2619
rect 1455 2589 1495 2597
rect 143 2551 588 2581
rect 1626 2564 1691 2565
rect 143 2548 566 2551
rect 143 2500 190 2548
rect 143 2482 153 2500
rect 171 2482 190 2500
rect 143 2478 190 2482
rect 1277 2539 1464 2563
rect 1495 2544 1888 2564
rect 1908 2544 1911 2564
rect 1495 2539 1911 2544
rect 144 2473 181 2478
rect 1277 2468 1314 2539
rect 1495 2538 1836 2539
rect 1429 2478 1460 2479
rect 1277 2448 1286 2468
rect 1306 2448 1314 2468
rect 1277 2438 1314 2448
rect 1373 2468 1460 2478
rect 1373 2448 1382 2468
rect 1402 2448 1460 2468
rect 1373 2439 1460 2448
rect 1373 2438 1410 2439
rect 132 2411 184 2413
rect 130 2407 563 2411
rect 130 2401 569 2407
rect 130 2383 151 2401
rect 169 2383 569 2401
rect 1429 2388 1460 2439
rect 1495 2468 1532 2538
rect 1798 2537 1835 2538
rect 1647 2478 1683 2479
rect 1495 2448 1504 2468
rect 1524 2448 1532 2468
rect 1495 2438 1532 2448
rect 1591 2468 1739 2478
rect 1839 2475 1935 2477
rect 1591 2448 1600 2468
rect 1620 2448 1710 2468
rect 1730 2448 1739 2468
rect 1591 2439 1739 2448
rect 1797 2468 1935 2475
rect 1797 2448 1806 2468
rect 1826 2448 1935 2468
rect 1797 2439 1935 2448
rect 1591 2438 1628 2439
rect 1321 2385 1362 2386
rect 130 2365 569 2383
rect 132 2176 184 2365
rect 530 2340 569 2365
rect 1213 2378 1362 2385
rect 1213 2358 1272 2378
rect 1292 2358 1331 2378
rect 1351 2358 1362 2378
rect 1213 2350 1362 2358
rect 1429 2381 1586 2388
rect 1429 2361 1549 2381
rect 1569 2361 1586 2381
rect 1429 2351 1586 2361
rect 1429 2350 1464 2351
rect 314 2315 501 2339
rect 530 2320 925 2340
rect 945 2320 948 2340
rect 1429 2329 1460 2350
rect 1647 2329 1683 2439
rect 1702 2438 1739 2439
rect 1798 2438 1835 2439
rect 1758 2379 1848 2385
rect 1758 2359 1767 2379
rect 1787 2377 1848 2379
rect 1787 2359 1812 2377
rect 1758 2357 1812 2359
rect 1832 2357 1848 2377
rect 1758 2351 1848 2357
rect 1272 2328 1309 2329
rect 530 2315 948 2320
rect 1271 2319 1309 2328
rect 314 2244 351 2315
rect 530 2314 873 2315
rect 530 2311 569 2314
rect 835 2313 872 2314
rect 466 2254 497 2255
rect 314 2224 323 2244
rect 343 2224 351 2244
rect 314 2214 351 2224
rect 410 2244 497 2254
rect 410 2224 419 2244
rect 439 2224 497 2244
rect 410 2215 497 2224
rect 410 2214 447 2215
rect 132 2158 148 2176
rect 166 2158 184 2176
rect 466 2164 497 2215
rect 532 2244 569 2311
rect 1271 2299 1280 2319
rect 1300 2299 1309 2319
rect 1271 2291 1309 2299
rect 1375 2323 1460 2329
rect 1490 2328 1527 2329
rect 1375 2303 1383 2323
rect 1403 2303 1460 2323
rect 1375 2295 1460 2303
rect 1489 2319 1527 2328
rect 1489 2299 1498 2319
rect 1518 2299 1527 2319
rect 1375 2294 1411 2295
rect 1489 2291 1527 2299
rect 1593 2327 1737 2329
rect 1593 2323 1653 2327
rect 1593 2303 1601 2323
rect 1621 2305 1653 2323
rect 1676 2323 1737 2327
rect 1676 2305 1709 2323
rect 1621 2303 1709 2305
rect 1729 2303 1737 2323
rect 1593 2295 1737 2303
rect 1593 2294 1629 2295
rect 1701 2294 1737 2295
rect 1803 2328 1840 2329
rect 1803 2327 1841 2328
rect 1803 2319 1867 2327
rect 1803 2299 1812 2319
rect 1832 2305 1867 2319
rect 1887 2305 1890 2325
rect 1832 2300 1890 2305
rect 1832 2299 1867 2300
rect 1272 2262 1309 2291
rect 1273 2260 1309 2262
rect 684 2254 720 2255
rect 532 2224 541 2244
rect 561 2224 569 2244
rect 532 2214 569 2224
rect 628 2244 776 2254
rect 876 2251 972 2253
rect 628 2224 637 2244
rect 657 2224 747 2244
rect 767 2224 776 2244
rect 628 2215 776 2224
rect 834 2244 972 2251
rect 834 2224 843 2244
rect 863 2224 972 2244
rect 1273 2238 1464 2260
rect 1490 2259 1527 2291
rect 1803 2287 1867 2299
rect 1490 2258 1765 2259
rect 1907 2258 1934 2439
rect 1490 2233 1934 2258
rect 2070 2264 2109 4079
rect 2411 4066 2444 4399
rect 2508 4431 2676 4432
rect 2802 4431 2842 4655
rect 3305 4659 3473 4660
rect 3714 4659 3749 4676
rect 4106 4666 4153 4677
rect 3305 4633 3749 4659
rect 3305 4631 3473 4633
rect 3669 4632 3749 4633
rect 3904 4632 3971 4658
rect 4110 4632 4153 4666
rect 3305 4453 3332 4631
rect 3372 4593 3436 4605
rect 3712 4601 3749 4632
rect 3930 4601 3967 4632
rect 4112 4607 4153 4632
rect 4544 4691 4585 4716
rect 4730 4691 4767 4722
rect 4948 4691 4985 4722
rect 5261 4718 5325 4730
rect 5365 4692 5392 4870
rect 4544 4657 4587 4691
rect 4726 4665 4793 4691
rect 4948 4690 5028 4691
rect 5224 4690 5392 4692
rect 4948 4664 5392 4690
rect 4544 4646 4591 4657
rect 4948 4647 4983 4664
rect 5224 4663 5392 4664
rect 5855 4668 5895 4892
rect 6021 4891 6189 4892
rect 6253 4924 6286 5257
rect 6588 5244 6627 7059
rect 6763 7065 7207 7090
rect 6763 6884 6790 7065
rect 6932 7064 7207 7065
rect 6830 7024 6894 7036
rect 7170 7032 7207 7064
rect 7233 7063 7424 7085
rect 7725 7079 7834 7099
rect 7854 7079 7863 7099
rect 7725 7072 7863 7079
rect 7921 7099 8069 7108
rect 7921 7079 7930 7099
rect 7950 7079 8040 7099
rect 8060 7079 8069 7099
rect 7725 7070 7821 7072
rect 7921 7069 8069 7079
rect 8128 7099 8165 7109
rect 8128 7079 8136 7099
rect 8156 7079 8165 7099
rect 7977 7068 8013 7069
rect 7388 7061 7424 7063
rect 7388 7032 7425 7061
rect 6830 7023 6865 7024
rect 6807 7018 6865 7023
rect 6807 6998 6810 7018
rect 6830 7004 6865 7018
rect 6885 7004 6894 7024
rect 6830 6996 6894 7004
rect 6856 6995 6894 6996
rect 6857 6994 6894 6995
rect 6960 7028 6996 7029
rect 7068 7028 7104 7029
rect 6960 7020 7104 7028
rect 6960 7000 6968 7020
rect 6988 7018 7076 7020
rect 6988 7000 7021 7018
rect 6960 6996 7021 7000
rect 7044 7000 7076 7018
rect 7096 7000 7104 7020
rect 7044 6996 7104 7000
rect 6960 6994 7104 6996
rect 7170 7024 7208 7032
rect 7286 7028 7322 7029
rect 7170 7004 7179 7024
rect 7199 7004 7208 7024
rect 7170 6995 7208 7004
rect 7237 7020 7322 7028
rect 7237 7000 7294 7020
rect 7314 7000 7322 7020
rect 7170 6994 7207 6995
rect 7237 6994 7322 7000
rect 7388 7024 7426 7032
rect 7388 7004 7397 7024
rect 7417 7004 7426 7024
rect 8128 7012 8165 7079
rect 8200 7108 8231 7159
rect 8513 7147 8531 7165
rect 8549 7147 8565 7165
rect 8250 7108 8287 7109
rect 8200 7099 8287 7108
rect 8200 7079 8258 7099
rect 8278 7079 8287 7099
rect 8200 7069 8287 7079
rect 8346 7099 8383 7109
rect 8346 7079 8354 7099
rect 8374 7079 8383 7099
rect 8200 7068 8231 7069
rect 7825 7009 7862 7010
rect 8128 7009 8167 7012
rect 7824 7008 8167 7009
rect 8346 7008 8383 7079
rect 7388 6995 7426 7004
rect 7749 7003 8167 7008
rect 7388 6994 7425 6995
rect 6849 6966 6939 6972
rect 6849 6946 6865 6966
rect 6885 6964 6939 6966
rect 6885 6946 6910 6964
rect 6849 6944 6910 6946
rect 6930 6944 6939 6964
rect 6849 6938 6939 6944
rect 6862 6884 6899 6885
rect 6958 6884 6995 6885
rect 7014 6884 7050 6994
rect 7237 6973 7268 6994
rect 7749 6983 7752 7003
rect 7772 6983 8167 7003
rect 8196 6984 8383 7008
rect 7233 6972 7268 6973
rect 7111 6962 7268 6972
rect 7111 6942 7128 6962
rect 7148 6942 7268 6962
rect 7111 6935 7268 6942
rect 7335 6965 7484 6973
rect 7335 6945 7346 6965
rect 7366 6945 7405 6965
rect 7425 6945 7484 6965
rect 7335 6938 7484 6945
rect 8128 6958 8167 6983
rect 8513 6958 8565 7147
rect 8128 6940 8567 6958
rect 7335 6937 7376 6938
rect 7069 6884 7106 6885
rect 6762 6875 6900 6884
rect 6762 6855 6871 6875
rect 6891 6855 6900 6875
rect 6762 6848 6900 6855
rect 6958 6875 7106 6884
rect 6958 6855 6967 6875
rect 6987 6855 7077 6875
rect 7097 6855 7106 6875
rect 6762 6846 6858 6848
rect 6958 6845 7106 6855
rect 7165 6875 7202 6885
rect 7165 6855 7173 6875
rect 7193 6855 7202 6875
rect 7014 6844 7050 6845
rect 6862 6785 6899 6786
rect 7165 6785 7202 6855
rect 7237 6884 7268 6935
rect 8128 6922 8528 6940
rect 8546 6922 8567 6940
rect 8128 6916 8567 6922
rect 8134 6912 8567 6916
rect 8513 6910 8565 6912
rect 7287 6884 7324 6885
rect 7237 6875 7324 6884
rect 7237 6855 7295 6875
rect 7315 6855 7324 6875
rect 7237 6845 7324 6855
rect 7383 6875 7420 6885
rect 7383 6855 7391 6875
rect 7411 6855 7420 6875
rect 7237 6844 7268 6845
rect 6861 6784 7202 6785
rect 7383 6784 7420 6855
rect 8516 6845 8553 6850
rect 6786 6779 7202 6784
rect 6786 6759 6789 6779
rect 6809 6759 7202 6779
rect 7233 6760 7420 6784
rect 8507 6841 8554 6845
rect 8507 6823 8526 6841
rect 8544 6823 8554 6841
rect 8507 6775 8554 6823
rect 8131 6772 8554 6775
rect 7006 6758 7071 6759
rect 8109 6742 8554 6772
rect 7202 6726 7242 6734
rect 7202 6704 7210 6726
rect 7234 6704 7242 6726
rect 6807 6475 6844 6481
rect 6807 6456 6815 6475
rect 6836 6456 6844 6475
rect 6807 6448 6844 6456
rect 6811 6115 6844 6448
rect 6908 6480 7076 6481
rect 7202 6480 7242 6704
rect 7705 6708 7873 6709
rect 8109 6708 8150 6742
rect 8507 6721 8554 6742
rect 7705 6698 8150 6708
rect 8222 6706 8365 6707
rect 7705 6682 8149 6698
rect 7705 6680 7873 6682
rect 8069 6681 8149 6682
rect 8222 6681 8367 6706
rect 8509 6681 8554 6721
rect 7705 6502 7732 6680
rect 7772 6642 7836 6654
rect 8112 6650 8149 6681
rect 8330 6650 8367 6681
rect 8512 6674 8554 6681
rect 7772 6641 7807 6642
rect 7749 6636 7807 6641
rect 7749 6616 7752 6636
rect 7772 6622 7807 6636
rect 7827 6622 7836 6642
rect 7772 6614 7836 6622
rect 7798 6613 7836 6614
rect 7799 6612 7836 6613
rect 7902 6646 7938 6647
rect 8010 6646 8046 6647
rect 7902 6638 8046 6646
rect 7902 6618 7910 6638
rect 7930 6634 8018 6638
rect 7930 6618 7974 6634
rect 7902 6614 7974 6618
rect 7994 6618 8018 6634
rect 8038 6618 8046 6638
rect 7994 6614 8046 6618
rect 7902 6612 8046 6614
rect 8112 6642 8150 6650
rect 8228 6646 8264 6647
rect 8112 6622 8121 6642
rect 8141 6622 8150 6642
rect 8112 6613 8150 6622
rect 8179 6638 8264 6646
rect 8179 6618 8236 6638
rect 8256 6618 8264 6638
rect 8112 6612 8149 6613
rect 8179 6612 8264 6618
rect 8330 6642 8368 6650
rect 8330 6622 8339 6642
rect 8359 6622 8368 6642
rect 8330 6613 8368 6622
rect 8512 6647 8555 6674
rect 8512 6629 8526 6647
rect 8544 6629 8555 6647
rect 8512 6621 8555 6629
rect 8517 6619 8555 6621
rect 8330 6612 8367 6613
rect 7791 6584 7881 6590
rect 7791 6564 7807 6584
rect 7827 6582 7881 6584
rect 7827 6564 7852 6582
rect 7791 6562 7852 6564
rect 7872 6562 7881 6582
rect 7791 6556 7881 6562
rect 7804 6502 7841 6503
rect 7900 6502 7937 6503
rect 7956 6502 7992 6612
rect 8179 6591 8210 6612
rect 8175 6590 8210 6591
rect 8053 6580 8210 6590
rect 8053 6560 8070 6580
rect 8090 6560 8210 6580
rect 8053 6553 8210 6560
rect 8277 6583 8426 6591
rect 8277 6563 8288 6583
rect 8308 6563 8347 6583
rect 8367 6563 8426 6583
rect 8277 6556 8426 6563
rect 8277 6555 8318 6556
rect 8514 6554 8551 6557
rect 8011 6502 8048 6503
rect 7704 6493 7842 6502
rect 6908 6454 7352 6480
rect 6908 6452 7076 6454
rect 6908 6274 6935 6452
rect 6975 6414 7039 6426
rect 7315 6422 7352 6454
rect 7378 6453 7569 6475
rect 7704 6473 7813 6493
rect 7833 6473 7842 6493
rect 7704 6466 7842 6473
rect 7900 6493 8048 6502
rect 7900 6473 7909 6493
rect 7929 6473 8019 6493
rect 8039 6473 8048 6493
rect 7704 6464 7800 6466
rect 7900 6463 8048 6473
rect 8107 6493 8144 6503
rect 8107 6473 8115 6493
rect 8135 6473 8144 6493
rect 7956 6462 7992 6463
rect 7533 6451 7569 6453
rect 7533 6422 7570 6451
rect 6975 6413 7010 6414
rect 6952 6408 7010 6413
rect 6952 6388 6955 6408
rect 6975 6394 7010 6408
rect 7030 6394 7039 6414
rect 6975 6388 7039 6394
rect 6952 6386 7039 6388
rect 6952 6382 6979 6386
rect 7001 6385 7039 6386
rect 7002 6384 7039 6385
rect 7105 6418 7141 6419
rect 7213 6418 7249 6419
rect 7105 6411 7249 6418
rect 7105 6410 7167 6411
rect 7105 6390 7113 6410
rect 7133 6393 7167 6410
rect 7186 6410 7249 6411
rect 7186 6393 7221 6410
rect 7133 6390 7221 6393
rect 7241 6390 7249 6410
rect 7105 6384 7249 6390
rect 7315 6414 7353 6422
rect 7431 6418 7467 6419
rect 7315 6394 7324 6414
rect 7344 6394 7353 6414
rect 7315 6385 7353 6394
rect 7382 6410 7467 6418
rect 7382 6390 7439 6410
rect 7459 6390 7467 6410
rect 7315 6384 7352 6385
rect 7382 6384 7467 6390
rect 7533 6414 7571 6422
rect 7533 6394 7542 6414
rect 7562 6394 7571 6414
rect 7804 6403 7841 6404
rect 8107 6403 8144 6473
rect 8179 6502 8210 6553
rect 8506 6548 8551 6554
rect 8506 6530 8524 6548
rect 8542 6530 8551 6548
rect 8506 6520 8551 6530
rect 8229 6502 8266 6503
rect 8179 6493 8266 6502
rect 8179 6473 8237 6493
rect 8257 6473 8266 6493
rect 8179 6463 8266 6473
rect 8325 6493 8362 6503
rect 8325 6473 8333 6493
rect 8353 6473 8362 6493
rect 8506 6478 8549 6520
rect 8412 6476 8549 6478
rect 8179 6462 8210 6463
rect 8325 6403 8362 6473
rect 7803 6402 8144 6403
rect 7533 6385 7571 6394
rect 7728 6397 8144 6402
rect 7533 6384 7570 6385
rect 6994 6356 7084 6362
rect 6994 6336 7010 6356
rect 7030 6354 7084 6356
rect 7030 6336 7055 6354
rect 6994 6334 7055 6336
rect 7075 6334 7084 6354
rect 6994 6328 7084 6334
rect 7007 6274 7044 6275
rect 7103 6274 7140 6275
rect 7159 6274 7195 6384
rect 7382 6363 7413 6384
rect 7728 6377 7731 6397
rect 7751 6377 8144 6397
rect 8328 6387 8362 6403
rect 8406 6455 8549 6476
rect 8104 6368 8144 6377
rect 8406 6368 8433 6455
rect 8506 6429 8549 6455
rect 8506 6411 8519 6429
rect 8537 6411 8549 6429
rect 8506 6400 8549 6411
rect 7378 6362 7413 6363
rect 7256 6352 7413 6362
rect 7256 6332 7273 6352
rect 7293 6332 7413 6352
rect 7256 6325 7413 6332
rect 7480 6355 7626 6363
rect 7480 6335 7491 6355
rect 7511 6335 7550 6355
rect 7570 6335 7626 6355
rect 8104 6351 8433 6368
rect 8104 6350 8144 6351
rect 7480 6328 7626 6335
rect 8501 6339 8541 6342
rect 8501 6333 8544 6339
rect 8126 6330 8544 6333
rect 7480 6327 7521 6328
rect 7214 6274 7251 6275
rect 6907 6265 7045 6274
rect 6907 6245 7016 6265
rect 7036 6245 7045 6265
rect 6907 6238 7045 6245
rect 7103 6265 7251 6274
rect 7103 6245 7112 6265
rect 7132 6245 7222 6265
rect 7242 6245 7251 6265
rect 6907 6236 7003 6238
rect 7103 6235 7251 6245
rect 7310 6265 7347 6275
rect 7310 6245 7318 6265
rect 7338 6245 7347 6265
rect 7159 6234 7195 6235
rect 7007 6175 7044 6176
rect 7310 6175 7347 6245
rect 7382 6274 7413 6325
rect 8126 6312 8517 6330
rect 8535 6312 8544 6330
rect 8126 6310 8544 6312
rect 8126 6302 8153 6310
rect 8394 6307 8544 6310
rect 7706 6296 7874 6297
rect 8125 6296 8153 6302
rect 7706 6280 8153 6296
rect 8501 6302 8544 6307
rect 7432 6274 7469 6275
rect 7382 6265 7469 6274
rect 7382 6245 7440 6265
rect 7460 6245 7469 6265
rect 7382 6235 7469 6245
rect 7528 6265 7565 6275
rect 7528 6245 7536 6265
rect 7556 6245 7565 6265
rect 7382 6234 7413 6235
rect 7006 6174 7347 6175
rect 7528 6174 7565 6245
rect 6931 6169 7347 6174
rect 6931 6149 6934 6169
rect 6954 6149 7347 6169
rect 7378 6150 7565 6174
rect 7706 6270 8150 6280
rect 7706 6268 7874 6270
rect 6806 6070 6848 6115
rect 7706 6090 7733 6268
rect 7773 6230 7837 6242
rect 8113 6238 8150 6270
rect 8176 6269 8367 6291
rect 8331 6267 8367 6269
rect 8331 6238 8368 6267
rect 8501 6246 8541 6302
rect 7773 6229 7808 6230
rect 7750 6224 7808 6229
rect 7750 6204 7753 6224
rect 7773 6210 7808 6224
rect 7828 6210 7837 6230
rect 7773 6202 7837 6210
rect 7799 6201 7837 6202
rect 7800 6200 7837 6201
rect 7903 6234 7939 6235
rect 8011 6234 8047 6235
rect 7903 6226 8047 6234
rect 7903 6206 7911 6226
rect 7931 6206 7966 6226
rect 7986 6206 8019 6226
rect 8039 6206 8047 6226
rect 7903 6200 8047 6206
rect 8113 6230 8151 6238
rect 8229 6234 8265 6235
rect 8113 6210 8122 6230
rect 8142 6210 8151 6230
rect 8113 6201 8151 6210
rect 8180 6226 8265 6234
rect 8180 6206 8237 6226
rect 8257 6206 8265 6226
rect 8113 6200 8150 6201
rect 8180 6200 8265 6206
rect 8331 6230 8369 6238
rect 8331 6210 8340 6230
rect 8360 6210 8369 6230
rect 8501 6228 8513 6246
rect 8531 6228 8541 6246
rect 8501 6218 8541 6228
rect 8331 6201 8369 6210
rect 8331 6200 8368 6201
rect 7792 6172 7882 6178
rect 7792 6152 7808 6172
rect 7828 6170 7882 6172
rect 7828 6152 7853 6170
rect 7792 6150 7853 6152
rect 7873 6150 7882 6170
rect 7792 6144 7882 6150
rect 7805 6090 7842 6091
rect 7901 6090 7938 6091
rect 7957 6090 7993 6200
rect 8180 6179 8211 6200
rect 8176 6178 8211 6179
rect 8054 6168 8211 6178
rect 8054 6148 8071 6168
rect 8091 6148 8211 6168
rect 8054 6141 8211 6148
rect 8278 6171 8427 6179
rect 8278 6151 8289 6171
rect 8309 6151 8348 6171
rect 8368 6151 8427 6171
rect 8278 6144 8427 6151
rect 8493 6147 8545 6165
rect 8278 6143 8319 6144
rect 8012 6090 8049 6091
rect 7705 6081 7843 6090
rect 7177 6070 7210 6072
rect 6806 6058 7253 6070
rect 6809 6044 7253 6058
rect 6809 6042 6977 6044
rect 6809 5864 6836 6042
rect 6876 6004 6940 6016
rect 7216 6012 7253 6044
rect 7279 6043 7470 6065
rect 7705 6061 7814 6081
rect 7834 6061 7843 6081
rect 7705 6054 7843 6061
rect 7901 6081 8049 6090
rect 7901 6061 7910 6081
rect 7930 6061 8020 6081
rect 8040 6061 8049 6081
rect 7705 6052 7801 6054
rect 7901 6051 8049 6061
rect 8108 6081 8145 6091
rect 8108 6061 8116 6081
rect 8136 6061 8145 6081
rect 7957 6050 7993 6051
rect 7434 6041 7470 6043
rect 7434 6012 7471 6041
rect 6876 6003 6911 6004
rect 6853 5998 6911 6003
rect 6853 5978 6856 5998
rect 6876 5984 6911 5998
rect 6931 5984 6940 6004
rect 6876 5976 6940 5984
rect 6902 5975 6940 5976
rect 6903 5974 6940 5975
rect 7006 6008 7042 6009
rect 7114 6008 7150 6009
rect 7006 6000 7150 6008
rect 7006 5980 7014 6000
rect 7034 5998 7122 6000
rect 7034 5980 7067 5998
rect 7006 5979 7067 5980
rect 7088 5980 7122 5998
rect 7142 5980 7150 6000
rect 7088 5979 7150 5980
rect 7006 5974 7150 5979
rect 7216 6004 7254 6012
rect 7332 6008 7368 6009
rect 7216 5984 7225 6004
rect 7245 5984 7254 6004
rect 7216 5975 7254 5984
rect 7283 6000 7368 6008
rect 7283 5980 7340 6000
rect 7360 5980 7368 6000
rect 7216 5974 7253 5975
rect 7283 5974 7368 5980
rect 7434 6004 7472 6012
rect 7434 5984 7443 6004
rect 7463 5984 7472 6004
rect 8108 5994 8145 6061
rect 8180 6090 8211 6141
rect 8493 6129 8511 6147
rect 8529 6129 8545 6147
rect 8230 6090 8267 6091
rect 8180 6081 8267 6090
rect 8180 6061 8238 6081
rect 8258 6061 8267 6081
rect 8180 6051 8267 6061
rect 8326 6081 8363 6091
rect 8326 6061 8334 6081
rect 8354 6061 8363 6081
rect 8180 6050 8211 6051
rect 7805 5991 7842 5992
rect 8108 5991 8147 5994
rect 7804 5990 8147 5991
rect 8326 5990 8363 6061
rect 7434 5975 7472 5984
rect 7729 5985 8147 5990
rect 7434 5974 7471 5975
rect 6895 5946 6985 5952
rect 6895 5926 6911 5946
rect 6931 5944 6985 5946
rect 6931 5926 6956 5944
rect 6895 5924 6956 5926
rect 6976 5924 6985 5944
rect 6895 5918 6985 5924
rect 6908 5864 6945 5865
rect 7004 5864 7041 5865
rect 7060 5864 7096 5974
rect 7283 5953 7314 5974
rect 7729 5965 7732 5985
rect 7752 5965 8147 5985
rect 8176 5966 8363 5990
rect 7279 5952 7314 5953
rect 7157 5942 7314 5952
rect 7157 5922 7174 5942
rect 7194 5922 7314 5942
rect 7157 5915 7314 5922
rect 7381 5945 7530 5953
rect 7381 5925 7392 5945
rect 7412 5925 7451 5945
rect 7471 5925 7530 5945
rect 7381 5918 7530 5925
rect 8108 5940 8147 5965
rect 8493 5940 8545 6129
rect 8108 5922 8547 5940
rect 7381 5917 7422 5918
rect 7115 5864 7152 5865
rect 6808 5855 6946 5864
rect 6808 5835 6917 5855
rect 6937 5835 6946 5855
rect 6808 5828 6946 5835
rect 7004 5855 7152 5864
rect 7004 5835 7013 5855
rect 7033 5835 7123 5855
rect 7143 5835 7152 5855
rect 6808 5826 6904 5828
rect 7004 5825 7152 5835
rect 7211 5855 7248 5865
rect 7211 5835 7219 5855
rect 7239 5835 7248 5855
rect 7060 5824 7096 5825
rect 6908 5765 6945 5766
rect 7211 5765 7248 5835
rect 7283 5864 7314 5915
rect 8108 5904 8508 5922
rect 8526 5904 8547 5922
rect 8108 5898 8547 5904
rect 8114 5894 8547 5898
rect 8493 5892 8545 5894
rect 7333 5864 7370 5865
rect 7283 5855 7370 5864
rect 7283 5835 7341 5855
rect 7361 5835 7370 5855
rect 7283 5825 7370 5835
rect 7429 5855 7466 5865
rect 7429 5835 7437 5855
rect 7457 5835 7466 5855
rect 7283 5824 7314 5825
rect 6907 5764 7248 5765
rect 7429 5764 7466 5835
rect 8496 5827 8533 5832
rect 8487 5823 8534 5827
rect 8487 5805 8506 5823
rect 8524 5805 8534 5823
rect 6832 5759 7248 5764
rect 6832 5739 6835 5759
rect 6855 5739 7248 5759
rect 7279 5740 7466 5764
rect 8091 5762 8131 5767
rect 8487 5762 8534 5805
rect 8091 5723 8534 5762
rect 7185 5708 7225 5716
rect 7185 5686 7193 5708
rect 7217 5686 7225 5708
rect 6891 5462 7059 5463
rect 7185 5462 7225 5686
rect 7688 5690 7856 5691
rect 8091 5690 8131 5723
rect 8487 5690 8534 5723
rect 7688 5689 8132 5690
rect 7688 5664 8133 5689
rect 7688 5662 7856 5664
rect 8052 5663 8133 5664
rect 8302 5663 8351 5689
rect 8487 5663 8536 5690
rect 7688 5484 7715 5662
rect 7755 5624 7819 5636
rect 8095 5632 8132 5663
rect 8313 5632 8350 5663
rect 8495 5638 8536 5663
rect 7755 5623 7790 5624
rect 7732 5618 7790 5623
rect 7732 5598 7735 5618
rect 7755 5604 7790 5618
rect 7810 5604 7819 5624
rect 7755 5596 7819 5604
rect 7781 5595 7819 5596
rect 7782 5594 7819 5595
rect 7885 5628 7921 5629
rect 7993 5628 8029 5629
rect 7885 5620 8029 5628
rect 7885 5600 7893 5620
rect 7913 5616 8001 5620
rect 7913 5600 7957 5616
rect 7885 5596 7957 5600
rect 7977 5600 8001 5616
rect 8021 5600 8029 5620
rect 7977 5596 8029 5600
rect 7885 5594 8029 5596
rect 8095 5624 8133 5632
rect 8211 5628 8247 5629
rect 8095 5604 8104 5624
rect 8124 5604 8133 5624
rect 8095 5595 8133 5604
rect 8162 5620 8247 5628
rect 8162 5600 8219 5620
rect 8239 5600 8247 5620
rect 8095 5594 8132 5595
rect 8162 5594 8247 5600
rect 8313 5624 8351 5632
rect 8313 5604 8322 5624
rect 8342 5604 8351 5624
rect 8313 5595 8351 5604
rect 8495 5629 8537 5638
rect 8495 5611 8509 5629
rect 8527 5611 8537 5629
rect 8495 5603 8537 5611
rect 8500 5601 8537 5603
rect 8313 5594 8350 5595
rect 7774 5566 7864 5572
rect 7774 5546 7790 5566
rect 7810 5564 7864 5566
rect 7810 5546 7835 5564
rect 7774 5544 7835 5546
rect 7855 5544 7864 5564
rect 7774 5538 7864 5544
rect 7787 5484 7824 5485
rect 7883 5484 7920 5485
rect 7939 5484 7975 5594
rect 8162 5573 8193 5594
rect 8158 5572 8193 5573
rect 8036 5562 8193 5572
rect 8036 5542 8053 5562
rect 8073 5542 8193 5562
rect 8036 5535 8193 5542
rect 8260 5565 8409 5573
rect 8260 5545 8271 5565
rect 8291 5545 8330 5565
rect 8350 5545 8409 5565
rect 8260 5538 8409 5545
rect 8260 5537 8301 5538
rect 8497 5536 8534 5539
rect 7994 5484 8031 5485
rect 7687 5475 7825 5484
rect 6891 5436 7335 5462
rect 6891 5434 7059 5436
rect 6891 5256 6918 5434
rect 6958 5396 7022 5408
rect 7298 5404 7335 5436
rect 7361 5435 7552 5457
rect 7687 5455 7796 5475
rect 7816 5455 7825 5475
rect 7687 5448 7825 5455
rect 7883 5475 8031 5484
rect 7883 5455 7892 5475
rect 7912 5455 8002 5475
rect 8022 5455 8031 5475
rect 7687 5446 7783 5448
rect 7883 5445 8031 5455
rect 8090 5475 8127 5485
rect 8090 5455 8098 5475
rect 8118 5455 8127 5475
rect 7939 5444 7975 5445
rect 7516 5433 7552 5435
rect 7516 5404 7553 5433
rect 6958 5395 6993 5396
rect 6935 5390 6993 5395
rect 6935 5370 6938 5390
rect 6958 5376 6993 5390
rect 7013 5376 7022 5396
rect 6958 5368 7022 5376
rect 6984 5367 7022 5368
rect 6985 5366 7022 5367
rect 7088 5400 7124 5401
rect 7196 5400 7232 5401
rect 7088 5392 7232 5400
rect 7088 5372 7096 5392
rect 7116 5391 7204 5392
rect 7116 5372 7151 5391
rect 7172 5372 7204 5391
rect 7224 5372 7232 5392
rect 7088 5366 7232 5372
rect 7298 5396 7336 5404
rect 7414 5400 7450 5401
rect 7298 5376 7307 5396
rect 7327 5376 7336 5396
rect 7298 5367 7336 5376
rect 7365 5392 7450 5400
rect 7365 5372 7422 5392
rect 7442 5372 7450 5392
rect 7298 5366 7335 5367
rect 7365 5366 7450 5372
rect 7516 5396 7554 5404
rect 7516 5376 7525 5396
rect 7545 5376 7554 5396
rect 7787 5385 7824 5386
rect 8090 5385 8127 5455
rect 8162 5484 8193 5535
rect 8489 5530 8534 5536
rect 8489 5512 8507 5530
rect 8525 5512 8534 5530
rect 8489 5502 8534 5512
rect 8212 5484 8249 5485
rect 8162 5475 8249 5484
rect 8162 5455 8220 5475
rect 8240 5455 8249 5475
rect 8162 5445 8249 5455
rect 8308 5475 8345 5485
rect 8308 5455 8316 5475
rect 8336 5455 8345 5475
rect 8489 5460 8532 5502
rect 8395 5458 8532 5460
rect 8162 5444 8193 5445
rect 8308 5385 8345 5455
rect 7786 5384 8127 5385
rect 7516 5367 7554 5376
rect 7711 5379 8127 5384
rect 7516 5366 7553 5367
rect 6977 5338 7067 5344
rect 6977 5318 6993 5338
rect 7013 5336 7067 5338
rect 7013 5318 7038 5336
rect 6977 5316 7038 5318
rect 7058 5316 7067 5336
rect 6977 5310 7067 5316
rect 6990 5256 7027 5257
rect 7086 5256 7123 5257
rect 7142 5256 7178 5366
rect 7365 5345 7396 5366
rect 7711 5359 7714 5379
rect 7734 5359 8127 5379
rect 8311 5369 8345 5385
rect 8389 5437 8532 5458
rect 8087 5350 8127 5359
rect 8389 5350 8416 5437
rect 8489 5411 8532 5437
rect 8489 5393 8502 5411
rect 8520 5393 8532 5411
rect 8489 5382 8532 5393
rect 7361 5344 7396 5345
rect 7239 5334 7396 5344
rect 7239 5314 7256 5334
rect 7276 5314 7396 5334
rect 7239 5307 7396 5314
rect 7463 5337 7612 5345
rect 7463 5317 7474 5337
rect 7494 5317 7533 5337
rect 7553 5317 7612 5337
rect 8087 5333 8416 5350
rect 8087 5332 8127 5333
rect 7463 5310 7612 5317
rect 8484 5321 8524 5324
rect 8484 5315 8527 5321
rect 8109 5312 8527 5315
rect 7463 5309 7504 5310
rect 7197 5256 7234 5257
rect 6890 5247 7028 5256
rect 6588 5072 6628 5244
rect 6890 5227 6999 5247
rect 7019 5227 7028 5247
rect 6890 5220 7028 5227
rect 7086 5247 7234 5256
rect 7086 5227 7095 5247
rect 7115 5227 7205 5247
rect 7225 5227 7234 5247
rect 6890 5218 6986 5220
rect 7086 5217 7234 5227
rect 7293 5247 7330 5257
rect 7293 5227 7301 5247
rect 7321 5227 7330 5247
rect 7142 5216 7178 5217
rect 6990 5157 7027 5158
rect 7293 5157 7330 5227
rect 7365 5256 7396 5307
rect 8109 5294 8500 5312
rect 8518 5294 8527 5312
rect 8109 5292 8527 5294
rect 8109 5284 8136 5292
rect 8377 5289 8527 5292
rect 7689 5278 7857 5279
rect 8108 5278 8136 5284
rect 7689 5262 8136 5278
rect 8484 5284 8527 5289
rect 7415 5256 7452 5257
rect 7365 5247 7452 5256
rect 7365 5227 7423 5247
rect 7443 5227 7452 5247
rect 7365 5217 7452 5227
rect 7511 5247 7548 5257
rect 7511 5227 7519 5247
rect 7539 5227 7548 5247
rect 7365 5216 7396 5217
rect 6989 5156 7330 5157
rect 7511 5156 7548 5227
rect 6914 5151 7330 5156
rect 6914 5131 6917 5151
rect 6937 5131 7330 5151
rect 7361 5132 7548 5156
rect 7689 5252 8133 5262
rect 7689 5250 7857 5252
rect 7689 5072 7716 5250
rect 7756 5212 7820 5224
rect 8096 5220 8133 5252
rect 8159 5251 8350 5273
rect 8314 5249 8350 5251
rect 8314 5220 8351 5249
rect 8484 5228 8524 5284
rect 7756 5211 7791 5212
rect 7733 5206 7791 5211
rect 7733 5186 7736 5206
rect 7756 5192 7791 5206
rect 7811 5192 7820 5212
rect 7756 5184 7820 5192
rect 7782 5183 7820 5184
rect 7783 5182 7820 5183
rect 7886 5216 7922 5217
rect 7994 5216 8030 5217
rect 7886 5208 8030 5216
rect 7886 5188 7894 5208
rect 7914 5188 7949 5208
rect 7969 5188 8002 5208
rect 8022 5188 8030 5208
rect 7886 5182 8030 5188
rect 8096 5212 8134 5220
rect 8212 5216 8248 5217
rect 8096 5192 8105 5212
rect 8125 5192 8134 5212
rect 8096 5183 8134 5192
rect 8163 5208 8248 5216
rect 8163 5188 8220 5208
rect 8240 5188 8248 5208
rect 8096 5182 8133 5183
rect 8163 5182 8248 5188
rect 8314 5212 8352 5220
rect 8314 5192 8323 5212
rect 8343 5192 8352 5212
rect 8484 5210 8496 5228
rect 8514 5210 8524 5228
rect 8484 5200 8524 5210
rect 8314 5183 8352 5192
rect 8314 5182 8351 5183
rect 7775 5154 7865 5160
rect 7775 5134 7791 5154
rect 7811 5152 7865 5154
rect 7811 5134 7836 5152
rect 7775 5132 7836 5134
rect 7856 5132 7865 5152
rect 7775 5126 7865 5132
rect 7788 5072 7825 5073
rect 7884 5072 7921 5073
rect 7940 5072 7976 5182
rect 8163 5161 8194 5182
rect 8159 5160 8194 5161
rect 8037 5150 8194 5160
rect 8037 5130 8054 5150
rect 8074 5130 8194 5150
rect 8037 5123 8194 5130
rect 8261 5153 8410 5161
rect 8261 5133 8272 5153
rect 8292 5133 8331 5153
rect 8351 5133 8410 5153
rect 8261 5126 8410 5133
rect 8476 5129 8528 5147
rect 8261 5125 8302 5126
rect 7995 5072 8032 5073
rect 6589 5057 6628 5072
rect 7688 5063 7826 5072
rect 6589 5056 6755 5057
rect 6881 5056 6921 5058
rect 6589 5030 7031 5056
rect 6589 5028 6755 5030
rect 6253 4916 6290 4924
rect 6253 4897 6261 4916
rect 6282 4897 6290 4916
rect 6253 4891 6290 4897
rect 6589 4850 6614 5028
rect 6654 4990 6718 5002
rect 6994 4998 7031 5030
rect 7057 5029 7248 5051
rect 7688 5043 7797 5063
rect 7817 5043 7826 5063
rect 7688 5036 7826 5043
rect 7884 5063 8032 5072
rect 7884 5043 7893 5063
rect 7913 5043 8003 5063
rect 8023 5043 8032 5063
rect 7688 5034 7784 5036
rect 7884 5033 8032 5043
rect 8091 5063 8128 5073
rect 8091 5043 8099 5063
rect 8119 5043 8128 5063
rect 7940 5032 7976 5033
rect 7212 5027 7248 5029
rect 7212 4998 7249 5027
rect 6654 4989 6689 4990
rect 6631 4984 6689 4989
rect 6631 4964 6634 4984
rect 6654 4970 6689 4984
rect 6709 4970 6718 4990
rect 6654 4962 6718 4970
rect 6680 4961 6718 4962
rect 6681 4960 6718 4961
rect 6784 4994 6820 4995
rect 6892 4994 6928 4995
rect 6784 4989 6928 4994
rect 6784 4986 6846 4989
rect 6784 4966 6792 4986
rect 6812 4966 6846 4986
rect 6784 4963 6846 4966
rect 6872 4986 6928 4989
rect 6872 4966 6900 4986
rect 6920 4966 6928 4986
rect 6872 4963 6928 4966
rect 6784 4960 6928 4963
rect 6994 4990 7032 4998
rect 7110 4994 7146 4995
rect 6994 4970 7003 4990
rect 7023 4970 7032 4990
rect 6994 4961 7032 4970
rect 7061 4986 7146 4994
rect 7061 4966 7118 4986
rect 7138 4966 7146 4986
rect 6994 4960 7031 4961
rect 7061 4960 7146 4966
rect 7212 4990 7250 4998
rect 7212 4970 7221 4990
rect 7241 4970 7250 4990
rect 8091 4976 8128 5043
rect 8163 5072 8194 5123
rect 8476 5111 8494 5129
rect 8512 5111 8528 5129
rect 8213 5072 8250 5073
rect 8163 5063 8250 5072
rect 8163 5043 8221 5063
rect 8241 5043 8250 5063
rect 8163 5033 8250 5043
rect 8309 5063 8346 5073
rect 8309 5043 8317 5063
rect 8337 5043 8346 5063
rect 8163 5032 8194 5033
rect 7788 4973 7825 4974
rect 8091 4973 8130 4976
rect 7787 4972 8130 4973
rect 8309 4972 8346 5043
rect 7212 4961 7250 4970
rect 7712 4967 8130 4972
rect 7212 4960 7249 4961
rect 6673 4932 6763 4938
rect 6673 4912 6689 4932
rect 6709 4930 6763 4932
rect 6709 4912 6734 4930
rect 6673 4910 6734 4912
rect 6754 4910 6763 4930
rect 6673 4904 6763 4910
rect 6686 4850 6723 4851
rect 6782 4850 6819 4851
rect 6838 4850 6874 4960
rect 7061 4939 7092 4960
rect 7712 4947 7715 4967
rect 7735 4947 8130 4967
rect 8159 4948 8346 4972
rect 7057 4938 7092 4939
rect 6935 4928 7092 4938
rect 6935 4908 6952 4928
rect 6972 4908 7092 4928
rect 6935 4901 7092 4908
rect 7159 4931 7308 4939
rect 7159 4911 7170 4931
rect 7190 4911 7229 4931
rect 7249 4911 7308 4931
rect 7159 4904 7308 4911
rect 8091 4922 8130 4947
rect 8476 4922 8528 5111
rect 8091 4904 8530 4922
rect 7159 4903 7200 4904
rect 6893 4850 6930 4851
rect 6589 4841 6724 4850
rect 6589 4821 6695 4841
rect 6715 4821 6724 4841
rect 6589 4814 6724 4821
rect 6782 4841 6930 4850
rect 6782 4821 6791 4841
rect 6811 4821 6901 4841
rect 6921 4821 6930 4841
rect 6589 4812 6682 4814
rect 6782 4811 6930 4821
rect 6989 4841 7026 4851
rect 6989 4821 6997 4841
rect 7017 4821 7026 4841
rect 6838 4810 6874 4811
rect 6686 4751 6723 4752
rect 6989 4751 7026 4821
rect 7061 4850 7092 4901
rect 8091 4886 8491 4904
rect 8509 4886 8530 4904
rect 8091 4880 8530 4886
rect 8097 4876 8530 4880
rect 8476 4874 8528 4876
rect 7111 4850 7148 4851
rect 7061 4841 7148 4850
rect 7061 4821 7119 4841
rect 7139 4821 7148 4841
rect 7061 4811 7148 4821
rect 7207 4841 7244 4851
rect 7207 4821 7215 4841
rect 7235 4821 7244 4841
rect 7061 4810 7092 4811
rect 6685 4750 7026 4751
rect 7207 4750 7244 4821
rect 8479 4809 8516 4814
rect 6610 4745 7026 4750
rect 6610 4725 6613 4745
rect 6633 4725 7026 4745
rect 7057 4726 7244 4750
rect 8470 4805 8517 4809
rect 8470 4787 8489 4805
rect 8507 4787 8517 4805
rect 8078 4728 8116 4729
rect 8470 4728 8517 4787
rect 6830 4724 6895 4725
rect 4945 4646 4983 4647
rect 4544 4608 4983 4646
rect 5855 4646 5863 4668
rect 5887 4646 5895 4668
rect 5855 4638 5895 4646
rect 7166 4690 7206 4698
rect 7166 4668 7174 4690
rect 7198 4668 7206 4690
rect 8078 4690 8517 4728
rect 8078 4689 8116 4690
rect 6166 4611 6231 4612
rect 3372 4592 3407 4593
rect 3349 4587 3407 4592
rect 3349 4567 3352 4587
rect 3372 4573 3407 4587
rect 3427 4573 3436 4593
rect 3372 4565 3436 4573
rect 3398 4564 3436 4565
rect 3399 4563 3436 4564
rect 3502 4597 3538 4598
rect 3610 4597 3646 4598
rect 3502 4589 3646 4597
rect 3502 4569 3510 4589
rect 3530 4585 3618 4589
rect 3530 4569 3574 4585
rect 3502 4565 3574 4569
rect 3594 4569 3618 4585
rect 3638 4569 3646 4589
rect 3594 4565 3646 4569
rect 3502 4563 3646 4565
rect 3712 4593 3750 4601
rect 3828 4597 3864 4598
rect 3712 4573 3721 4593
rect 3741 4573 3750 4593
rect 3712 4564 3750 4573
rect 3779 4589 3864 4597
rect 3779 4569 3836 4589
rect 3856 4569 3864 4589
rect 3712 4563 3749 4564
rect 3779 4563 3864 4569
rect 3930 4593 3968 4601
rect 3930 4573 3939 4593
rect 3959 4573 3968 4593
rect 3930 4564 3968 4573
rect 4112 4598 4154 4607
rect 4112 4580 4126 4598
rect 4144 4580 4154 4598
rect 4112 4572 4154 4580
rect 4117 4570 4154 4572
rect 3930 4563 3967 4564
rect 3391 4535 3481 4541
rect 3391 4515 3407 4535
rect 3427 4533 3481 4535
rect 3427 4515 3452 4533
rect 3391 4513 3452 4515
rect 3472 4513 3481 4533
rect 3391 4507 3481 4513
rect 3404 4453 3441 4454
rect 3500 4453 3537 4454
rect 3556 4453 3592 4563
rect 3779 4542 3810 4563
rect 4544 4549 4591 4608
rect 4945 4607 4983 4608
rect 3775 4541 3810 4542
rect 3653 4531 3810 4541
rect 3653 4511 3670 4531
rect 3690 4511 3810 4531
rect 3653 4504 3810 4511
rect 3877 4534 4026 4542
rect 3877 4514 3888 4534
rect 3908 4514 3947 4534
rect 3967 4514 4026 4534
rect 4544 4531 4554 4549
rect 4572 4531 4591 4549
rect 4544 4527 4591 4531
rect 5817 4586 6004 4610
rect 6035 4591 6428 4611
rect 6448 4591 6451 4611
rect 6035 4586 6451 4591
rect 4545 4522 4582 4527
rect 3877 4507 4026 4514
rect 5817 4515 5854 4586
rect 6035 4585 6376 4586
rect 5969 4525 6000 4526
rect 3877 4506 3918 4507
rect 4114 4505 4151 4508
rect 3611 4453 3648 4454
rect 3304 4444 3442 4453
rect 2508 4405 2952 4431
rect 2508 4403 2676 4405
rect 2508 4225 2535 4403
rect 2575 4365 2639 4377
rect 2915 4373 2952 4405
rect 2978 4404 3169 4426
rect 3304 4424 3413 4444
rect 3433 4424 3442 4444
rect 3304 4417 3442 4424
rect 3500 4444 3648 4453
rect 3500 4424 3509 4444
rect 3529 4424 3619 4444
rect 3639 4424 3648 4444
rect 3304 4415 3400 4417
rect 3500 4414 3648 4424
rect 3707 4444 3744 4454
rect 3707 4424 3715 4444
rect 3735 4424 3744 4444
rect 3556 4413 3592 4414
rect 3133 4402 3169 4404
rect 3133 4373 3170 4402
rect 2575 4364 2610 4365
rect 2552 4359 2610 4364
rect 2552 4339 2555 4359
rect 2575 4345 2610 4359
rect 2630 4345 2639 4365
rect 2575 4339 2639 4345
rect 2552 4337 2639 4339
rect 2552 4333 2579 4337
rect 2601 4336 2639 4337
rect 2602 4335 2639 4336
rect 2705 4369 2741 4370
rect 2813 4369 2849 4370
rect 2705 4362 2849 4369
rect 2705 4361 2767 4362
rect 2705 4341 2713 4361
rect 2733 4344 2767 4361
rect 2786 4361 2849 4362
rect 2786 4344 2821 4361
rect 2733 4341 2821 4344
rect 2841 4341 2849 4361
rect 2705 4335 2849 4341
rect 2915 4365 2953 4373
rect 3031 4369 3067 4370
rect 2915 4345 2924 4365
rect 2944 4345 2953 4365
rect 2915 4336 2953 4345
rect 2982 4361 3067 4369
rect 2982 4341 3039 4361
rect 3059 4341 3067 4361
rect 2915 4335 2952 4336
rect 2982 4335 3067 4341
rect 3133 4365 3171 4373
rect 3133 4345 3142 4365
rect 3162 4345 3171 4365
rect 3404 4354 3441 4355
rect 3707 4354 3744 4424
rect 3779 4453 3810 4504
rect 4106 4499 4151 4505
rect 4106 4481 4124 4499
rect 4142 4481 4151 4499
rect 5817 4495 5826 4515
rect 5846 4495 5854 4515
rect 5817 4485 5854 4495
rect 5913 4515 6000 4525
rect 5913 4495 5922 4515
rect 5942 4495 6000 4515
rect 5913 4486 6000 4495
rect 5913 4485 5950 4486
rect 4106 4471 4151 4481
rect 3829 4453 3866 4454
rect 3779 4444 3866 4453
rect 3779 4424 3837 4444
rect 3857 4424 3866 4444
rect 3779 4414 3866 4424
rect 3925 4444 3962 4454
rect 3925 4424 3933 4444
rect 3953 4424 3962 4444
rect 4106 4429 4149 4471
rect 4533 4460 4585 4462
rect 4012 4427 4149 4429
rect 3779 4413 3810 4414
rect 3925 4354 3962 4424
rect 3403 4353 3744 4354
rect 3133 4336 3171 4345
rect 3328 4348 3744 4353
rect 3133 4335 3170 4336
rect 2594 4307 2684 4313
rect 2594 4287 2610 4307
rect 2630 4305 2684 4307
rect 2630 4287 2655 4305
rect 2594 4285 2655 4287
rect 2675 4285 2684 4305
rect 2594 4279 2684 4285
rect 2607 4225 2644 4226
rect 2703 4225 2740 4226
rect 2759 4225 2795 4335
rect 2982 4314 3013 4335
rect 3328 4328 3331 4348
rect 3351 4328 3744 4348
rect 3928 4338 3962 4354
rect 4006 4406 4149 4427
rect 4531 4456 4964 4460
rect 4531 4450 4970 4456
rect 4531 4432 4552 4450
rect 4570 4432 4970 4450
rect 5969 4435 6000 4486
rect 6035 4515 6072 4585
rect 6338 4584 6375 4585
rect 6187 4525 6223 4526
rect 6035 4495 6044 4515
rect 6064 4495 6072 4515
rect 6035 4485 6072 4495
rect 6131 4515 6279 4525
rect 6379 4522 6475 4524
rect 6131 4495 6140 4515
rect 6160 4495 6250 4515
rect 6270 4495 6279 4515
rect 6131 4486 6279 4495
rect 6337 4515 6475 4522
rect 6337 4495 6346 4515
rect 6366 4495 6475 4515
rect 6337 4486 6475 4495
rect 6131 4485 6168 4486
rect 5861 4432 5902 4433
rect 4531 4414 4970 4432
rect 3704 4319 3744 4328
rect 4006 4319 4033 4406
rect 4106 4380 4149 4406
rect 4106 4362 4119 4380
rect 4137 4362 4149 4380
rect 4106 4351 4149 4362
rect 2978 4313 3013 4314
rect 2856 4303 3013 4313
rect 2856 4283 2873 4303
rect 2893 4283 3013 4303
rect 2856 4276 3013 4283
rect 3080 4306 3226 4314
rect 3080 4286 3091 4306
rect 3111 4286 3150 4306
rect 3170 4286 3226 4306
rect 3704 4302 4033 4319
rect 3704 4301 3744 4302
rect 3080 4279 3226 4286
rect 4101 4290 4141 4293
rect 4101 4284 4144 4290
rect 3726 4281 4144 4284
rect 3080 4278 3121 4279
rect 2814 4225 2851 4226
rect 2507 4216 2645 4225
rect 2507 4196 2616 4216
rect 2636 4196 2645 4216
rect 2507 4189 2645 4196
rect 2703 4216 2851 4225
rect 2703 4196 2712 4216
rect 2732 4196 2822 4216
rect 2842 4196 2851 4216
rect 2507 4187 2603 4189
rect 2703 4186 2851 4196
rect 2910 4216 2947 4226
rect 2910 4196 2918 4216
rect 2938 4196 2947 4216
rect 2759 4185 2795 4186
rect 2607 4126 2644 4127
rect 2910 4126 2947 4196
rect 2982 4225 3013 4276
rect 3726 4263 4117 4281
rect 4135 4263 4144 4281
rect 3726 4261 4144 4263
rect 3726 4253 3753 4261
rect 3994 4258 4144 4261
rect 3306 4247 3474 4248
rect 3725 4247 3753 4253
rect 3306 4231 3753 4247
rect 4101 4253 4144 4258
rect 3032 4225 3069 4226
rect 2982 4216 3069 4225
rect 2982 4196 3040 4216
rect 3060 4196 3069 4216
rect 2982 4186 3069 4196
rect 3128 4216 3165 4226
rect 3128 4196 3136 4216
rect 3156 4196 3165 4216
rect 2982 4185 3013 4186
rect 2606 4125 2947 4126
rect 3128 4125 3165 4196
rect 2531 4120 2947 4125
rect 2531 4100 2534 4120
rect 2554 4100 2947 4120
rect 2978 4101 3165 4125
rect 3306 4221 3750 4231
rect 3306 4219 3474 4221
rect 2340 4026 2384 4027
rect 2340 4020 2385 4026
rect 2340 4002 2352 4020
rect 2374 4002 2385 4020
rect 2406 4021 2448 4066
rect 3306 4041 3333 4219
rect 3373 4181 3437 4193
rect 3713 4189 3750 4221
rect 3776 4220 3967 4242
rect 3931 4218 3967 4220
rect 3931 4189 3968 4218
rect 4101 4197 4141 4253
rect 3373 4180 3408 4181
rect 3350 4175 3408 4180
rect 3350 4155 3353 4175
rect 3373 4161 3408 4175
rect 3428 4161 3437 4181
rect 3373 4153 3437 4161
rect 3399 4152 3437 4153
rect 3400 4151 3437 4152
rect 3503 4185 3539 4186
rect 3611 4185 3647 4186
rect 3503 4177 3647 4185
rect 3503 4157 3511 4177
rect 3531 4157 3566 4177
rect 3586 4157 3619 4177
rect 3639 4157 3647 4177
rect 3503 4151 3647 4157
rect 3713 4181 3751 4189
rect 3829 4185 3865 4186
rect 3713 4161 3722 4181
rect 3742 4161 3751 4181
rect 3713 4152 3751 4161
rect 3780 4177 3865 4185
rect 3780 4157 3837 4177
rect 3857 4157 3865 4177
rect 3713 4151 3750 4152
rect 3780 4151 3865 4157
rect 3931 4181 3969 4189
rect 3931 4161 3940 4181
rect 3960 4161 3969 4181
rect 4101 4179 4113 4197
rect 4131 4179 4141 4197
rect 4533 4225 4585 4414
rect 4931 4389 4970 4414
rect 5753 4425 5902 4432
rect 5753 4405 5812 4425
rect 5832 4405 5871 4425
rect 5891 4405 5902 4425
rect 5753 4397 5902 4405
rect 5969 4428 6126 4435
rect 5969 4408 6089 4428
rect 6109 4408 6126 4428
rect 5969 4398 6126 4408
rect 5969 4397 6004 4398
rect 4715 4364 4902 4388
rect 4931 4369 5326 4389
rect 5346 4369 5349 4389
rect 5969 4376 6000 4397
rect 6187 4376 6223 4486
rect 6242 4485 6279 4486
rect 6338 4485 6375 4486
rect 6298 4426 6388 4432
rect 6298 4406 6307 4426
rect 6327 4424 6388 4426
rect 6327 4406 6352 4424
rect 6298 4404 6352 4406
rect 6372 4404 6388 4424
rect 6298 4398 6388 4404
rect 5812 4375 5849 4376
rect 4931 4364 5349 4369
rect 5811 4366 5849 4375
rect 4715 4293 4752 4364
rect 4931 4363 5274 4364
rect 4931 4360 4970 4363
rect 5236 4362 5273 4363
rect 4867 4303 4898 4304
rect 4715 4273 4724 4293
rect 4744 4273 4752 4293
rect 4715 4263 4752 4273
rect 4811 4293 4898 4303
rect 4811 4273 4820 4293
rect 4840 4273 4898 4293
rect 4811 4264 4898 4273
rect 4811 4263 4848 4264
rect 4533 4207 4549 4225
rect 4567 4207 4585 4225
rect 4867 4213 4898 4264
rect 4933 4293 4970 4360
rect 5811 4346 5820 4366
rect 5840 4346 5849 4366
rect 5811 4338 5849 4346
rect 5915 4370 6000 4376
rect 6030 4375 6067 4376
rect 5915 4350 5923 4370
rect 5943 4350 6000 4370
rect 5915 4342 6000 4350
rect 6029 4366 6067 4375
rect 6029 4346 6038 4366
rect 6058 4346 6067 4366
rect 5915 4341 5951 4342
rect 6029 4338 6067 4346
rect 6133 4370 6277 4376
rect 6133 4350 6141 4370
rect 6161 4364 6249 4370
rect 6161 4350 6190 4364
rect 6133 4342 6190 4350
rect 6133 4341 6169 4342
rect 6213 4350 6249 4364
rect 6269 4350 6277 4370
rect 6213 4342 6277 4350
rect 6241 4341 6277 4342
rect 6343 4375 6380 4376
rect 6343 4374 6381 4375
rect 6343 4366 6407 4374
rect 6343 4346 6352 4366
rect 6372 4352 6407 4366
rect 6427 4352 6430 4372
rect 6372 4347 6430 4352
rect 6372 4346 6407 4347
rect 5812 4309 5849 4338
rect 5813 4307 5849 4309
rect 5085 4303 5121 4304
rect 4933 4273 4942 4293
rect 4962 4273 4970 4293
rect 4933 4263 4970 4273
rect 5029 4293 5177 4303
rect 5277 4300 5373 4302
rect 5029 4273 5038 4293
rect 5058 4273 5148 4293
rect 5168 4273 5177 4293
rect 5029 4264 5177 4273
rect 5235 4293 5373 4300
rect 5235 4273 5244 4293
rect 5264 4273 5373 4293
rect 5813 4285 6004 4307
rect 6030 4306 6067 4338
rect 6343 4334 6407 4346
rect 6447 4308 6474 4486
rect 6771 4439 6808 4445
rect 6771 4420 6779 4439
rect 6800 4420 6808 4439
rect 6771 4412 6808 4420
rect 6306 4306 6474 4308
rect 6030 4280 6474 4306
rect 6140 4278 6180 4280
rect 6306 4279 6474 4280
rect 5235 4264 5373 4273
rect 6433 4274 6474 4279
rect 5029 4263 5066 4264
rect 4759 4210 4800 4211
rect 4533 4189 4585 4207
rect 4651 4203 4800 4210
rect 4101 4169 4141 4179
rect 4651 4183 4710 4203
rect 4730 4183 4769 4203
rect 4789 4183 4800 4203
rect 4651 4175 4800 4183
rect 4867 4206 5024 4213
rect 4867 4186 4987 4206
rect 5007 4186 5024 4206
rect 4867 4176 5024 4186
rect 4867 4175 4902 4176
rect 3931 4152 3969 4161
rect 4867 4154 4898 4175
rect 5085 4154 5121 4264
rect 5140 4263 5177 4264
rect 5236 4263 5273 4264
rect 5196 4204 5286 4210
rect 5196 4184 5205 4204
rect 5225 4202 5286 4204
rect 5225 4184 5250 4202
rect 5196 4182 5250 4184
rect 5270 4182 5286 4202
rect 5196 4176 5286 4182
rect 4710 4153 4747 4154
rect 3931 4151 3968 4152
rect 3392 4123 3482 4129
rect 3392 4103 3408 4123
rect 3428 4121 3482 4123
rect 3428 4103 3453 4121
rect 3392 4101 3453 4103
rect 3473 4101 3482 4121
rect 3392 4095 3482 4101
rect 3405 4041 3442 4042
rect 3501 4041 3538 4042
rect 3557 4041 3593 4151
rect 3780 4130 3811 4151
rect 4709 4144 4747 4153
rect 3776 4129 3811 4130
rect 3654 4119 3811 4129
rect 3654 4099 3671 4119
rect 3691 4099 3811 4119
rect 3654 4092 3811 4099
rect 3878 4122 4027 4130
rect 3878 4102 3889 4122
rect 3909 4102 3948 4122
rect 3968 4102 4027 4122
rect 4537 4126 4577 4136
rect 3878 4095 4027 4102
rect 4093 4098 4145 4116
rect 3878 4094 3919 4095
rect 3612 4041 3649 4042
rect 3305 4032 3443 4041
rect 2777 4021 2810 4023
rect 2406 4009 2853 4021
rect 2340 3972 2385 4002
rect 2357 3026 2385 3972
rect 2409 3995 2853 4009
rect 2409 3993 2577 3995
rect 2409 3815 2436 3993
rect 2476 3955 2540 3967
rect 2816 3963 2853 3995
rect 2879 3994 3070 4016
rect 3305 4012 3414 4032
rect 3434 4012 3443 4032
rect 3305 4005 3443 4012
rect 3501 4032 3649 4041
rect 3501 4012 3510 4032
rect 3530 4012 3620 4032
rect 3640 4012 3649 4032
rect 3305 4003 3401 4005
rect 3501 4002 3649 4012
rect 3708 4032 3745 4042
rect 3708 4012 3716 4032
rect 3736 4012 3745 4032
rect 3557 4001 3593 4002
rect 3034 3992 3070 3994
rect 3034 3963 3071 3992
rect 2476 3954 2511 3955
rect 2453 3949 2511 3954
rect 2453 3929 2456 3949
rect 2476 3935 2511 3949
rect 2531 3935 2540 3955
rect 2476 3927 2540 3935
rect 2502 3926 2540 3927
rect 2503 3925 2540 3926
rect 2606 3959 2642 3960
rect 2714 3959 2750 3960
rect 2606 3953 2750 3959
rect 2606 3951 2667 3953
rect 2606 3931 2614 3951
rect 2634 3936 2667 3951
rect 2686 3951 2750 3953
rect 2686 3936 2722 3951
rect 2634 3931 2722 3936
rect 2742 3931 2750 3951
rect 2606 3925 2750 3931
rect 2816 3955 2854 3963
rect 2932 3959 2968 3960
rect 2816 3935 2825 3955
rect 2845 3935 2854 3955
rect 2816 3926 2854 3935
rect 2883 3951 2968 3959
rect 2883 3931 2940 3951
rect 2960 3931 2968 3951
rect 2816 3925 2853 3926
rect 2883 3925 2968 3931
rect 3034 3955 3072 3963
rect 3034 3935 3043 3955
rect 3063 3935 3072 3955
rect 3708 3945 3745 4012
rect 3780 4041 3811 4092
rect 4093 4080 4111 4098
rect 4129 4080 4145 4098
rect 3830 4041 3867 4042
rect 3780 4032 3867 4041
rect 3780 4012 3838 4032
rect 3858 4012 3867 4032
rect 3780 4002 3867 4012
rect 3926 4032 3963 4042
rect 3926 4012 3934 4032
rect 3954 4012 3963 4032
rect 3780 4001 3811 4002
rect 3405 3942 3442 3943
rect 3708 3942 3747 3945
rect 3404 3941 3747 3942
rect 3926 3941 3963 4012
rect 3034 3926 3072 3935
rect 3329 3936 3747 3941
rect 3034 3925 3071 3926
rect 2495 3897 2585 3903
rect 2495 3877 2511 3897
rect 2531 3895 2585 3897
rect 2531 3877 2556 3895
rect 2495 3875 2556 3877
rect 2576 3875 2585 3895
rect 2495 3869 2585 3875
rect 2508 3815 2545 3816
rect 2604 3815 2641 3816
rect 2660 3815 2696 3925
rect 2883 3904 2914 3925
rect 3329 3916 3332 3936
rect 3352 3916 3747 3936
rect 3776 3917 3963 3941
rect 2879 3903 2914 3904
rect 2757 3893 2914 3903
rect 2757 3873 2774 3893
rect 2794 3873 2914 3893
rect 2757 3866 2914 3873
rect 2981 3896 3130 3904
rect 2981 3876 2992 3896
rect 3012 3876 3051 3896
rect 3071 3876 3130 3896
rect 2981 3869 3130 3876
rect 3708 3891 3747 3916
rect 4093 3891 4145 4080
rect 4537 4108 4547 4126
rect 4565 4108 4577 4126
rect 4709 4124 4718 4144
rect 4738 4124 4747 4144
rect 4709 4116 4747 4124
rect 4813 4148 4898 4154
rect 4928 4153 4965 4154
rect 4813 4128 4821 4148
rect 4841 4128 4898 4148
rect 4813 4120 4898 4128
rect 4927 4144 4965 4153
rect 4927 4124 4936 4144
rect 4956 4124 4965 4144
rect 4813 4119 4849 4120
rect 4927 4116 4965 4124
rect 5031 4148 5175 4154
rect 5031 4128 5039 4148
rect 5059 4128 5092 4148
rect 5112 4128 5147 4148
rect 5167 4128 5175 4148
rect 5031 4120 5175 4128
rect 5031 4119 5067 4120
rect 5139 4119 5175 4120
rect 5241 4153 5278 4154
rect 5241 4152 5279 4153
rect 5241 4144 5305 4152
rect 5241 4124 5250 4144
rect 5270 4130 5305 4144
rect 5325 4130 5328 4150
rect 5270 4125 5328 4130
rect 5270 4124 5305 4125
rect 4537 4052 4577 4108
rect 4710 4087 4747 4116
rect 4711 4085 4747 4087
rect 4711 4063 4902 4085
rect 4928 4084 4965 4116
rect 5241 4112 5305 4124
rect 5345 4086 5372 4264
rect 5204 4084 5372 4086
rect 4928 4074 5372 4084
rect 5513 4180 5700 4204
rect 5731 4185 6124 4205
rect 6144 4185 6147 4205
rect 5731 4180 6147 4185
rect 5513 4109 5550 4180
rect 5731 4179 6072 4180
rect 5665 4119 5696 4120
rect 5513 4089 5522 4109
rect 5542 4089 5550 4109
rect 5513 4079 5550 4089
rect 5609 4109 5696 4119
rect 5609 4089 5618 4109
rect 5638 4089 5696 4109
rect 5609 4080 5696 4089
rect 5609 4079 5646 4080
rect 4534 4047 4577 4052
rect 4925 4058 5372 4074
rect 4925 4052 4953 4058
rect 5204 4057 5372 4058
rect 4534 4044 4684 4047
rect 4925 4044 4952 4052
rect 4534 4042 4952 4044
rect 4534 4024 4543 4042
rect 4561 4024 4952 4042
rect 5665 4029 5696 4080
rect 5731 4109 5768 4179
rect 6034 4178 6071 4179
rect 5883 4119 5919 4120
rect 5731 4089 5740 4109
rect 5760 4089 5768 4109
rect 5731 4079 5768 4089
rect 5827 4109 5975 4119
rect 6075 4116 6171 4118
rect 5827 4089 5836 4109
rect 5856 4089 5946 4109
rect 5966 4089 5975 4109
rect 5827 4080 5975 4089
rect 6033 4109 6171 4116
rect 6033 4089 6042 4109
rect 6062 4089 6171 4109
rect 6433 4092 6473 4274
rect 6033 4080 6171 4089
rect 5827 4079 5864 4080
rect 5557 4026 5598 4027
rect 4534 4021 4952 4024
rect 4534 4015 4577 4021
rect 4537 4012 4577 4015
rect 5449 4019 5598 4026
rect 4934 4003 4974 4004
rect 4645 3986 4974 4003
rect 5449 3999 5508 4019
rect 5528 3999 5567 4019
rect 5587 3999 5598 4019
rect 5449 3991 5598 3999
rect 5665 4022 5822 4029
rect 5665 4002 5785 4022
rect 5805 4002 5822 4022
rect 5665 3992 5822 4002
rect 5665 3991 5700 3992
rect 4529 3943 4572 3954
rect 4529 3925 4541 3943
rect 4559 3925 4572 3943
rect 4529 3899 4572 3925
rect 4645 3899 4672 3986
rect 4934 3977 4974 3986
rect 3708 3873 4147 3891
rect 2981 3868 3022 3869
rect 2715 3815 2752 3816
rect 2408 3806 2546 3815
rect 2408 3786 2517 3806
rect 2537 3786 2546 3806
rect 2408 3779 2546 3786
rect 2604 3806 2752 3815
rect 2604 3786 2613 3806
rect 2633 3786 2723 3806
rect 2743 3786 2752 3806
rect 2408 3777 2504 3779
rect 2604 3776 2752 3786
rect 2811 3806 2848 3816
rect 2811 3786 2819 3806
rect 2839 3786 2848 3806
rect 2660 3775 2696 3776
rect 2508 3716 2545 3717
rect 2811 3716 2848 3786
rect 2883 3815 2914 3866
rect 3708 3855 4108 3873
rect 4126 3855 4147 3873
rect 3708 3849 4147 3855
rect 3714 3845 4147 3849
rect 4529 3878 4672 3899
rect 4716 3951 4750 3967
rect 4934 3957 5327 3977
rect 5347 3957 5350 3977
rect 5665 3970 5696 3991
rect 5883 3970 5919 4080
rect 5938 4079 5975 4080
rect 6034 4079 6071 4080
rect 5994 4020 6084 4026
rect 5994 4000 6003 4020
rect 6023 4018 6084 4020
rect 6023 4000 6048 4018
rect 5994 3998 6048 4000
rect 6068 3998 6084 4018
rect 5994 3992 6084 3998
rect 5508 3969 5545 3970
rect 4934 3952 5350 3957
rect 5507 3960 5545 3969
rect 4934 3951 5275 3952
rect 4716 3881 4753 3951
rect 4868 3891 4899 3892
rect 4529 3876 4666 3878
rect 4093 3843 4145 3845
rect 4529 3834 4572 3876
rect 4716 3861 4725 3881
rect 4745 3861 4753 3881
rect 4716 3851 4753 3861
rect 4812 3881 4899 3891
rect 4812 3861 4821 3881
rect 4841 3861 4899 3881
rect 4812 3852 4899 3861
rect 4812 3851 4849 3852
rect 4527 3824 4572 3834
rect 2933 3815 2970 3816
rect 2883 3806 2970 3815
rect 2883 3786 2941 3806
rect 2961 3786 2970 3806
rect 2883 3776 2970 3786
rect 3029 3806 3066 3816
rect 3029 3786 3037 3806
rect 3057 3786 3066 3806
rect 4527 3806 4536 3824
rect 4554 3806 4572 3824
rect 4527 3800 4572 3806
rect 4868 3801 4899 3852
rect 4934 3881 4971 3951
rect 5237 3950 5274 3951
rect 5507 3940 5516 3960
rect 5536 3940 5545 3960
rect 5507 3932 5545 3940
rect 5611 3964 5696 3970
rect 5726 3969 5763 3970
rect 5611 3944 5619 3964
rect 5639 3944 5696 3964
rect 5611 3936 5696 3944
rect 5725 3960 5763 3969
rect 5725 3940 5734 3960
rect 5754 3940 5763 3960
rect 5611 3935 5647 3936
rect 5725 3932 5763 3940
rect 5829 3964 5973 3970
rect 5829 3944 5837 3964
rect 5857 3945 5889 3964
rect 5910 3945 5945 3964
rect 5857 3944 5945 3945
rect 5965 3944 5973 3964
rect 5829 3936 5973 3944
rect 5829 3935 5865 3936
rect 5937 3935 5973 3936
rect 6039 3969 6076 3970
rect 6039 3968 6077 3969
rect 6039 3960 6103 3968
rect 6039 3940 6048 3960
rect 6068 3946 6103 3960
rect 6123 3946 6126 3966
rect 6068 3941 6126 3946
rect 6068 3940 6103 3941
rect 5508 3903 5545 3932
rect 5509 3901 5545 3903
rect 5086 3891 5122 3892
rect 4934 3861 4943 3881
rect 4963 3861 4971 3881
rect 4934 3851 4971 3861
rect 5030 3881 5178 3891
rect 5278 3888 5374 3890
rect 5030 3861 5039 3881
rect 5059 3861 5149 3881
rect 5169 3861 5178 3881
rect 5030 3852 5178 3861
rect 5236 3881 5374 3888
rect 5236 3861 5245 3881
rect 5265 3861 5374 3881
rect 5509 3879 5700 3901
rect 5726 3900 5763 3932
rect 6039 3928 6103 3940
rect 6143 3902 6170 4080
rect 6002 3900 6170 3902
rect 5726 3874 6170 3900
rect 5236 3852 5374 3861
rect 5030 3851 5067 3852
rect 4527 3797 4564 3800
rect 4760 3798 4801 3799
rect 2883 3775 2914 3776
rect 2507 3715 2848 3716
rect 3029 3715 3066 3786
rect 4652 3791 4801 3798
rect 4096 3778 4133 3783
rect 4087 3774 4134 3778
rect 4087 3756 4106 3774
rect 4124 3756 4134 3774
rect 4652 3771 4711 3791
rect 4731 3771 4770 3791
rect 4790 3771 4801 3791
rect 4652 3763 4801 3771
rect 4868 3794 5025 3801
rect 4868 3774 4988 3794
rect 5008 3774 5025 3794
rect 4868 3764 5025 3774
rect 4868 3763 4903 3764
rect 2432 3710 2848 3715
rect 2432 3690 2435 3710
rect 2455 3690 2848 3710
rect 2879 3691 3066 3715
rect 3691 3713 3731 3718
rect 4087 3713 4134 3756
rect 4868 3742 4899 3763
rect 5086 3742 5122 3852
rect 5141 3851 5178 3852
rect 5237 3851 5274 3852
rect 5197 3792 5287 3798
rect 5197 3772 5206 3792
rect 5226 3790 5287 3792
rect 5226 3772 5251 3790
rect 5197 3770 5251 3772
rect 5271 3770 5287 3790
rect 5197 3764 5287 3770
rect 4711 3741 4748 3742
rect 3691 3674 4134 3713
rect 4524 3733 4561 3735
rect 4524 3725 4566 3733
rect 4524 3707 4534 3725
rect 4552 3707 4566 3725
rect 4524 3698 4566 3707
rect 4710 3732 4748 3741
rect 4710 3712 4719 3732
rect 4739 3712 4748 3732
rect 4710 3704 4748 3712
rect 4814 3736 4899 3742
rect 4929 3741 4966 3742
rect 4814 3716 4822 3736
rect 4842 3716 4899 3736
rect 4814 3708 4899 3716
rect 4928 3732 4966 3741
rect 4928 3712 4937 3732
rect 4957 3712 4966 3732
rect 4814 3707 4850 3708
rect 4928 3704 4966 3712
rect 5032 3740 5176 3742
rect 5032 3736 5084 3740
rect 5032 3716 5040 3736
rect 5060 3720 5084 3736
rect 5104 3736 5176 3740
rect 5104 3720 5148 3736
rect 5060 3716 5148 3720
rect 5168 3716 5176 3736
rect 5032 3708 5176 3716
rect 5032 3707 5068 3708
rect 5140 3707 5176 3708
rect 5242 3741 5279 3742
rect 5242 3740 5280 3741
rect 5242 3732 5306 3740
rect 5242 3712 5251 3732
rect 5271 3718 5306 3732
rect 5326 3718 5329 3738
rect 5271 3713 5329 3718
rect 5271 3712 5306 3713
rect 2785 3659 2825 3667
rect 2785 3637 2793 3659
rect 2817 3637 2825 3659
rect 2491 3413 2659 3414
rect 2785 3413 2825 3637
rect 3288 3641 3456 3642
rect 3691 3641 3731 3674
rect 4087 3641 4134 3674
rect 4525 3673 4566 3698
rect 4711 3673 4748 3704
rect 4929 3673 4966 3704
rect 5242 3700 5306 3712
rect 5346 3674 5373 3852
rect 4525 3646 4574 3673
rect 4710 3647 4759 3673
rect 4928 3672 5009 3673
rect 5205 3672 5373 3674
rect 4928 3647 5373 3672
rect 4929 3646 5373 3647
rect 3288 3640 3732 3641
rect 3288 3615 3733 3640
rect 3288 3613 3456 3615
rect 3652 3614 3733 3615
rect 3902 3614 3951 3640
rect 4087 3614 4136 3641
rect 3288 3435 3315 3613
rect 3355 3575 3419 3587
rect 3695 3583 3732 3614
rect 3913 3583 3950 3614
rect 4095 3589 4136 3614
rect 4527 3613 4574 3646
rect 4930 3613 4970 3646
rect 5205 3645 5373 3646
rect 5836 3650 5876 3874
rect 6002 3873 6170 3874
rect 5836 3628 5844 3650
rect 5868 3628 5876 3650
rect 5836 3620 5876 3628
rect 3355 3574 3390 3575
rect 3332 3569 3390 3574
rect 3332 3549 3335 3569
rect 3355 3555 3390 3569
rect 3410 3555 3419 3575
rect 3355 3547 3419 3555
rect 3381 3546 3419 3547
rect 3382 3545 3419 3546
rect 3485 3579 3521 3580
rect 3593 3579 3629 3580
rect 3485 3571 3629 3579
rect 3485 3551 3493 3571
rect 3513 3567 3601 3571
rect 3513 3551 3557 3567
rect 3485 3547 3557 3551
rect 3577 3551 3601 3567
rect 3621 3551 3629 3571
rect 3577 3547 3629 3551
rect 3485 3545 3629 3547
rect 3695 3575 3733 3583
rect 3811 3579 3847 3580
rect 3695 3555 3704 3575
rect 3724 3555 3733 3575
rect 3695 3546 3733 3555
rect 3762 3571 3847 3579
rect 3762 3551 3819 3571
rect 3839 3551 3847 3571
rect 3695 3545 3732 3546
rect 3762 3545 3847 3551
rect 3913 3575 3951 3583
rect 3913 3555 3922 3575
rect 3942 3555 3951 3575
rect 3913 3546 3951 3555
rect 4095 3580 4137 3589
rect 4095 3562 4109 3580
rect 4127 3562 4137 3580
rect 4095 3554 4137 3562
rect 4100 3552 4137 3554
rect 4527 3574 4970 3613
rect 3913 3545 3950 3546
rect 3374 3517 3464 3523
rect 3374 3497 3390 3517
rect 3410 3515 3464 3517
rect 3410 3497 3435 3515
rect 3374 3495 3435 3497
rect 3455 3495 3464 3515
rect 3374 3489 3464 3495
rect 3387 3435 3424 3436
rect 3483 3435 3520 3436
rect 3539 3435 3575 3545
rect 3762 3524 3793 3545
rect 4527 3531 4574 3574
rect 4930 3569 4970 3574
rect 5595 3572 5782 3596
rect 5813 3577 6206 3597
rect 6226 3577 6229 3597
rect 5813 3572 6229 3577
rect 3758 3523 3793 3524
rect 3636 3513 3793 3523
rect 3636 3493 3653 3513
rect 3673 3493 3793 3513
rect 3636 3486 3793 3493
rect 3860 3516 4009 3524
rect 3860 3496 3871 3516
rect 3891 3496 3930 3516
rect 3950 3496 4009 3516
rect 4527 3513 4537 3531
rect 4555 3513 4574 3531
rect 4527 3509 4574 3513
rect 4528 3504 4565 3509
rect 3860 3489 4009 3496
rect 5595 3501 5632 3572
rect 5813 3571 6154 3572
rect 5747 3511 5778 3512
rect 3860 3488 3901 3489
rect 4097 3487 4134 3490
rect 3594 3435 3631 3436
rect 3287 3426 3425 3435
rect 2491 3387 2935 3413
rect 2491 3385 2659 3387
rect 2491 3207 2518 3385
rect 2558 3347 2622 3359
rect 2898 3355 2935 3387
rect 2961 3386 3152 3408
rect 3287 3406 3396 3426
rect 3416 3406 3425 3426
rect 3287 3399 3425 3406
rect 3483 3426 3631 3435
rect 3483 3406 3492 3426
rect 3512 3406 3602 3426
rect 3622 3406 3631 3426
rect 3287 3397 3383 3399
rect 3483 3396 3631 3406
rect 3690 3426 3727 3436
rect 3690 3406 3698 3426
rect 3718 3406 3727 3426
rect 3539 3395 3575 3396
rect 3116 3384 3152 3386
rect 3116 3355 3153 3384
rect 2558 3346 2593 3347
rect 2535 3341 2593 3346
rect 2535 3321 2538 3341
rect 2558 3327 2593 3341
rect 2613 3327 2622 3347
rect 2558 3319 2622 3327
rect 2584 3318 2622 3319
rect 2585 3317 2622 3318
rect 2688 3351 2724 3352
rect 2796 3351 2832 3352
rect 2688 3343 2832 3351
rect 2688 3323 2696 3343
rect 2716 3342 2804 3343
rect 2716 3323 2751 3342
rect 2772 3323 2804 3342
rect 2824 3323 2832 3343
rect 2688 3317 2832 3323
rect 2898 3347 2936 3355
rect 3014 3351 3050 3352
rect 2898 3327 2907 3347
rect 2927 3327 2936 3347
rect 2898 3318 2936 3327
rect 2965 3343 3050 3351
rect 2965 3323 3022 3343
rect 3042 3323 3050 3343
rect 2898 3317 2935 3318
rect 2965 3317 3050 3323
rect 3116 3347 3154 3355
rect 3116 3327 3125 3347
rect 3145 3327 3154 3347
rect 3387 3336 3424 3337
rect 3690 3336 3727 3406
rect 3762 3435 3793 3486
rect 4089 3481 4134 3487
rect 4089 3463 4107 3481
rect 4125 3463 4134 3481
rect 5595 3481 5604 3501
rect 5624 3481 5632 3501
rect 5595 3471 5632 3481
rect 5691 3501 5778 3511
rect 5691 3481 5700 3501
rect 5720 3481 5778 3501
rect 5691 3472 5778 3481
rect 5691 3471 5728 3472
rect 4089 3453 4134 3463
rect 3812 3435 3849 3436
rect 3762 3426 3849 3435
rect 3762 3406 3820 3426
rect 3840 3406 3849 3426
rect 3762 3396 3849 3406
rect 3908 3426 3945 3436
rect 3908 3406 3916 3426
rect 3936 3406 3945 3426
rect 4089 3411 4132 3453
rect 4516 3442 4568 3444
rect 3995 3409 4132 3411
rect 3762 3395 3793 3396
rect 3908 3336 3945 3406
rect 3386 3335 3727 3336
rect 3116 3318 3154 3327
rect 3311 3330 3727 3335
rect 3116 3317 3153 3318
rect 2577 3289 2667 3295
rect 2577 3269 2593 3289
rect 2613 3287 2667 3289
rect 2613 3269 2638 3287
rect 2577 3267 2638 3269
rect 2658 3267 2667 3287
rect 2577 3261 2667 3267
rect 2590 3207 2627 3208
rect 2686 3207 2723 3208
rect 2742 3207 2778 3317
rect 2965 3296 2996 3317
rect 3311 3310 3314 3330
rect 3334 3310 3727 3330
rect 3911 3320 3945 3336
rect 3989 3388 4132 3409
rect 4514 3438 4947 3442
rect 4514 3432 4953 3438
rect 4514 3414 4535 3432
rect 4553 3414 4953 3432
rect 5747 3421 5778 3472
rect 5813 3501 5850 3571
rect 6116 3570 6153 3571
rect 5965 3511 6001 3512
rect 5813 3481 5822 3501
rect 5842 3481 5850 3501
rect 5813 3471 5850 3481
rect 5909 3501 6057 3511
rect 6157 3508 6253 3510
rect 5909 3481 5918 3501
rect 5938 3481 6028 3501
rect 6048 3481 6057 3501
rect 5909 3472 6057 3481
rect 6115 3501 6253 3508
rect 6115 3481 6124 3501
rect 6144 3481 6253 3501
rect 6115 3472 6253 3481
rect 5909 3471 5946 3472
rect 5639 3418 5680 3419
rect 4514 3396 4953 3414
rect 3687 3301 3727 3310
rect 3989 3301 4016 3388
rect 4089 3362 4132 3388
rect 4089 3344 4102 3362
rect 4120 3344 4132 3362
rect 4089 3333 4132 3344
rect 2961 3295 2996 3296
rect 2839 3285 2996 3295
rect 2839 3265 2856 3285
rect 2876 3265 2996 3285
rect 2839 3258 2996 3265
rect 3063 3288 3212 3296
rect 3063 3268 3074 3288
rect 3094 3268 3133 3288
rect 3153 3268 3212 3288
rect 3687 3284 4016 3301
rect 3687 3283 3727 3284
rect 3063 3261 3212 3268
rect 4084 3272 4124 3275
rect 4084 3266 4127 3272
rect 3709 3263 4127 3266
rect 3063 3260 3104 3261
rect 2797 3207 2834 3208
rect 2490 3198 2628 3207
rect 2490 3178 2599 3198
rect 2619 3178 2628 3198
rect 2490 3171 2628 3178
rect 2686 3198 2834 3207
rect 2686 3178 2695 3198
rect 2715 3178 2805 3198
rect 2825 3178 2834 3198
rect 2490 3169 2586 3171
rect 2686 3168 2834 3178
rect 2893 3198 2930 3208
rect 2893 3178 2901 3198
rect 2921 3178 2930 3198
rect 2742 3167 2778 3168
rect 2590 3108 2627 3109
rect 2893 3108 2930 3178
rect 2965 3207 2996 3258
rect 3709 3245 4100 3263
rect 4118 3245 4127 3263
rect 3709 3243 4127 3245
rect 3709 3235 3736 3243
rect 3977 3240 4127 3243
rect 3289 3229 3457 3230
rect 3708 3229 3736 3235
rect 3289 3213 3736 3229
rect 4084 3235 4127 3240
rect 3015 3207 3052 3208
rect 2965 3198 3052 3207
rect 2965 3178 3023 3198
rect 3043 3178 3052 3198
rect 2965 3168 3052 3178
rect 3111 3198 3148 3208
rect 3111 3178 3119 3198
rect 3139 3178 3148 3198
rect 2965 3167 2996 3168
rect 2589 3107 2930 3108
rect 3111 3107 3148 3178
rect 2514 3102 2930 3107
rect 2514 3082 2517 3102
rect 2537 3082 2930 3102
rect 2961 3083 3148 3107
rect 3289 3203 3733 3213
rect 3289 3201 3457 3203
rect 2356 3008 2385 3026
rect 3289 3023 3316 3201
rect 3356 3163 3420 3175
rect 3696 3171 3733 3203
rect 3759 3202 3950 3224
rect 3914 3200 3950 3202
rect 3914 3171 3951 3200
rect 4084 3179 4124 3235
rect 3356 3162 3391 3163
rect 3333 3157 3391 3162
rect 3333 3137 3336 3157
rect 3356 3143 3391 3157
rect 3411 3143 3420 3163
rect 3356 3135 3420 3143
rect 3382 3134 3420 3135
rect 3383 3133 3420 3134
rect 3486 3167 3522 3168
rect 3594 3167 3630 3168
rect 3486 3159 3630 3167
rect 3486 3139 3494 3159
rect 3514 3139 3549 3159
rect 3569 3139 3602 3159
rect 3622 3139 3630 3159
rect 3486 3133 3630 3139
rect 3696 3163 3734 3171
rect 3812 3167 3848 3168
rect 3696 3143 3705 3163
rect 3725 3143 3734 3163
rect 3696 3134 3734 3143
rect 3763 3159 3848 3167
rect 3763 3139 3820 3159
rect 3840 3139 3848 3159
rect 3696 3133 3733 3134
rect 3763 3133 3848 3139
rect 3914 3163 3952 3171
rect 3914 3143 3923 3163
rect 3943 3143 3952 3163
rect 4084 3161 4096 3179
rect 4114 3161 4124 3179
rect 4516 3207 4568 3396
rect 4914 3371 4953 3396
rect 5531 3411 5680 3418
rect 5531 3391 5590 3411
rect 5610 3391 5649 3411
rect 5669 3391 5680 3411
rect 5531 3383 5680 3391
rect 5747 3414 5904 3421
rect 5747 3394 5867 3414
rect 5887 3394 5904 3414
rect 5747 3384 5904 3394
rect 5747 3383 5782 3384
rect 4698 3346 4885 3370
rect 4914 3351 5309 3371
rect 5329 3351 5332 3371
rect 5747 3362 5778 3383
rect 5965 3362 6001 3472
rect 6020 3471 6057 3472
rect 6116 3471 6153 3472
rect 6076 3412 6166 3418
rect 6076 3392 6085 3412
rect 6105 3410 6166 3412
rect 6105 3392 6130 3410
rect 6076 3390 6130 3392
rect 6150 3390 6166 3410
rect 6076 3384 6166 3390
rect 5590 3361 5627 3362
rect 4914 3346 5332 3351
rect 5589 3352 5627 3361
rect 4698 3275 4735 3346
rect 4914 3345 5257 3346
rect 4914 3342 4953 3345
rect 5219 3344 5256 3345
rect 4850 3285 4881 3286
rect 4698 3255 4707 3275
rect 4727 3255 4735 3275
rect 4698 3245 4735 3255
rect 4794 3275 4881 3285
rect 4794 3255 4803 3275
rect 4823 3255 4881 3275
rect 4794 3246 4881 3255
rect 4794 3245 4831 3246
rect 4516 3189 4532 3207
rect 4550 3189 4568 3207
rect 4850 3195 4881 3246
rect 4916 3275 4953 3342
rect 5589 3332 5598 3352
rect 5618 3332 5627 3352
rect 5589 3324 5627 3332
rect 5693 3356 5778 3362
rect 5808 3361 5845 3362
rect 5693 3336 5701 3356
rect 5721 3336 5778 3356
rect 5693 3328 5778 3336
rect 5807 3352 5845 3361
rect 5807 3332 5816 3352
rect 5836 3332 5845 3352
rect 5693 3327 5729 3328
rect 5807 3324 5845 3332
rect 5911 3357 6055 3362
rect 5911 3356 5973 3357
rect 5911 3336 5919 3356
rect 5939 3338 5973 3356
rect 5994 3356 6055 3357
rect 5994 3338 6027 3356
rect 5939 3336 6027 3338
rect 6047 3336 6055 3356
rect 5911 3328 6055 3336
rect 5911 3327 5947 3328
rect 6019 3327 6055 3328
rect 6121 3361 6158 3362
rect 6121 3360 6159 3361
rect 6121 3352 6185 3360
rect 6121 3332 6130 3352
rect 6150 3338 6185 3352
rect 6205 3338 6208 3358
rect 6150 3333 6208 3338
rect 6150 3332 6185 3333
rect 5590 3295 5627 3324
rect 5591 3293 5627 3295
rect 5068 3285 5104 3286
rect 4916 3255 4925 3275
rect 4945 3255 4953 3275
rect 4916 3245 4953 3255
rect 5012 3275 5160 3285
rect 5260 3282 5356 3284
rect 5012 3255 5021 3275
rect 5041 3255 5131 3275
rect 5151 3255 5160 3275
rect 5012 3246 5160 3255
rect 5218 3275 5356 3282
rect 5218 3255 5227 3275
rect 5247 3255 5356 3275
rect 5591 3271 5782 3293
rect 5808 3292 5845 3324
rect 6121 3320 6185 3332
rect 6225 3294 6252 3472
rect 6084 3292 6252 3294
rect 5808 3278 6252 3292
rect 5808 3266 6255 3278
rect 5851 3264 5884 3266
rect 5218 3246 5356 3255
rect 5012 3245 5049 3246
rect 4742 3192 4783 3193
rect 4516 3171 4568 3189
rect 4634 3185 4783 3192
rect 4084 3151 4124 3161
rect 4634 3165 4693 3185
rect 4713 3165 4752 3185
rect 4772 3165 4783 3185
rect 4634 3157 4783 3165
rect 4850 3188 5007 3195
rect 4850 3168 4970 3188
rect 4990 3168 5007 3188
rect 4850 3158 5007 3168
rect 4850 3157 4885 3158
rect 3914 3134 3952 3143
rect 4850 3136 4881 3157
rect 5068 3136 5104 3246
rect 5123 3245 5160 3246
rect 5219 3245 5256 3246
rect 5179 3186 5269 3192
rect 5179 3166 5188 3186
rect 5208 3184 5269 3186
rect 5208 3166 5233 3184
rect 5179 3164 5233 3166
rect 5253 3164 5269 3184
rect 5179 3158 5269 3164
rect 4693 3135 4730 3136
rect 3914 3133 3951 3134
rect 3375 3105 3465 3111
rect 3375 3085 3391 3105
rect 3411 3103 3465 3105
rect 3411 3085 3436 3103
rect 3375 3083 3436 3085
rect 3456 3083 3465 3103
rect 3375 3077 3465 3083
rect 3388 3023 3425 3024
rect 3484 3023 3521 3024
rect 3540 3023 3576 3133
rect 3763 3112 3794 3133
rect 4692 3126 4730 3135
rect 3759 3111 3794 3112
rect 3637 3101 3794 3111
rect 3637 3081 3654 3101
rect 3674 3081 3794 3101
rect 3637 3074 3794 3081
rect 3861 3104 4010 3112
rect 3861 3084 3872 3104
rect 3892 3084 3931 3104
rect 3951 3084 4010 3104
rect 4520 3108 4560 3118
rect 3861 3077 4010 3084
rect 4076 3080 4128 3098
rect 3861 3076 3902 3077
rect 3595 3023 3632 3024
rect 2326 3006 2385 3008
rect 3288 3014 3426 3023
rect 2326 3005 2494 3006
rect 2620 3005 2660 3007
rect 2326 2979 2770 3005
rect 2326 2977 2494 2979
rect 2326 2975 2407 2977
rect 2326 2799 2353 2975
rect 2393 2939 2457 2951
rect 2733 2947 2770 2979
rect 2796 2978 2987 3000
rect 3288 2994 3397 3014
rect 3417 2994 3426 3014
rect 3288 2987 3426 2994
rect 3484 3014 3632 3023
rect 3484 2994 3493 3014
rect 3513 2994 3603 3014
rect 3623 2994 3632 3014
rect 3288 2985 3384 2987
rect 3484 2984 3632 2994
rect 3691 3014 3728 3024
rect 3691 2994 3699 3014
rect 3719 2994 3728 3014
rect 3540 2983 3576 2984
rect 2951 2976 2987 2978
rect 2951 2947 2988 2976
rect 2393 2938 2428 2939
rect 2370 2933 2428 2938
rect 2370 2913 2373 2933
rect 2393 2919 2428 2933
rect 2448 2919 2457 2939
rect 2393 2911 2457 2919
rect 2419 2910 2457 2911
rect 2420 2909 2457 2910
rect 2523 2943 2559 2944
rect 2631 2943 2667 2944
rect 2523 2935 2667 2943
rect 2523 2915 2531 2935
rect 2551 2934 2639 2935
rect 2551 2916 2586 2934
rect 2604 2916 2639 2934
rect 2551 2915 2639 2916
rect 2659 2915 2667 2935
rect 2523 2909 2667 2915
rect 2733 2939 2771 2947
rect 2849 2943 2885 2944
rect 2733 2919 2742 2939
rect 2762 2919 2771 2939
rect 2733 2910 2771 2919
rect 2800 2935 2885 2943
rect 2800 2915 2857 2935
rect 2877 2915 2885 2935
rect 2733 2909 2770 2910
rect 2800 2909 2885 2915
rect 2951 2939 2989 2947
rect 2951 2919 2960 2939
rect 2980 2919 2989 2939
rect 3691 2927 3728 2994
rect 3763 3023 3794 3074
rect 4076 3062 4094 3080
rect 4112 3062 4128 3080
rect 3813 3023 3850 3024
rect 3763 3014 3850 3023
rect 3763 2994 3821 3014
rect 3841 2994 3850 3014
rect 3763 2984 3850 2994
rect 3909 3014 3946 3024
rect 3909 2994 3917 3014
rect 3937 2994 3946 3014
rect 3763 2983 3794 2984
rect 3388 2924 3425 2925
rect 3691 2924 3730 2927
rect 3387 2923 3730 2924
rect 3909 2923 3946 2994
rect 2951 2910 2989 2919
rect 3312 2918 3730 2923
rect 2951 2909 2988 2910
rect 2412 2881 2502 2887
rect 2412 2861 2428 2881
rect 2448 2879 2502 2881
rect 2448 2861 2473 2879
rect 2412 2859 2473 2861
rect 2493 2859 2502 2879
rect 2412 2853 2502 2859
rect 2425 2799 2462 2800
rect 2521 2799 2558 2800
rect 2577 2799 2613 2909
rect 2800 2888 2831 2909
rect 3312 2898 3315 2918
rect 3335 2898 3730 2918
rect 3759 2899 3946 2923
rect 2796 2887 2831 2888
rect 2674 2877 2831 2887
rect 2674 2857 2691 2877
rect 2711 2857 2831 2877
rect 2674 2850 2831 2857
rect 2898 2880 3047 2888
rect 2898 2860 2909 2880
rect 2929 2860 2968 2880
rect 2988 2860 3047 2880
rect 2898 2853 3047 2860
rect 3691 2873 3730 2898
rect 4076 2873 4128 3062
rect 4520 3090 4530 3108
rect 4548 3090 4560 3108
rect 4692 3106 4701 3126
rect 4721 3106 4730 3126
rect 4692 3098 4730 3106
rect 4796 3130 4881 3136
rect 4911 3135 4948 3136
rect 4796 3110 4804 3130
rect 4824 3110 4881 3130
rect 4796 3102 4881 3110
rect 4910 3126 4948 3135
rect 4910 3106 4919 3126
rect 4939 3106 4948 3126
rect 4796 3101 4832 3102
rect 4910 3098 4948 3106
rect 5014 3130 5158 3136
rect 5014 3110 5022 3130
rect 5042 3110 5075 3130
rect 5095 3110 5130 3130
rect 5150 3110 5158 3130
rect 5014 3102 5158 3110
rect 5014 3101 5050 3102
rect 5122 3101 5158 3102
rect 5224 3135 5261 3136
rect 5224 3134 5262 3135
rect 5224 3126 5288 3134
rect 5224 3106 5233 3126
rect 5253 3112 5288 3126
rect 5308 3112 5311 3132
rect 5253 3107 5311 3112
rect 5253 3106 5288 3107
rect 4520 3034 4560 3090
rect 4693 3069 4730 3098
rect 4694 3067 4730 3069
rect 4694 3045 4885 3067
rect 4911 3066 4948 3098
rect 5224 3094 5288 3106
rect 5328 3068 5355 3246
rect 6213 3221 6255 3266
rect 5187 3066 5355 3068
rect 4911 3056 5355 3066
rect 5496 3162 5683 3186
rect 5714 3167 6107 3187
rect 6127 3167 6130 3187
rect 5714 3162 6130 3167
rect 5496 3091 5533 3162
rect 5714 3161 6055 3162
rect 5648 3101 5679 3102
rect 5496 3071 5505 3091
rect 5525 3071 5533 3091
rect 5496 3061 5533 3071
rect 5592 3091 5679 3101
rect 5592 3071 5601 3091
rect 5621 3071 5679 3091
rect 5592 3062 5679 3071
rect 5592 3061 5629 3062
rect 4517 3029 4560 3034
rect 4908 3040 5355 3056
rect 4908 3034 4936 3040
rect 5187 3039 5355 3040
rect 4517 3026 4667 3029
rect 4908 3026 4935 3034
rect 4517 3024 4935 3026
rect 4517 3006 4526 3024
rect 4544 3006 4935 3024
rect 5648 3011 5679 3062
rect 5714 3091 5751 3161
rect 6017 3160 6054 3161
rect 5866 3101 5902 3102
rect 5714 3071 5723 3091
rect 5743 3071 5751 3091
rect 5714 3061 5751 3071
rect 5810 3091 5958 3101
rect 6058 3098 6154 3100
rect 5810 3071 5819 3091
rect 5839 3071 5929 3091
rect 5949 3071 5958 3091
rect 5810 3062 5958 3071
rect 6016 3091 6154 3098
rect 6016 3071 6025 3091
rect 6045 3071 6154 3091
rect 6016 3062 6154 3071
rect 5810 3061 5847 3062
rect 5540 3008 5581 3009
rect 4517 3003 4935 3006
rect 4517 2997 4560 3003
rect 4520 2994 4560 2997
rect 5435 3001 5581 3008
rect 4917 2985 4957 2986
rect 4628 2968 4957 2985
rect 5435 2981 5491 3001
rect 5511 2981 5550 3001
rect 5570 2981 5581 3001
rect 5435 2973 5581 2981
rect 5648 3004 5805 3011
rect 5648 2984 5768 3004
rect 5788 2984 5805 3004
rect 5648 2974 5805 2984
rect 5648 2973 5683 2974
rect 4512 2925 4555 2936
rect 4512 2907 4524 2925
rect 4542 2907 4555 2925
rect 4512 2881 4555 2907
rect 4628 2881 4655 2968
rect 4917 2959 4957 2968
rect 3691 2855 4130 2873
rect 2898 2852 2939 2853
rect 2632 2799 2669 2800
rect 2325 2790 2463 2799
rect 2325 2770 2434 2790
rect 2454 2770 2463 2790
rect 2325 2763 2463 2770
rect 2521 2790 2669 2799
rect 2521 2770 2530 2790
rect 2550 2770 2640 2790
rect 2660 2770 2669 2790
rect 2325 2761 2421 2763
rect 2521 2760 2669 2770
rect 2728 2790 2765 2800
rect 2728 2770 2736 2790
rect 2756 2770 2765 2790
rect 2577 2759 2613 2760
rect 2425 2700 2462 2701
rect 2728 2700 2765 2770
rect 2800 2799 2831 2850
rect 3691 2837 4091 2855
rect 4109 2837 4130 2855
rect 3691 2831 4130 2837
rect 3697 2827 4130 2831
rect 4512 2860 4655 2881
rect 4699 2933 4733 2949
rect 4917 2939 5310 2959
rect 5330 2939 5333 2959
rect 5648 2952 5679 2973
rect 5866 2952 5902 3062
rect 5921 3061 5958 3062
rect 6017 3061 6054 3062
rect 5977 3002 6067 3008
rect 5977 2982 5986 3002
rect 6006 3000 6067 3002
rect 6006 2982 6031 3000
rect 5977 2980 6031 2982
rect 6051 2980 6067 3000
rect 5977 2974 6067 2980
rect 5491 2951 5528 2952
rect 4917 2934 5333 2939
rect 5490 2942 5528 2951
rect 4917 2933 5258 2934
rect 4699 2863 4736 2933
rect 4851 2873 4882 2874
rect 4512 2858 4649 2860
rect 4076 2825 4128 2827
rect 4512 2816 4555 2858
rect 4699 2843 4708 2863
rect 4728 2843 4736 2863
rect 4699 2833 4736 2843
rect 4795 2863 4882 2873
rect 4795 2843 4804 2863
rect 4824 2843 4882 2863
rect 4795 2834 4882 2843
rect 4795 2833 4832 2834
rect 4510 2806 4555 2816
rect 2850 2799 2887 2800
rect 2800 2790 2887 2799
rect 2800 2770 2858 2790
rect 2878 2770 2887 2790
rect 2800 2760 2887 2770
rect 2946 2790 2983 2800
rect 2946 2770 2954 2790
rect 2974 2770 2983 2790
rect 4510 2788 4519 2806
rect 4537 2788 4555 2806
rect 4510 2782 4555 2788
rect 4851 2783 4882 2834
rect 4917 2863 4954 2933
rect 5220 2932 5257 2933
rect 5490 2922 5499 2942
rect 5519 2922 5528 2942
rect 5490 2914 5528 2922
rect 5594 2946 5679 2952
rect 5709 2951 5746 2952
rect 5594 2926 5602 2946
rect 5622 2926 5679 2946
rect 5594 2918 5679 2926
rect 5708 2942 5746 2951
rect 5708 2922 5717 2942
rect 5737 2922 5746 2942
rect 5594 2917 5630 2918
rect 5708 2914 5746 2922
rect 5812 2946 5956 2952
rect 5812 2926 5820 2946
rect 5840 2943 5928 2946
rect 5840 2926 5875 2943
rect 5812 2925 5875 2926
rect 5894 2926 5928 2943
rect 5948 2926 5956 2946
rect 5894 2925 5956 2926
rect 5812 2918 5956 2925
rect 5812 2917 5848 2918
rect 5920 2917 5956 2918
rect 6022 2951 6059 2952
rect 6022 2950 6060 2951
rect 6082 2950 6109 2954
rect 6022 2948 6109 2950
rect 6022 2942 6086 2948
rect 6022 2922 6031 2942
rect 6051 2928 6086 2942
rect 6106 2928 6109 2948
rect 6051 2923 6109 2928
rect 6051 2922 6086 2923
rect 5491 2885 5528 2914
rect 5492 2883 5528 2885
rect 5069 2873 5105 2874
rect 4917 2843 4926 2863
rect 4946 2843 4954 2863
rect 4917 2833 4954 2843
rect 5013 2863 5161 2873
rect 5261 2870 5357 2872
rect 5013 2843 5022 2863
rect 5042 2843 5132 2863
rect 5152 2843 5161 2863
rect 5013 2834 5161 2843
rect 5219 2863 5357 2870
rect 5219 2843 5228 2863
rect 5248 2843 5357 2863
rect 5492 2861 5683 2883
rect 5709 2882 5746 2914
rect 6022 2910 6086 2922
rect 6126 2884 6153 3062
rect 5985 2882 6153 2884
rect 5709 2856 6153 2882
rect 5219 2834 5357 2843
rect 5013 2833 5050 2834
rect 4510 2779 4547 2782
rect 4743 2780 4784 2781
rect 2800 2759 2831 2760
rect 2424 2699 2765 2700
rect 2946 2699 2983 2770
rect 4635 2773 4784 2780
rect 4079 2760 4116 2765
rect 2349 2694 2765 2699
rect 2349 2674 2352 2694
rect 2372 2674 2765 2694
rect 2796 2675 2983 2699
rect 4070 2756 4117 2760
rect 4070 2738 4089 2756
rect 4107 2738 4117 2756
rect 4635 2753 4694 2773
rect 4714 2753 4753 2773
rect 4773 2753 4784 2773
rect 4635 2745 4784 2753
rect 4851 2776 5008 2783
rect 4851 2756 4971 2776
rect 4991 2756 5008 2776
rect 4851 2746 5008 2756
rect 4851 2745 4886 2746
rect 4070 2690 4117 2738
rect 4851 2724 4882 2745
rect 5069 2724 5105 2834
rect 5124 2833 5161 2834
rect 5220 2833 5257 2834
rect 5180 2774 5270 2780
rect 5180 2754 5189 2774
rect 5209 2772 5270 2774
rect 5209 2754 5234 2772
rect 5180 2752 5234 2754
rect 5254 2752 5270 2772
rect 5180 2746 5270 2752
rect 4694 2723 4731 2724
rect 3694 2687 4117 2690
rect 2569 2673 2634 2674
rect 3672 2657 4117 2687
rect 4506 2715 4544 2717
rect 4506 2707 4549 2715
rect 4506 2689 4517 2707
rect 4535 2689 4549 2707
rect 4506 2662 4549 2689
rect 4693 2714 4731 2723
rect 4693 2694 4702 2714
rect 4722 2694 4731 2714
rect 4693 2686 4731 2694
rect 4797 2718 4882 2724
rect 4912 2723 4949 2724
rect 4797 2698 4805 2718
rect 4825 2698 4882 2718
rect 4797 2690 4882 2698
rect 4911 2714 4949 2723
rect 4911 2694 4920 2714
rect 4940 2694 4949 2714
rect 4797 2689 4833 2690
rect 4911 2686 4949 2694
rect 5015 2722 5159 2724
rect 5015 2718 5067 2722
rect 5015 2698 5023 2718
rect 5043 2702 5067 2718
rect 5087 2718 5159 2722
rect 5087 2702 5131 2718
rect 5043 2698 5131 2702
rect 5151 2698 5159 2718
rect 5015 2690 5159 2698
rect 5015 2689 5051 2690
rect 5123 2689 5159 2690
rect 5225 2723 5262 2724
rect 5225 2722 5263 2723
rect 5225 2714 5289 2722
rect 5225 2694 5234 2714
rect 5254 2700 5289 2714
rect 5309 2700 5312 2720
rect 5254 2695 5312 2700
rect 5254 2694 5289 2695
rect 2765 2641 2805 2649
rect 2765 2619 2773 2641
rect 2797 2619 2805 2641
rect 2370 2390 2407 2396
rect 2370 2371 2378 2390
rect 2399 2371 2407 2390
rect 2370 2363 2407 2371
rect 2070 2242 2077 2264
rect 2101 2242 2109 2264
rect 2070 2236 2109 2242
rect 1600 2231 1640 2233
rect 1766 2232 1934 2233
rect 1868 2231 1905 2232
rect 834 2215 972 2224
rect 628 2214 665 2215
rect 358 2161 399 2162
rect 132 2140 184 2158
rect 250 2154 399 2161
rect 250 2134 309 2154
rect 329 2134 368 2154
rect 388 2134 399 2154
rect 250 2126 399 2134
rect 466 2157 623 2164
rect 466 2137 586 2157
rect 606 2137 623 2157
rect 466 2127 623 2137
rect 466 2126 501 2127
rect 466 2105 497 2126
rect 684 2105 720 2215
rect 739 2214 776 2215
rect 835 2214 872 2215
rect 795 2155 885 2161
rect 795 2135 804 2155
rect 824 2153 885 2155
rect 824 2135 849 2153
rect 795 2133 849 2135
rect 869 2133 885 2153
rect 795 2127 885 2133
rect 309 2104 346 2105
rect 308 2095 346 2104
rect 136 2077 176 2087
rect 136 2059 146 2077
rect 164 2059 176 2077
rect 308 2075 317 2095
rect 337 2075 346 2095
rect 308 2067 346 2075
rect 412 2099 497 2105
rect 527 2104 564 2105
rect 412 2079 420 2099
rect 440 2079 497 2099
rect 412 2071 497 2079
rect 526 2095 564 2104
rect 526 2075 535 2095
rect 555 2075 564 2095
rect 412 2070 448 2071
rect 526 2067 564 2075
rect 630 2099 774 2105
rect 630 2079 638 2099
rect 658 2079 691 2099
rect 711 2079 746 2099
rect 766 2079 774 2099
rect 630 2071 774 2079
rect 630 2070 666 2071
rect 738 2070 774 2071
rect 840 2104 877 2105
rect 840 2103 878 2104
rect 840 2095 904 2103
rect 840 2075 849 2095
rect 869 2081 904 2095
rect 924 2081 927 2101
rect 869 2076 927 2081
rect 869 2075 904 2076
rect 136 2003 176 2059
rect 309 2038 346 2067
rect 310 2036 346 2038
rect 310 2014 501 2036
rect 527 2035 564 2067
rect 840 2063 904 2075
rect 944 2037 971 2215
rect 803 2035 971 2037
rect 527 2025 971 2035
rect 1112 2131 1299 2155
rect 1330 2136 1723 2156
rect 1743 2136 1746 2156
rect 1330 2131 1746 2136
rect 1112 2060 1149 2131
rect 1330 2130 1671 2131
rect 1264 2070 1295 2071
rect 1112 2040 1121 2060
rect 1141 2040 1149 2060
rect 1112 2030 1149 2040
rect 1208 2060 1295 2070
rect 1208 2040 1217 2060
rect 1237 2040 1295 2060
rect 1208 2031 1295 2040
rect 1208 2030 1245 2031
rect 133 1998 176 2003
rect 524 2009 971 2025
rect 524 2003 552 2009
rect 803 2008 971 2009
rect 133 1995 283 1998
rect 524 1995 551 2003
rect 133 1993 551 1995
rect 133 1975 142 1993
rect 160 1975 551 1993
rect 1264 1980 1295 2031
rect 1330 2060 1367 2130
rect 1633 2129 1670 2130
rect 1871 2072 1904 2231
rect 1482 2070 1518 2071
rect 1330 2040 1339 2060
rect 1359 2040 1367 2060
rect 1330 2030 1367 2040
rect 1426 2060 1574 2070
rect 1674 2067 1770 2069
rect 1426 2040 1435 2060
rect 1455 2040 1545 2060
rect 1565 2040 1574 2060
rect 1426 2031 1574 2040
rect 1632 2060 1770 2067
rect 1632 2040 1641 2060
rect 1661 2040 1770 2060
rect 1871 2068 1907 2072
rect 1871 2050 1880 2068
rect 1902 2050 1907 2068
rect 1871 2044 1907 2050
rect 1632 2031 1770 2040
rect 1426 2030 1463 2031
rect 1156 1977 1197 1978
rect 133 1972 551 1975
rect 133 1966 176 1972
rect 136 1963 176 1966
rect 1048 1970 1197 1977
rect 533 1954 573 1955
rect 244 1937 573 1954
rect 1048 1950 1107 1970
rect 1127 1950 1166 1970
rect 1186 1950 1197 1970
rect 1048 1942 1197 1950
rect 1264 1973 1421 1980
rect 1264 1953 1384 1973
rect 1404 1953 1421 1973
rect 1264 1943 1421 1953
rect 1264 1942 1299 1943
rect 128 1894 171 1905
rect 128 1876 140 1894
rect 158 1876 171 1894
rect 128 1850 171 1876
rect 244 1850 271 1937
rect 533 1928 573 1937
rect 128 1829 271 1850
rect 315 1902 349 1918
rect 533 1908 926 1928
rect 946 1908 949 1928
rect 1264 1921 1295 1942
rect 1482 1921 1518 2031
rect 1537 2030 1574 2031
rect 1633 2030 1670 2031
rect 1593 1971 1683 1977
rect 1593 1951 1602 1971
rect 1622 1969 1683 1971
rect 1622 1951 1647 1969
rect 1593 1949 1647 1951
rect 1667 1949 1683 1969
rect 1593 1943 1683 1949
rect 1107 1920 1144 1921
rect 533 1903 949 1908
rect 1106 1911 1144 1920
rect 533 1902 874 1903
rect 315 1832 352 1902
rect 467 1842 498 1843
rect 128 1827 265 1829
rect 128 1785 171 1827
rect 315 1812 324 1832
rect 344 1812 352 1832
rect 315 1802 352 1812
rect 411 1832 498 1842
rect 411 1812 420 1832
rect 440 1812 498 1832
rect 411 1803 498 1812
rect 411 1802 448 1803
rect 126 1775 171 1785
rect 126 1757 135 1775
rect 153 1757 171 1775
rect 126 1751 171 1757
rect 467 1752 498 1803
rect 533 1832 570 1902
rect 836 1901 873 1902
rect 1106 1891 1115 1911
rect 1135 1891 1144 1911
rect 1106 1883 1144 1891
rect 1210 1915 1295 1921
rect 1325 1920 1362 1921
rect 1210 1895 1218 1915
rect 1238 1895 1295 1915
rect 1210 1887 1295 1895
rect 1324 1911 1362 1920
rect 1324 1891 1333 1911
rect 1353 1891 1362 1911
rect 1210 1886 1246 1887
rect 1324 1883 1362 1891
rect 1428 1915 1572 1921
rect 1428 1895 1436 1915
rect 1456 1896 1488 1915
rect 1509 1896 1544 1915
rect 1456 1895 1544 1896
rect 1564 1895 1572 1915
rect 1428 1887 1572 1895
rect 1428 1886 1464 1887
rect 1536 1886 1572 1887
rect 1638 1920 1675 1921
rect 1638 1919 1676 1920
rect 1638 1911 1702 1919
rect 1638 1891 1647 1911
rect 1667 1897 1702 1911
rect 1722 1897 1725 1917
rect 1667 1892 1725 1897
rect 1667 1891 1702 1892
rect 1107 1854 1144 1883
rect 1108 1852 1144 1854
rect 685 1842 721 1843
rect 533 1812 542 1832
rect 562 1812 570 1832
rect 533 1802 570 1812
rect 629 1832 777 1842
rect 877 1839 973 1841
rect 629 1812 638 1832
rect 658 1812 748 1832
rect 768 1812 777 1832
rect 629 1803 777 1812
rect 835 1832 973 1839
rect 835 1812 844 1832
rect 864 1812 973 1832
rect 1108 1830 1299 1852
rect 1325 1851 1362 1883
rect 1638 1879 1702 1891
rect 1742 1853 1769 2031
rect 2374 2030 2407 2363
rect 2471 2395 2639 2396
rect 2765 2395 2805 2619
rect 3268 2623 3436 2624
rect 3672 2623 3713 2657
rect 4070 2636 4117 2657
rect 3268 2613 3713 2623
rect 3785 2621 3928 2622
rect 3268 2597 3712 2613
rect 3268 2595 3436 2597
rect 3632 2596 3712 2597
rect 3785 2596 3930 2621
rect 4072 2596 4117 2636
rect 3268 2417 3295 2595
rect 3335 2557 3399 2569
rect 3675 2565 3712 2596
rect 3893 2565 3930 2596
rect 4075 2589 4117 2596
rect 4507 2655 4549 2662
rect 4694 2655 4731 2686
rect 4912 2655 4949 2686
rect 5225 2682 5289 2694
rect 5329 2656 5356 2834
rect 4507 2615 4552 2655
rect 4694 2630 4839 2655
rect 4912 2654 4992 2655
rect 5188 2654 5356 2656
rect 4912 2638 5356 2654
rect 4696 2629 4839 2630
rect 4911 2628 5356 2638
rect 4507 2594 4554 2615
rect 4911 2594 4952 2628
rect 5188 2627 5356 2628
rect 5819 2632 5859 2856
rect 5985 2855 6153 2856
rect 6217 2888 6250 3221
rect 6217 2880 6254 2888
rect 6217 2861 6225 2880
rect 6246 2861 6254 2880
rect 6217 2855 6254 2861
rect 5819 2610 5827 2632
rect 5851 2610 5859 2632
rect 5819 2602 5859 2610
rect 3335 2556 3370 2557
rect 3312 2551 3370 2556
rect 3312 2531 3315 2551
rect 3335 2537 3370 2551
rect 3390 2537 3399 2557
rect 3335 2529 3399 2537
rect 3361 2528 3399 2529
rect 3362 2527 3399 2528
rect 3465 2561 3501 2562
rect 3573 2561 3609 2562
rect 3465 2553 3609 2561
rect 3465 2533 3473 2553
rect 3493 2549 3581 2553
rect 3493 2533 3537 2549
rect 3465 2529 3537 2533
rect 3557 2533 3581 2549
rect 3601 2533 3609 2553
rect 3557 2529 3609 2533
rect 3465 2527 3609 2529
rect 3675 2557 3713 2565
rect 3791 2561 3827 2562
rect 3675 2537 3684 2557
rect 3704 2537 3713 2557
rect 3675 2528 3713 2537
rect 3742 2553 3827 2561
rect 3742 2533 3799 2553
rect 3819 2533 3827 2553
rect 3675 2527 3712 2528
rect 3742 2527 3827 2533
rect 3893 2557 3931 2565
rect 3893 2537 3902 2557
rect 3922 2537 3931 2557
rect 3893 2528 3931 2537
rect 4075 2562 4118 2589
rect 4075 2544 4089 2562
rect 4107 2544 4118 2562
rect 4075 2536 4118 2544
rect 4080 2534 4118 2536
rect 4507 2564 4952 2594
rect 5990 2577 6055 2578
rect 4507 2561 4930 2564
rect 3893 2527 3930 2528
rect 3354 2499 3444 2505
rect 3354 2479 3370 2499
rect 3390 2497 3444 2499
rect 3390 2479 3415 2497
rect 3354 2477 3415 2479
rect 3435 2477 3444 2497
rect 3354 2471 3444 2477
rect 3367 2417 3404 2418
rect 3463 2417 3500 2418
rect 3519 2417 3555 2527
rect 3742 2506 3773 2527
rect 4507 2513 4554 2561
rect 3738 2505 3773 2506
rect 3616 2495 3773 2505
rect 3616 2475 3633 2495
rect 3653 2475 3773 2495
rect 3616 2468 3773 2475
rect 3840 2498 3989 2506
rect 3840 2478 3851 2498
rect 3871 2478 3910 2498
rect 3930 2478 3989 2498
rect 4507 2495 4517 2513
rect 4535 2495 4554 2513
rect 4507 2491 4554 2495
rect 5641 2552 5828 2576
rect 5859 2557 6252 2577
rect 6272 2557 6275 2577
rect 5859 2552 6275 2557
rect 4508 2486 4545 2491
rect 3840 2471 3989 2478
rect 5641 2481 5678 2552
rect 5859 2551 6200 2552
rect 5793 2491 5824 2492
rect 3840 2470 3881 2471
rect 4077 2469 4114 2472
rect 3574 2417 3611 2418
rect 3267 2408 3405 2417
rect 2471 2369 2915 2395
rect 2471 2367 2639 2369
rect 2471 2189 2498 2367
rect 2538 2329 2602 2341
rect 2878 2337 2915 2369
rect 2941 2368 3132 2390
rect 3267 2388 3376 2408
rect 3396 2388 3405 2408
rect 3267 2381 3405 2388
rect 3463 2408 3611 2417
rect 3463 2388 3472 2408
rect 3492 2388 3582 2408
rect 3602 2388 3611 2408
rect 3267 2379 3363 2381
rect 3463 2378 3611 2388
rect 3670 2408 3707 2418
rect 3670 2388 3678 2408
rect 3698 2388 3707 2408
rect 3519 2377 3555 2378
rect 3096 2366 3132 2368
rect 3096 2337 3133 2366
rect 2538 2328 2573 2329
rect 2515 2323 2573 2328
rect 2515 2303 2518 2323
rect 2538 2309 2573 2323
rect 2593 2309 2602 2329
rect 2538 2303 2602 2309
rect 2515 2301 2602 2303
rect 2515 2297 2542 2301
rect 2564 2300 2602 2301
rect 2565 2299 2602 2300
rect 2668 2333 2704 2334
rect 2776 2333 2812 2334
rect 2668 2326 2812 2333
rect 2668 2325 2730 2326
rect 2668 2305 2676 2325
rect 2696 2308 2730 2325
rect 2749 2325 2812 2326
rect 2749 2308 2784 2325
rect 2696 2305 2784 2308
rect 2804 2305 2812 2325
rect 2668 2299 2812 2305
rect 2878 2329 2916 2337
rect 2994 2333 3030 2334
rect 2878 2309 2887 2329
rect 2907 2309 2916 2329
rect 2878 2300 2916 2309
rect 2945 2325 3030 2333
rect 2945 2305 3002 2325
rect 3022 2305 3030 2325
rect 2878 2299 2915 2300
rect 2945 2299 3030 2305
rect 3096 2329 3134 2337
rect 3096 2309 3105 2329
rect 3125 2309 3134 2329
rect 3367 2318 3404 2319
rect 3670 2318 3707 2388
rect 3742 2417 3773 2468
rect 4069 2463 4114 2469
rect 4069 2445 4087 2463
rect 4105 2445 4114 2463
rect 5641 2461 5650 2481
rect 5670 2461 5678 2481
rect 5641 2451 5678 2461
rect 5737 2481 5824 2491
rect 5737 2461 5746 2481
rect 5766 2461 5824 2481
rect 5737 2452 5824 2461
rect 5737 2451 5774 2452
rect 4069 2435 4114 2445
rect 3792 2417 3829 2418
rect 3742 2408 3829 2417
rect 3742 2388 3800 2408
rect 3820 2388 3829 2408
rect 3742 2378 3829 2388
rect 3888 2408 3925 2418
rect 3888 2388 3896 2408
rect 3916 2388 3925 2408
rect 4069 2393 4112 2435
rect 4496 2424 4548 2426
rect 3975 2391 4112 2393
rect 3742 2377 3773 2378
rect 3888 2318 3925 2388
rect 3366 2317 3707 2318
rect 3096 2300 3134 2309
rect 3291 2312 3707 2317
rect 3096 2299 3133 2300
rect 2557 2271 2647 2277
rect 2557 2251 2573 2271
rect 2593 2269 2647 2271
rect 2593 2251 2618 2269
rect 2557 2249 2618 2251
rect 2638 2249 2647 2269
rect 2557 2243 2647 2249
rect 2570 2189 2607 2190
rect 2666 2189 2703 2190
rect 2722 2189 2758 2299
rect 2945 2278 2976 2299
rect 3291 2292 3294 2312
rect 3314 2292 3707 2312
rect 3891 2302 3925 2318
rect 3969 2370 4112 2391
rect 4494 2420 4927 2424
rect 4494 2414 4933 2420
rect 4494 2396 4515 2414
rect 4533 2396 4933 2414
rect 5793 2401 5824 2452
rect 5859 2481 5896 2551
rect 6162 2550 6199 2551
rect 6011 2491 6047 2492
rect 5859 2461 5868 2481
rect 5888 2461 5896 2481
rect 5859 2451 5896 2461
rect 5955 2481 6103 2491
rect 6203 2488 6299 2490
rect 5955 2461 5964 2481
rect 5984 2461 6074 2481
rect 6094 2461 6103 2481
rect 5955 2452 6103 2461
rect 6161 2481 6299 2488
rect 6161 2461 6170 2481
rect 6190 2461 6299 2481
rect 6161 2452 6299 2461
rect 5955 2451 5992 2452
rect 5685 2398 5726 2399
rect 4494 2378 4933 2396
rect 3667 2283 3707 2292
rect 3969 2283 3996 2370
rect 4069 2344 4112 2370
rect 4069 2326 4082 2344
rect 4100 2326 4112 2344
rect 4069 2315 4112 2326
rect 2941 2277 2976 2278
rect 2819 2267 2976 2277
rect 2819 2247 2836 2267
rect 2856 2247 2976 2267
rect 2819 2240 2976 2247
rect 3043 2270 3189 2278
rect 3043 2250 3054 2270
rect 3074 2250 3113 2270
rect 3133 2250 3189 2270
rect 3667 2266 3996 2283
rect 3667 2265 3707 2266
rect 3043 2243 3189 2250
rect 4064 2254 4104 2257
rect 4064 2248 4107 2254
rect 3689 2245 4107 2248
rect 3043 2242 3084 2243
rect 2777 2189 2814 2190
rect 2470 2180 2608 2189
rect 2470 2160 2579 2180
rect 2599 2160 2608 2180
rect 2470 2153 2608 2160
rect 2666 2180 2814 2189
rect 2666 2160 2675 2180
rect 2695 2160 2785 2180
rect 2805 2160 2814 2180
rect 2470 2151 2566 2153
rect 2666 2150 2814 2160
rect 2873 2180 2910 2190
rect 2873 2160 2881 2180
rect 2901 2160 2910 2180
rect 2722 2149 2758 2150
rect 2570 2090 2607 2091
rect 2873 2090 2910 2160
rect 2945 2189 2976 2240
rect 3689 2227 4080 2245
rect 4098 2227 4107 2245
rect 3689 2225 4107 2227
rect 3689 2217 3716 2225
rect 3957 2222 4107 2225
rect 3269 2211 3437 2212
rect 3688 2211 3716 2217
rect 3269 2195 3716 2211
rect 4064 2217 4107 2222
rect 2995 2189 3032 2190
rect 2945 2180 3032 2189
rect 2945 2160 3003 2180
rect 3023 2160 3032 2180
rect 2945 2150 3032 2160
rect 3091 2180 3128 2190
rect 3091 2160 3099 2180
rect 3119 2160 3128 2180
rect 2945 2149 2976 2150
rect 2569 2089 2910 2090
rect 3091 2089 3128 2160
rect 2494 2084 2910 2089
rect 2494 2064 2497 2084
rect 2517 2064 2910 2084
rect 2941 2065 3128 2089
rect 3269 2185 3713 2195
rect 3269 2183 3437 2185
rect 2369 1985 2411 2030
rect 3269 2005 3296 2183
rect 3336 2145 3400 2157
rect 3676 2153 3713 2185
rect 3739 2184 3930 2206
rect 3894 2182 3930 2184
rect 3894 2153 3931 2182
rect 4064 2161 4104 2217
rect 3336 2144 3371 2145
rect 3313 2139 3371 2144
rect 3313 2119 3316 2139
rect 3336 2125 3371 2139
rect 3391 2125 3400 2145
rect 3336 2117 3400 2125
rect 3362 2116 3400 2117
rect 3363 2115 3400 2116
rect 3466 2149 3502 2150
rect 3574 2149 3610 2150
rect 3466 2141 3610 2149
rect 3466 2121 3474 2141
rect 3494 2121 3529 2141
rect 3549 2121 3582 2141
rect 3602 2121 3610 2141
rect 3466 2115 3610 2121
rect 3676 2145 3714 2153
rect 3792 2149 3828 2150
rect 3676 2125 3685 2145
rect 3705 2125 3714 2145
rect 3676 2116 3714 2125
rect 3743 2141 3828 2149
rect 3743 2121 3800 2141
rect 3820 2121 3828 2141
rect 3676 2115 3713 2116
rect 3743 2115 3828 2121
rect 3894 2145 3932 2153
rect 3894 2125 3903 2145
rect 3923 2125 3932 2145
rect 4064 2143 4076 2161
rect 4094 2143 4104 2161
rect 4496 2189 4548 2378
rect 4894 2353 4933 2378
rect 5577 2391 5726 2398
rect 5577 2371 5636 2391
rect 5656 2371 5695 2391
rect 5715 2371 5726 2391
rect 5577 2363 5726 2371
rect 5793 2394 5950 2401
rect 5793 2374 5913 2394
rect 5933 2374 5950 2394
rect 5793 2364 5950 2374
rect 5793 2363 5828 2364
rect 4678 2328 4865 2352
rect 4894 2333 5289 2353
rect 5309 2333 5312 2353
rect 5793 2342 5824 2363
rect 6011 2342 6047 2452
rect 6066 2451 6103 2452
rect 6162 2451 6199 2452
rect 6122 2392 6212 2398
rect 6122 2372 6131 2392
rect 6151 2390 6212 2392
rect 6151 2372 6176 2390
rect 6122 2370 6176 2372
rect 6196 2370 6212 2390
rect 6122 2364 6212 2370
rect 5636 2341 5673 2342
rect 4894 2328 5312 2333
rect 5635 2332 5673 2341
rect 4678 2257 4715 2328
rect 4894 2327 5237 2328
rect 4894 2324 4933 2327
rect 5199 2326 5236 2327
rect 4830 2267 4861 2268
rect 4678 2237 4687 2257
rect 4707 2237 4715 2257
rect 4678 2227 4715 2237
rect 4774 2257 4861 2267
rect 4774 2237 4783 2257
rect 4803 2237 4861 2257
rect 4774 2228 4861 2237
rect 4774 2227 4811 2228
rect 4496 2171 4512 2189
rect 4530 2171 4548 2189
rect 4830 2177 4861 2228
rect 4896 2257 4933 2324
rect 5635 2312 5644 2332
rect 5664 2312 5673 2332
rect 5635 2304 5673 2312
rect 5739 2336 5824 2342
rect 5854 2341 5891 2342
rect 5739 2316 5747 2336
rect 5767 2316 5824 2336
rect 5739 2308 5824 2316
rect 5853 2332 5891 2341
rect 5853 2312 5862 2332
rect 5882 2312 5891 2332
rect 5739 2307 5775 2308
rect 5853 2304 5891 2312
rect 5957 2340 6101 2342
rect 5957 2336 6017 2340
rect 5957 2316 5965 2336
rect 5985 2318 6017 2336
rect 6040 2336 6101 2340
rect 6040 2318 6073 2336
rect 5985 2316 6073 2318
rect 6093 2316 6101 2336
rect 5957 2308 6101 2316
rect 5957 2307 5993 2308
rect 6065 2307 6101 2308
rect 6167 2341 6204 2342
rect 6167 2340 6205 2341
rect 6167 2332 6231 2340
rect 6167 2312 6176 2332
rect 6196 2318 6231 2332
rect 6251 2318 6254 2338
rect 6196 2313 6254 2318
rect 6196 2312 6231 2313
rect 5636 2275 5673 2304
rect 5637 2273 5673 2275
rect 5048 2267 5084 2268
rect 4896 2237 4905 2257
rect 4925 2237 4933 2257
rect 4896 2227 4933 2237
rect 4992 2257 5140 2267
rect 5240 2264 5336 2266
rect 4992 2237 5001 2257
rect 5021 2237 5111 2257
rect 5131 2237 5140 2257
rect 4992 2228 5140 2237
rect 5198 2257 5336 2264
rect 5198 2237 5207 2257
rect 5227 2237 5336 2257
rect 5637 2251 5828 2273
rect 5854 2272 5891 2304
rect 6167 2300 6231 2312
rect 5854 2271 6129 2272
rect 6271 2271 6298 2452
rect 5854 2246 6298 2271
rect 6434 2277 6473 4092
rect 6775 4079 6808 4412
rect 6872 4444 7040 4445
rect 7166 4444 7206 4668
rect 7669 4672 7837 4673
rect 8078 4672 8113 4689
rect 8470 4679 8517 4690
rect 7669 4646 8113 4672
rect 7669 4644 7837 4646
rect 8033 4645 8113 4646
rect 8268 4645 8335 4671
rect 8474 4645 8517 4679
rect 7669 4466 7696 4644
rect 7736 4606 7800 4618
rect 8076 4614 8113 4645
rect 8294 4614 8331 4645
rect 8476 4620 8517 4645
rect 7736 4605 7771 4606
rect 7713 4600 7771 4605
rect 7713 4580 7716 4600
rect 7736 4586 7771 4600
rect 7791 4586 7800 4606
rect 7736 4578 7800 4586
rect 7762 4577 7800 4578
rect 7763 4576 7800 4577
rect 7866 4610 7902 4611
rect 7974 4610 8010 4611
rect 7866 4602 8010 4610
rect 7866 4582 7874 4602
rect 7894 4598 7982 4602
rect 7894 4582 7938 4598
rect 7866 4578 7938 4582
rect 7958 4582 7982 4598
rect 8002 4582 8010 4602
rect 7958 4578 8010 4582
rect 7866 4576 8010 4578
rect 8076 4606 8114 4614
rect 8192 4610 8228 4611
rect 8076 4586 8085 4606
rect 8105 4586 8114 4606
rect 8076 4577 8114 4586
rect 8143 4602 8228 4610
rect 8143 4582 8200 4602
rect 8220 4582 8228 4602
rect 8076 4576 8113 4577
rect 8143 4576 8228 4582
rect 8294 4606 8332 4614
rect 8294 4586 8303 4606
rect 8323 4586 8332 4606
rect 8294 4577 8332 4586
rect 8476 4611 8518 4620
rect 8476 4593 8490 4611
rect 8508 4593 8518 4611
rect 8476 4585 8518 4593
rect 8481 4583 8518 4585
rect 8294 4576 8331 4577
rect 7755 4548 7845 4554
rect 7755 4528 7771 4548
rect 7791 4546 7845 4548
rect 7791 4528 7816 4546
rect 7755 4526 7816 4528
rect 7836 4526 7845 4546
rect 7755 4520 7845 4526
rect 7768 4466 7805 4467
rect 7864 4466 7901 4467
rect 7920 4466 7956 4576
rect 8143 4555 8174 4576
rect 8139 4554 8174 4555
rect 8017 4544 8174 4554
rect 8017 4524 8034 4544
rect 8054 4524 8174 4544
rect 8017 4517 8174 4524
rect 8241 4547 8390 4555
rect 8241 4527 8252 4547
rect 8272 4527 8311 4547
rect 8331 4527 8390 4547
rect 8241 4520 8390 4527
rect 8241 4519 8282 4520
rect 8478 4518 8515 4521
rect 7975 4466 8012 4467
rect 7668 4457 7806 4466
rect 6872 4418 7316 4444
rect 6872 4416 7040 4418
rect 6872 4238 6899 4416
rect 6939 4378 7003 4390
rect 7279 4386 7316 4418
rect 7342 4417 7533 4439
rect 7668 4437 7777 4457
rect 7797 4437 7806 4457
rect 7668 4430 7806 4437
rect 7864 4457 8012 4466
rect 7864 4437 7873 4457
rect 7893 4437 7983 4457
rect 8003 4437 8012 4457
rect 7668 4428 7764 4430
rect 7864 4427 8012 4437
rect 8071 4457 8108 4467
rect 8071 4437 8079 4457
rect 8099 4437 8108 4457
rect 7920 4426 7956 4427
rect 7497 4415 7533 4417
rect 7497 4386 7534 4415
rect 6939 4377 6974 4378
rect 6916 4372 6974 4377
rect 6916 4352 6919 4372
rect 6939 4358 6974 4372
rect 6994 4358 7003 4378
rect 6939 4352 7003 4358
rect 6916 4350 7003 4352
rect 6916 4346 6943 4350
rect 6965 4349 7003 4350
rect 6966 4348 7003 4349
rect 7069 4382 7105 4383
rect 7177 4382 7213 4383
rect 7069 4375 7213 4382
rect 7069 4374 7131 4375
rect 7069 4354 7077 4374
rect 7097 4357 7131 4374
rect 7150 4374 7213 4375
rect 7150 4357 7185 4374
rect 7097 4354 7185 4357
rect 7205 4354 7213 4374
rect 7069 4348 7213 4354
rect 7279 4378 7317 4386
rect 7395 4382 7431 4383
rect 7279 4358 7288 4378
rect 7308 4358 7317 4378
rect 7279 4349 7317 4358
rect 7346 4374 7431 4382
rect 7346 4354 7403 4374
rect 7423 4354 7431 4374
rect 7279 4348 7316 4349
rect 7346 4348 7431 4354
rect 7497 4378 7535 4386
rect 7497 4358 7506 4378
rect 7526 4358 7535 4378
rect 7768 4367 7805 4368
rect 8071 4367 8108 4437
rect 8143 4466 8174 4517
rect 8470 4512 8515 4518
rect 8470 4494 8488 4512
rect 8506 4494 8515 4512
rect 8470 4484 8515 4494
rect 8193 4466 8230 4467
rect 8143 4457 8230 4466
rect 8143 4437 8201 4457
rect 8221 4437 8230 4457
rect 8143 4427 8230 4437
rect 8289 4457 8326 4467
rect 8289 4437 8297 4457
rect 8317 4437 8326 4457
rect 8470 4442 8513 4484
rect 8376 4440 8513 4442
rect 8143 4426 8174 4427
rect 8289 4367 8326 4437
rect 7767 4366 8108 4367
rect 7497 4349 7535 4358
rect 7692 4361 8108 4366
rect 7497 4348 7534 4349
rect 6958 4320 7048 4326
rect 6958 4300 6974 4320
rect 6994 4318 7048 4320
rect 6994 4300 7019 4318
rect 6958 4298 7019 4300
rect 7039 4298 7048 4318
rect 6958 4292 7048 4298
rect 6971 4238 7008 4239
rect 7067 4238 7104 4239
rect 7123 4238 7159 4348
rect 7346 4327 7377 4348
rect 7692 4341 7695 4361
rect 7715 4341 8108 4361
rect 8292 4351 8326 4367
rect 8370 4419 8513 4440
rect 8068 4332 8108 4341
rect 8370 4332 8397 4419
rect 8470 4393 8513 4419
rect 8470 4375 8483 4393
rect 8501 4375 8513 4393
rect 8470 4364 8513 4375
rect 7342 4326 7377 4327
rect 7220 4316 7377 4326
rect 7220 4296 7237 4316
rect 7257 4296 7377 4316
rect 7220 4289 7377 4296
rect 7444 4319 7590 4327
rect 7444 4299 7455 4319
rect 7475 4299 7514 4319
rect 7534 4299 7590 4319
rect 8068 4315 8397 4332
rect 8068 4314 8108 4315
rect 7444 4292 7590 4299
rect 8465 4303 8505 4306
rect 8465 4297 8508 4303
rect 8090 4294 8508 4297
rect 7444 4291 7485 4292
rect 7178 4238 7215 4239
rect 6871 4229 7009 4238
rect 6871 4209 6980 4229
rect 7000 4209 7009 4229
rect 6871 4202 7009 4209
rect 7067 4229 7215 4238
rect 7067 4209 7076 4229
rect 7096 4209 7186 4229
rect 7206 4209 7215 4229
rect 6871 4200 6967 4202
rect 7067 4199 7215 4209
rect 7274 4229 7311 4239
rect 7274 4209 7282 4229
rect 7302 4209 7311 4229
rect 7123 4198 7159 4199
rect 6971 4139 7008 4140
rect 7274 4139 7311 4209
rect 7346 4238 7377 4289
rect 8090 4276 8481 4294
rect 8499 4276 8508 4294
rect 8090 4274 8508 4276
rect 8090 4266 8117 4274
rect 8358 4271 8508 4274
rect 7670 4260 7838 4261
rect 8089 4260 8117 4266
rect 7670 4244 8117 4260
rect 8465 4266 8508 4271
rect 7396 4238 7433 4239
rect 7346 4229 7433 4238
rect 7346 4209 7404 4229
rect 7424 4209 7433 4229
rect 7346 4199 7433 4209
rect 7492 4229 7529 4239
rect 7492 4209 7500 4229
rect 7520 4209 7529 4229
rect 7346 4198 7377 4199
rect 6970 4138 7311 4139
rect 7492 4138 7529 4209
rect 6895 4133 7311 4138
rect 6895 4113 6898 4133
rect 6918 4113 7311 4133
rect 7342 4114 7529 4138
rect 7670 4234 8114 4244
rect 7670 4232 7838 4234
rect 6704 4039 6748 4040
rect 6704 4033 6749 4039
rect 6704 4015 6716 4033
rect 6738 4015 6749 4033
rect 6770 4034 6812 4079
rect 7670 4054 7697 4232
rect 7737 4194 7801 4206
rect 8077 4202 8114 4234
rect 8140 4233 8331 4255
rect 8295 4231 8331 4233
rect 8295 4202 8332 4231
rect 8465 4210 8505 4266
rect 7737 4193 7772 4194
rect 7714 4188 7772 4193
rect 7714 4168 7717 4188
rect 7737 4174 7772 4188
rect 7792 4174 7801 4194
rect 7737 4166 7801 4174
rect 7763 4165 7801 4166
rect 7764 4164 7801 4165
rect 7867 4198 7903 4199
rect 7975 4198 8011 4199
rect 7867 4190 8011 4198
rect 7867 4170 7875 4190
rect 7895 4170 7930 4190
rect 7950 4170 7983 4190
rect 8003 4170 8011 4190
rect 7867 4164 8011 4170
rect 8077 4194 8115 4202
rect 8193 4198 8229 4199
rect 8077 4174 8086 4194
rect 8106 4174 8115 4194
rect 8077 4165 8115 4174
rect 8144 4190 8229 4198
rect 8144 4170 8201 4190
rect 8221 4170 8229 4190
rect 8077 4164 8114 4165
rect 8144 4164 8229 4170
rect 8295 4194 8333 4202
rect 8295 4174 8304 4194
rect 8324 4174 8333 4194
rect 8465 4192 8477 4210
rect 8495 4192 8505 4210
rect 8465 4182 8505 4192
rect 8295 4165 8333 4174
rect 8295 4164 8332 4165
rect 7756 4136 7846 4142
rect 7756 4116 7772 4136
rect 7792 4134 7846 4136
rect 7792 4116 7817 4134
rect 7756 4114 7817 4116
rect 7837 4114 7846 4134
rect 7756 4108 7846 4114
rect 7769 4054 7806 4055
rect 7865 4054 7902 4055
rect 7921 4054 7957 4164
rect 8144 4143 8175 4164
rect 8140 4142 8175 4143
rect 8018 4132 8175 4142
rect 8018 4112 8035 4132
rect 8055 4112 8175 4132
rect 8018 4105 8175 4112
rect 8242 4135 8391 4143
rect 8242 4115 8253 4135
rect 8273 4115 8312 4135
rect 8332 4115 8391 4135
rect 8242 4108 8391 4115
rect 8457 4111 8509 4129
rect 8242 4107 8283 4108
rect 7976 4054 8013 4055
rect 7669 4045 7807 4054
rect 7141 4034 7174 4036
rect 6770 4022 7217 4034
rect 6704 3985 6749 4015
rect 6721 3039 6749 3985
rect 6773 4008 7217 4022
rect 6773 4006 6941 4008
rect 6773 3828 6800 4006
rect 6840 3968 6904 3980
rect 7180 3976 7217 4008
rect 7243 4007 7434 4029
rect 7669 4025 7778 4045
rect 7798 4025 7807 4045
rect 7669 4018 7807 4025
rect 7865 4045 8013 4054
rect 7865 4025 7874 4045
rect 7894 4025 7984 4045
rect 8004 4025 8013 4045
rect 7669 4016 7765 4018
rect 7865 4015 8013 4025
rect 8072 4045 8109 4055
rect 8072 4025 8080 4045
rect 8100 4025 8109 4045
rect 7921 4014 7957 4015
rect 7398 4005 7434 4007
rect 7398 3976 7435 4005
rect 6840 3967 6875 3968
rect 6817 3962 6875 3967
rect 6817 3942 6820 3962
rect 6840 3948 6875 3962
rect 6895 3948 6904 3968
rect 6840 3940 6904 3948
rect 6866 3939 6904 3940
rect 6867 3938 6904 3939
rect 6970 3972 7006 3973
rect 7078 3972 7114 3973
rect 6970 3966 7114 3972
rect 6970 3964 7031 3966
rect 6970 3944 6978 3964
rect 6998 3949 7031 3964
rect 7050 3964 7114 3966
rect 7050 3949 7086 3964
rect 6998 3944 7086 3949
rect 7106 3944 7114 3964
rect 6970 3938 7114 3944
rect 7180 3968 7218 3976
rect 7296 3972 7332 3973
rect 7180 3948 7189 3968
rect 7209 3948 7218 3968
rect 7180 3939 7218 3948
rect 7247 3964 7332 3972
rect 7247 3944 7304 3964
rect 7324 3944 7332 3964
rect 7180 3938 7217 3939
rect 7247 3938 7332 3944
rect 7398 3968 7436 3976
rect 7398 3948 7407 3968
rect 7427 3948 7436 3968
rect 8072 3958 8109 4025
rect 8144 4054 8175 4105
rect 8457 4093 8475 4111
rect 8493 4093 8509 4111
rect 8194 4054 8231 4055
rect 8144 4045 8231 4054
rect 8144 4025 8202 4045
rect 8222 4025 8231 4045
rect 8144 4015 8231 4025
rect 8290 4045 8327 4055
rect 8290 4025 8298 4045
rect 8318 4025 8327 4045
rect 8144 4014 8175 4015
rect 7769 3955 7806 3956
rect 8072 3955 8111 3958
rect 7768 3954 8111 3955
rect 8290 3954 8327 4025
rect 7398 3939 7436 3948
rect 7693 3949 8111 3954
rect 7398 3938 7435 3939
rect 6859 3910 6949 3916
rect 6859 3890 6875 3910
rect 6895 3908 6949 3910
rect 6895 3890 6920 3908
rect 6859 3888 6920 3890
rect 6940 3888 6949 3908
rect 6859 3882 6949 3888
rect 6872 3828 6909 3829
rect 6968 3828 7005 3829
rect 7024 3828 7060 3938
rect 7247 3917 7278 3938
rect 7693 3929 7696 3949
rect 7716 3929 8111 3949
rect 8140 3930 8327 3954
rect 7243 3916 7278 3917
rect 7121 3906 7278 3916
rect 7121 3886 7138 3906
rect 7158 3886 7278 3906
rect 7121 3879 7278 3886
rect 7345 3909 7494 3917
rect 7345 3889 7356 3909
rect 7376 3889 7415 3909
rect 7435 3889 7494 3909
rect 7345 3882 7494 3889
rect 8072 3904 8111 3929
rect 8457 3904 8509 4093
rect 8072 3886 8511 3904
rect 7345 3881 7386 3882
rect 7079 3828 7116 3829
rect 6772 3819 6910 3828
rect 6772 3799 6881 3819
rect 6901 3799 6910 3819
rect 6772 3792 6910 3799
rect 6968 3819 7116 3828
rect 6968 3799 6977 3819
rect 6997 3799 7087 3819
rect 7107 3799 7116 3819
rect 6772 3790 6868 3792
rect 6968 3789 7116 3799
rect 7175 3819 7212 3829
rect 7175 3799 7183 3819
rect 7203 3799 7212 3819
rect 7024 3788 7060 3789
rect 6872 3729 6909 3730
rect 7175 3729 7212 3799
rect 7247 3828 7278 3879
rect 8072 3868 8472 3886
rect 8490 3868 8511 3886
rect 8072 3862 8511 3868
rect 8078 3858 8511 3862
rect 8457 3856 8509 3858
rect 7297 3828 7334 3829
rect 7247 3819 7334 3828
rect 7247 3799 7305 3819
rect 7325 3799 7334 3819
rect 7247 3789 7334 3799
rect 7393 3819 7430 3829
rect 7393 3799 7401 3819
rect 7421 3799 7430 3819
rect 7247 3788 7278 3789
rect 6871 3728 7212 3729
rect 7393 3728 7430 3799
rect 8460 3791 8497 3796
rect 8451 3787 8498 3791
rect 8451 3769 8470 3787
rect 8488 3769 8498 3787
rect 6796 3723 7212 3728
rect 6796 3703 6799 3723
rect 6819 3703 7212 3723
rect 7243 3704 7430 3728
rect 8055 3726 8095 3731
rect 8451 3726 8498 3769
rect 8055 3687 8498 3726
rect 7149 3672 7189 3680
rect 7149 3650 7157 3672
rect 7181 3650 7189 3672
rect 6855 3426 7023 3427
rect 7149 3426 7189 3650
rect 7652 3654 7820 3655
rect 8055 3654 8095 3687
rect 8451 3654 8498 3687
rect 7652 3653 8096 3654
rect 7652 3628 8097 3653
rect 7652 3626 7820 3628
rect 8016 3627 8097 3628
rect 8266 3627 8315 3653
rect 8451 3627 8500 3654
rect 7652 3448 7679 3626
rect 7719 3588 7783 3600
rect 8059 3596 8096 3627
rect 8277 3596 8314 3627
rect 8459 3602 8500 3627
rect 7719 3587 7754 3588
rect 7696 3582 7754 3587
rect 7696 3562 7699 3582
rect 7719 3568 7754 3582
rect 7774 3568 7783 3588
rect 7719 3560 7783 3568
rect 7745 3559 7783 3560
rect 7746 3558 7783 3559
rect 7849 3592 7885 3593
rect 7957 3592 7993 3593
rect 7849 3584 7993 3592
rect 7849 3564 7857 3584
rect 7877 3580 7965 3584
rect 7877 3564 7921 3580
rect 7849 3560 7921 3564
rect 7941 3564 7965 3580
rect 7985 3564 7993 3584
rect 7941 3560 7993 3564
rect 7849 3558 7993 3560
rect 8059 3588 8097 3596
rect 8175 3592 8211 3593
rect 8059 3568 8068 3588
rect 8088 3568 8097 3588
rect 8059 3559 8097 3568
rect 8126 3584 8211 3592
rect 8126 3564 8183 3584
rect 8203 3564 8211 3584
rect 8059 3558 8096 3559
rect 8126 3558 8211 3564
rect 8277 3588 8315 3596
rect 8277 3568 8286 3588
rect 8306 3568 8315 3588
rect 8277 3559 8315 3568
rect 8459 3593 8501 3602
rect 8459 3575 8473 3593
rect 8491 3575 8501 3593
rect 8459 3567 8501 3575
rect 8464 3565 8501 3567
rect 8277 3558 8314 3559
rect 7738 3530 7828 3536
rect 7738 3510 7754 3530
rect 7774 3528 7828 3530
rect 7774 3510 7799 3528
rect 7738 3508 7799 3510
rect 7819 3508 7828 3528
rect 7738 3502 7828 3508
rect 7751 3448 7788 3449
rect 7847 3448 7884 3449
rect 7903 3448 7939 3558
rect 8126 3537 8157 3558
rect 8122 3536 8157 3537
rect 8000 3526 8157 3536
rect 8000 3506 8017 3526
rect 8037 3506 8157 3526
rect 8000 3499 8157 3506
rect 8224 3529 8373 3537
rect 8224 3509 8235 3529
rect 8255 3509 8294 3529
rect 8314 3509 8373 3529
rect 8224 3502 8373 3509
rect 8224 3501 8265 3502
rect 8461 3500 8498 3503
rect 7958 3448 7995 3449
rect 7651 3439 7789 3448
rect 6855 3400 7299 3426
rect 6855 3398 7023 3400
rect 6855 3220 6882 3398
rect 6922 3360 6986 3372
rect 7262 3368 7299 3400
rect 7325 3399 7516 3421
rect 7651 3419 7760 3439
rect 7780 3419 7789 3439
rect 7651 3412 7789 3419
rect 7847 3439 7995 3448
rect 7847 3419 7856 3439
rect 7876 3419 7966 3439
rect 7986 3419 7995 3439
rect 7651 3410 7747 3412
rect 7847 3409 7995 3419
rect 8054 3439 8091 3449
rect 8054 3419 8062 3439
rect 8082 3419 8091 3439
rect 7903 3408 7939 3409
rect 7480 3397 7516 3399
rect 7480 3368 7517 3397
rect 6922 3359 6957 3360
rect 6899 3354 6957 3359
rect 6899 3334 6902 3354
rect 6922 3340 6957 3354
rect 6977 3340 6986 3360
rect 6922 3332 6986 3340
rect 6948 3331 6986 3332
rect 6949 3330 6986 3331
rect 7052 3364 7088 3365
rect 7160 3364 7196 3365
rect 7052 3356 7196 3364
rect 7052 3336 7060 3356
rect 7080 3355 7168 3356
rect 7080 3336 7115 3355
rect 7136 3336 7168 3355
rect 7188 3336 7196 3356
rect 7052 3330 7196 3336
rect 7262 3360 7300 3368
rect 7378 3364 7414 3365
rect 7262 3340 7271 3360
rect 7291 3340 7300 3360
rect 7262 3331 7300 3340
rect 7329 3356 7414 3364
rect 7329 3336 7386 3356
rect 7406 3336 7414 3356
rect 7262 3330 7299 3331
rect 7329 3330 7414 3336
rect 7480 3360 7518 3368
rect 7480 3340 7489 3360
rect 7509 3340 7518 3360
rect 7751 3349 7788 3350
rect 8054 3349 8091 3419
rect 8126 3448 8157 3499
rect 8453 3494 8498 3500
rect 8453 3476 8471 3494
rect 8489 3476 8498 3494
rect 8453 3466 8498 3476
rect 8176 3448 8213 3449
rect 8126 3439 8213 3448
rect 8126 3419 8184 3439
rect 8204 3419 8213 3439
rect 8126 3409 8213 3419
rect 8272 3439 8309 3449
rect 8272 3419 8280 3439
rect 8300 3419 8309 3439
rect 8453 3424 8496 3466
rect 8359 3422 8496 3424
rect 8126 3408 8157 3409
rect 8272 3349 8309 3419
rect 7750 3348 8091 3349
rect 7480 3331 7518 3340
rect 7675 3343 8091 3348
rect 7480 3330 7517 3331
rect 6941 3302 7031 3308
rect 6941 3282 6957 3302
rect 6977 3300 7031 3302
rect 6977 3282 7002 3300
rect 6941 3280 7002 3282
rect 7022 3280 7031 3300
rect 6941 3274 7031 3280
rect 6954 3220 6991 3221
rect 7050 3220 7087 3221
rect 7106 3220 7142 3330
rect 7329 3309 7360 3330
rect 7675 3323 7678 3343
rect 7698 3323 8091 3343
rect 8275 3333 8309 3349
rect 8353 3401 8496 3422
rect 8051 3314 8091 3323
rect 8353 3314 8380 3401
rect 8453 3375 8496 3401
rect 8453 3357 8466 3375
rect 8484 3357 8496 3375
rect 8453 3346 8496 3357
rect 7325 3308 7360 3309
rect 7203 3298 7360 3308
rect 7203 3278 7220 3298
rect 7240 3278 7360 3298
rect 7203 3271 7360 3278
rect 7427 3301 7576 3309
rect 7427 3281 7438 3301
rect 7458 3281 7497 3301
rect 7517 3281 7576 3301
rect 8051 3297 8380 3314
rect 8051 3296 8091 3297
rect 7427 3274 7576 3281
rect 8448 3285 8488 3288
rect 8448 3279 8491 3285
rect 8073 3276 8491 3279
rect 7427 3273 7468 3274
rect 7161 3220 7198 3221
rect 6854 3211 6992 3220
rect 6854 3191 6963 3211
rect 6983 3191 6992 3211
rect 6854 3184 6992 3191
rect 7050 3211 7198 3220
rect 7050 3191 7059 3211
rect 7079 3191 7169 3211
rect 7189 3191 7198 3211
rect 6854 3182 6950 3184
rect 7050 3181 7198 3191
rect 7257 3211 7294 3221
rect 7257 3191 7265 3211
rect 7285 3191 7294 3211
rect 7106 3180 7142 3181
rect 6954 3121 6991 3122
rect 7257 3121 7294 3191
rect 7329 3220 7360 3271
rect 8073 3258 8464 3276
rect 8482 3258 8491 3276
rect 8073 3256 8491 3258
rect 8073 3248 8100 3256
rect 8341 3253 8491 3256
rect 7653 3242 7821 3243
rect 8072 3242 8100 3248
rect 7653 3226 8100 3242
rect 8448 3248 8491 3253
rect 7379 3220 7416 3221
rect 7329 3211 7416 3220
rect 7329 3191 7387 3211
rect 7407 3191 7416 3211
rect 7329 3181 7416 3191
rect 7475 3211 7512 3221
rect 7475 3191 7483 3211
rect 7503 3191 7512 3211
rect 7329 3180 7360 3181
rect 6953 3120 7294 3121
rect 7475 3120 7512 3191
rect 6878 3115 7294 3120
rect 6878 3095 6881 3115
rect 6901 3095 7294 3115
rect 7325 3096 7512 3120
rect 7653 3216 8097 3226
rect 7653 3214 7821 3216
rect 6720 3021 6749 3039
rect 7653 3036 7680 3214
rect 7720 3176 7784 3188
rect 8060 3184 8097 3216
rect 8123 3215 8314 3237
rect 8278 3213 8314 3215
rect 8278 3184 8315 3213
rect 8448 3192 8488 3248
rect 7720 3175 7755 3176
rect 7697 3170 7755 3175
rect 7697 3150 7700 3170
rect 7720 3156 7755 3170
rect 7775 3156 7784 3176
rect 7720 3148 7784 3156
rect 7746 3147 7784 3148
rect 7747 3146 7784 3147
rect 7850 3180 7886 3181
rect 7958 3180 7994 3181
rect 7850 3172 7994 3180
rect 7850 3152 7858 3172
rect 7878 3152 7913 3172
rect 7933 3152 7966 3172
rect 7986 3152 7994 3172
rect 7850 3146 7994 3152
rect 8060 3176 8098 3184
rect 8176 3180 8212 3181
rect 8060 3156 8069 3176
rect 8089 3156 8098 3176
rect 8060 3147 8098 3156
rect 8127 3172 8212 3180
rect 8127 3152 8184 3172
rect 8204 3152 8212 3172
rect 8060 3146 8097 3147
rect 8127 3146 8212 3152
rect 8278 3176 8316 3184
rect 8278 3156 8287 3176
rect 8307 3156 8316 3176
rect 8448 3174 8460 3192
rect 8478 3174 8488 3192
rect 8448 3164 8488 3174
rect 8278 3147 8316 3156
rect 8278 3146 8315 3147
rect 7739 3118 7829 3124
rect 7739 3098 7755 3118
rect 7775 3116 7829 3118
rect 7775 3098 7800 3116
rect 7739 3096 7800 3098
rect 7820 3096 7829 3116
rect 7739 3090 7829 3096
rect 7752 3036 7789 3037
rect 7848 3036 7885 3037
rect 7904 3036 7940 3146
rect 8127 3125 8158 3146
rect 8123 3124 8158 3125
rect 8001 3114 8158 3124
rect 8001 3094 8018 3114
rect 8038 3094 8158 3114
rect 8001 3087 8158 3094
rect 8225 3117 8374 3125
rect 8225 3097 8236 3117
rect 8256 3097 8295 3117
rect 8315 3097 8374 3117
rect 8225 3090 8374 3097
rect 8440 3093 8492 3111
rect 8225 3089 8266 3090
rect 7959 3036 7996 3037
rect 6690 3019 6749 3021
rect 7652 3027 7790 3036
rect 6690 3018 6858 3019
rect 6984 3018 7024 3020
rect 6690 2992 7134 3018
rect 6690 2990 6858 2992
rect 6690 2988 6771 2990
rect 6690 2812 6717 2988
rect 6757 2952 6821 2964
rect 7097 2960 7134 2992
rect 7160 2991 7351 3013
rect 7652 3007 7761 3027
rect 7781 3007 7790 3027
rect 7652 3000 7790 3007
rect 7848 3027 7996 3036
rect 7848 3007 7857 3027
rect 7877 3007 7967 3027
rect 7987 3007 7996 3027
rect 7652 2998 7748 3000
rect 7848 2997 7996 3007
rect 8055 3027 8092 3037
rect 8055 3007 8063 3027
rect 8083 3007 8092 3027
rect 7904 2996 7940 2997
rect 7315 2989 7351 2991
rect 7315 2960 7352 2989
rect 6757 2951 6792 2952
rect 6734 2946 6792 2951
rect 6734 2926 6737 2946
rect 6757 2932 6792 2946
rect 6812 2932 6821 2952
rect 6757 2924 6821 2932
rect 6783 2923 6821 2924
rect 6784 2922 6821 2923
rect 6887 2956 6923 2957
rect 6995 2956 7031 2957
rect 6887 2948 7031 2956
rect 6887 2928 6895 2948
rect 6915 2947 7003 2948
rect 6915 2929 6950 2947
rect 6968 2929 7003 2947
rect 6915 2928 7003 2929
rect 7023 2928 7031 2948
rect 6887 2922 7031 2928
rect 7097 2952 7135 2960
rect 7213 2956 7249 2957
rect 7097 2932 7106 2952
rect 7126 2932 7135 2952
rect 7097 2923 7135 2932
rect 7164 2948 7249 2956
rect 7164 2928 7221 2948
rect 7241 2928 7249 2948
rect 7097 2922 7134 2923
rect 7164 2922 7249 2928
rect 7315 2952 7353 2960
rect 7315 2932 7324 2952
rect 7344 2932 7353 2952
rect 8055 2940 8092 3007
rect 8127 3036 8158 3087
rect 8440 3075 8458 3093
rect 8476 3075 8492 3093
rect 8177 3036 8214 3037
rect 8127 3027 8214 3036
rect 8127 3007 8185 3027
rect 8205 3007 8214 3027
rect 8127 2997 8214 3007
rect 8273 3027 8310 3037
rect 8273 3007 8281 3027
rect 8301 3007 8310 3027
rect 8127 2996 8158 2997
rect 7752 2937 7789 2938
rect 8055 2937 8094 2940
rect 7751 2936 8094 2937
rect 8273 2936 8310 3007
rect 7315 2923 7353 2932
rect 7676 2931 8094 2936
rect 7315 2922 7352 2923
rect 6776 2894 6866 2900
rect 6776 2874 6792 2894
rect 6812 2892 6866 2894
rect 6812 2874 6837 2892
rect 6776 2872 6837 2874
rect 6857 2872 6866 2892
rect 6776 2866 6866 2872
rect 6789 2812 6826 2813
rect 6885 2812 6922 2813
rect 6941 2812 6977 2922
rect 7164 2901 7195 2922
rect 7676 2911 7679 2931
rect 7699 2911 8094 2931
rect 8123 2912 8310 2936
rect 7160 2900 7195 2901
rect 7038 2890 7195 2900
rect 7038 2870 7055 2890
rect 7075 2870 7195 2890
rect 7038 2863 7195 2870
rect 7262 2893 7411 2901
rect 7262 2873 7273 2893
rect 7293 2873 7332 2893
rect 7352 2873 7411 2893
rect 7262 2866 7411 2873
rect 8055 2886 8094 2911
rect 8440 2886 8492 3075
rect 8055 2868 8494 2886
rect 7262 2865 7303 2866
rect 6996 2812 7033 2813
rect 6689 2803 6827 2812
rect 6689 2783 6798 2803
rect 6818 2783 6827 2803
rect 6689 2776 6827 2783
rect 6885 2803 7033 2812
rect 6885 2783 6894 2803
rect 6914 2783 7004 2803
rect 7024 2783 7033 2803
rect 6689 2774 6785 2776
rect 6885 2773 7033 2783
rect 7092 2803 7129 2813
rect 7092 2783 7100 2803
rect 7120 2783 7129 2803
rect 6941 2772 6977 2773
rect 6789 2713 6826 2714
rect 7092 2713 7129 2783
rect 7164 2812 7195 2863
rect 8055 2850 8455 2868
rect 8473 2850 8494 2868
rect 8055 2844 8494 2850
rect 8061 2840 8494 2844
rect 8440 2838 8492 2840
rect 7214 2812 7251 2813
rect 7164 2803 7251 2812
rect 7164 2783 7222 2803
rect 7242 2783 7251 2803
rect 7164 2773 7251 2783
rect 7310 2803 7347 2813
rect 7310 2783 7318 2803
rect 7338 2783 7347 2803
rect 7164 2772 7195 2773
rect 6788 2712 7129 2713
rect 7310 2712 7347 2783
rect 8443 2773 8480 2778
rect 6713 2707 7129 2712
rect 6713 2687 6716 2707
rect 6736 2687 7129 2707
rect 7160 2688 7347 2712
rect 8434 2769 8481 2773
rect 8434 2751 8453 2769
rect 8471 2751 8481 2769
rect 8434 2703 8481 2751
rect 8058 2700 8481 2703
rect 6933 2686 6998 2687
rect 8036 2670 8481 2700
rect 7129 2654 7169 2662
rect 7129 2632 7137 2654
rect 7161 2632 7169 2654
rect 6734 2403 6771 2409
rect 6734 2384 6742 2403
rect 6763 2384 6771 2403
rect 6734 2376 6771 2384
rect 6434 2255 6441 2277
rect 6465 2255 6473 2277
rect 6434 2249 6473 2255
rect 5964 2244 6004 2246
rect 6130 2245 6298 2246
rect 6232 2244 6269 2245
rect 5198 2228 5336 2237
rect 4992 2227 5029 2228
rect 4722 2174 4763 2175
rect 4496 2153 4548 2171
rect 4614 2167 4763 2174
rect 4064 2133 4104 2143
rect 4614 2147 4673 2167
rect 4693 2147 4732 2167
rect 4752 2147 4763 2167
rect 4614 2139 4763 2147
rect 4830 2170 4987 2177
rect 4830 2150 4950 2170
rect 4970 2150 4987 2170
rect 4830 2140 4987 2150
rect 4830 2139 4865 2140
rect 3894 2116 3932 2125
rect 4830 2118 4861 2139
rect 5048 2118 5084 2228
rect 5103 2227 5140 2228
rect 5199 2227 5236 2228
rect 5159 2168 5249 2174
rect 5159 2148 5168 2168
rect 5188 2166 5249 2168
rect 5188 2148 5213 2166
rect 5159 2146 5213 2148
rect 5233 2146 5249 2166
rect 5159 2140 5249 2146
rect 4673 2117 4710 2118
rect 3894 2115 3931 2116
rect 3355 2087 3445 2093
rect 3355 2067 3371 2087
rect 3391 2085 3445 2087
rect 3391 2067 3416 2085
rect 3355 2065 3416 2067
rect 3436 2065 3445 2085
rect 3355 2059 3445 2065
rect 3368 2005 3405 2006
rect 3464 2005 3501 2006
rect 3520 2005 3556 2115
rect 3743 2094 3774 2115
rect 4672 2108 4710 2117
rect 3739 2093 3774 2094
rect 3617 2083 3774 2093
rect 3617 2063 3634 2083
rect 3654 2063 3774 2083
rect 3617 2056 3774 2063
rect 3841 2086 3990 2094
rect 3841 2066 3852 2086
rect 3872 2066 3911 2086
rect 3931 2066 3990 2086
rect 4500 2090 4540 2100
rect 3841 2059 3990 2066
rect 4056 2062 4108 2080
rect 3841 2058 3882 2059
rect 3575 2005 3612 2006
rect 3268 1996 3406 2005
rect 2740 1985 2773 1987
rect 2369 1973 2816 1985
rect 1601 1851 1769 1853
rect 1325 1825 1769 1851
rect 835 1803 973 1812
rect 629 1802 666 1803
rect 126 1748 163 1751
rect 359 1749 400 1750
rect 251 1742 400 1749
rect 251 1722 310 1742
rect 330 1722 369 1742
rect 389 1722 400 1742
rect 251 1714 400 1722
rect 467 1745 624 1752
rect 467 1725 587 1745
rect 607 1725 624 1745
rect 467 1715 624 1725
rect 467 1714 502 1715
rect 467 1693 498 1714
rect 685 1693 721 1803
rect 740 1802 777 1803
rect 836 1802 873 1803
rect 796 1743 886 1749
rect 796 1723 805 1743
rect 825 1741 886 1743
rect 825 1723 850 1741
rect 796 1721 850 1723
rect 870 1721 886 1741
rect 796 1715 886 1721
rect 310 1692 347 1693
rect 123 1684 160 1686
rect 123 1676 165 1684
rect 123 1658 133 1676
rect 151 1658 165 1676
rect 123 1649 165 1658
rect 309 1683 347 1692
rect 309 1663 318 1683
rect 338 1663 347 1683
rect 309 1655 347 1663
rect 413 1687 498 1693
rect 528 1692 565 1693
rect 413 1667 421 1687
rect 441 1667 498 1687
rect 413 1659 498 1667
rect 527 1683 565 1692
rect 527 1663 536 1683
rect 556 1663 565 1683
rect 413 1658 449 1659
rect 527 1655 565 1663
rect 631 1691 775 1693
rect 631 1687 683 1691
rect 631 1667 639 1687
rect 659 1671 683 1687
rect 703 1687 775 1691
rect 703 1671 747 1687
rect 659 1667 747 1671
rect 767 1667 775 1687
rect 631 1659 775 1667
rect 631 1658 667 1659
rect 739 1658 775 1659
rect 841 1692 878 1693
rect 841 1691 879 1692
rect 841 1683 905 1691
rect 841 1663 850 1683
rect 870 1669 905 1683
rect 925 1669 928 1689
rect 870 1664 928 1669
rect 870 1663 905 1664
rect 124 1624 165 1649
rect 310 1624 347 1655
rect 528 1624 565 1655
rect 841 1651 905 1663
rect 945 1625 972 1803
rect 124 1597 173 1624
rect 309 1598 358 1624
rect 527 1623 608 1624
rect 804 1623 972 1625
rect 527 1598 972 1623
rect 528 1597 972 1598
rect 126 1564 173 1597
rect 529 1564 569 1597
rect 804 1596 972 1597
rect 1435 1601 1475 1825
rect 1601 1824 1769 1825
rect 2372 1959 2816 1973
rect 2372 1957 2540 1959
rect 2372 1779 2399 1957
rect 2439 1919 2503 1931
rect 2779 1927 2816 1959
rect 2842 1958 3033 1980
rect 3268 1976 3377 1996
rect 3397 1976 3406 1996
rect 3268 1969 3406 1976
rect 3464 1996 3612 2005
rect 3464 1976 3473 1996
rect 3493 1976 3583 1996
rect 3603 1976 3612 1996
rect 3268 1967 3364 1969
rect 3464 1966 3612 1976
rect 3671 1996 3708 2006
rect 3671 1976 3679 1996
rect 3699 1976 3708 1996
rect 3520 1965 3556 1966
rect 2997 1956 3033 1958
rect 2997 1927 3034 1956
rect 2439 1918 2474 1919
rect 2416 1913 2474 1918
rect 2416 1893 2419 1913
rect 2439 1899 2474 1913
rect 2494 1899 2503 1919
rect 2439 1891 2503 1899
rect 2465 1890 2503 1891
rect 2466 1889 2503 1890
rect 2569 1923 2605 1924
rect 2677 1923 2713 1924
rect 2569 1915 2713 1923
rect 2569 1895 2577 1915
rect 2597 1913 2685 1915
rect 2597 1895 2630 1913
rect 2569 1894 2630 1895
rect 2651 1895 2685 1913
rect 2705 1895 2713 1915
rect 2651 1894 2713 1895
rect 2569 1889 2713 1894
rect 2779 1919 2817 1927
rect 2895 1923 2931 1924
rect 2779 1899 2788 1919
rect 2808 1899 2817 1919
rect 2779 1890 2817 1899
rect 2846 1915 2931 1923
rect 2846 1895 2903 1915
rect 2923 1895 2931 1915
rect 2779 1889 2816 1890
rect 2846 1889 2931 1895
rect 2997 1919 3035 1927
rect 2997 1899 3006 1919
rect 3026 1899 3035 1919
rect 3671 1909 3708 1976
rect 3743 2005 3774 2056
rect 4056 2044 4074 2062
rect 4092 2044 4108 2062
rect 3793 2005 3830 2006
rect 3743 1996 3830 2005
rect 3743 1976 3801 1996
rect 3821 1976 3830 1996
rect 3743 1966 3830 1976
rect 3889 1996 3926 2006
rect 3889 1976 3897 1996
rect 3917 1976 3926 1996
rect 3743 1965 3774 1966
rect 3368 1906 3405 1907
rect 3671 1906 3710 1909
rect 3367 1905 3710 1906
rect 3889 1905 3926 1976
rect 2997 1890 3035 1899
rect 3292 1900 3710 1905
rect 2997 1889 3034 1890
rect 2458 1861 2548 1867
rect 2458 1841 2474 1861
rect 2494 1859 2548 1861
rect 2494 1841 2519 1859
rect 2458 1839 2519 1841
rect 2539 1839 2548 1859
rect 2458 1833 2548 1839
rect 2471 1779 2508 1780
rect 2567 1779 2604 1780
rect 2623 1779 2659 1889
rect 2846 1868 2877 1889
rect 3292 1880 3295 1900
rect 3315 1880 3710 1900
rect 3739 1881 3926 1905
rect 2842 1867 2877 1868
rect 2720 1857 2877 1867
rect 2720 1837 2737 1857
rect 2757 1837 2877 1857
rect 2720 1830 2877 1837
rect 2944 1860 3093 1868
rect 2944 1840 2955 1860
rect 2975 1840 3014 1860
rect 3034 1840 3093 1860
rect 2944 1833 3093 1840
rect 3671 1855 3710 1880
rect 4056 1855 4108 2044
rect 4500 2072 4510 2090
rect 4528 2072 4540 2090
rect 4672 2088 4681 2108
rect 4701 2088 4710 2108
rect 4672 2080 4710 2088
rect 4776 2112 4861 2118
rect 4891 2117 4928 2118
rect 4776 2092 4784 2112
rect 4804 2092 4861 2112
rect 4776 2084 4861 2092
rect 4890 2108 4928 2117
rect 4890 2088 4899 2108
rect 4919 2088 4928 2108
rect 4776 2083 4812 2084
rect 4890 2080 4928 2088
rect 4994 2112 5138 2118
rect 4994 2092 5002 2112
rect 5022 2092 5055 2112
rect 5075 2092 5110 2112
rect 5130 2092 5138 2112
rect 4994 2084 5138 2092
rect 4994 2083 5030 2084
rect 5102 2083 5138 2084
rect 5204 2117 5241 2118
rect 5204 2116 5242 2117
rect 5204 2108 5268 2116
rect 5204 2088 5213 2108
rect 5233 2094 5268 2108
rect 5288 2094 5291 2114
rect 5233 2089 5291 2094
rect 5233 2088 5268 2089
rect 4500 2016 4540 2072
rect 4673 2051 4710 2080
rect 4674 2049 4710 2051
rect 4674 2027 4865 2049
rect 4891 2048 4928 2080
rect 5204 2076 5268 2088
rect 5308 2050 5335 2228
rect 5167 2048 5335 2050
rect 4891 2038 5335 2048
rect 5476 2144 5663 2168
rect 5694 2149 6087 2169
rect 6107 2149 6110 2169
rect 5694 2144 6110 2149
rect 5476 2073 5513 2144
rect 5694 2143 6035 2144
rect 5628 2083 5659 2084
rect 5476 2053 5485 2073
rect 5505 2053 5513 2073
rect 5476 2043 5513 2053
rect 5572 2073 5659 2083
rect 5572 2053 5581 2073
rect 5601 2053 5659 2073
rect 5572 2044 5659 2053
rect 5572 2043 5609 2044
rect 4497 2011 4540 2016
rect 4888 2022 5335 2038
rect 4888 2016 4916 2022
rect 5167 2021 5335 2022
rect 4497 2008 4647 2011
rect 4888 2008 4915 2016
rect 4497 2006 4915 2008
rect 4497 1988 4506 2006
rect 4524 1988 4915 2006
rect 5628 1993 5659 2044
rect 5694 2073 5731 2143
rect 5997 2142 6034 2143
rect 6235 2085 6268 2244
rect 5846 2083 5882 2084
rect 5694 2053 5703 2073
rect 5723 2053 5731 2073
rect 5694 2043 5731 2053
rect 5790 2073 5938 2083
rect 6038 2080 6134 2082
rect 5790 2053 5799 2073
rect 5819 2053 5909 2073
rect 5929 2053 5938 2073
rect 5790 2044 5938 2053
rect 5996 2073 6134 2080
rect 5996 2053 6005 2073
rect 6025 2053 6134 2073
rect 6235 2081 6271 2085
rect 6235 2063 6244 2081
rect 6266 2063 6271 2081
rect 6235 2057 6271 2063
rect 5996 2044 6134 2053
rect 5790 2043 5827 2044
rect 5520 1990 5561 1991
rect 4497 1985 4915 1988
rect 4497 1979 4540 1985
rect 4500 1976 4540 1979
rect 5412 1983 5561 1990
rect 4897 1967 4937 1968
rect 4608 1950 4937 1967
rect 5412 1963 5471 1983
rect 5491 1963 5530 1983
rect 5550 1963 5561 1983
rect 5412 1955 5561 1963
rect 5628 1986 5785 1993
rect 5628 1966 5748 1986
rect 5768 1966 5785 1986
rect 5628 1956 5785 1966
rect 5628 1955 5663 1956
rect 4492 1907 4535 1918
rect 4492 1889 4504 1907
rect 4522 1889 4535 1907
rect 4492 1863 4535 1889
rect 4608 1863 4635 1950
rect 4897 1941 4937 1950
rect 3671 1837 4110 1855
rect 2944 1832 2985 1833
rect 2678 1779 2715 1780
rect 2371 1770 2509 1779
rect 2371 1750 2480 1770
rect 2500 1750 2509 1770
rect 2371 1743 2509 1750
rect 2567 1770 2715 1779
rect 2567 1750 2576 1770
rect 2596 1750 2686 1770
rect 2706 1750 2715 1770
rect 2371 1741 2467 1743
rect 2567 1740 2715 1750
rect 2774 1770 2811 1780
rect 2774 1750 2782 1770
rect 2802 1750 2811 1770
rect 2623 1739 2659 1740
rect 2471 1680 2508 1681
rect 2774 1680 2811 1750
rect 2846 1779 2877 1830
rect 3671 1819 4071 1837
rect 4089 1819 4110 1837
rect 3671 1813 4110 1819
rect 3677 1809 4110 1813
rect 4492 1842 4635 1863
rect 4679 1915 4713 1931
rect 4897 1921 5290 1941
rect 5310 1921 5313 1941
rect 5628 1934 5659 1955
rect 5846 1934 5882 2044
rect 5901 2043 5938 2044
rect 5997 2043 6034 2044
rect 5957 1984 6047 1990
rect 5957 1964 5966 1984
rect 5986 1982 6047 1984
rect 5986 1964 6011 1982
rect 5957 1962 6011 1964
rect 6031 1962 6047 1982
rect 5957 1956 6047 1962
rect 5471 1933 5508 1934
rect 4897 1916 5313 1921
rect 5470 1924 5508 1933
rect 4897 1915 5238 1916
rect 4679 1845 4716 1915
rect 4831 1855 4862 1856
rect 4492 1840 4629 1842
rect 4056 1807 4108 1809
rect 4492 1798 4535 1840
rect 4679 1825 4688 1845
rect 4708 1825 4716 1845
rect 4679 1815 4716 1825
rect 4775 1845 4862 1855
rect 4775 1825 4784 1845
rect 4804 1825 4862 1845
rect 4775 1816 4862 1825
rect 4775 1815 4812 1816
rect 4490 1788 4535 1798
rect 2896 1779 2933 1780
rect 2846 1770 2933 1779
rect 2846 1750 2904 1770
rect 2924 1750 2933 1770
rect 2846 1740 2933 1750
rect 2992 1770 3029 1780
rect 2992 1750 3000 1770
rect 3020 1750 3029 1770
rect 4490 1770 4499 1788
rect 4517 1770 4535 1788
rect 4490 1764 4535 1770
rect 4831 1765 4862 1816
rect 4897 1845 4934 1915
rect 5200 1914 5237 1915
rect 5470 1904 5479 1924
rect 5499 1904 5508 1924
rect 5470 1896 5508 1904
rect 5574 1928 5659 1934
rect 5689 1933 5726 1934
rect 5574 1908 5582 1928
rect 5602 1908 5659 1928
rect 5574 1900 5659 1908
rect 5688 1924 5726 1933
rect 5688 1904 5697 1924
rect 5717 1904 5726 1924
rect 5574 1899 5610 1900
rect 5688 1896 5726 1904
rect 5792 1928 5936 1934
rect 5792 1908 5800 1928
rect 5820 1909 5852 1928
rect 5873 1909 5908 1928
rect 5820 1908 5908 1909
rect 5928 1908 5936 1928
rect 5792 1900 5936 1908
rect 5792 1899 5828 1900
rect 5900 1899 5936 1900
rect 6002 1933 6039 1934
rect 6002 1932 6040 1933
rect 6002 1924 6066 1932
rect 6002 1904 6011 1924
rect 6031 1910 6066 1924
rect 6086 1910 6089 1930
rect 6031 1905 6089 1910
rect 6031 1904 6066 1905
rect 5471 1867 5508 1896
rect 5472 1865 5508 1867
rect 5049 1855 5085 1856
rect 4897 1825 4906 1845
rect 4926 1825 4934 1845
rect 4897 1815 4934 1825
rect 4993 1845 5141 1855
rect 5241 1852 5337 1854
rect 4993 1825 5002 1845
rect 5022 1825 5112 1845
rect 5132 1825 5141 1845
rect 4993 1816 5141 1825
rect 5199 1845 5337 1852
rect 5199 1825 5208 1845
rect 5228 1825 5337 1845
rect 5472 1843 5663 1865
rect 5689 1864 5726 1896
rect 6002 1892 6066 1904
rect 6106 1866 6133 2044
rect 6738 2043 6771 2376
rect 6835 2408 7003 2409
rect 7129 2408 7169 2632
rect 7632 2636 7800 2637
rect 8036 2636 8077 2670
rect 8434 2649 8481 2670
rect 7632 2626 8077 2636
rect 8149 2634 8292 2635
rect 7632 2610 8076 2626
rect 7632 2608 7800 2610
rect 7996 2609 8076 2610
rect 8149 2609 8294 2634
rect 8436 2609 8481 2649
rect 7632 2430 7659 2608
rect 7699 2570 7763 2582
rect 8039 2578 8076 2609
rect 8257 2578 8294 2609
rect 8439 2602 8481 2609
rect 7699 2569 7734 2570
rect 7676 2564 7734 2569
rect 7676 2544 7679 2564
rect 7699 2550 7734 2564
rect 7754 2550 7763 2570
rect 7699 2542 7763 2550
rect 7725 2541 7763 2542
rect 7726 2540 7763 2541
rect 7829 2574 7865 2575
rect 7937 2574 7973 2575
rect 7829 2566 7973 2574
rect 7829 2546 7837 2566
rect 7857 2562 7945 2566
rect 7857 2546 7901 2562
rect 7829 2542 7901 2546
rect 7921 2546 7945 2562
rect 7965 2546 7973 2566
rect 7921 2542 7973 2546
rect 7829 2540 7973 2542
rect 8039 2570 8077 2578
rect 8155 2574 8191 2575
rect 8039 2550 8048 2570
rect 8068 2550 8077 2570
rect 8039 2541 8077 2550
rect 8106 2566 8191 2574
rect 8106 2546 8163 2566
rect 8183 2546 8191 2566
rect 8039 2540 8076 2541
rect 8106 2540 8191 2546
rect 8257 2570 8295 2578
rect 8257 2550 8266 2570
rect 8286 2550 8295 2570
rect 8257 2541 8295 2550
rect 8439 2575 8482 2602
rect 8439 2557 8453 2575
rect 8471 2557 8482 2575
rect 8439 2549 8482 2557
rect 8444 2547 8482 2549
rect 8257 2540 8294 2541
rect 7718 2512 7808 2518
rect 7718 2492 7734 2512
rect 7754 2510 7808 2512
rect 7754 2492 7779 2510
rect 7718 2490 7779 2492
rect 7799 2490 7808 2510
rect 7718 2484 7808 2490
rect 7731 2430 7768 2431
rect 7827 2430 7864 2431
rect 7883 2430 7919 2540
rect 8106 2519 8137 2540
rect 8102 2518 8137 2519
rect 7980 2508 8137 2518
rect 7980 2488 7997 2508
rect 8017 2488 8137 2508
rect 7980 2481 8137 2488
rect 8204 2511 8353 2519
rect 8204 2491 8215 2511
rect 8235 2491 8274 2511
rect 8294 2491 8353 2511
rect 8204 2484 8353 2491
rect 8204 2483 8245 2484
rect 8441 2482 8478 2485
rect 7938 2430 7975 2431
rect 7631 2421 7769 2430
rect 6835 2382 7279 2408
rect 6835 2380 7003 2382
rect 6835 2202 6862 2380
rect 6902 2342 6966 2354
rect 7242 2350 7279 2382
rect 7305 2381 7496 2403
rect 7631 2401 7740 2421
rect 7760 2401 7769 2421
rect 7631 2394 7769 2401
rect 7827 2421 7975 2430
rect 7827 2401 7836 2421
rect 7856 2401 7946 2421
rect 7966 2401 7975 2421
rect 7631 2392 7727 2394
rect 7827 2391 7975 2401
rect 8034 2421 8071 2431
rect 8034 2401 8042 2421
rect 8062 2401 8071 2421
rect 7883 2390 7919 2391
rect 7460 2379 7496 2381
rect 7460 2350 7497 2379
rect 6902 2341 6937 2342
rect 6879 2336 6937 2341
rect 6879 2316 6882 2336
rect 6902 2322 6937 2336
rect 6957 2322 6966 2342
rect 6902 2316 6966 2322
rect 6879 2314 6966 2316
rect 6879 2310 6906 2314
rect 6928 2313 6966 2314
rect 6929 2312 6966 2313
rect 7032 2346 7068 2347
rect 7140 2346 7176 2347
rect 7032 2339 7176 2346
rect 7032 2338 7094 2339
rect 7032 2318 7040 2338
rect 7060 2321 7094 2338
rect 7113 2338 7176 2339
rect 7113 2321 7148 2338
rect 7060 2318 7148 2321
rect 7168 2318 7176 2338
rect 7032 2312 7176 2318
rect 7242 2342 7280 2350
rect 7358 2346 7394 2347
rect 7242 2322 7251 2342
rect 7271 2322 7280 2342
rect 7242 2313 7280 2322
rect 7309 2338 7394 2346
rect 7309 2318 7366 2338
rect 7386 2318 7394 2338
rect 7242 2312 7279 2313
rect 7309 2312 7394 2318
rect 7460 2342 7498 2350
rect 7460 2322 7469 2342
rect 7489 2322 7498 2342
rect 7731 2331 7768 2332
rect 8034 2331 8071 2401
rect 8106 2430 8137 2481
rect 8433 2476 8478 2482
rect 8433 2458 8451 2476
rect 8469 2458 8478 2476
rect 8433 2448 8478 2458
rect 8156 2430 8193 2431
rect 8106 2421 8193 2430
rect 8106 2401 8164 2421
rect 8184 2401 8193 2421
rect 8106 2391 8193 2401
rect 8252 2421 8289 2431
rect 8252 2401 8260 2421
rect 8280 2401 8289 2421
rect 8433 2406 8476 2448
rect 8339 2404 8476 2406
rect 8106 2390 8137 2391
rect 8252 2331 8289 2401
rect 7730 2330 8071 2331
rect 7460 2313 7498 2322
rect 7655 2325 8071 2330
rect 7460 2312 7497 2313
rect 6921 2284 7011 2290
rect 6921 2264 6937 2284
rect 6957 2282 7011 2284
rect 6957 2264 6982 2282
rect 6921 2262 6982 2264
rect 7002 2262 7011 2282
rect 6921 2256 7011 2262
rect 6934 2202 6971 2203
rect 7030 2202 7067 2203
rect 7086 2202 7122 2312
rect 7309 2291 7340 2312
rect 7655 2305 7658 2325
rect 7678 2305 8071 2325
rect 8255 2315 8289 2331
rect 8333 2383 8476 2404
rect 8031 2296 8071 2305
rect 8333 2296 8360 2383
rect 8433 2357 8476 2383
rect 8433 2339 8446 2357
rect 8464 2339 8476 2357
rect 8433 2328 8476 2339
rect 7305 2290 7340 2291
rect 7183 2280 7340 2290
rect 7183 2260 7200 2280
rect 7220 2260 7340 2280
rect 7183 2253 7340 2260
rect 7407 2283 7553 2291
rect 7407 2263 7418 2283
rect 7438 2263 7477 2283
rect 7497 2263 7553 2283
rect 8031 2279 8360 2296
rect 8031 2278 8071 2279
rect 7407 2256 7553 2263
rect 8428 2267 8468 2270
rect 8428 2261 8471 2267
rect 8053 2258 8471 2261
rect 7407 2255 7448 2256
rect 7141 2202 7178 2203
rect 6834 2193 6972 2202
rect 6834 2173 6943 2193
rect 6963 2173 6972 2193
rect 6834 2166 6972 2173
rect 7030 2193 7178 2202
rect 7030 2173 7039 2193
rect 7059 2173 7149 2193
rect 7169 2173 7178 2193
rect 6834 2164 6930 2166
rect 7030 2163 7178 2173
rect 7237 2193 7274 2203
rect 7237 2173 7245 2193
rect 7265 2173 7274 2193
rect 7086 2162 7122 2163
rect 6934 2103 6971 2104
rect 7237 2103 7274 2173
rect 7309 2202 7340 2253
rect 8053 2240 8444 2258
rect 8462 2240 8471 2258
rect 8053 2238 8471 2240
rect 8053 2230 8080 2238
rect 8321 2235 8471 2238
rect 7633 2224 7801 2225
rect 8052 2224 8080 2230
rect 7633 2208 8080 2224
rect 8428 2230 8471 2235
rect 7359 2202 7396 2203
rect 7309 2193 7396 2202
rect 7309 2173 7367 2193
rect 7387 2173 7396 2193
rect 7309 2163 7396 2173
rect 7455 2193 7492 2203
rect 7455 2173 7463 2193
rect 7483 2173 7492 2193
rect 7309 2162 7340 2163
rect 6933 2102 7274 2103
rect 7455 2102 7492 2173
rect 6858 2097 7274 2102
rect 6858 2077 6861 2097
rect 6881 2077 7274 2097
rect 7305 2078 7492 2102
rect 7633 2198 8077 2208
rect 7633 2196 7801 2198
rect 6733 1998 6775 2043
rect 7633 2018 7660 2196
rect 7700 2158 7764 2170
rect 8040 2166 8077 2198
rect 8103 2197 8294 2219
rect 8258 2195 8294 2197
rect 8258 2166 8295 2195
rect 8428 2174 8468 2230
rect 7700 2157 7735 2158
rect 7677 2152 7735 2157
rect 7677 2132 7680 2152
rect 7700 2138 7735 2152
rect 7755 2138 7764 2158
rect 7700 2130 7764 2138
rect 7726 2129 7764 2130
rect 7727 2128 7764 2129
rect 7830 2162 7866 2163
rect 7938 2162 7974 2163
rect 7830 2154 7974 2162
rect 7830 2134 7838 2154
rect 7858 2134 7893 2154
rect 7913 2134 7946 2154
rect 7966 2134 7974 2154
rect 7830 2128 7974 2134
rect 8040 2158 8078 2166
rect 8156 2162 8192 2163
rect 8040 2138 8049 2158
rect 8069 2138 8078 2158
rect 8040 2129 8078 2138
rect 8107 2154 8192 2162
rect 8107 2134 8164 2154
rect 8184 2134 8192 2154
rect 8040 2128 8077 2129
rect 8107 2128 8192 2134
rect 8258 2158 8296 2166
rect 8258 2138 8267 2158
rect 8287 2138 8296 2158
rect 8428 2156 8440 2174
rect 8458 2156 8468 2174
rect 8428 2146 8468 2156
rect 8258 2129 8296 2138
rect 8258 2128 8295 2129
rect 7719 2100 7809 2106
rect 7719 2080 7735 2100
rect 7755 2098 7809 2100
rect 7755 2080 7780 2098
rect 7719 2078 7780 2080
rect 7800 2078 7809 2098
rect 7719 2072 7809 2078
rect 7732 2018 7769 2019
rect 7828 2018 7865 2019
rect 7884 2018 7920 2128
rect 8107 2107 8138 2128
rect 8103 2106 8138 2107
rect 7981 2096 8138 2106
rect 7981 2076 7998 2096
rect 8018 2076 8138 2096
rect 7981 2069 8138 2076
rect 8205 2099 8354 2107
rect 8205 2079 8216 2099
rect 8236 2079 8275 2099
rect 8295 2079 8354 2099
rect 8205 2072 8354 2079
rect 8420 2075 8472 2093
rect 8205 2071 8246 2072
rect 7939 2018 7976 2019
rect 7632 2009 7770 2018
rect 7104 1998 7137 2000
rect 6733 1986 7180 1998
rect 5965 1864 6133 1866
rect 5689 1838 6133 1864
rect 5199 1816 5337 1825
rect 4993 1815 5030 1816
rect 4490 1761 4527 1764
rect 4723 1762 4764 1763
rect 2846 1739 2877 1740
rect 2470 1679 2811 1680
rect 2992 1679 3029 1750
rect 4615 1755 4764 1762
rect 4059 1742 4096 1747
rect 4050 1738 4097 1742
rect 4050 1720 4069 1738
rect 4087 1720 4097 1738
rect 4615 1735 4674 1755
rect 4694 1735 4733 1755
rect 4753 1735 4764 1755
rect 4615 1727 4764 1735
rect 4831 1758 4988 1765
rect 4831 1738 4951 1758
rect 4971 1738 4988 1758
rect 4831 1728 4988 1738
rect 4831 1727 4866 1728
rect 2395 1674 2811 1679
rect 2395 1654 2398 1674
rect 2418 1654 2811 1674
rect 2842 1655 3029 1679
rect 3654 1677 3694 1682
rect 4050 1677 4097 1720
rect 4831 1706 4862 1727
rect 5049 1706 5085 1816
rect 5104 1815 5141 1816
rect 5200 1815 5237 1816
rect 5160 1756 5250 1762
rect 5160 1736 5169 1756
rect 5189 1754 5250 1756
rect 5189 1736 5214 1754
rect 5160 1734 5214 1736
rect 5234 1734 5250 1754
rect 5160 1728 5250 1734
rect 4674 1705 4711 1706
rect 3654 1638 4097 1677
rect 4487 1697 4524 1699
rect 4487 1689 4529 1697
rect 4487 1671 4497 1689
rect 4515 1671 4529 1689
rect 4487 1662 4529 1671
rect 4673 1696 4711 1705
rect 4673 1676 4682 1696
rect 4702 1676 4711 1696
rect 4673 1668 4711 1676
rect 4777 1700 4862 1706
rect 4892 1705 4929 1706
rect 4777 1680 4785 1700
rect 4805 1680 4862 1700
rect 4777 1672 4862 1680
rect 4891 1696 4929 1705
rect 4891 1676 4900 1696
rect 4920 1676 4929 1696
rect 4777 1671 4813 1672
rect 4891 1668 4929 1676
rect 4995 1704 5139 1706
rect 4995 1700 5047 1704
rect 4995 1680 5003 1700
rect 5023 1684 5047 1700
rect 5067 1700 5139 1704
rect 5067 1684 5111 1700
rect 5023 1680 5111 1684
rect 5131 1680 5139 1700
rect 4995 1672 5139 1680
rect 4995 1671 5031 1672
rect 5103 1671 5139 1672
rect 5205 1705 5242 1706
rect 5205 1704 5243 1705
rect 5205 1696 5269 1704
rect 5205 1676 5214 1696
rect 5234 1682 5269 1696
rect 5289 1682 5292 1702
rect 5234 1677 5292 1682
rect 5234 1676 5269 1677
rect 1435 1579 1443 1601
rect 1467 1579 1475 1601
rect 1435 1571 1475 1579
rect 2748 1623 2788 1631
rect 2748 1601 2756 1623
rect 2780 1601 2788 1623
rect 126 1525 569 1564
rect 126 1482 173 1525
rect 529 1520 569 1525
rect 1194 1523 1381 1547
rect 1412 1528 1805 1548
rect 1825 1528 1828 1548
rect 1412 1523 1828 1528
rect 126 1464 136 1482
rect 154 1464 173 1482
rect 126 1460 173 1464
rect 127 1455 164 1460
rect 1194 1452 1231 1523
rect 1412 1522 1753 1523
rect 1346 1462 1377 1463
rect 1194 1432 1203 1452
rect 1223 1432 1231 1452
rect 1194 1422 1231 1432
rect 1290 1452 1377 1462
rect 1290 1432 1299 1452
rect 1319 1432 1377 1452
rect 1290 1423 1377 1432
rect 1290 1422 1327 1423
rect 115 1393 167 1395
rect 113 1389 546 1393
rect 113 1383 552 1389
rect 113 1365 134 1383
rect 152 1365 552 1383
rect 1346 1372 1377 1423
rect 1412 1452 1449 1522
rect 1715 1521 1752 1522
rect 1564 1462 1600 1463
rect 1412 1432 1421 1452
rect 1441 1432 1449 1452
rect 1412 1422 1449 1432
rect 1508 1452 1656 1462
rect 1756 1459 1852 1461
rect 1508 1432 1517 1452
rect 1537 1432 1627 1452
rect 1647 1432 1656 1452
rect 1508 1423 1656 1432
rect 1714 1452 1852 1459
rect 1714 1432 1723 1452
rect 1743 1432 1852 1452
rect 1714 1423 1852 1432
rect 1508 1422 1545 1423
rect 1238 1369 1279 1370
rect 113 1347 552 1365
rect 115 1158 167 1347
rect 513 1322 552 1347
rect 1130 1362 1279 1369
rect 1130 1342 1189 1362
rect 1209 1342 1248 1362
rect 1268 1342 1279 1362
rect 1130 1334 1279 1342
rect 1346 1365 1503 1372
rect 1346 1345 1466 1365
rect 1486 1345 1503 1365
rect 1346 1335 1503 1345
rect 1346 1334 1381 1335
rect 297 1297 484 1321
rect 513 1302 908 1322
rect 928 1302 931 1322
rect 1346 1313 1377 1334
rect 1564 1313 1600 1423
rect 1619 1422 1656 1423
rect 1715 1422 1752 1423
rect 1675 1363 1765 1369
rect 1675 1343 1684 1363
rect 1704 1361 1765 1363
rect 1704 1343 1729 1361
rect 1675 1341 1729 1343
rect 1749 1341 1765 1361
rect 1675 1335 1765 1341
rect 1189 1312 1226 1313
rect 513 1297 931 1302
rect 1188 1303 1226 1312
rect 297 1226 334 1297
rect 513 1296 856 1297
rect 513 1293 552 1296
rect 818 1295 855 1296
rect 449 1236 480 1237
rect 297 1206 306 1226
rect 326 1206 334 1226
rect 297 1196 334 1206
rect 393 1226 480 1236
rect 393 1206 402 1226
rect 422 1206 480 1226
rect 393 1197 480 1206
rect 393 1196 430 1197
rect 115 1140 131 1158
rect 149 1140 167 1158
rect 449 1146 480 1197
rect 515 1226 552 1293
rect 1188 1283 1197 1303
rect 1217 1283 1226 1303
rect 1188 1275 1226 1283
rect 1292 1307 1377 1313
rect 1407 1312 1444 1313
rect 1292 1287 1300 1307
rect 1320 1287 1377 1307
rect 1292 1279 1377 1287
rect 1406 1303 1444 1312
rect 1406 1283 1415 1303
rect 1435 1283 1444 1303
rect 1292 1278 1328 1279
rect 1406 1275 1444 1283
rect 1510 1307 1654 1313
rect 1510 1287 1518 1307
rect 1538 1302 1626 1307
rect 1538 1287 1574 1302
rect 1510 1285 1574 1287
rect 1593 1287 1626 1302
rect 1646 1287 1654 1307
rect 1593 1285 1654 1287
rect 1510 1279 1654 1285
rect 1510 1278 1546 1279
rect 1618 1278 1654 1279
rect 1720 1312 1757 1313
rect 1720 1311 1758 1312
rect 1720 1303 1784 1311
rect 1720 1283 1729 1303
rect 1749 1289 1784 1303
rect 1804 1289 1807 1309
rect 1749 1284 1807 1289
rect 1749 1283 1784 1284
rect 1189 1246 1226 1275
rect 1190 1244 1226 1246
rect 667 1236 703 1237
rect 515 1206 524 1226
rect 544 1206 552 1226
rect 515 1196 552 1206
rect 611 1226 759 1236
rect 859 1233 955 1235
rect 611 1206 620 1226
rect 640 1206 730 1226
rect 750 1206 759 1226
rect 611 1197 759 1206
rect 817 1226 955 1233
rect 817 1206 826 1226
rect 846 1206 955 1226
rect 1190 1222 1381 1244
rect 1407 1243 1444 1275
rect 1720 1271 1784 1283
rect 1824 1245 1851 1423
rect 1683 1243 1851 1245
rect 1407 1229 1851 1243
rect 2454 1377 2622 1378
rect 2748 1377 2788 1601
rect 3251 1605 3419 1606
rect 3654 1605 3694 1638
rect 4050 1605 4097 1638
rect 4488 1637 4529 1662
rect 4674 1637 4711 1668
rect 4892 1637 4929 1668
rect 5205 1664 5269 1676
rect 5309 1638 5336 1816
rect 4488 1610 4537 1637
rect 4673 1611 4722 1637
rect 4891 1636 4972 1637
rect 5168 1636 5336 1638
rect 4891 1611 5336 1636
rect 4892 1610 5336 1611
rect 3251 1604 3695 1605
rect 3251 1579 3696 1604
rect 3251 1577 3419 1579
rect 3615 1578 3696 1579
rect 3865 1578 3914 1604
rect 4050 1578 4099 1605
rect 3251 1399 3278 1577
rect 3318 1539 3382 1551
rect 3658 1547 3695 1578
rect 3876 1547 3913 1578
rect 4058 1553 4099 1578
rect 4490 1577 4537 1610
rect 4893 1577 4933 1610
rect 5168 1609 5336 1610
rect 5799 1614 5839 1838
rect 5965 1837 6133 1838
rect 6736 1972 7180 1986
rect 6736 1970 6904 1972
rect 6736 1792 6763 1970
rect 6803 1932 6867 1944
rect 7143 1940 7180 1972
rect 7206 1971 7397 1993
rect 7632 1989 7741 2009
rect 7761 1989 7770 2009
rect 7632 1982 7770 1989
rect 7828 2009 7976 2018
rect 7828 1989 7837 2009
rect 7857 1989 7947 2009
rect 7967 1989 7976 2009
rect 7632 1980 7728 1982
rect 7828 1979 7976 1989
rect 8035 2009 8072 2019
rect 8035 1989 8043 2009
rect 8063 1989 8072 2009
rect 7884 1978 7920 1979
rect 7361 1969 7397 1971
rect 7361 1940 7398 1969
rect 6803 1931 6838 1932
rect 6780 1926 6838 1931
rect 6780 1906 6783 1926
rect 6803 1912 6838 1926
rect 6858 1912 6867 1932
rect 6803 1904 6867 1912
rect 6829 1903 6867 1904
rect 6830 1902 6867 1903
rect 6933 1936 6969 1937
rect 7041 1936 7077 1937
rect 6933 1928 7077 1936
rect 6933 1908 6941 1928
rect 6961 1926 7049 1928
rect 6961 1908 6994 1926
rect 6933 1907 6994 1908
rect 7015 1908 7049 1926
rect 7069 1908 7077 1928
rect 7015 1907 7077 1908
rect 6933 1902 7077 1907
rect 7143 1932 7181 1940
rect 7259 1936 7295 1937
rect 7143 1912 7152 1932
rect 7172 1912 7181 1932
rect 7143 1903 7181 1912
rect 7210 1928 7295 1936
rect 7210 1908 7267 1928
rect 7287 1908 7295 1928
rect 7143 1902 7180 1903
rect 7210 1902 7295 1908
rect 7361 1932 7399 1940
rect 7361 1912 7370 1932
rect 7390 1912 7399 1932
rect 8035 1922 8072 1989
rect 8107 2018 8138 2069
rect 8420 2057 8438 2075
rect 8456 2057 8472 2075
rect 8157 2018 8194 2019
rect 8107 2009 8194 2018
rect 8107 1989 8165 2009
rect 8185 1989 8194 2009
rect 8107 1979 8194 1989
rect 8253 2009 8290 2019
rect 8253 1989 8261 2009
rect 8281 1989 8290 2009
rect 8107 1978 8138 1979
rect 7732 1919 7769 1920
rect 8035 1919 8074 1922
rect 7731 1918 8074 1919
rect 8253 1918 8290 1989
rect 7361 1903 7399 1912
rect 7656 1913 8074 1918
rect 7361 1902 7398 1903
rect 6822 1874 6912 1880
rect 6822 1854 6838 1874
rect 6858 1872 6912 1874
rect 6858 1854 6883 1872
rect 6822 1852 6883 1854
rect 6903 1852 6912 1872
rect 6822 1846 6912 1852
rect 6835 1792 6872 1793
rect 6931 1792 6968 1793
rect 6987 1792 7023 1902
rect 7210 1881 7241 1902
rect 7656 1893 7659 1913
rect 7679 1893 8074 1913
rect 8103 1894 8290 1918
rect 7206 1880 7241 1881
rect 7084 1870 7241 1880
rect 7084 1850 7101 1870
rect 7121 1850 7241 1870
rect 7084 1843 7241 1850
rect 7308 1873 7457 1881
rect 7308 1853 7319 1873
rect 7339 1853 7378 1873
rect 7398 1853 7457 1873
rect 7308 1846 7457 1853
rect 8035 1868 8074 1893
rect 8420 1868 8472 2057
rect 8035 1850 8474 1868
rect 7308 1845 7349 1846
rect 7042 1792 7079 1793
rect 6735 1783 6873 1792
rect 6735 1763 6844 1783
rect 6864 1763 6873 1783
rect 6735 1756 6873 1763
rect 6931 1783 7079 1792
rect 6931 1763 6940 1783
rect 6960 1763 7050 1783
rect 7070 1763 7079 1783
rect 6735 1754 6831 1756
rect 6931 1753 7079 1763
rect 7138 1783 7175 1793
rect 7138 1763 7146 1783
rect 7166 1763 7175 1783
rect 6987 1752 7023 1753
rect 6835 1693 6872 1694
rect 7138 1693 7175 1763
rect 7210 1792 7241 1843
rect 8035 1832 8435 1850
rect 8453 1832 8474 1850
rect 8035 1826 8474 1832
rect 8041 1822 8474 1826
rect 8420 1820 8472 1822
rect 7260 1792 7297 1793
rect 7210 1783 7297 1792
rect 7210 1763 7268 1783
rect 7288 1763 7297 1783
rect 7210 1753 7297 1763
rect 7356 1783 7393 1793
rect 7356 1763 7364 1783
rect 7384 1763 7393 1783
rect 7210 1752 7241 1753
rect 6834 1692 7175 1693
rect 7356 1692 7393 1763
rect 8423 1755 8460 1760
rect 8414 1751 8461 1755
rect 8414 1733 8433 1751
rect 8451 1733 8461 1751
rect 6759 1687 7175 1692
rect 6759 1667 6762 1687
rect 6782 1667 7175 1687
rect 7206 1668 7393 1692
rect 8018 1690 8058 1695
rect 8414 1690 8461 1733
rect 8018 1651 8461 1690
rect 5799 1592 5807 1614
rect 5831 1592 5839 1614
rect 5799 1584 5839 1592
rect 7112 1636 7152 1644
rect 7112 1614 7120 1636
rect 7144 1614 7152 1636
rect 3318 1538 3353 1539
rect 3295 1533 3353 1538
rect 3295 1513 3298 1533
rect 3318 1519 3353 1533
rect 3373 1519 3382 1539
rect 3318 1511 3382 1519
rect 3344 1510 3382 1511
rect 3345 1509 3382 1510
rect 3448 1543 3484 1544
rect 3556 1543 3592 1544
rect 3448 1535 3592 1543
rect 3448 1515 3456 1535
rect 3476 1531 3564 1535
rect 3476 1515 3520 1531
rect 3448 1511 3520 1515
rect 3540 1515 3564 1531
rect 3584 1515 3592 1535
rect 3540 1511 3592 1515
rect 3448 1509 3592 1511
rect 3658 1539 3696 1547
rect 3774 1543 3810 1544
rect 3658 1519 3667 1539
rect 3687 1519 3696 1539
rect 3658 1510 3696 1519
rect 3725 1535 3810 1543
rect 3725 1515 3782 1535
rect 3802 1515 3810 1535
rect 3658 1509 3695 1510
rect 3725 1509 3810 1515
rect 3876 1539 3914 1547
rect 3876 1519 3885 1539
rect 3905 1519 3914 1539
rect 3876 1510 3914 1519
rect 4058 1544 4100 1553
rect 4058 1526 4072 1544
rect 4090 1526 4100 1544
rect 4058 1518 4100 1526
rect 4063 1516 4100 1518
rect 4490 1538 4933 1577
rect 3876 1509 3913 1510
rect 3337 1481 3427 1487
rect 3337 1461 3353 1481
rect 3373 1479 3427 1481
rect 3373 1461 3398 1479
rect 3337 1459 3398 1461
rect 3418 1459 3427 1479
rect 3337 1453 3427 1459
rect 3350 1399 3387 1400
rect 3446 1399 3483 1400
rect 3502 1399 3538 1509
rect 3725 1488 3756 1509
rect 4490 1495 4537 1538
rect 4893 1533 4933 1538
rect 5558 1536 5745 1560
rect 5776 1541 6169 1561
rect 6189 1541 6192 1561
rect 5776 1536 6192 1541
rect 3721 1487 3756 1488
rect 3599 1477 3756 1487
rect 3599 1457 3616 1477
rect 3636 1457 3756 1477
rect 3599 1450 3756 1457
rect 3823 1480 3972 1488
rect 3823 1460 3834 1480
rect 3854 1460 3893 1480
rect 3913 1460 3972 1480
rect 4490 1477 4500 1495
rect 4518 1477 4537 1495
rect 4490 1473 4537 1477
rect 4491 1468 4528 1473
rect 3823 1453 3972 1460
rect 5558 1465 5595 1536
rect 5776 1535 6117 1536
rect 5710 1475 5741 1476
rect 3823 1452 3864 1453
rect 4060 1451 4097 1454
rect 3557 1399 3594 1400
rect 3250 1390 3388 1399
rect 2454 1351 2898 1377
rect 2454 1349 2622 1351
rect 1407 1217 1854 1229
rect 1450 1215 1483 1217
rect 817 1197 955 1206
rect 611 1196 648 1197
rect 341 1143 382 1144
rect 115 1122 167 1140
rect 233 1136 382 1143
rect 233 1116 292 1136
rect 312 1116 351 1136
rect 371 1116 382 1136
rect 233 1108 382 1116
rect 449 1139 606 1146
rect 449 1119 569 1139
rect 589 1119 606 1139
rect 449 1109 606 1119
rect 449 1108 484 1109
rect 449 1087 480 1108
rect 667 1087 703 1197
rect 722 1196 759 1197
rect 818 1196 855 1197
rect 778 1137 868 1143
rect 778 1117 787 1137
rect 807 1135 868 1137
rect 807 1117 832 1135
rect 778 1115 832 1117
rect 852 1115 868 1135
rect 778 1109 868 1115
rect 292 1086 329 1087
rect 291 1077 329 1086
rect 119 1059 159 1069
rect 119 1041 129 1059
rect 147 1041 159 1059
rect 291 1057 300 1077
rect 320 1057 329 1077
rect 291 1049 329 1057
rect 395 1081 480 1087
rect 510 1086 547 1087
rect 395 1061 403 1081
rect 423 1061 480 1081
rect 395 1053 480 1061
rect 509 1077 547 1086
rect 509 1057 518 1077
rect 538 1057 547 1077
rect 395 1052 431 1053
rect 509 1049 547 1057
rect 613 1081 757 1087
rect 613 1061 621 1081
rect 641 1061 674 1081
rect 694 1061 729 1081
rect 749 1061 757 1081
rect 613 1053 757 1061
rect 613 1052 649 1053
rect 721 1052 757 1053
rect 823 1086 860 1087
rect 823 1085 861 1086
rect 823 1077 887 1085
rect 823 1057 832 1077
rect 852 1063 887 1077
rect 907 1063 910 1083
rect 852 1058 910 1063
rect 852 1057 887 1058
rect 119 985 159 1041
rect 292 1020 329 1049
rect 293 1018 329 1020
rect 293 996 484 1018
rect 510 1017 547 1049
rect 823 1045 887 1057
rect 927 1019 954 1197
rect 1812 1172 1854 1217
rect 786 1017 954 1019
rect 510 1007 954 1017
rect 1095 1113 1282 1137
rect 1313 1118 1706 1138
rect 1726 1118 1729 1138
rect 1313 1113 1729 1118
rect 1095 1042 1132 1113
rect 1313 1112 1654 1113
rect 1247 1052 1278 1053
rect 1095 1022 1104 1042
rect 1124 1022 1132 1042
rect 1095 1012 1132 1022
rect 1191 1042 1278 1052
rect 1191 1022 1200 1042
rect 1220 1022 1278 1042
rect 1191 1013 1278 1022
rect 1191 1012 1228 1013
rect 116 980 159 985
rect 507 991 954 1007
rect 507 985 535 991
rect 786 990 954 991
rect 116 977 266 980
rect 507 977 534 985
rect 116 975 534 977
rect 116 957 125 975
rect 143 957 534 975
rect 1247 962 1278 1013
rect 1313 1042 1350 1112
rect 1616 1111 1653 1112
rect 1465 1052 1501 1053
rect 1313 1022 1322 1042
rect 1342 1022 1350 1042
rect 1313 1012 1350 1022
rect 1409 1042 1557 1052
rect 1657 1049 1753 1051
rect 1409 1022 1418 1042
rect 1438 1022 1528 1042
rect 1548 1022 1557 1042
rect 1409 1013 1557 1022
rect 1615 1042 1753 1049
rect 1615 1022 1624 1042
rect 1644 1022 1753 1042
rect 1615 1013 1753 1022
rect 1409 1012 1446 1013
rect 1139 959 1180 960
rect 116 954 534 957
rect 116 948 159 954
rect 119 945 159 948
rect 1034 952 1180 959
rect 516 936 556 937
rect 227 919 556 936
rect 1034 932 1090 952
rect 1110 932 1149 952
rect 1169 932 1180 952
rect 1034 924 1180 932
rect 1247 955 1404 962
rect 1247 935 1367 955
rect 1387 935 1404 955
rect 1247 925 1404 935
rect 1247 924 1282 925
rect 111 876 154 887
rect 111 858 123 876
rect 141 858 154 876
rect 111 832 154 858
rect 227 832 254 919
rect 516 910 556 919
rect 111 811 254 832
rect 298 884 332 900
rect 516 890 909 910
rect 929 890 932 910
rect 1247 903 1278 924
rect 1465 903 1501 1013
rect 1520 1012 1557 1013
rect 1616 1012 1653 1013
rect 1576 953 1666 959
rect 1576 933 1585 953
rect 1605 951 1666 953
rect 1605 933 1630 951
rect 1576 931 1630 933
rect 1650 931 1666 951
rect 1576 925 1666 931
rect 1090 902 1127 903
rect 516 885 932 890
rect 1089 893 1127 902
rect 516 884 857 885
rect 298 814 335 884
rect 450 824 481 825
rect 111 809 248 811
rect 111 767 154 809
rect 298 794 307 814
rect 327 794 335 814
rect 298 784 335 794
rect 394 814 481 824
rect 394 794 403 814
rect 423 794 481 814
rect 394 785 481 794
rect 394 784 431 785
rect 109 757 154 767
rect 109 739 118 757
rect 136 739 154 757
rect 109 733 154 739
rect 450 734 481 785
rect 516 814 553 884
rect 819 883 856 884
rect 1089 873 1098 893
rect 1118 873 1127 893
rect 1089 865 1127 873
rect 1193 897 1278 903
rect 1308 902 1345 903
rect 1193 877 1201 897
rect 1221 877 1278 897
rect 1193 869 1278 877
rect 1307 893 1345 902
rect 1307 873 1316 893
rect 1336 873 1345 893
rect 1193 868 1229 869
rect 1307 865 1345 873
rect 1411 897 1555 903
rect 1411 877 1419 897
rect 1439 894 1527 897
rect 1439 877 1474 894
rect 1411 876 1474 877
rect 1493 877 1527 894
rect 1547 877 1555 897
rect 1493 876 1555 877
rect 1411 869 1555 876
rect 1411 868 1447 869
rect 1519 868 1555 869
rect 1621 902 1658 903
rect 1621 901 1659 902
rect 1681 901 1708 905
rect 1621 899 1708 901
rect 1621 893 1685 899
rect 1621 873 1630 893
rect 1650 879 1685 893
rect 1705 879 1708 899
rect 1650 874 1708 879
rect 1650 873 1685 874
rect 1090 836 1127 865
rect 1091 834 1127 836
rect 668 824 704 825
rect 516 794 525 814
rect 545 794 553 814
rect 516 784 553 794
rect 612 814 760 824
rect 860 821 956 823
rect 612 794 621 814
rect 641 794 731 814
rect 751 794 760 814
rect 612 785 760 794
rect 818 814 956 821
rect 818 794 827 814
rect 847 794 956 814
rect 1091 812 1282 834
rect 1308 833 1345 865
rect 1621 861 1685 873
rect 1725 835 1752 1013
rect 1584 833 1752 835
rect 1308 807 1752 833
rect 818 785 956 794
rect 612 784 649 785
rect 109 730 146 733
rect 342 731 383 732
rect 234 724 383 731
rect 234 704 293 724
rect 313 704 352 724
rect 372 704 383 724
rect 234 696 383 704
rect 450 727 607 734
rect 450 707 570 727
rect 590 707 607 727
rect 450 697 607 707
rect 450 696 485 697
rect 450 675 481 696
rect 668 675 704 785
rect 723 784 760 785
rect 819 784 856 785
rect 779 725 869 731
rect 779 705 788 725
rect 808 723 869 725
rect 808 705 833 723
rect 779 703 833 705
rect 853 703 869 723
rect 779 697 869 703
rect 293 674 330 675
rect 106 666 143 668
rect 106 658 148 666
rect 106 640 116 658
rect 134 640 148 658
rect 106 631 148 640
rect 292 665 330 674
rect 292 645 301 665
rect 321 645 330 665
rect 292 637 330 645
rect 396 669 481 675
rect 511 674 548 675
rect 396 649 404 669
rect 424 649 481 669
rect 396 641 481 649
rect 510 665 548 674
rect 510 645 519 665
rect 539 645 548 665
rect 396 640 432 641
rect 510 637 548 645
rect 614 673 758 675
rect 614 669 666 673
rect 614 649 622 669
rect 642 653 666 669
rect 686 669 758 673
rect 686 653 730 669
rect 642 649 730 653
rect 750 649 758 669
rect 614 641 758 649
rect 614 640 650 641
rect 722 640 758 641
rect 824 674 861 675
rect 824 673 862 674
rect 824 665 888 673
rect 824 645 833 665
rect 853 651 888 665
rect 908 651 911 671
rect 853 646 911 651
rect 853 645 888 646
rect 107 606 148 631
rect 293 606 330 637
rect 511 615 548 637
rect 824 633 888 645
rect 506 606 548 615
rect 928 607 955 785
rect 107 594 152 606
rect 103 536 152 594
rect 293 580 355 606
rect 506 605 591 606
rect 787 605 955 607
rect 506 579 955 605
rect 506 536 545 579
rect 787 578 955 579
rect 1418 583 1458 807
rect 1584 806 1752 807
rect 1816 839 1849 1172
rect 2454 1171 2481 1349
rect 2521 1311 2585 1323
rect 2861 1319 2898 1351
rect 2924 1350 3115 1372
rect 3250 1370 3359 1390
rect 3379 1370 3388 1390
rect 3250 1363 3388 1370
rect 3446 1390 3594 1399
rect 3446 1370 3455 1390
rect 3475 1370 3565 1390
rect 3585 1370 3594 1390
rect 3250 1361 3346 1363
rect 3446 1360 3594 1370
rect 3653 1390 3690 1400
rect 3653 1370 3661 1390
rect 3681 1370 3690 1390
rect 3502 1359 3538 1360
rect 3079 1348 3115 1350
rect 3079 1319 3116 1348
rect 2521 1310 2556 1311
rect 2498 1305 2556 1310
rect 2498 1285 2501 1305
rect 2521 1291 2556 1305
rect 2576 1291 2585 1311
rect 2521 1283 2585 1291
rect 2547 1282 2585 1283
rect 2548 1281 2585 1282
rect 2651 1315 2687 1316
rect 2759 1315 2795 1316
rect 2651 1307 2795 1315
rect 2651 1287 2659 1307
rect 2679 1306 2767 1307
rect 2679 1287 2714 1306
rect 2735 1287 2767 1306
rect 2787 1287 2795 1307
rect 2651 1281 2795 1287
rect 2861 1311 2899 1319
rect 2977 1315 3013 1316
rect 2861 1291 2870 1311
rect 2890 1291 2899 1311
rect 2861 1282 2899 1291
rect 2928 1307 3013 1315
rect 2928 1287 2985 1307
rect 3005 1287 3013 1307
rect 2861 1281 2898 1282
rect 2928 1281 3013 1287
rect 3079 1311 3117 1319
rect 3079 1291 3088 1311
rect 3108 1291 3117 1311
rect 3350 1300 3387 1301
rect 3653 1300 3690 1370
rect 3725 1399 3756 1450
rect 4052 1445 4097 1451
rect 4052 1427 4070 1445
rect 4088 1427 4097 1445
rect 5558 1445 5567 1465
rect 5587 1445 5595 1465
rect 5558 1435 5595 1445
rect 5654 1465 5741 1475
rect 5654 1445 5663 1465
rect 5683 1445 5741 1465
rect 5654 1436 5741 1445
rect 5654 1435 5691 1436
rect 4052 1417 4097 1427
rect 3775 1399 3812 1400
rect 3725 1390 3812 1399
rect 3725 1370 3783 1390
rect 3803 1370 3812 1390
rect 3725 1360 3812 1370
rect 3871 1390 3908 1400
rect 3871 1370 3879 1390
rect 3899 1370 3908 1390
rect 4052 1375 4095 1417
rect 4479 1406 4531 1408
rect 3958 1373 4095 1375
rect 3725 1359 3756 1360
rect 3871 1300 3908 1370
rect 3349 1299 3690 1300
rect 3079 1282 3117 1291
rect 3274 1294 3690 1299
rect 3079 1281 3116 1282
rect 2540 1253 2630 1259
rect 2540 1233 2556 1253
rect 2576 1251 2630 1253
rect 2576 1233 2601 1251
rect 2540 1231 2601 1233
rect 2621 1231 2630 1251
rect 2540 1225 2630 1231
rect 2553 1171 2590 1172
rect 2649 1171 2686 1172
rect 2705 1171 2741 1281
rect 2928 1260 2959 1281
rect 3274 1274 3277 1294
rect 3297 1274 3690 1294
rect 3874 1284 3908 1300
rect 3952 1352 4095 1373
rect 4477 1402 4910 1406
rect 4477 1396 4916 1402
rect 4477 1378 4498 1396
rect 4516 1378 4916 1396
rect 5710 1385 5741 1436
rect 5776 1465 5813 1535
rect 6079 1534 6116 1535
rect 5928 1475 5964 1476
rect 5776 1445 5785 1465
rect 5805 1445 5813 1465
rect 5776 1435 5813 1445
rect 5872 1465 6020 1475
rect 6120 1472 6216 1474
rect 5872 1445 5881 1465
rect 5901 1445 5991 1465
rect 6011 1445 6020 1465
rect 5872 1436 6020 1445
rect 6078 1465 6216 1472
rect 6078 1445 6087 1465
rect 6107 1445 6216 1465
rect 6078 1436 6216 1445
rect 5872 1435 5909 1436
rect 5602 1382 5643 1383
rect 4477 1360 4916 1378
rect 3650 1265 3690 1274
rect 3952 1265 3979 1352
rect 4052 1326 4095 1352
rect 4052 1308 4065 1326
rect 4083 1308 4095 1326
rect 4052 1297 4095 1308
rect 2924 1259 2959 1260
rect 2802 1249 2959 1259
rect 2802 1229 2819 1249
rect 2839 1229 2959 1249
rect 2802 1222 2959 1229
rect 3026 1252 3175 1260
rect 3026 1232 3037 1252
rect 3057 1232 3096 1252
rect 3116 1232 3175 1252
rect 3650 1248 3979 1265
rect 3650 1247 3690 1248
rect 3026 1225 3175 1232
rect 4047 1236 4087 1239
rect 4047 1230 4090 1236
rect 3672 1227 4090 1230
rect 3026 1224 3067 1225
rect 2760 1171 2797 1172
rect 2453 1162 2591 1171
rect 2453 1142 2562 1162
rect 2582 1142 2591 1162
rect 2453 1135 2591 1142
rect 2649 1162 2797 1171
rect 2649 1142 2658 1162
rect 2678 1142 2768 1162
rect 2788 1142 2797 1162
rect 2453 1133 2549 1135
rect 2649 1132 2797 1142
rect 2856 1162 2893 1172
rect 2856 1142 2864 1162
rect 2884 1142 2893 1162
rect 2705 1131 2741 1132
rect 2553 1072 2590 1073
rect 2856 1072 2893 1142
rect 2928 1171 2959 1222
rect 3672 1209 4063 1227
rect 4081 1209 4090 1227
rect 3672 1207 4090 1209
rect 3672 1199 3699 1207
rect 3940 1204 4090 1207
rect 3252 1193 3420 1194
rect 3671 1193 3699 1199
rect 3252 1177 3699 1193
rect 4047 1199 4090 1204
rect 2978 1171 3015 1172
rect 2928 1162 3015 1171
rect 2928 1142 2986 1162
rect 3006 1142 3015 1162
rect 2928 1132 3015 1142
rect 3074 1162 3111 1172
rect 3074 1142 3082 1162
rect 3102 1142 3111 1162
rect 2928 1131 2959 1132
rect 2552 1071 2893 1072
rect 3074 1071 3111 1142
rect 2477 1066 2893 1071
rect 2477 1046 2480 1066
rect 2500 1046 2893 1066
rect 2924 1047 3111 1071
rect 3252 1167 3696 1177
rect 3252 1165 3420 1167
rect 3252 987 3279 1165
rect 3319 1127 3383 1139
rect 3659 1135 3696 1167
rect 3722 1166 3913 1188
rect 3877 1164 3913 1166
rect 3877 1135 3914 1164
rect 4047 1143 4087 1199
rect 3319 1126 3354 1127
rect 3296 1121 3354 1126
rect 3296 1101 3299 1121
rect 3319 1107 3354 1121
rect 3374 1107 3383 1127
rect 3319 1099 3383 1107
rect 3345 1098 3383 1099
rect 3346 1097 3383 1098
rect 3449 1131 3485 1132
rect 3557 1131 3593 1132
rect 3449 1123 3593 1131
rect 3449 1103 3457 1123
rect 3477 1103 3512 1123
rect 3532 1103 3565 1123
rect 3585 1103 3593 1123
rect 3449 1097 3593 1103
rect 3659 1127 3697 1135
rect 3775 1131 3811 1132
rect 3659 1107 3668 1127
rect 3688 1107 3697 1127
rect 3659 1098 3697 1107
rect 3726 1123 3811 1131
rect 3726 1103 3783 1123
rect 3803 1103 3811 1123
rect 3659 1097 3696 1098
rect 3726 1097 3811 1103
rect 3877 1127 3915 1135
rect 3877 1107 3886 1127
rect 3906 1107 3915 1127
rect 4047 1125 4059 1143
rect 4077 1125 4087 1143
rect 4479 1171 4531 1360
rect 4877 1335 4916 1360
rect 5494 1375 5643 1382
rect 5494 1355 5553 1375
rect 5573 1355 5612 1375
rect 5632 1355 5643 1375
rect 5494 1347 5643 1355
rect 5710 1378 5867 1385
rect 5710 1358 5830 1378
rect 5850 1358 5867 1378
rect 5710 1348 5867 1358
rect 5710 1347 5745 1348
rect 4661 1310 4848 1334
rect 4877 1315 5272 1335
rect 5292 1315 5295 1335
rect 5710 1326 5741 1347
rect 5928 1326 5964 1436
rect 5983 1435 6020 1436
rect 6079 1435 6116 1436
rect 6039 1376 6129 1382
rect 6039 1356 6048 1376
rect 6068 1374 6129 1376
rect 6068 1356 6093 1374
rect 6039 1354 6093 1356
rect 6113 1354 6129 1374
rect 6039 1348 6129 1354
rect 5553 1325 5590 1326
rect 4877 1310 5295 1315
rect 5552 1316 5590 1325
rect 4661 1239 4698 1310
rect 4877 1309 5220 1310
rect 4877 1306 4916 1309
rect 5182 1308 5219 1309
rect 4813 1249 4844 1250
rect 4661 1219 4670 1239
rect 4690 1219 4698 1239
rect 4661 1209 4698 1219
rect 4757 1239 4844 1249
rect 4757 1219 4766 1239
rect 4786 1219 4844 1239
rect 4757 1210 4844 1219
rect 4757 1209 4794 1210
rect 4479 1153 4495 1171
rect 4513 1153 4531 1171
rect 4813 1159 4844 1210
rect 4879 1239 4916 1306
rect 5552 1296 5561 1316
rect 5581 1296 5590 1316
rect 5552 1288 5590 1296
rect 5656 1320 5741 1326
rect 5771 1325 5808 1326
rect 5656 1300 5664 1320
rect 5684 1300 5741 1320
rect 5656 1292 5741 1300
rect 5770 1316 5808 1325
rect 5770 1296 5779 1316
rect 5799 1296 5808 1316
rect 5656 1291 5692 1292
rect 5770 1288 5808 1296
rect 5874 1320 6018 1326
rect 5874 1300 5882 1320
rect 5902 1315 5990 1320
rect 5902 1300 5938 1315
rect 5874 1298 5938 1300
rect 5957 1300 5990 1315
rect 6010 1300 6018 1320
rect 5957 1298 6018 1300
rect 5874 1292 6018 1298
rect 5874 1291 5910 1292
rect 5982 1291 6018 1292
rect 6084 1325 6121 1326
rect 6084 1324 6122 1325
rect 6084 1316 6148 1324
rect 6084 1296 6093 1316
rect 6113 1302 6148 1316
rect 6168 1302 6171 1322
rect 6113 1297 6171 1302
rect 6113 1296 6148 1297
rect 5553 1259 5590 1288
rect 5554 1257 5590 1259
rect 5031 1249 5067 1250
rect 4879 1219 4888 1239
rect 4908 1219 4916 1239
rect 4879 1209 4916 1219
rect 4975 1239 5123 1249
rect 5223 1246 5319 1248
rect 4975 1219 4984 1239
rect 5004 1219 5094 1239
rect 5114 1219 5123 1239
rect 4975 1210 5123 1219
rect 5181 1239 5319 1246
rect 5181 1219 5190 1239
rect 5210 1219 5319 1239
rect 5554 1235 5745 1257
rect 5771 1256 5808 1288
rect 6084 1284 6148 1296
rect 6188 1258 6215 1436
rect 6047 1256 6215 1258
rect 5771 1242 6215 1256
rect 6818 1390 6986 1391
rect 7112 1390 7152 1614
rect 7615 1618 7783 1619
rect 8018 1618 8058 1651
rect 8414 1618 8461 1651
rect 7615 1617 8059 1618
rect 7615 1592 8060 1617
rect 7615 1590 7783 1592
rect 7979 1591 8060 1592
rect 8229 1591 8278 1617
rect 8414 1591 8463 1618
rect 7615 1412 7642 1590
rect 7682 1552 7746 1564
rect 8022 1560 8059 1591
rect 8240 1560 8277 1591
rect 8422 1566 8463 1591
rect 7682 1551 7717 1552
rect 7659 1546 7717 1551
rect 7659 1526 7662 1546
rect 7682 1532 7717 1546
rect 7737 1532 7746 1552
rect 7682 1524 7746 1532
rect 7708 1523 7746 1524
rect 7709 1522 7746 1523
rect 7812 1556 7848 1557
rect 7920 1556 7956 1557
rect 7812 1548 7956 1556
rect 7812 1528 7820 1548
rect 7840 1544 7928 1548
rect 7840 1528 7884 1544
rect 7812 1524 7884 1528
rect 7904 1528 7928 1544
rect 7948 1528 7956 1548
rect 7904 1524 7956 1528
rect 7812 1522 7956 1524
rect 8022 1552 8060 1560
rect 8138 1556 8174 1557
rect 8022 1532 8031 1552
rect 8051 1532 8060 1552
rect 8022 1523 8060 1532
rect 8089 1548 8174 1556
rect 8089 1528 8146 1548
rect 8166 1528 8174 1548
rect 8022 1522 8059 1523
rect 8089 1522 8174 1528
rect 8240 1552 8278 1560
rect 8240 1532 8249 1552
rect 8269 1532 8278 1552
rect 8240 1523 8278 1532
rect 8422 1557 8464 1566
rect 8422 1539 8436 1557
rect 8454 1539 8464 1557
rect 8422 1531 8464 1539
rect 8427 1529 8464 1531
rect 8240 1522 8277 1523
rect 7701 1494 7791 1500
rect 7701 1474 7717 1494
rect 7737 1492 7791 1494
rect 7737 1474 7762 1492
rect 7701 1472 7762 1474
rect 7782 1472 7791 1492
rect 7701 1466 7791 1472
rect 7714 1412 7751 1413
rect 7810 1412 7847 1413
rect 7866 1412 7902 1522
rect 8089 1501 8120 1522
rect 8085 1500 8120 1501
rect 7963 1490 8120 1500
rect 7963 1470 7980 1490
rect 8000 1470 8120 1490
rect 7963 1463 8120 1470
rect 8187 1493 8336 1501
rect 8187 1473 8198 1493
rect 8218 1473 8257 1493
rect 8277 1473 8336 1493
rect 8187 1466 8336 1473
rect 8187 1465 8228 1466
rect 8424 1464 8461 1467
rect 7921 1412 7958 1413
rect 7614 1403 7752 1412
rect 6818 1364 7262 1390
rect 6818 1362 6986 1364
rect 5771 1230 6218 1242
rect 5814 1228 5847 1230
rect 5181 1210 5319 1219
rect 4975 1209 5012 1210
rect 4705 1156 4746 1157
rect 4479 1135 4531 1153
rect 4597 1149 4746 1156
rect 4047 1115 4087 1125
rect 4597 1129 4656 1149
rect 4676 1129 4715 1149
rect 4735 1129 4746 1149
rect 4597 1121 4746 1129
rect 4813 1152 4970 1159
rect 4813 1132 4933 1152
rect 4953 1132 4970 1152
rect 4813 1122 4970 1132
rect 4813 1121 4848 1122
rect 3877 1098 3915 1107
rect 4813 1100 4844 1121
rect 5031 1100 5067 1210
rect 5086 1209 5123 1210
rect 5182 1209 5219 1210
rect 5142 1150 5232 1156
rect 5142 1130 5151 1150
rect 5171 1148 5232 1150
rect 5171 1130 5196 1148
rect 5142 1128 5196 1130
rect 5216 1128 5232 1148
rect 5142 1122 5232 1128
rect 4656 1099 4693 1100
rect 3877 1097 3914 1098
rect 3338 1069 3428 1075
rect 3338 1049 3354 1069
rect 3374 1067 3428 1069
rect 3374 1049 3399 1067
rect 3338 1047 3399 1049
rect 3419 1047 3428 1067
rect 3338 1041 3428 1047
rect 3351 987 3388 988
rect 3447 987 3484 988
rect 3503 987 3539 1097
rect 3726 1076 3757 1097
rect 4655 1090 4693 1099
rect 3722 1075 3757 1076
rect 3600 1065 3757 1075
rect 3600 1045 3617 1065
rect 3637 1045 3757 1065
rect 3600 1038 3757 1045
rect 3824 1068 3973 1076
rect 3824 1048 3835 1068
rect 3855 1048 3894 1068
rect 3914 1048 3973 1068
rect 4483 1072 4523 1082
rect 3824 1041 3973 1048
rect 4039 1044 4091 1062
rect 3824 1040 3865 1041
rect 3558 987 3595 988
rect 3251 978 3389 987
rect 3251 958 3360 978
rect 3380 958 3389 978
rect 3251 951 3389 958
rect 3447 978 3595 987
rect 3447 958 3456 978
rect 3476 958 3566 978
rect 3586 958 3595 978
rect 3251 949 3347 951
rect 3447 948 3595 958
rect 3654 978 3691 988
rect 3654 958 3662 978
rect 3682 958 3691 978
rect 3503 947 3539 948
rect 3654 891 3691 958
rect 3726 987 3757 1038
rect 4039 1026 4057 1044
rect 4075 1026 4091 1044
rect 3776 987 3813 988
rect 3726 978 3813 987
rect 3726 958 3784 978
rect 3804 958 3813 978
rect 3726 948 3813 958
rect 3872 978 3909 988
rect 3872 958 3880 978
rect 3900 958 3909 978
rect 3726 947 3757 948
rect 3351 888 3388 889
rect 3654 888 3693 891
rect 3350 887 3693 888
rect 3872 887 3909 958
rect 3275 882 3693 887
rect 3275 862 3278 882
rect 3298 862 3693 882
rect 3722 863 3909 887
rect 1816 831 1853 839
rect 1816 812 1824 831
rect 1845 812 1853 831
rect 1816 806 1853 812
rect 3654 837 3693 862
rect 4039 837 4091 1026
rect 4483 1054 4493 1072
rect 4511 1054 4523 1072
rect 4655 1070 4664 1090
rect 4684 1070 4693 1090
rect 4655 1062 4693 1070
rect 4759 1094 4844 1100
rect 4874 1099 4911 1100
rect 4759 1074 4767 1094
rect 4787 1074 4844 1094
rect 4759 1066 4844 1074
rect 4873 1090 4911 1099
rect 4873 1070 4882 1090
rect 4902 1070 4911 1090
rect 4759 1065 4795 1066
rect 4873 1062 4911 1070
rect 4977 1094 5121 1100
rect 4977 1074 4985 1094
rect 5005 1074 5038 1094
rect 5058 1074 5093 1094
rect 5113 1074 5121 1094
rect 4977 1066 5121 1074
rect 4977 1065 5013 1066
rect 5085 1065 5121 1066
rect 5187 1099 5224 1100
rect 5187 1098 5225 1099
rect 5187 1090 5251 1098
rect 5187 1070 5196 1090
rect 5216 1076 5251 1090
rect 5271 1076 5274 1096
rect 5216 1071 5274 1076
rect 5216 1070 5251 1071
rect 4483 998 4523 1054
rect 4656 1033 4693 1062
rect 4657 1031 4693 1033
rect 4657 1009 4848 1031
rect 4874 1030 4911 1062
rect 5187 1058 5251 1070
rect 5291 1032 5318 1210
rect 6176 1185 6218 1230
rect 5150 1030 5318 1032
rect 4874 1020 5318 1030
rect 5459 1126 5646 1150
rect 5677 1131 6070 1151
rect 6090 1131 6093 1151
rect 5677 1126 6093 1131
rect 5459 1055 5496 1126
rect 5677 1125 6018 1126
rect 5611 1065 5642 1066
rect 5459 1035 5468 1055
rect 5488 1035 5496 1055
rect 5459 1025 5496 1035
rect 5555 1055 5642 1065
rect 5555 1035 5564 1055
rect 5584 1035 5642 1055
rect 5555 1026 5642 1035
rect 5555 1025 5592 1026
rect 4480 993 4523 998
rect 4871 1004 5318 1020
rect 4871 998 4899 1004
rect 5150 1003 5318 1004
rect 4480 990 4630 993
rect 4871 990 4898 998
rect 4480 988 4898 990
rect 4480 970 4489 988
rect 4507 970 4898 988
rect 5611 975 5642 1026
rect 5677 1055 5714 1125
rect 5980 1124 6017 1125
rect 5829 1065 5865 1066
rect 5677 1035 5686 1055
rect 5706 1035 5714 1055
rect 5677 1025 5714 1035
rect 5773 1055 5921 1065
rect 6021 1062 6117 1064
rect 5773 1035 5782 1055
rect 5802 1035 5892 1055
rect 5912 1035 5921 1055
rect 5773 1026 5921 1035
rect 5979 1055 6117 1062
rect 5979 1035 5988 1055
rect 6008 1035 6117 1055
rect 5979 1026 6117 1035
rect 5773 1025 5810 1026
rect 5503 972 5544 973
rect 4480 967 4898 970
rect 4480 961 4523 967
rect 4483 958 4523 961
rect 5398 965 5544 972
rect 4880 949 4920 950
rect 4591 932 4920 949
rect 5398 945 5454 965
rect 5474 945 5513 965
rect 5533 945 5544 965
rect 5398 937 5544 945
rect 5611 968 5768 975
rect 5611 948 5731 968
rect 5751 948 5768 968
rect 5611 938 5768 948
rect 5611 937 5646 938
rect 4475 889 4518 900
rect 4475 871 4487 889
rect 4505 871 4518 889
rect 4475 845 4518 871
rect 4591 845 4618 932
rect 4880 923 4920 932
rect 3654 819 4093 837
rect 3654 801 4054 819
rect 4072 801 4093 819
rect 3654 795 4093 801
rect 3660 791 4093 795
rect 4475 824 4618 845
rect 4662 897 4696 913
rect 4880 903 5273 923
rect 5293 903 5296 923
rect 5611 916 5642 937
rect 5829 916 5865 1026
rect 5884 1025 5921 1026
rect 5980 1025 6017 1026
rect 5940 966 6030 972
rect 5940 946 5949 966
rect 5969 964 6030 966
rect 5969 946 5994 964
rect 5940 944 5994 946
rect 6014 944 6030 964
rect 5940 938 6030 944
rect 5454 915 5491 916
rect 4880 898 5296 903
rect 5453 906 5491 915
rect 4880 897 5221 898
rect 4662 827 4699 897
rect 4814 837 4845 838
rect 4475 822 4612 824
rect 4039 789 4091 791
rect 4475 780 4518 822
rect 4662 807 4671 827
rect 4691 807 4699 827
rect 4662 797 4699 807
rect 4758 827 4845 837
rect 4758 807 4767 827
rect 4787 807 4845 827
rect 4758 798 4845 807
rect 4758 797 4795 798
rect 4473 770 4518 780
rect 4473 752 4482 770
rect 4500 752 4518 770
rect 4473 746 4518 752
rect 4814 747 4845 798
rect 4880 827 4917 897
rect 5183 896 5220 897
rect 5453 886 5462 906
rect 5482 886 5491 906
rect 5453 878 5491 886
rect 5557 910 5642 916
rect 5672 915 5709 916
rect 5557 890 5565 910
rect 5585 890 5642 910
rect 5557 882 5642 890
rect 5671 906 5709 915
rect 5671 886 5680 906
rect 5700 886 5709 906
rect 5557 881 5593 882
rect 5671 878 5709 886
rect 5775 910 5919 916
rect 5775 890 5783 910
rect 5803 907 5891 910
rect 5803 890 5838 907
rect 5775 889 5838 890
rect 5857 890 5891 907
rect 5911 890 5919 910
rect 5857 889 5919 890
rect 5775 882 5919 889
rect 5775 881 5811 882
rect 5883 881 5919 882
rect 5985 915 6022 916
rect 5985 914 6023 915
rect 6045 914 6072 918
rect 5985 912 6072 914
rect 5985 906 6049 912
rect 5985 886 5994 906
rect 6014 892 6049 906
rect 6069 892 6072 912
rect 6014 887 6072 892
rect 6014 886 6049 887
rect 5454 849 5491 878
rect 5455 847 5491 849
rect 5032 837 5068 838
rect 4880 807 4889 827
rect 4909 807 4917 827
rect 4880 797 4917 807
rect 4976 827 5124 837
rect 5224 834 5320 836
rect 4976 807 4985 827
rect 5005 807 5095 827
rect 5115 807 5124 827
rect 4976 798 5124 807
rect 5182 827 5320 834
rect 5182 807 5191 827
rect 5211 807 5320 827
rect 5455 825 5646 847
rect 5672 846 5709 878
rect 5985 874 6049 886
rect 6089 848 6116 1026
rect 5948 846 6116 848
rect 5672 820 6116 846
rect 5182 798 5320 807
rect 4976 797 5013 798
rect 4473 743 4510 746
rect 4706 744 4747 745
rect 4598 737 4747 744
rect 4042 724 4079 729
rect 4033 720 4080 724
rect 4033 702 4052 720
rect 4070 702 4080 720
rect 4598 717 4657 737
rect 4677 717 4716 737
rect 4736 717 4747 737
rect 4598 709 4747 717
rect 4814 740 4971 747
rect 4814 720 4934 740
rect 4954 720 4971 740
rect 4814 710 4971 720
rect 4814 709 4849 710
rect 4033 639 4080 702
rect 4814 688 4845 709
rect 5032 688 5068 798
rect 5087 797 5124 798
rect 5183 797 5220 798
rect 5143 738 5233 744
rect 5143 718 5152 738
rect 5172 736 5233 738
rect 5172 718 5197 736
rect 5143 716 5197 718
rect 5217 716 5233 736
rect 5143 710 5233 716
rect 4657 687 4694 688
rect 4470 679 4507 681
rect 4470 671 4512 679
rect 4470 653 4480 671
rect 4498 653 4512 671
rect 4470 644 4512 653
rect 4656 678 4694 687
rect 4656 658 4665 678
rect 4685 658 4694 678
rect 4656 650 4694 658
rect 4760 682 4845 688
rect 4875 687 4912 688
rect 4760 662 4768 682
rect 4788 662 4845 682
rect 4760 654 4845 662
rect 4874 678 4912 687
rect 4874 658 4883 678
rect 4903 658 4912 678
rect 4760 653 4796 654
rect 4874 650 4912 658
rect 4978 686 5122 688
rect 4978 682 5030 686
rect 4978 662 4986 682
rect 5006 666 5030 682
rect 5050 682 5122 686
rect 5050 666 5094 682
rect 5006 662 5094 666
rect 5114 662 5122 682
rect 4978 654 5122 662
rect 4978 653 5014 654
rect 5086 653 5122 654
rect 5188 687 5225 688
rect 5188 686 5226 687
rect 5188 678 5252 686
rect 5188 658 5197 678
rect 5217 664 5252 678
rect 5272 664 5275 684
rect 5217 659 5275 664
rect 5217 658 5252 659
rect 4033 624 4083 639
rect 4033 599 4047 624
rect 4079 599 4083 624
rect 4471 619 4512 644
rect 4657 619 4694 650
rect 4875 628 4912 650
rect 5188 646 5252 658
rect 4870 619 4912 628
rect 5292 620 5319 798
rect 4471 607 4516 619
rect 4033 586 4080 599
rect 1418 561 1426 583
rect 1450 561 1458 583
rect 1418 553 1458 561
rect 4467 549 4516 607
rect 4657 593 4719 619
rect 4870 618 4955 619
rect 5151 618 5319 620
rect 4870 592 5319 618
rect 4870 549 4909 592
rect 5151 591 5319 592
rect 5782 596 5822 820
rect 5948 819 6116 820
rect 6180 852 6213 1185
rect 6818 1184 6845 1362
rect 6885 1324 6949 1336
rect 7225 1332 7262 1364
rect 7288 1363 7479 1385
rect 7614 1383 7723 1403
rect 7743 1383 7752 1403
rect 7614 1376 7752 1383
rect 7810 1403 7958 1412
rect 7810 1383 7819 1403
rect 7839 1383 7929 1403
rect 7949 1383 7958 1403
rect 7614 1374 7710 1376
rect 7810 1373 7958 1383
rect 8017 1403 8054 1413
rect 8017 1383 8025 1403
rect 8045 1383 8054 1403
rect 7866 1372 7902 1373
rect 7443 1361 7479 1363
rect 7443 1332 7480 1361
rect 6885 1323 6920 1324
rect 6862 1318 6920 1323
rect 6862 1298 6865 1318
rect 6885 1304 6920 1318
rect 6940 1304 6949 1324
rect 6885 1296 6949 1304
rect 6911 1295 6949 1296
rect 6912 1294 6949 1295
rect 7015 1328 7051 1329
rect 7123 1328 7159 1329
rect 7015 1320 7159 1328
rect 7015 1300 7023 1320
rect 7043 1319 7131 1320
rect 7043 1300 7078 1319
rect 7099 1300 7131 1319
rect 7151 1300 7159 1320
rect 7015 1294 7159 1300
rect 7225 1324 7263 1332
rect 7341 1328 7377 1329
rect 7225 1304 7234 1324
rect 7254 1304 7263 1324
rect 7225 1295 7263 1304
rect 7292 1320 7377 1328
rect 7292 1300 7349 1320
rect 7369 1300 7377 1320
rect 7225 1294 7262 1295
rect 7292 1294 7377 1300
rect 7443 1324 7481 1332
rect 7443 1304 7452 1324
rect 7472 1304 7481 1324
rect 7714 1313 7751 1314
rect 8017 1313 8054 1383
rect 8089 1412 8120 1463
rect 8416 1458 8461 1464
rect 8416 1440 8434 1458
rect 8452 1440 8461 1458
rect 8416 1430 8461 1440
rect 8139 1412 8176 1413
rect 8089 1403 8176 1412
rect 8089 1383 8147 1403
rect 8167 1383 8176 1403
rect 8089 1373 8176 1383
rect 8235 1403 8272 1413
rect 8235 1383 8243 1403
rect 8263 1383 8272 1403
rect 8416 1388 8459 1430
rect 8322 1386 8459 1388
rect 8089 1372 8120 1373
rect 8235 1313 8272 1383
rect 7713 1312 8054 1313
rect 7443 1295 7481 1304
rect 7638 1307 8054 1312
rect 7443 1294 7480 1295
rect 6904 1266 6994 1272
rect 6904 1246 6920 1266
rect 6940 1264 6994 1266
rect 6940 1246 6965 1264
rect 6904 1244 6965 1246
rect 6985 1244 6994 1264
rect 6904 1238 6994 1244
rect 6917 1184 6954 1185
rect 7013 1184 7050 1185
rect 7069 1184 7105 1294
rect 7292 1273 7323 1294
rect 7638 1287 7641 1307
rect 7661 1287 8054 1307
rect 8238 1297 8272 1313
rect 8316 1365 8459 1386
rect 8014 1278 8054 1287
rect 8316 1278 8343 1365
rect 8416 1339 8459 1365
rect 8416 1321 8429 1339
rect 8447 1321 8459 1339
rect 8416 1310 8459 1321
rect 7288 1272 7323 1273
rect 7166 1262 7323 1272
rect 7166 1242 7183 1262
rect 7203 1242 7323 1262
rect 7166 1235 7323 1242
rect 7390 1265 7539 1273
rect 7390 1245 7401 1265
rect 7421 1245 7460 1265
rect 7480 1245 7539 1265
rect 8014 1261 8343 1278
rect 8014 1260 8054 1261
rect 7390 1238 7539 1245
rect 8411 1249 8451 1252
rect 8411 1243 8454 1249
rect 8036 1240 8454 1243
rect 7390 1237 7431 1238
rect 7124 1184 7161 1185
rect 6817 1175 6955 1184
rect 6817 1155 6926 1175
rect 6946 1155 6955 1175
rect 6817 1148 6955 1155
rect 7013 1175 7161 1184
rect 7013 1155 7022 1175
rect 7042 1155 7132 1175
rect 7152 1155 7161 1175
rect 6817 1146 6913 1148
rect 7013 1145 7161 1155
rect 7220 1175 7257 1185
rect 7220 1155 7228 1175
rect 7248 1155 7257 1175
rect 7069 1144 7105 1145
rect 6917 1085 6954 1086
rect 7220 1085 7257 1155
rect 7292 1184 7323 1235
rect 8036 1222 8427 1240
rect 8445 1222 8454 1240
rect 8036 1220 8454 1222
rect 8036 1212 8063 1220
rect 8304 1217 8454 1220
rect 7616 1206 7784 1207
rect 8035 1206 8063 1212
rect 7616 1190 8063 1206
rect 8411 1212 8454 1217
rect 7342 1184 7379 1185
rect 7292 1175 7379 1184
rect 7292 1155 7350 1175
rect 7370 1155 7379 1175
rect 7292 1145 7379 1155
rect 7438 1175 7475 1185
rect 7438 1155 7446 1175
rect 7466 1155 7475 1175
rect 7292 1144 7323 1145
rect 6916 1084 7257 1085
rect 7438 1084 7475 1155
rect 6841 1079 7257 1084
rect 6841 1059 6844 1079
rect 6864 1059 7257 1079
rect 7288 1060 7475 1084
rect 7616 1180 8060 1190
rect 7616 1178 7784 1180
rect 7616 1000 7643 1178
rect 7683 1140 7747 1152
rect 8023 1148 8060 1180
rect 8086 1179 8277 1201
rect 8241 1177 8277 1179
rect 8241 1148 8278 1177
rect 8411 1156 8451 1212
rect 7683 1139 7718 1140
rect 7660 1134 7718 1139
rect 7660 1114 7663 1134
rect 7683 1120 7718 1134
rect 7738 1120 7747 1140
rect 7683 1112 7747 1120
rect 7709 1111 7747 1112
rect 7710 1110 7747 1111
rect 7813 1144 7849 1145
rect 7921 1144 7957 1145
rect 7813 1136 7957 1144
rect 7813 1116 7821 1136
rect 7841 1116 7876 1136
rect 7896 1116 7929 1136
rect 7949 1116 7957 1136
rect 7813 1110 7957 1116
rect 8023 1140 8061 1148
rect 8139 1144 8175 1145
rect 8023 1120 8032 1140
rect 8052 1120 8061 1140
rect 8023 1111 8061 1120
rect 8090 1136 8175 1144
rect 8090 1116 8147 1136
rect 8167 1116 8175 1136
rect 8023 1110 8060 1111
rect 8090 1110 8175 1116
rect 8241 1140 8279 1148
rect 8241 1120 8250 1140
rect 8270 1120 8279 1140
rect 8411 1138 8423 1156
rect 8441 1138 8451 1156
rect 8411 1128 8451 1138
rect 8241 1111 8279 1120
rect 8241 1110 8278 1111
rect 7702 1082 7792 1088
rect 7702 1062 7718 1082
rect 7738 1080 7792 1082
rect 7738 1062 7763 1080
rect 7702 1060 7763 1062
rect 7783 1060 7792 1080
rect 7702 1054 7792 1060
rect 7715 1000 7752 1001
rect 7811 1000 7848 1001
rect 7867 1000 7903 1110
rect 8090 1089 8121 1110
rect 8086 1088 8121 1089
rect 7964 1078 8121 1088
rect 7964 1058 7981 1078
rect 8001 1058 8121 1078
rect 7964 1051 8121 1058
rect 8188 1081 8337 1089
rect 8188 1061 8199 1081
rect 8219 1061 8258 1081
rect 8278 1061 8337 1081
rect 8188 1054 8337 1061
rect 8403 1057 8455 1075
rect 8188 1053 8229 1054
rect 7922 1000 7959 1001
rect 7615 991 7753 1000
rect 7615 971 7724 991
rect 7744 971 7753 991
rect 7615 964 7753 971
rect 7811 991 7959 1000
rect 7811 971 7820 991
rect 7840 971 7930 991
rect 7950 971 7959 991
rect 7615 962 7711 964
rect 7811 961 7959 971
rect 8018 991 8055 1001
rect 8018 971 8026 991
rect 8046 971 8055 991
rect 7867 960 7903 961
rect 8018 904 8055 971
rect 8090 1000 8121 1051
rect 8403 1039 8421 1057
rect 8439 1039 8455 1057
rect 8140 1000 8177 1001
rect 8090 991 8177 1000
rect 8090 971 8148 991
rect 8168 971 8177 991
rect 8090 961 8177 971
rect 8236 991 8273 1001
rect 8236 971 8244 991
rect 8264 971 8273 991
rect 8090 960 8121 961
rect 7715 901 7752 902
rect 8018 901 8057 904
rect 7714 900 8057 901
rect 8236 900 8273 971
rect 7639 895 8057 900
rect 7639 875 7642 895
rect 7662 875 8057 895
rect 8086 876 8273 900
rect 6180 844 6217 852
rect 6180 825 6188 844
rect 6209 825 6217 844
rect 6180 819 6217 825
rect 8018 850 8057 875
rect 8403 850 8455 1039
rect 8018 832 8457 850
rect 8018 814 8418 832
rect 8436 814 8457 832
rect 8018 808 8457 814
rect 8024 804 8457 808
rect 8403 802 8455 804
rect 8406 737 8443 742
rect 8397 733 8444 737
rect 8397 715 8416 733
rect 8434 715 8444 733
rect 8397 652 8444 715
rect 8397 637 8447 652
rect 8397 612 8411 637
rect 8443 612 8447 637
rect 8397 599 8444 612
rect 5782 574 5790 596
rect 5814 574 5822 596
rect 5782 566 5822 574
rect 101 509 506 536
rect 542 509 545 536
rect 4465 522 4870 549
rect 4906 522 4909 549
rect 4465 518 4909 522
rect 4465 517 4891 518
rect 101 505 545 509
rect 101 504 527 505
rect 6224 347 6289 348
rect 1860 334 1925 335
rect 1511 309 1698 333
rect 1729 313 2122 334
rect 2143 313 2145 334
rect 1729 309 2145 313
rect 5875 322 6062 346
rect 6093 326 6486 347
rect 6507 326 6509 347
rect 6093 322 6509 326
rect 1511 238 1548 309
rect 1729 308 2070 309
rect 1663 248 1694 249
rect 1511 218 1520 238
rect 1540 218 1548 238
rect 1511 208 1548 218
rect 1607 238 1694 248
rect 1607 218 1616 238
rect 1636 218 1694 238
rect 1607 209 1694 218
rect 1607 208 1644 209
rect 1663 158 1694 209
rect 1729 238 1766 308
rect 2032 307 2069 308
rect 4349 260 4414 261
rect 1881 248 1917 249
rect 1729 218 1738 238
rect 1758 218 1766 238
rect 1729 208 1766 218
rect 1825 238 1973 248
rect 2073 245 2234 247
rect 1825 218 1834 238
rect 1854 218 1944 238
rect 1964 218 1973 238
rect 1825 209 1973 218
rect 2031 240 2234 245
rect 2031 238 2204 240
rect 2031 218 2040 238
rect 2060 220 2204 238
rect 2224 220 2234 240
rect 2060 218 2234 220
rect 2031 211 2234 218
rect 4000 235 4187 259
rect 4218 239 4611 260
rect 4632 239 4634 260
rect 4218 235 4634 239
rect 5875 251 5912 322
rect 6093 321 6434 322
rect 6027 261 6058 262
rect 2031 209 2169 211
rect 1825 208 1862 209
rect 1555 155 1596 156
rect 1447 148 1596 155
rect 1447 128 1506 148
rect 1526 128 1565 148
rect 1585 128 1596 148
rect 1447 120 1596 128
rect 1663 151 1820 158
rect 1663 131 1783 151
rect 1803 131 1820 151
rect 1663 121 1820 131
rect 1663 120 1698 121
rect 1663 99 1694 120
rect 1881 99 1917 209
rect 1936 208 1973 209
rect 2032 208 2069 209
rect 1992 149 2082 155
rect 1992 129 2001 149
rect 2021 147 2082 149
rect 2021 129 2046 147
rect 1992 127 2046 129
rect 2066 127 2082 147
rect 1992 121 2082 127
rect 1506 98 1543 99
rect 1505 89 1543 98
rect 1505 69 1514 89
rect 1534 69 1543 89
rect 1505 61 1543 69
rect 1609 93 1694 99
rect 1724 98 1761 99
rect 1609 73 1617 93
rect 1637 73 1694 93
rect 1609 65 1694 73
rect 1723 89 1761 98
rect 1723 69 1732 89
rect 1752 69 1761 89
rect 1609 64 1645 65
rect 1723 61 1761 69
rect 1827 94 1971 99
rect 1827 93 1888 94
rect 1827 73 1835 93
rect 1855 73 1888 93
rect 1827 70 1888 73
rect 1911 93 1971 94
rect 1911 73 1943 93
rect 1963 73 1971 93
rect 1911 70 1971 73
rect 1827 65 1971 70
rect 1827 64 1863 65
rect 1935 64 1971 65
rect 2037 98 2074 99
rect 2037 97 2075 98
rect 2037 89 2101 97
rect 2037 69 2046 89
rect 2066 75 2101 89
rect 2121 75 2124 95
rect 2066 70 2124 75
rect 2066 69 2101 70
rect 1506 32 1543 61
rect 1507 30 1543 32
rect 1507 8 1698 30
rect 1724 29 1761 61
rect 2037 57 2101 69
rect 2141 31 2168 209
rect 4000 164 4037 235
rect 4218 234 4559 235
rect 4152 174 4183 175
rect 4000 144 4009 164
rect 4029 144 4037 164
rect 4000 134 4037 144
rect 4096 164 4183 174
rect 4096 144 4105 164
rect 4125 144 4183 164
rect 4096 135 4183 144
rect 4096 134 4133 135
rect 4152 84 4183 135
rect 4218 164 4255 234
rect 4521 233 4558 234
rect 5875 231 5884 251
rect 5904 231 5912 251
rect 5875 221 5912 231
rect 5971 251 6058 261
rect 5971 231 5980 251
rect 6000 231 6058 251
rect 5971 222 6058 231
rect 5971 221 6008 222
rect 4370 174 4406 175
rect 4218 144 4227 164
rect 4247 144 4255 164
rect 4218 134 4255 144
rect 4314 164 4462 174
rect 4562 171 4684 173
rect 4314 144 4323 164
rect 4343 144 4433 164
rect 4453 144 4462 164
rect 4314 135 4462 144
rect 4520 169 4684 171
rect 6027 171 6058 222
rect 6093 251 6130 321
rect 6396 320 6433 321
rect 6245 261 6281 262
rect 6093 231 6102 251
rect 6122 231 6130 251
rect 6093 221 6130 231
rect 6189 251 6337 261
rect 6437 258 6598 260
rect 6189 231 6198 251
rect 6218 231 6308 251
rect 6328 231 6337 251
rect 6189 222 6337 231
rect 6395 253 6598 258
rect 6395 251 6568 253
rect 6395 231 6404 251
rect 6424 233 6568 251
rect 6588 233 6598 253
rect 6424 231 6598 233
rect 6395 224 6598 231
rect 6395 222 6533 224
rect 6189 221 6226 222
rect 4520 166 4723 169
rect 5919 168 5960 169
rect 4520 164 4693 166
rect 4520 144 4529 164
rect 4549 146 4693 164
rect 4713 146 4723 166
rect 4549 144 4723 146
rect 4520 137 4723 144
rect 5811 161 5960 168
rect 5811 141 5870 161
rect 5890 141 5929 161
rect 5949 141 5960 161
rect 4520 135 4658 137
rect 4314 134 4351 135
rect 4044 81 4085 82
rect 3936 74 4085 81
rect 3936 54 3995 74
rect 4015 54 4054 74
rect 4074 54 4085 74
rect 3936 46 4085 54
rect 4152 77 4309 84
rect 4152 57 4272 77
rect 4292 57 4309 77
rect 4152 47 4309 57
rect 4152 46 4187 47
rect 2000 29 2168 31
rect 1724 3 2168 29
rect 4152 25 4183 46
rect 4370 25 4406 135
rect 4425 134 4462 135
rect 4521 134 4558 135
rect 4481 75 4571 81
rect 4481 55 4490 75
rect 4510 73 4571 75
rect 4510 55 4535 73
rect 4481 53 4535 55
rect 4555 53 4571 73
rect 4481 47 4571 53
rect 3995 24 4032 25
rect 1834 0 1874 3
rect 2000 2 2168 3
rect 3994 15 4032 24
rect 3994 -5 4003 15
rect 4023 -5 4032 15
rect 3994 -13 4032 -5
rect 4098 19 4183 25
rect 4213 24 4250 25
rect 4098 -1 4106 19
rect 4126 -1 4183 19
rect 4098 -9 4183 -1
rect 4212 15 4250 24
rect 4212 -5 4221 15
rect 4241 -5 4250 15
rect 4098 -10 4134 -9
rect 4212 -13 4250 -5
rect 4316 19 4460 25
rect 4316 -1 4324 19
rect 4344 -1 4432 19
rect 4452 -1 4460 19
rect 4316 -9 4460 -1
rect 4316 -10 4352 -9
rect 4424 -10 4460 -9
rect 4526 24 4563 25
rect 4526 23 4564 24
rect 4526 15 4590 23
rect 4526 -5 4535 15
rect 4555 1 4590 15
rect 4610 1 4613 21
rect 4555 -4 4613 1
rect 4555 -5 4590 -4
rect 3995 -42 4032 -13
rect 3996 -44 4032 -42
rect 3996 -66 4187 -44
rect 4213 -45 4250 -13
rect 4526 -17 4590 -5
rect 4630 -43 4657 135
rect 5811 133 5960 141
rect 6027 164 6184 171
rect 6027 144 6147 164
rect 6167 144 6184 164
rect 6027 134 6184 144
rect 6027 133 6062 134
rect 6027 112 6058 133
rect 6245 112 6281 222
rect 6300 221 6337 222
rect 6396 221 6433 222
rect 6356 162 6446 168
rect 6356 142 6365 162
rect 6385 160 6446 162
rect 6385 142 6410 160
rect 6356 140 6410 142
rect 6430 140 6446 160
rect 6356 134 6446 140
rect 5870 111 5907 112
rect 5869 102 5907 111
rect 5869 82 5878 102
rect 5898 82 5907 102
rect 5869 74 5907 82
rect 5973 106 6058 112
rect 6088 111 6125 112
rect 5973 86 5981 106
rect 6001 86 6058 106
rect 5973 78 6058 86
rect 6087 102 6125 111
rect 6087 82 6096 102
rect 6116 82 6125 102
rect 5973 77 6009 78
rect 6087 74 6125 82
rect 6191 108 6335 112
rect 6191 106 6255 108
rect 6191 86 6199 106
rect 6219 86 6255 106
rect 6191 84 6255 86
rect 6278 106 6335 108
rect 6278 86 6307 106
rect 6327 86 6335 106
rect 6278 84 6335 86
rect 6191 78 6335 84
rect 6191 77 6227 78
rect 6299 77 6335 78
rect 6401 111 6438 112
rect 6401 110 6439 111
rect 6401 102 6465 110
rect 6401 82 6410 102
rect 6430 88 6465 102
rect 6485 88 6488 108
rect 6430 83 6488 88
rect 6430 82 6465 83
rect 5870 45 5907 74
rect 5871 43 5907 45
rect 5871 21 6062 43
rect 6088 42 6125 74
rect 6401 70 6465 82
rect 6505 44 6532 222
rect 6364 42 6532 44
rect 6088 16 6532 42
rect 6198 13 6238 16
rect 6364 15 6532 16
rect 4489 -45 4657 -43
rect 4213 -71 4657 -45
rect 4323 -74 4363 -71
rect 4489 -72 4657 -71
<< viali >>
rect 2883 8727 2907 8749
rect 2488 8479 2509 8498
rect 1035 8428 1055 8448
rect 419 8242 439 8262
rect 959 8241 979 8261
rect 801 8187 821 8207
rect 1014 8189 1034 8209
rect 1833 8244 1853 8264
rect 1217 8058 1237 8078
rect 1036 8016 1056 8036
rect 1757 8057 1777 8077
rect 1598 8004 1619 8023
rect 1812 8005 1832 8025
rect 7247 8740 7271 8762
rect 3425 8639 3445 8659
rect 3647 8637 3667 8657
rect 3480 8587 3500 8607
rect 4020 8586 4040 8606
rect 2628 8411 2648 8431
rect 2840 8416 2859 8434
rect 2683 8359 2703 8379
rect 3404 8400 3424 8420
rect 3223 8358 3243 8378
rect 2607 8172 2627 8192
rect 3426 8227 3446 8247
rect 3639 8229 3659 8249
rect 6852 8492 6873 8511
rect 5399 8441 5419 8461
rect 4783 8255 4803 8275
rect 5323 8254 5343 8274
rect 3481 8175 3501 8195
rect 4021 8174 4041 8194
rect 420 7830 440 7850
rect 960 7829 980 7849
rect 793 7779 813 7799
rect 1015 7777 1035 7797
rect 2529 8001 2549 8021
rect 2740 8008 2759 8025
rect 2584 7949 2604 7969
rect 3405 7988 3425 8008
rect 3124 7948 3144 7968
rect 5165 8200 5185 8220
rect 5378 8202 5398 8222
rect 6197 8257 6217 8277
rect 5581 8071 5601 8091
rect 5400 8029 5420 8049
rect 6121 8070 6141 8090
rect 5962 8017 5983 8036
rect 6176 8018 6196 8038
rect 7789 8652 7809 8672
rect 8011 8650 8031 8670
rect 7844 8600 7864 8620
rect 8384 8599 8404 8619
rect 6992 8424 7012 8444
rect 7204 8429 7223 8447
rect 7047 8372 7067 8392
rect 7768 8413 7788 8433
rect 7587 8371 7607 8391
rect 6971 8185 6991 8205
rect 7790 8240 7810 8260
rect 8003 8242 8023 8262
rect 7845 8188 7865 8208
rect 8385 8187 8405 8207
rect 4784 7843 4804 7863
rect 2508 7762 2528 7782
rect 5324 7842 5344 7862
rect 5157 7792 5177 7812
rect 5379 7790 5399 7810
rect 1553 7687 1577 7709
rect 2866 7709 2890 7731
rect 1915 7636 1935 7656
rect 1299 7450 1319 7470
rect 1018 7410 1038 7430
rect 1839 7449 1859 7469
rect 1682 7397 1703 7416
rect 1894 7397 1914 7417
rect 6893 8014 6913 8034
rect 7104 8021 7123 8038
rect 6948 7962 6968 7982
rect 7769 8001 7789 8021
rect 7488 7961 7508 7981
rect 6872 7775 6892 7795
rect 5917 7700 5941 7722
rect 7230 7722 7254 7744
rect 3408 7621 3428 7641
rect 3630 7619 3650 7639
rect 3463 7569 3483 7589
rect 6279 7649 6299 7669
rect 4003 7568 4023 7588
rect 402 7224 422 7244
rect 942 7223 962 7243
rect 784 7169 804 7189
rect 997 7171 1017 7191
rect 1816 7226 1836 7246
rect 1200 7040 1220 7060
rect 1019 6998 1039 7018
rect 1740 7039 1760 7059
rect 1584 6984 1603 7002
rect 1795 6987 1815 7007
rect 403 6812 423 6832
rect 943 6811 963 6831
rect 776 6761 796 6781
rect 998 6759 1018 6779
rect 2611 7393 2631 7413
rect 2824 7395 2845 7414
rect 2666 7341 2686 7361
rect 3387 7382 3407 7402
rect 3206 7340 3226 7360
rect 2431 7242 2453 7260
rect 2590 7154 2610 7174
rect 3409 7209 3429 7229
rect 3622 7211 3642 7231
rect 5663 7463 5683 7483
rect 5382 7423 5402 7443
rect 6203 7462 6223 7482
rect 6046 7410 6067 7429
rect 6258 7410 6278 7430
rect 7772 7634 7792 7654
rect 7994 7632 8014 7652
rect 7827 7582 7847 7602
rect 8367 7581 8387 7601
rect 4766 7237 4786 7257
rect 5306 7236 5326 7256
rect 3464 7157 3484 7177
rect 4004 7156 4024 7176
rect 2232 7046 2256 7068
rect 1934 6920 1955 6939
rect 1536 6669 1560 6691
rect 1961 6616 1981 6636
rect 1345 6430 1365 6450
rect 998 6392 1018 6412
rect 1885 6429 1905 6449
rect 1729 6376 1747 6394
rect 1940 6377 1960 6397
rect 382 6206 402 6226
rect 922 6205 942 6225
rect 764 6151 784 6171
rect 977 6153 997 6173
rect 1796 6208 1816 6228
rect 1180 6022 1200 6042
rect 999 5980 1019 6000
rect 1720 6021 1740 6041
rect 1561 5968 1582 5987
rect 1775 5969 1795 5989
rect 383 5794 403 5814
rect 923 5793 943 5813
rect 756 5743 776 5763
rect 978 5741 998 5761
rect 1516 5651 1540 5673
rect 1878 5600 1898 5620
rect 1262 5414 1282 5434
rect 981 5374 1001 5394
rect 1802 5413 1822 5433
rect 1647 5357 1666 5374
rect 1857 5361 1877 5381
rect 365 5188 385 5208
rect 905 5187 925 5207
rect 747 5133 767 5153
rect 960 5135 980 5155
rect 1959 5290 1981 5308
rect 1779 5190 1799 5210
rect 1163 5004 1183 5024
rect 982 4962 1002 4982
rect 1703 5003 1723 5023
rect 1547 4948 1566 4966
rect 1758 4951 1778 4971
rect 366 4776 386 4796
rect 906 4775 926 4795
rect 739 4725 759 4745
rect 961 4723 981 4743
rect 2446 6985 2466 7005
rect 2657 6983 2680 7005
rect 2501 6933 2521 6953
rect 3388 6970 3408 6990
rect 3041 6932 3061 6952
rect 5148 7182 5168 7202
rect 5361 7184 5381 7204
rect 6180 7239 6200 7259
rect 5564 7053 5584 7073
rect 5383 7011 5403 7031
rect 6104 7052 6124 7072
rect 5948 6997 5967 7015
rect 6159 7000 6179 7020
rect 2425 6746 2445 6766
rect 4767 6825 4787 6845
rect 5307 6824 5327 6844
rect 5140 6774 5160 6794
rect 5362 6772 5382 6792
rect 2846 6691 2870 6713
rect 2451 6443 2472 6462
rect 6975 7406 6995 7426
rect 7188 7408 7209 7427
rect 7030 7354 7050 7374
rect 7751 7395 7771 7415
rect 7570 7353 7590 7373
rect 6795 7255 6817 7273
rect 6954 7167 6974 7187
rect 7773 7222 7793 7242
rect 7986 7224 8006 7244
rect 7828 7170 7848 7190
rect 8368 7169 8388 7189
rect 6596 7059 6620 7081
rect 6298 6933 6319 6952
rect 5900 6682 5924 6704
rect 3388 6603 3408 6623
rect 3610 6601 3630 6621
rect 3443 6551 3463 6571
rect 3983 6550 4003 6570
rect 6325 6629 6345 6649
rect 2591 6375 2611 6395
rect 2803 6380 2822 6398
rect 2646 6323 2666 6343
rect 3367 6364 3387 6384
rect 3186 6322 3206 6342
rect 2570 6136 2590 6156
rect 3389 6191 3409 6211
rect 3602 6193 3622 6213
rect 5709 6443 5729 6463
rect 5362 6405 5382 6425
rect 6249 6442 6269 6462
rect 6093 6389 6111 6407
rect 6304 6390 6324 6410
rect 4746 6219 4766 6239
rect 5286 6218 5306 6238
rect 3444 6139 3464 6159
rect 3984 6138 4004 6158
rect 2492 5965 2512 5985
rect 2703 5966 2724 5985
rect 2547 5913 2567 5933
rect 3368 5952 3388 5972
rect 3087 5912 3107 5932
rect 5128 6164 5148 6184
rect 5341 6166 5361 6186
rect 6160 6221 6180 6241
rect 5544 6035 5564 6055
rect 5363 5993 5383 6013
rect 6084 6034 6104 6054
rect 5925 5981 5946 6000
rect 6139 5982 6159 6002
rect 4747 5807 4767 5827
rect 2471 5726 2491 5746
rect 5287 5806 5307 5826
rect 5120 5756 5140 5776
rect 5342 5754 5362 5774
rect 2829 5673 2853 5695
rect 5880 5664 5904 5686
rect 3371 5585 3391 5605
rect 3593 5583 3613 5603
rect 3426 5533 3446 5553
rect 6242 5613 6262 5633
rect 3966 5532 3986 5552
rect 2574 5357 2594 5377
rect 2787 5359 2808 5378
rect 2629 5305 2649 5325
rect 3350 5346 3370 5366
rect 3169 5304 3189 5324
rect 2553 5118 2573 5138
rect 3372 5173 3392 5193
rect 3585 5175 3605 5195
rect 5626 5427 5646 5447
rect 5345 5387 5365 5407
rect 6166 5426 6186 5446
rect 6011 5370 6030 5387
rect 6221 5374 6241 5394
rect 4729 5201 4749 5221
rect 5269 5200 5289 5220
rect 3427 5121 3447 5141
rect 3967 5120 3987 5140
rect 1897 4884 1918 4903
rect 2270 4951 2290 4971
rect 2482 4950 2508 4976
rect 2325 4899 2345 4919
rect 3351 4934 3371 4954
rect 2865 4898 2885 4918
rect 5111 5146 5131 5166
rect 5324 5148 5344 5168
rect 6323 5303 6345 5321
rect 6143 5203 6163 5223
rect 5527 5017 5547 5037
rect 5346 4975 5366 4995
rect 6067 5016 6087 5036
rect 5911 4961 5930 4979
rect 6122 4964 6142 4984
rect 2249 4712 2269 4732
rect 4730 4789 4750 4809
rect 5270 4788 5290 4808
rect 5103 4738 5123 4758
rect 5325 4736 5345 4756
rect 1499 4633 1523 4655
rect 2810 4655 2834 4677
rect 2064 4578 2084 4598
rect 1448 4392 1468 4412
rect 962 4356 982 4376
rect 1988 4391 2008 4411
rect 1826 4328 1849 4351
rect 2043 4339 2063 4359
rect 2415 4407 2436 4426
rect 346 4170 366 4190
rect 886 4169 906 4189
rect 728 4115 748 4135
rect 941 4117 961 4137
rect 1760 4172 1780 4192
rect 1144 3986 1164 4006
rect 963 3944 983 3964
rect 1684 3985 1704 4005
rect 1525 3932 1546 3951
rect 1739 3933 1759 3953
rect 347 3758 367 3778
rect 887 3757 907 3777
rect 720 3707 740 3727
rect 942 3705 962 3725
rect 1480 3615 1504 3637
rect 1842 3564 1862 3584
rect 1226 3378 1246 3398
rect 945 3338 965 3358
rect 1766 3377 1786 3397
rect 1609 3325 1630 3344
rect 1821 3325 1841 3345
rect 329 3152 349 3172
rect 869 3151 889 3171
rect 711 3097 731 3117
rect 924 3099 944 3119
rect 1743 3154 1763 3174
rect 1127 2968 1147 2988
rect 946 2926 966 2946
rect 1667 2967 1687 2987
rect 1511 2912 1530 2930
rect 1722 2915 1742 2935
rect 330 2740 350 2760
rect 870 2739 890 2759
rect 703 2689 723 2709
rect 925 2687 945 2707
rect 1861 2848 1882 2867
rect 1463 2597 1487 2619
rect 1888 2544 1908 2564
rect 1272 2358 1292 2378
rect 925 2320 945 2340
rect 1812 2357 1832 2377
rect 1653 2305 1676 2327
rect 1867 2305 1887 2325
rect 6810 6998 6830 7018
rect 7021 6996 7044 7018
rect 6865 6946 6885 6966
rect 7752 6983 7772 7003
rect 7405 6945 7425 6965
rect 6789 6759 6809 6779
rect 7210 6704 7234 6726
rect 6815 6456 6836 6475
rect 7752 6616 7772 6636
rect 7974 6614 7994 6634
rect 7807 6564 7827 6584
rect 8347 6563 8367 6583
rect 6955 6388 6975 6408
rect 7167 6393 7186 6411
rect 7010 6336 7030 6356
rect 7731 6377 7751 6397
rect 7550 6335 7570 6355
rect 6934 6149 6954 6169
rect 7753 6204 7773 6224
rect 7966 6206 7986 6226
rect 7808 6152 7828 6172
rect 8348 6151 8368 6171
rect 6856 5978 6876 5998
rect 7067 5979 7088 5998
rect 6911 5926 6931 5946
rect 7732 5965 7752 5985
rect 7451 5925 7471 5945
rect 6835 5739 6855 5759
rect 7193 5686 7217 5708
rect 7735 5598 7755 5618
rect 7957 5596 7977 5616
rect 7790 5546 7810 5566
rect 8330 5545 8350 5565
rect 6938 5370 6958 5390
rect 7151 5372 7172 5391
rect 6993 5318 7013 5338
rect 7714 5359 7734 5379
rect 7533 5317 7553 5337
rect 6917 5131 6937 5151
rect 7736 5186 7756 5206
rect 7949 5188 7969 5208
rect 7791 5134 7811 5154
rect 8331 5133 8351 5153
rect 6261 4897 6282 4916
rect 6634 4964 6654 4984
rect 6846 4963 6872 4989
rect 6689 4912 6709 4932
rect 7715 4947 7735 4967
rect 7229 4911 7249 4931
rect 6613 4725 6633 4745
rect 5863 4646 5887 4668
rect 7174 4668 7198 4690
rect 3352 4567 3372 4587
rect 3574 4565 3594 4585
rect 3407 4515 3427 4535
rect 3947 4514 3967 4534
rect 6428 4591 6448 4611
rect 2555 4339 2575 4359
rect 2767 4344 2786 4362
rect 2610 4287 2630 4307
rect 3331 4328 3351 4348
rect 3150 4286 3170 4306
rect 2534 4100 2554 4120
rect 2352 4002 2374 4020
rect 3353 4155 3373 4175
rect 3566 4157 3586 4177
rect 5812 4405 5832 4425
rect 5326 4369 5346 4389
rect 6352 4404 6372 4424
rect 6190 4341 6213 4364
rect 6407 4352 6427 4372
rect 6779 4420 6800 4439
rect 4710 4183 4730 4203
rect 5250 4182 5270 4202
rect 3408 4103 3428 4123
rect 3948 4102 3968 4122
rect 2456 3929 2476 3949
rect 2667 3936 2686 3953
rect 2511 3877 2531 3897
rect 3332 3916 3352 3936
rect 3051 3876 3071 3896
rect 5092 4128 5112 4148
rect 5305 4130 5325 4150
rect 6124 4185 6144 4205
rect 5508 3999 5528 4019
rect 5327 3957 5347 3977
rect 6048 3998 6068 4018
rect 5889 3945 5910 3964
rect 6103 3946 6123 3966
rect 4711 3771 4731 3791
rect 2435 3690 2455 3710
rect 5251 3770 5271 3790
rect 5084 3720 5104 3740
rect 5306 3718 5326 3738
rect 2793 3637 2817 3659
rect 5844 3628 5868 3650
rect 3335 3549 3355 3569
rect 3557 3547 3577 3567
rect 3390 3497 3410 3517
rect 6206 3577 6226 3597
rect 3930 3496 3950 3516
rect 2538 3321 2558 3341
rect 2751 3323 2772 3342
rect 2593 3269 2613 3289
rect 3314 3310 3334 3330
rect 3133 3268 3153 3288
rect 2517 3082 2537 3102
rect 3336 3137 3356 3157
rect 3549 3139 3569 3159
rect 5590 3391 5610 3411
rect 5309 3351 5329 3371
rect 6130 3390 6150 3410
rect 5973 3338 5994 3357
rect 6185 3338 6205 3358
rect 4693 3165 4713 3185
rect 5233 3164 5253 3184
rect 3391 3085 3411 3105
rect 3931 3084 3951 3104
rect 2373 2913 2393 2933
rect 2586 2916 2604 2934
rect 2428 2861 2448 2881
rect 3315 2898 3335 2918
rect 2968 2860 2988 2880
rect 5075 3110 5095 3130
rect 5288 3112 5308 3132
rect 6107 3167 6127 3187
rect 5491 2981 5511 3001
rect 5310 2939 5330 2959
rect 6031 2980 6051 3000
rect 5875 2925 5894 2943
rect 6086 2928 6106 2948
rect 2352 2674 2372 2694
rect 4694 2753 4714 2773
rect 5234 2752 5254 2772
rect 5067 2702 5087 2722
rect 5289 2700 5309 2720
rect 2773 2619 2797 2641
rect 2378 2371 2399 2390
rect 2077 2242 2101 2264
rect 309 2134 329 2154
rect 849 2133 869 2153
rect 691 2079 711 2099
rect 904 2081 924 2101
rect 1723 2136 1743 2156
rect 1880 2050 1902 2068
rect 1107 1950 1127 1970
rect 926 1908 946 1928
rect 1647 1949 1667 1969
rect 1488 1896 1509 1915
rect 1702 1897 1722 1917
rect 6225 2861 6246 2880
rect 5827 2610 5851 2632
rect 3315 2531 3335 2551
rect 3537 2529 3557 2549
rect 3370 2479 3390 2499
rect 3910 2478 3930 2498
rect 6252 2557 6272 2577
rect 2518 2303 2538 2323
rect 2730 2308 2749 2326
rect 2573 2251 2593 2271
rect 3294 2292 3314 2312
rect 3113 2250 3133 2270
rect 2497 2064 2517 2084
rect 3316 2119 3336 2139
rect 3529 2121 3549 2141
rect 5636 2371 5656 2391
rect 5289 2333 5309 2353
rect 6176 2370 6196 2390
rect 6017 2318 6040 2340
rect 6231 2318 6251 2338
rect 7716 4580 7736 4600
rect 7938 4578 7958 4598
rect 7771 4528 7791 4548
rect 8311 4527 8331 4547
rect 6919 4352 6939 4372
rect 7131 4357 7150 4375
rect 6974 4300 6994 4320
rect 7695 4341 7715 4361
rect 7514 4299 7534 4319
rect 6898 4113 6918 4133
rect 6716 4015 6738 4033
rect 7717 4168 7737 4188
rect 7930 4170 7950 4190
rect 7772 4116 7792 4136
rect 8312 4115 8332 4135
rect 6820 3942 6840 3962
rect 7031 3949 7050 3966
rect 6875 3890 6895 3910
rect 7696 3929 7716 3949
rect 7415 3889 7435 3909
rect 6799 3703 6819 3723
rect 7157 3650 7181 3672
rect 7699 3562 7719 3582
rect 7921 3560 7941 3580
rect 7754 3510 7774 3530
rect 8294 3509 8314 3529
rect 6902 3334 6922 3354
rect 7115 3336 7136 3355
rect 6957 3282 6977 3302
rect 7678 3323 7698 3343
rect 7497 3281 7517 3301
rect 6881 3095 6901 3115
rect 7700 3150 7720 3170
rect 7913 3152 7933 3172
rect 7755 3098 7775 3118
rect 8295 3097 8315 3117
rect 6737 2926 6757 2946
rect 6950 2929 6968 2947
rect 6792 2874 6812 2894
rect 7679 2911 7699 2931
rect 7332 2873 7352 2893
rect 6716 2687 6736 2707
rect 7137 2632 7161 2654
rect 6742 2384 6763 2403
rect 6441 2255 6465 2277
rect 4673 2147 4693 2167
rect 5213 2146 5233 2166
rect 3371 2067 3391 2087
rect 3911 2066 3931 2086
rect 310 1722 330 1742
rect 850 1721 870 1741
rect 683 1671 703 1691
rect 905 1669 925 1689
rect 2419 1893 2439 1913
rect 2630 1894 2651 1913
rect 2474 1841 2494 1861
rect 3295 1880 3315 1900
rect 3014 1840 3034 1860
rect 5055 2092 5075 2112
rect 5268 2094 5288 2114
rect 6087 2149 6107 2169
rect 6244 2063 6266 2081
rect 5471 1963 5491 1983
rect 5290 1921 5310 1941
rect 6011 1962 6031 1982
rect 5852 1909 5873 1928
rect 6066 1910 6086 1930
rect 7679 2544 7699 2564
rect 7901 2542 7921 2562
rect 7734 2492 7754 2512
rect 8274 2491 8294 2511
rect 6882 2316 6902 2336
rect 7094 2321 7113 2339
rect 6937 2264 6957 2284
rect 7658 2305 7678 2325
rect 7477 2263 7497 2283
rect 6861 2077 6881 2097
rect 7680 2132 7700 2152
rect 7893 2134 7913 2154
rect 7735 2080 7755 2100
rect 8275 2079 8295 2099
rect 4674 1735 4694 1755
rect 2398 1654 2418 1674
rect 5214 1734 5234 1754
rect 5047 1684 5067 1704
rect 5269 1682 5289 1702
rect 1443 1579 1467 1601
rect 2756 1601 2780 1623
rect 1805 1528 1825 1548
rect 1189 1342 1209 1362
rect 908 1302 928 1322
rect 1729 1341 1749 1361
rect 1574 1285 1593 1302
rect 1784 1289 1804 1309
rect 6783 1906 6803 1926
rect 6994 1907 7015 1926
rect 6838 1854 6858 1874
rect 7659 1893 7679 1913
rect 7378 1853 7398 1873
rect 6762 1667 6782 1687
rect 5807 1592 5831 1614
rect 7120 1614 7144 1636
rect 3298 1513 3318 1533
rect 3520 1511 3540 1531
rect 3353 1461 3373 1481
rect 6169 1541 6189 1561
rect 3893 1460 3913 1480
rect 292 1116 312 1136
rect 832 1115 852 1135
rect 674 1061 694 1081
rect 887 1063 907 1083
rect 1706 1118 1726 1138
rect 1090 932 1110 952
rect 909 890 929 910
rect 1630 931 1650 951
rect 1474 876 1493 894
rect 1685 879 1705 899
rect 293 704 313 724
rect 833 703 853 723
rect 666 653 686 673
rect 888 651 908 671
rect 2501 1285 2521 1305
rect 2714 1287 2735 1306
rect 2556 1233 2576 1253
rect 3277 1274 3297 1294
rect 3096 1232 3116 1252
rect 2480 1046 2500 1066
rect 3299 1101 3319 1121
rect 3512 1103 3532 1123
rect 5553 1355 5573 1375
rect 5272 1315 5292 1335
rect 6093 1354 6113 1374
rect 5938 1298 5957 1315
rect 6148 1302 6168 1322
rect 7662 1526 7682 1546
rect 7884 1524 7904 1544
rect 7717 1474 7737 1494
rect 8257 1473 8277 1493
rect 4656 1129 4676 1149
rect 5196 1128 5216 1148
rect 3354 1049 3374 1069
rect 3894 1048 3914 1068
rect 3278 862 3298 882
rect 1824 812 1845 831
rect 5038 1074 5058 1094
rect 5251 1076 5271 1096
rect 6070 1131 6090 1151
rect 5454 945 5474 965
rect 5273 903 5293 923
rect 5994 944 6014 964
rect 5838 889 5857 907
rect 6049 892 6069 912
rect 4657 717 4677 737
rect 5197 716 5217 736
rect 5030 666 5050 686
rect 5252 664 5272 684
rect 4047 599 4079 624
rect 1426 561 1450 583
rect 6865 1298 6885 1318
rect 7078 1300 7099 1319
rect 6920 1246 6940 1266
rect 7641 1287 7661 1307
rect 7460 1245 7480 1265
rect 6844 1059 6864 1079
rect 7663 1114 7683 1134
rect 7876 1116 7896 1136
rect 7718 1062 7738 1082
rect 8258 1061 8278 1081
rect 7642 875 7662 895
rect 6188 825 6209 844
rect 8411 612 8443 637
rect 5790 574 5814 596
rect 506 509 542 536
rect 4870 522 4906 549
rect 2122 313 2143 334
rect 6486 326 6507 347
rect 2204 220 2224 240
rect 4611 239 4632 260
rect 1506 128 1526 148
rect 2046 127 2066 147
rect 1888 70 1911 94
rect 2101 75 2121 95
rect 6568 233 6588 253
rect 4693 146 4713 166
rect 5870 141 5890 161
rect 3995 54 4015 74
rect 4535 53 4555 73
rect 4590 1 4610 21
rect 6410 140 6430 160
rect 6255 84 6278 108
rect 6465 88 6485 108
<< metal1 >>
rect 7751 8770 8037 8771
rect 7236 8762 8039 8770
rect 3387 8757 3673 8758
rect 2872 8749 3675 8757
rect 2872 8732 2883 8749
rect 2873 8727 2883 8732
rect 2907 8732 3675 8749
rect 7236 8745 7247 8762
rect 2907 8727 2912 8732
rect 2873 8714 2912 8727
rect 3417 8666 3452 8667
rect 3396 8659 3452 8666
rect 3396 8639 3425 8659
rect 3445 8639 3452 8659
rect 3396 8634 3452 8639
rect 3636 8657 3675 8732
rect 7237 8740 7247 8745
rect 7271 8745 8039 8762
rect 7271 8740 7276 8745
rect 7237 8727 7276 8740
rect 7781 8679 7816 8680
rect 3636 8637 3647 8657
rect 3667 8637 3675 8657
rect 2480 8498 2862 8503
rect 2480 8479 2488 8498
rect 2509 8479 2862 8498
rect 2480 8471 2862 8479
rect 1031 8453 1063 8454
rect 1028 8448 1063 8453
rect 1028 8428 1035 8448
rect 1055 8428 1063 8448
rect 2833 8441 2862 8471
rect 2620 8438 2655 8439
rect 1028 8420 1063 8428
rect 410 8262 995 8270
rect 410 8242 419 8262
rect 439 8261 995 8262
rect 439 8242 959 8261
rect 410 8241 959 8242
rect 979 8241 995 8261
rect 410 8235 995 8241
rect 1029 8214 1063 8420
rect 2599 8431 2655 8438
rect 2599 8411 2628 8431
rect 2648 8411 2655 8431
rect 2599 8406 2655 8411
rect 2832 8434 2866 8441
rect 2832 8416 2840 8434
rect 2859 8416 2866 8434
rect 2832 8408 2866 8416
rect 3396 8428 3430 8634
rect 3636 8633 3675 8637
rect 7760 8672 7816 8679
rect 7760 8652 7789 8672
rect 7809 8652 7816 8672
rect 7760 8647 7816 8652
rect 8000 8670 8039 8745
rect 8000 8650 8011 8670
rect 8031 8650 8039 8670
rect 3464 8607 4049 8613
rect 3464 8587 3480 8607
rect 3500 8606 4049 8607
rect 3500 8587 4020 8606
rect 3464 8586 4020 8587
rect 4040 8586 4049 8606
rect 3464 8578 4049 8586
rect 6844 8511 7226 8516
rect 6844 8492 6852 8511
rect 6873 8492 7226 8511
rect 6844 8484 7226 8492
rect 5395 8466 5427 8467
rect 5392 8461 5427 8466
rect 5392 8441 5399 8461
rect 5419 8441 5427 8461
rect 7197 8454 7226 8484
rect 6984 8451 7019 8452
rect 5392 8433 5427 8441
rect 3396 8420 3431 8428
rect 793 8207 828 8214
rect 793 8187 801 8207
rect 821 8187 828 8207
rect 793 8114 828 8187
rect 1007 8209 1063 8214
rect 1007 8189 1014 8209
rect 1034 8189 1063 8209
rect 1007 8182 1063 8189
rect 1098 8316 1128 8318
rect 1827 8316 1860 8317
rect 1098 8290 1861 8316
rect 1007 8181 1042 8182
rect 1098 8115 1128 8290
rect 1827 8269 1861 8290
rect 1826 8264 1861 8269
rect 1826 8244 1833 8264
rect 1853 8244 1861 8264
rect 1826 8236 1861 8244
rect 1093 8114 1128 8115
rect 792 8087 1128 8114
rect 1098 8086 1128 8087
rect 1208 8078 1793 8086
rect 1208 8058 1217 8078
rect 1237 8077 1793 8078
rect 1237 8058 1757 8077
rect 1208 8057 1757 8058
rect 1777 8057 1793 8077
rect 1208 8051 1793 8057
rect 1032 8041 1064 8042
rect 1029 8036 1064 8041
rect 1029 8016 1036 8036
rect 1056 8016 1064 8036
rect 1827 8030 1861 8236
rect 2599 8200 2633 8406
rect 3396 8400 3404 8420
rect 3424 8400 3431 8420
rect 3396 8395 3431 8400
rect 3396 8394 3428 8395
rect 2667 8379 3252 8385
rect 2667 8359 2683 8379
rect 2703 8378 3252 8379
rect 2703 8359 3223 8378
rect 2667 8358 3223 8359
rect 3243 8358 3252 8378
rect 2667 8350 3252 8358
rect 3332 8349 3362 8350
rect 3332 8322 3668 8349
rect 3332 8321 3367 8322
rect 2599 8192 2634 8200
rect 2599 8172 2607 8192
rect 2627 8172 2634 8192
rect 2599 8167 2634 8172
rect 2599 8146 2633 8167
rect 3332 8146 3362 8321
rect 3418 8254 3453 8255
rect 2599 8120 3362 8146
rect 2600 8119 2633 8120
rect 3332 8118 3362 8120
rect 3397 8247 3453 8254
rect 3397 8227 3426 8247
rect 3446 8227 3453 8247
rect 3397 8222 3453 8227
rect 3632 8249 3667 8322
rect 3632 8229 3639 8249
rect 3659 8229 3667 8249
rect 4774 8275 5359 8283
rect 4774 8255 4783 8275
rect 4803 8274 5359 8275
rect 4803 8255 5323 8274
rect 4774 8254 5323 8255
rect 5343 8254 5359 8274
rect 4774 8248 5359 8254
rect 3632 8222 3667 8229
rect 5393 8227 5427 8433
rect 6963 8444 7019 8451
rect 6963 8424 6992 8444
rect 7012 8424 7019 8444
rect 6963 8419 7019 8424
rect 7196 8447 7230 8454
rect 7196 8429 7204 8447
rect 7223 8429 7230 8447
rect 7196 8421 7230 8429
rect 7760 8441 7794 8647
rect 8000 8646 8039 8650
rect 7828 8620 8413 8626
rect 7828 8600 7844 8620
rect 7864 8619 8413 8620
rect 7864 8600 8384 8619
rect 7828 8599 8384 8600
rect 8404 8599 8413 8619
rect 7828 8591 8413 8599
rect 7760 8433 7795 8441
rect 1029 8008 1064 8016
rect 411 7850 996 7858
rect 411 7830 420 7850
rect 440 7849 996 7850
rect 440 7830 960 7849
rect 411 7829 960 7830
rect 980 7829 996 7849
rect 411 7823 996 7829
rect 785 7799 824 7803
rect 1030 7802 1064 8008
rect 1593 8023 1628 8029
rect 1593 8004 1598 8023
rect 1619 8004 1628 8023
rect 1593 7995 1628 8004
rect 1805 8025 1861 8030
rect 1805 8005 1812 8025
rect 1832 8005 1861 8025
rect 1805 7998 1861 8005
rect 2428 8069 2762 8097
rect 1805 7997 1840 7998
rect 1597 7927 1626 7995
rect 1597 7893 1943 7927
rect 785 7779 793 7799
rect 813 7779 824 7799
rect 785 7704 824 7779
rect 1008 7797 1064 7802
rect 1008 7777 1015 7797
rect 1035 7777 1064 7797
rect 1008 7770 1064 7777
rect 1008 7769 1043 7770
rect 1548 7709 1587 7722
rect 1548 7704 1553 7709
rect 785 7687 1553 7704
rect 1577 7704 1587 7709
rect 1577 7687 1588 7704
rect 785 7679 1588 7687
rect 787 7678 1073 7679
rect 1904 7656 1943 7893
rect 1904 7644 1915 7656
rect 1908 7636 1915 7644
rect 1935 7636 1943 7656
rect 1908 7628 1943 7636
rect 1290 7470 1875 7478
rect 1290 7450 1299 7470
rect 1319 7469 1875 7470
rect 1319 7450 1839 7469
rect 1290 7449 1839 7450
rect 1859 7449 1875 7469
rect 1290 7443 1875 7449
rect 1014 7435 1046 7436
rect 1011 7430 1046 7435
rect 1011 7410 1018 7430
rect 1038 7410 1046 7430
rect 1909 7422 1943 7628
rect 1011 7402 1046 7410
rect 393 7244 978 7252
rect 393 7224 402 7244
rect 422 7243 978 7244
rect 422 7224 942 7243
rect 393 7223 942 7224
rect 962 7223 978 7243
rect 393 7217 978 7223
rect 1012 7196 1046 7402
rect 1677 7416 1708 7422
rect 1677 7397 1682 7416
rect 1703 7397 1708 7416
rect 1677 7355 1708 7397
rect 1887 7417 1943 7422
rect 1887 7397 1894 7417
rect 1914 7397 1943 7417
rect 1887 7390 1943 7397
rect 1887 7389 1922 7390
rect 1677 7327 2016 7355
rect 776 7189 811 7196
rect 776 7169 784 7189
rect 804 7169 811 7189
rect 776 7096 811 7169
rect 990 7191 1046 7196
rect 990 7171 997 7191
rect 1017 7171 1046 7191
rect 990 7164 1046 7171
rect 1081 7298 1111 7300
rect 1810 7298 1843 7299
rect 1081 7272 1844 7298
rect 990 7163 1025 7164
rect 1081 7097 1111 7272
rect 1810 7251 1844 7272
rect 1809 7246 1844 7251
rect 1809 7226 1816 7246
rect 1836 7226 1844 7246
rect 1809 7218 1844 7226
rect 1076 7096 1111 7097
rect 775 7069 1111 7096
rect 1081 7068 1111 7069
rect 1191 7060 1776 7068
rect 1191 7040 1200 7060
rect 1220 7059 1776 7060
rect 1220 7040 1740 7059
rect 1191 7039 1740 7040
rect 1760 7039 1776 7059
rect 1191 7033 1776 7039
rect 1015 7023 1047 7024
rect 1012 7018 1047 7023
rect 1012 6998 1019 7018
rect 1039 6998 1047 7018
rect 1810 7012 1844 7218
rect 1012 6990 1047 6998
rect 394 6832 979 6840
rect 394 6812 403 6832
rect 423 6831 979 6832
rect 423 6812 943 6831
rect 394 6811 943 6812
rect 963 6811 979 6831
rect 394 6805 979 6811
rect 768 6781 807 6785
rect 1013 6784 1047 6990
rect 1577 7002 1611 7010
rect 1577 6984 1584 7002
rect 1603 6984 1611 7002
rect 1577 6977 1611 6984
rect 1788 7007 1844 7012
rect 1788 6987 1795 7007
rect 1815 6987 1844 7007
rect 1788 6980 1844 6987
rect 1788 6979 1823 6980
rect 1581 6947 1610 6977
rect 1581 6939 1963 6947
rect 1581 6920 1934 6939
rect 1955 6920 1963 6939
rect 1581 6915 1963 6920
rect 768 6761 776 6781
rect 796 6761 807 6781
rect 768 6686 807 6761
rect 991 6779 1047 6784
rect 991 6759 998 6779
rect 1018 6759 1047 6779
rect 991 6752 1047 6759
rect 991 6751 1026 6752
rect 1531 6691 1570 6704
rect 1531 6686 1536 6691
rect 768 6669 1536 6686
rect 1560 6686 1570 6691
rect 1560 6669 1571 6686
rect 768 6661 1571 6669
rect 770 6660 1056 6661
rect 1987 6642 2016 7327
rect 2428 7260 2460 8069
rect 2736 8034 2762 8069
rect 2521 8028 2556 8029
rect 2500 8021 2556 8028
rect 2500 8001 2529 8021
rect 2549 8001 2556 8021
rect 2500 7996 2556 8001
rect 2732 8025 2768 8034
rect 2732 8008 2740 8025
rect 2759 8008 2768 8025
rect 2732 7999 2768 8008
rect 3397 8016 3431 8222
rect 5157 8220 5192 8227
rect 3465 8195 4050 8201
rect 3465 8175 3481 8195
rect 3501 8194 4050 8195
rect 3501 8175 4021 8194
rect 3465 8174 4021 8175
rect 4041 8174 4050 8194
rect 3465 8166 4050 8174
rect 5157 8200 5165 8220
rect 5185 8200 5192 8220
rect 5157 8127 5192 8200
rect 5371 8222 5427 8227
rect 5371 8202 5378 8222
rect 5398 8202 5427 8222
rect 5371 8195 5427 8202
rect 5462 8329 5492 8331
rect 6191 8329 6224 8330
rect 5462 8303 6225 8329
rect 5371 8194 5406 8195
rect 5462 8128 5492 8303
rect 6191 8282 6225 8303
rect 6190 8277 6225 8282
rect 6190 8257 6197 8277
rect 6217 8257 6225 8277
rect 6190 8249 6225 8257
rect 5457 8127 5492 8128
rect 5156 8100 5492 8127
rect 5462 8099 5492 8100
rect 5572 8091 6157 8099
rect 5572 8071 5581 8091
rect 5601 8090 6157 8091
rect 5601 8071 6121 8090
rect 5572 8070 6121 8071
rect 6141 8070 6157 8090
rect 5572 8064 6157 8070
rect 5396 8054 5428 8055
rect 5393 8049 5428 8054
rect 5393 8029 5400 8049
rect 5420 8029 5428 8049
rect 6191 8043 6225 8249
rect 6963 8213 6997 8419
rect 7760 8413 7768 8433
rect 7788 8413 7795 8433
rect 7760 8408 7795 8413
rect 7760 8407 7792 8408
rect 7031 8392 7616 8398
rect 7031 8372 7047 8392
rect 7067 8391 7616 8392
rect 7067 8372 7587 8391
rect 7031 8371 7587 8372
rect 7607 8371 7616 8391
rect 7031 8363 7616 8371
rect 7696 8362 7726 8363
rect 7696 8335 8032 8362
rect 7696 8334 7731 8335
rect 6963 8205 6998 8213
rect 6963 8185 6971 8205
rect 6991 8185 6998 8205
rect 6963 8180 6998 8185
rect 6963 8159 6997 8180
rect 7696 8159 7726 8334
rect 7782 8267 7817 8268
rect 6963 8133 7726 8159
rect 6964 8132 6997 8133
rect 7696 8131 7726 8133
rect 7761 8260 7817 8267
rect 7761 8240 7790 8260
rect 7810 8240 7817 8260
rect 7761 8235 7817 8240
rect 7996 8262 8031 8335
rect 7996 8242 8003 8262
rect 8023 8242 8031 8262
rect 7996 8235 8031 8242
rect 5393 8021 5428 8029
rect 3397 8008 3432 8016
rect 2500 7790 2534 7996
rect 3397 7988 3405 8008
rect 3425 7988 3432 8008
rect 3397 7983 3432 7988
rect 3397 7982 3429 7983
rect 2568 7969 3153 7975
rect 2568 7949 2584 7969
rect 2604 7968 3153 7969
rect 2604 7949 3124 7968
rect 2568 7948 3124 7949
rect 3144 7948 3153 7968
rect 2568 7940 3153 7948
rect 4775 7863 5360 7871
rect 4775 7843 4784 7863
rect 4804 7862 5360 7863
rect 4804 7843 5324 7862
rect 4775 7842 5324 7843
rect 5344 7842 5360 7862
rect 4775 7836 5360 7842
rect 5149 7812 5188 7816
rect 5394 7815 5428 8021
rect 5957 8036 5992 8042
rect 5957 8017 5962 8036
rect 5983 8017 5992 8036
rect 5957 8008 5992 8017
rect 6169 8038 6225 8043
rect 6169 8018 6176 8038
rect 6196 8018 6225 8038
rect 6169 8011 6225 8018
rect 6792 8082 7126 8110
rect 6169 8010 6204 8011
rect 5961 7940 5990 8008
rect 5961 7906 6307 7940
rect 5149 7792 5157 7812
rect 5177 7792 5188 7812
rect 2500 7782 2535 7790
rect 2500 7762 2508 7782
rect 2528 7774 2535 7782
rect 2528 7762 2539 7774
rect 2500 7525 2539 7762
rect 3370 7739 3656 7740
rect 2855 7731 3658 7739
rect 2855 7714 2866 7731
rect 2856 7709 2866 7714
rect 2890 7714 3658 7731
rect 2890 7709 2895 7714
rect 2856 7696 2895 7709
rect 3400 7648 3435 7649
rect 3379 7641 3435 7648
rect 3379 7621 3408 7641
rect 3428 7621 3435 7641
rect 3379 7616 3435 7621
rect 3619 7639 3658 7714
rect 5149 7717 5188 7792
rect 5372 7810 5428 7815
rect 5372 7790 5379 7810
rect 5399 7790 5428 7810
rect 5372 7783 5428 7790
rect 5372 7782 5407 7783
rect 5912 7722 5951 7735
rect 5912 7717 5917 7722
rect 5149 7700 5917 7717
rect 5941 7717 5951 7722
rect 5941 7700 5952 7717
rect 5149 7692 5952 7700
rect 5151 7691 5437 7692
rect 6268 7669 6307 7906
rect 6268 7657 6279 7669
rect 6272 7649 6279 7657
rect 6299 7649 6307 7669
rect 6272 7641 6307 7649
rect 3619 7619 3630 7639
rect 3650 7619 3658 7639
rect 2500 7491 2846 7525
rect 2817 7423 2846 7491
rect 2603 7420 2638 7421
rect 2428 7242 2431 7260
rect 2453 7242 2460 7260
rect 2428 7230 2460 7242
rect 2582 7413 2638 7420
rect 2582 7393 2611 7413
rect 2631 7393 2638 7413
rect 2582 7388 2638 7393
rect 2815 7414 2850 7423
rect 2815 7395 2824 7414
rect 2845 7395 2850 7414
rect 2815 7389 2850 7395
rect 3379 7410 3413 7616
rect 3619 7615 3658 7619
rect 3447 7589 4032 7595
rect 3447 7569 3463 7589
rect 3483 7588 4032 7589
rect 3483 7569 4003 7588
rect 3447 7568 4003 7569
rect 4023 7568 4032 7588
rect 3447 7560 4032 7568
rect 5654 7483 6239 7491
rect 5654 7463 5663 7483
rect 5683 7482 6239 7483
rect 5683 7463 6203 7482
rect 5654 7462 6203 7463
rect 6223 7462 6239 7482
rect 5654 7456 6239 7462
rect 5378 7448 5410 7449
rect 5375 7443 5410 7448
rect 5375 7423 5382 7443
rect 5402 7423 5410 7443
rect 6273 7435 6307 7641
rect 5375 7415 5410 7423
rect 3379 7402 3414 7410
rect 2582 7182 2616 7388
rect 3379 7382 3387 7402
rect 3407 7382 3414 7402
rect 3379 7377 3414 7382
rect 3379 7376 3411 7377
rect 2650 7361 3235 7367
rect 2650 7341 2666 7361
rect 2686 7360 3235 7361
rect 2686 7341 3206 7360
rect 2650 7340 3206 7341
rect 3226 7340 3235 7360
rect 2650 7332 3235 7340
rect 3315 7331 3345 7332
rect 3315 7304 3651 7331
rect 3315 7303 3350 7304
rect 2582 7174 2617 7182
rect 2582 7154 2590 7174
rect 2610 7154 2617 7174
rect 2582 7149 2617 7154
rect 2582 7128 2616 7149
rect 3315 7128 3345 7303
rect 3401 7236 3436 7237
rect 2582 7102 3345 7128
rect 2583 7101 2616 7102
rect 3315 7100 3345 7102
rect 3380 7229 3436 7236
rect 3380 7209 3409 7229
rect 3429 7209 3436 7229
rect 3380 7204 3436 7209
rect 3615 7231 3650 7304
rect 3615 7211 3622 7231
rect 3642 7211 3650 7231
rect 4757 7257 5342 7265
rect 4757 7237 4766 7257
rect 4786 7256 5342 7257
rect 4786 7237 5306 7256
rect 4757 7236 5306 7237
rect 5326 7236 5342 7256
rect 4757 7230 5342 7236
rect 3615 7204 3650 7211
rect 5376 7209 5410 7415
rect 6041 7429 6072 7435
rect 6041 7410 6046 7429
rect 6067 7410 6072 7429
rect 6041 7368 6072 7410
rect 6251 7430 6307 7435
rect 6251 7410 6258 7430
rect 6278 7410 6307 7430
rect 6251 7403 6307 7410
rect 6251 7402 6286 7403
rect 6041 7340 6380 7368
rect 2220 7068 2683 7076
rect 2220 7046 2232 7068
rect 2256 7046 2683 7068
rect 2220 7045 2683 7046
rect 2222 7033 2261 7045
rect 2656 7014 2683 7045
rect 2438 7012 2473 7013
rect 2417 7005 2473 7012
rect 2417 6985 2446 7005
rect 2466 6985 2473 7005
rect 2417 6980 2473 6985
rect 2652 7005 2685 7014
rect 2652 6983 2657 7005
rect 2680 6983 2685 7005
rect 2417 6774 2451 6980
rect 2652 6977 2685 6983
rect 3380 6998 3414 7204
rect 5140 7202 5175 7209
rect 3448 7177 4033 7183
rect 3448 7157 3464 7177
rect 3484 7176 4033 7177
rect 3484 7157 4004 7176
rect 3448 7156 4004 7157
rect 4024 7156 4033 7176
rect 3448 7148 4033 7156
rect 5140 7182 5148 7202
rect 5168 7182 5175 7202
rect 5140 7109 5175 7182
rect 5354 7204 5410 7209
rect 5354 7184 5361 7204
rect 5381 7184 5410 7204
rect 5354 7177 5410 7184
rect 5445 7311 5475 7313
rect 6174 7311 6207 7312
rect 5445 7285 6208 7311
rect 5354 7176 5389 7177
rect 5445 7110 5475 7285
rect 6174 7264 6208 7285
rect 6173 7259 6208 7264
rect 6173 7239 6180 7259
rect 6200 7239 6208 7259
rect 6173 7231 6208 7239
rect 5440 7109 5475 7110
rect 5139 7082 5475 7109
rect 5445 7081 5475 7082
rect 5555 7073 6140 7081
rect 5555 7053 5564 7073
rect 5584 7072 6140 7073
rect 5584 7053 6104 7072
rect 5555 7052 6104 7053
rect 6124 7052 6140 7072
rect 5555 7046 6140 7052
rect 5379 7036 5411 7037
rect 5376 7031 5411 7036
rect 5376 7011 5383 7031
rect 5403 7011 5411 7031
rect 6174 7025 6208 7231
rect 5376 7003 5411 7011
rect 3380 6990 3415 6998
rect 3380 6970 3388 6990
rect 3408 6970 3415 6990
rect 3380 6965 3415 6970
rect 3380 6964 3412 6965
rect 2485 6953 3070 6959
rect 2485 6933 2501 6953
rect 2521 6952 3070 6953
rect 2521 6933 3041 6952
rect 2485 6932 3041 6933
rect 3061 6932 3070 6952
rect 2485 6924 3070 6932
rect 4758 6845 5343 6853
rect 4758 6825 4767 6845
rect 4787 6844 5343 6845
rect 4787 6825 5307 6844
rect 4758 6824 5307 6825
rect 5327 6824 5343 6844
rect 4758 6818 5343 6824
rect 5132 6794 5171 6798
rect 5377 6797 5411 7003
rect 5941 7015 5975 7023
rect 5941 6997 5948 7015
rect 5967 6997 5975 7015
rect 5941 6990 5975 6997
rect 6152 7020 6208 7025
rect 6152 7000 6159 7020
rect 6179 7000 6208 7020
rect 6152 6993 6208 7000
rect 6152 6992 6187 6993
rect 5945 6960 5974 6990
rect 5945 6952 6327 6960
rect 5945 6933 6298 6952
rect 6319 6933 6327 6952
rect 5945 6928 6327 6933
rect 5132 6774 5140 6794
rect 5160 6774 5171 6794
rect 2417 6773 2452 6774
rect 2385 6766 2452 6773
rect 2385 6746 2425 6766
rect 2445 6746 2452 6766
rect 2385 6743 2452 6746
rect 2385 6740 2450 6743
rect 1956 6639 2021 6642
rect 1954 6636 2021 6639
rect 1954 6616 1961 6636
rect 1981 6616 2021 6636
rect 1954 6609 2021 6616
rect 1954 6608 1989 6609
rect 1336 6450 1921 6458
rect 1336 6430 1345 6450
rect 1365 6449 1921 6450
rect 1365 6430 1885 6449
rect 1336 6429 1885 6430
rect 1905 6429 1921 6449
rect 1336 6423 1921 6429
rect 994 6417 1026 6418
rect 991 6412 1026 6417
rect 991 6392 998 6412
rect 1018 6392 1026 6412
rect 991 6384 1026 6392
rect 373 6226 958 6234
rect 373 6206 382 6226
rect 402 6225 958 6226
rect 402 6206 922 6225
rect 373 6205 922 6206
rect 942 6205 958 6225
rect 373 6199 958 6205
rect 992 6178 1026 6384
rect 1719 6394 1760 6405
rect 1955 6402 1989 6608
rect 1719 6376 1729 6394
rect 1747 6376 1760 6394
rect 1719 6368 1760 6376
rect 1933 6397 1989 6402
rect 1933 6377 1940 6397
rect 1960 6377 1989 6397
rect 1933 6370 1989 6377
rect 1933 6369 1968 6370
rect 1728 6338 1754 6368
rect 1728 6337 2066 6338
rect 1728 6301 2082 6337
rect 756 6171 791 6178
rect 756 6151 764 6171
rect 784 6151 791 6171
rect 756 6078 791 6151
rect 970 6173 1026 6178
rect 970 6153 977 6173
rect 997 6153 1026 6173
rect 970 6146 1026 6153
rect 1061 6280 1091 6282
rect 1790 6280 1823 6281
rect 1061 6254 1824 6280
rect 970 6145 1005 6146
rect 1061 6079 1091 6254
rect 1790 6233 1824 6254
rect 1789 6228 1824 6233
rect 1789 6208 1796 6228
rect 1816 6208 1824 6228
rect 1789 6200 1824 6208
rect 1056 6078 1091 6079
rect 755 6051 1091 6078
rect 1061 6050 1091 6051
rect 1171 6042 1756 6050
rect 1171 6022 1180 6042
rect 1200 6041 1756 6042
rect 1200 6022 1720 6041
rect 1171 6021 1720 6022
rect 1740 6021 1756 6041
rect 1171 6015 1756 6021
rect 995 6005 1027 6006
rect 992 6000 1027 6005
rect 992 5980 999 6000
rect 1019 5980 1027 6000
rect 1790 5994 1824 6200
rect 992 5972 1027 5980
rect 374 5814 959 5822
rect 374 5794 383 5814
rect 403 5813 959 5814
rect 403 5794 923 5813
rect 374 5793 923 5794
rect 943 5793 959 5813
rect 374 5787 959 5793
rect 748 5763 787 5767
rect 993 5766 1027 5972
rect 1556 5987 1591 5993
rect 1556 5968 1561 5987
rect 1582 5968 1591 5987
rect 1556 5959 1591 5968
rect 1768 5989 1824 5994
rect 1768 5969 1775 5989
rect 1795 5969 1824 5989
rect 1768 5962 1824 5969
rect 1768 5961 1803 5962
rect 1560 5891 1589 5959
rect 1560 5857 1906 5891
rect 748 5743 756 5763
rect 776 5743 787 5763
rect 748 5668 787 5743
rect 971 5761 1027 5766
rect 971 5741 978 5761
rect 998 5741 1027 5761
rect 971 5734 1027 5741
rect 971 5733 1006 5734
rect 1511 5673 1550 5686
rect 1511 5668 1516 5673
rect 748 5651 1516 5668
rect 1540 5668 1550 5673
rect 1540 5651 1551 5668
rect 748 5643 1551 5651
rect 750 5642 1036 5643
rect 1867 5620 1906 5857
rect 1867 5608 1878 5620
rect 1871 5600 1878 5608
rect 1898 5600 1906 5620
rect 1871 5592 1906 5600
rect 1253 5434 1838 5442
rect 1253 5414 1262 5434
rect 1282 5433 1838 5434
rect 1282 5414 1802 5433
rect 1253 5413 1802 5414
rect 1822 5413 1838 5433
rect 1253 5407 1838 5413
rect 977 5399 1009 5400
rect 974 5394 1009 5399
rect 974 5374 981 5394
rect 1001 5374 1009 5394
rect 1872 5386 1906 5592
rect 974 5366 1009 5374
rect 356 5208 941 5216
rect 356 5188 365 5208
rect 385 5207 941 5208
rect 385 5188 905 5207
rect 356 5187 905 5188
rect 925 5187 941 5207
rect 356 5181 941 5187
rect 975 5160 1009 5366
rect 1638 5374 1674 5383
rect 1638 5357 1647 5374
rect 1666 5357 1674 5374
rect 1638 5348 1674 5357
rect 1850 5381 1906 5386
rect 1850 5361 1857 5381
rect 1877 5361 1906 5381
rect 1850 5354 1906 5361
rect 1850 5353 1885 5354
rect 1644 5313 1670 5348
rect 1952 5313 1984 5314
rect 1644 5308 1984 5313
rect 1644 5290 1959 5308
rect 1981 5290 1984 5308
rect 1644 5285 1984 5290
rect 1952 5284 1984 5285
rect 739 5153 774 5160
rect 739 5133 747 5153
rect 767 5133 774 5153
rect 739 5060 774 5133
rect 953 5155 1009 5160
rect 953 5135 960 5155
rect 980 5135 1009 5155
rect 953 5128 1009 5135
rect 1044 5262 1074 5264
rect 1773 5262 1806 5263
rect 1044 5236 1807 5262
rect 953 5127 988 5128
rect 1044 5061 1074 5236
rect 1773 5215 1807 5236
rect 1772 5210 1807 5215
rect 1772 5190 1779 5210
rect 1799 5190 1807 5210
rect 1772 5182 1807 5190
rect 1039 5060 1074 5061
rect 738 5033 1074 5060
rect 1044 5032 1074 5033
rect 1154 5024 1739 5032
rect 1154 5004 1163 5024
rect 1183 5023 1739 5024
rect 1183 5004 1703 5023
rect 1154 5003 1703 5004
rect 1723 5003 1739 5023
rect 1154 4997 1739 5003
rect 978 4987 1010 4988
rect 975 4982 1010 4987
rect 975 4962 982 4982
rect 1002 4962 1010 4982
rect 1773 4976 1807 5182
rect 975 4954 1010 4962
rect 357 4796 942 4804
rect 357 4776 366 4796
rect 386 4795 942 4796
rect 386 4776 906 4795
rect 357 4775 906 4776
rect 926 4775 942 4795
rect 357 4769 942 4775
rect 731 4745 770 4749
rect 976 4748 1010 4954
rect 1540 4966 1574 4974
rect 1540 4948 1547 4966
rect 1566 4948 1574 4966
rect 1540 4941 1574 4948
rect 1751 4971 1807 4976
rect 1751 4951 1758 4971
rect 1778 4951 1807 4971
rect 1751 4944 1807 4951
rect 1751 4943 1786 4944
rect 1544 4911 1573 4941
rect 1544 4903 1926 4911
rect 1544 4884 1897 4903
rect 1918 4884 1926 4903
rect 1544 4879 1926 4884
rect 731 4725 739 4745
rect 759 4725 770 4745
rect 731 4650 770 4725
rect 954 4743 1010 4748
rect 954 4723 961 4743
rect 981 4723 1010 4743
rect 954 4716 1010 4723
rect 954 4715 989 4716
rect 1494 4655 1533 4668
rect 1494 4650 1499 4655
rect 731 4633 1499 4650
rect 1523 4650 1533 4655
rect 1523 4633 1534 4650
rect 731 4625 1534 4633
rect 733 4624 1019 4625
rect 2055 4601 2082 6301
rect 2390 6055 2419 6740
rect 3350 6721 3636 6722
rect 2835 6713 3638 6721
rect 2835 6696 2846 6713
rect 2836 6691 2846 6696
rect 2870 6696 3638 6713
rect 2870 6691 2875 6696
rect 2836 6678 2875 6691
rect 3380 6630 3415 6631
rect 3359 6623 3415 6630
rect 3359 6603 3388 6623
rect 3408 6603 3415 6623
rect 3359 6598 3415 6603
rect 3599 6621 3638 6696
rect 5132 6699 5171 6774
rect 5355 6792 5411 6797
rect 5355 6772 5362 6792
rect 5382 6772 5411 6792
rect 5355 6765 5411 6772
rect 5355 6764 5390 6765
rect 5895 6704 5934 6717
rect 5895 6699 5900 6704
rect 5132 6682 5900 6699
rect 5924 6699 5934 6704
rect 5924 6682 5935 6699
rect 5132 6674 5935 6682
rect 5134 6673 5420 6674
rect 6351 6655 6380 7340
rect 6792 7273 6824 8082
rect 7100 8047 7126 8082
rect 6885 8041 6920 8042
rect 6864 8034 6920 8041
rect 6864 8014 6893 8034
rect 6913 8014 6920 8034
rect 6864 8009 6920 8014
rect 7096 8038 7132 8047
rect 7096 8021 7104 8038
rect 7123 8021 7132 8038
rect 7096 8012 7132 8021
rect 7761 8029 7795 8235
rect 7829 8208 8414 8214
rect 7829 8188 7845 8208
rect 7865 8207 8414 8208
rect 7865 8188 8385 8207
rect 7829 8187 8385 8188
rect 8405 8187 8414 8207
rect 7829 8179 8414 8187
rect 7761 8021 7796 8029
rect 6864 7803 6898 8009
rect 7761 8001 7769 8021
rect 7789 8001 7796 8021
rect 7761 7996 7796 8001
rect 7761 7995 7793 7996
rect 6932 7982 7517 7988
rect 6932 7962 6948 7982
rect 6968 7981 7517 7982
rect 6968 7962 7488 7981
rect 6932 7961 7488 7962
rect 7508 7961 7517 7981
rect 6932 7953 7517 7961
rect 6864 7795 6899 7803
rect 6864 7775 6872 7795
rect 6892 7787 6899 7795
rect 6892 7775 6903 7787
rect 6864 7538 6903 7775
rect 7734 7752 8020 7753
rect 7219 7744 8022 7752
rect 7219 7727 7230 7744
rect 7220 7722 7230 7727
rect 7254 7727 8022 7744
rect 7254 7722 7259 7727
rect 7220 7709 7259 7722
rect 7764 7661 7799 7662
rect 7743 7654 7799 7661
rect 7743 7634 7772 7654
rect 7792 7634 7799 7654
rect 7743 7629 7799 7634
rect 7983 7652 8022 7727
rect 7983 7632 7994 7652
rect 8014 7632 8022 7652
rect 6864 7504 7210 7538
rect 7181 7436 7210 7504
rect 6967 7433 7002 7434
rect 6792 7255 6795 7273
rect 6817 7255 6824 7273
rect 6792 7243 6824 7255
rect 6946 7426 7002 7433
rect 6946 7406 6975 7426
rect 6995 7406 7002 7426
rect 6946 7401 7002 7406
rect 7179 7427 7214 7436
rect 7179 7408 7188 7427
rect 7209 7408 7214 7427
rect 7179 7402 7214 7408
rect 7743 7423 7777 7629
rect 7983 7628 8022 7632
rect 7811 7602 8396 7608
rect 7811 7582 7827 7602
rect 7847 7601 8396 7602
rect 7847 7582 8367 7601
rect 7811 7581 8367 7582
rect 8387 7581 8396 7601
rect 7811 7573 8396 7581
rect 7743 7415 7778 7423
rect 6946 7195 6980 7401
rect 7743 7395 7751 7415
rect 7771 7395 7778 7415
rect 7743 7390 7778 7395
rect 7743 7389 7775 7390
rect 7014 7374 7599 7380
rect 7014 7354 7030 7374
rect 7050 7373 7599 7374
rect 7050 7354 7570 7373
rect 7014 7353 7570 7354
rect 7590 7353 7599 7373
rect 7014 7345 7599 7353
rect 7679 7344 7709 7345
rect 7679 7317 8015 7344
rect 7679 7316 7714 7317
rect 6946 7187 6981 7195
rect 6946 7167 6954 7187
rect 6974 7167 6981 7187
rect 6946 7162 6981 7167
rect 6946 7141 6980 7162
rect 7679 7141 7709 7316
rect 7765 7249 7800 7250
rect 6946 7115 7709 7141
rect 6947 7114 6980 7115
rect 7679 7113 7709 7115
rect 7744 7242 7800 7249
rect 7744 7222 7773 7242
rect 7793 7222 7800 7242
rect 7744 7217 7800 7222
rect 7979 7244 8014 7317
rect 7979 7224 7986 7244
rect 8006 7224 8014 7244
rect 7979 7217 8014 7224
rect 6584 7081 7047 7089
rect 6584 7059 6596 7081
rect 6620 7059 7047 7081
rect 6584 7058 7047 7059
rect 6586 7046 6625 7058
rect 7020 7027 7047 7058
rect 6802 7025 6837 7026
rect 6781 7018 6837 7025
rect 6781 6998 6810 7018
rect 6830 6998 6837 7018
rect 6781 6993 6837 6998
rect 7016 7018 7049 7027
rect 7016 6996 7021 7018
rect 7044 6996 7049 7018
rect 6781 6787 6815 6993
rect 7016 6990 7049 6996
rect 7744 7011 7778 7217
rect 7812 7190 8397 7196
rect 7812 7170 7828 7190
rect 7848 7189 8397 7190
rect 7848 7170 8368 7189
rect 7812 7169 8368 7170
rect 8388 7169 8397 7189
rect 7812 7161 8397 7169
rect 7744 7003 7779 7011
rect 7744 6983 7752 7003
rect 7772 6983 7779 7003
rect 7744 6978 7779 6983
rect 7744 6977 7776 6978
rect 6849 6966 7434 6972
rect 6849 6946 6865 6966
rect 6885 6965 7434 6966
rect 6885 6946 7405 6965
rect 6849 6945 7405 6946
rect 7425 6945 7434 6965
rect 6849 6937 7434 6945
rect 6781 6786 6816 6787
rect 6749 6779 6816 6786
rect 6749 6759 6789 6779
rect 6809 6759 6816 6779
rect 6749 6756 6816 6759
rect 6749 6753 6814 6756
rect 6320 6652 6385 6655
rect 6318 6649 6385 6652
rect 6318 6629 6325 6649
rect 6345 6629 6385 6649
rect 6318 6622 6385 6629
rect 6318 6621 6353 6622
rect 3599 6601 3610 6621
rect 3630 6601 3638 6621
rect 2443 6462 2825 6467
rect 2443 6443 2451 6462
rect 2472 6443 2825 6462
rect 2443 6435 2825 6443
rect 2796 6405 2825 6435
rect 2583 6402 2618 6403
rect 2562 6395 2618 6402
rect 2562 6375 2591 6395
rect 2611 6375 2618 6395
rect 2562 6370 2618 6375
rect 2795 6398 2829 6405
rect 2795 6380 2803 6398
rect 2822 6380 2829 6398
rect 2795 6372 2829 6380
rect 3359 6392 3393 6598
rect 3599 6597 3638 6601
rect 3427 6571 4012 6577
rect 3427 6551 3443 6571
rect 3463 6570 4012 6571
rect 3463 6551 3983 6570
rect 3427 6550 3983 6551
rect 4003 6550 4012 6570
rect 3427 6542 4012 6550
rect 5700 6463 6285 6471
rect 5700 6443 5709 6463
rect 5729 6462 6285 6463
rect 5729 6443 6249 6462
rect 5700 6442 6249 6443
rect 6269 6442 6285 6462
rect 5700 6436 6285 6442
rect 5358 6430 5390 6431
rect 5355 6425 5390 6430
rect 5355 6405 5362 6425
rect 5382 6405 5390 6425
rect 5355 6397 5390 6405
rect 3359 6384 3394 6392
rect 2562 6164 2596 6370
rect 3359 6364 3367 6384
rect 3387 6364 3394 6384
rect 3359 6359 3394 6364
rect 3359 6358 3391 6359
rect 2630 6343 3215 6349
rect 2630 6323 2646 6343
rect 2666 6342 3215 6343
rect 2666 6323 3186 6342
rect 2630 6322 3186 6323
rect 3206 6322 3215 6342
rect 2630 6314 3215 6322
rect 3295 6313 3325 6314
rect 3295 6286 3631 6313
rect 3295 6285 3330 6286
rect 2562 6156 2597 6164
rect 2562 6136 2570 6156
rect 2590 6136 2597 6156
rect 2562 6131 2597 6136
rect 2562 6110 2596 6131
rect 3295 6110 3325 6285
rect 3381 6218 3416 6219
rect 2562 6084 3325 6110
rect 2563 6083 2596 6084
rect 3295 6082 3325 6084
rect 3360 6211 3416 6218
rect 3360 6191 3389 6211
rect 3409 6191 3416 6211
rect 3360 6186 3416 6191
rect 3595 6213 3630 6286
rect 3595 6193 3602 6213
rect 3622 6193 3630 6213
rect 4737 6239 5322 6247
rect 4737 6219 4746 6239
rect 4766 6238 5322 6239
rect 4766 6219 5286 6238
rect 4737 6218 5286 6219
rect 5306 6218 5322 6238
rect 4737 6212 5322 6218
rect 3595 6186 3630 6193
rect 5356 6191 5390 6397
rect 6083 6407 6124 6418
rect 6319 6415 6353 6621
rect 6083 6389 6093 6407
rect 6111 6389 6124 6407
rect 6083 6381 6124 6389
rect 6297 6410 6353 6415
rect 6297 6390 6304 6410
rect 6324 6390 6353 6410
rect 6297 6383 6353 6390
rect 6297 6382 6332 6383
rect 6092 6351 6118 6381
rect 6092 6350 6430 6351
rect 6092 6314 6446 6350
rect 2390 6027 2729 6055
rect 2484 5992 2519 5993
rect 2463 5985 2519 5992
rect 2463 5965 2492 5985
rect 2512 5965 2519 5985
rect 2463 5960 2519 5965
rect 2698 5985 2729 6027
rect 2698 5966 2703 5985
rect 2724 5966 2729 5985
rect 2698 5960 2729 5966
rect 3360 5980 3394 6186
rect 5120 6184 5155 6191
rect 3428 6159 4013 6165
rect 3428 6139 3444 6159
rect 3464 6158 4013 6159
rect 3464 6139 3984 6158
rect 3428 6138 3984 6139
rect 4004 6138 4013 6158
rect 3428 6130 4013 6138
rect 5120 6164 5128 6184
rect 5148 6164 5155 6184
rect 5120 6091 5155 6164
rect 5334 6186 5390 6191
rect 5334 6166 5341 6186
rect 5361 6166 5390 6186
rect 5334 6159 5390 6166
rect 5425 6293 5455 6295
rect 6154 6293 6187 6294
rect 5425 6267 6188 6293
rect 5334 6158 5369 6159
rect 5425 6092 5455 6267
rect 6154 6246 6188 6267
rect 6153 6241 6188 6246
rect 6153 6221 6160 6241
rect 6180 6221 6188 6241
rect 6153 6213 6188 6221
rect 5420 6091 5455 6092
rect 5119 6064 5455 6091
rect 5425 6063 5455 6064
rect 5535 6055 6120 6063
rect 5535 6035 5544 6055
rect 5564 6054 6120 6055
rect 5564 6035 6084 6054
rect 5535 6034 6084 6035
rect 6104 6034 6120 6054
rect 5535 6028 6120 6034
rect 5359 6018 5391 6019
rect 5356 6013 5391 6018
rect 5356 5993 5363 6013
rect 5383 5993 5391 6013
rect 6154 6007 6188 6213
rect 5356 5985 5391 5993
rect 3360 5972 3395 5980
rect 2463 5754 2497 5960
rect 3360 5952 3368 5972
rect 3388 5952 3395 5972
rect 3360 5947 3395 5952
rect 3360 5946 3392 5947
rect 2531 5933 3116 5939
rect 2531 5913 2547 5933
rect 2567 5932 3116 5933
rect 2567 5913 3087 5932
rect 2531 5912 3087 5913
rect 3107 5912 3116 5932
rect 2531 5904 3116 5912
rect 4738 5827 5323 5835
rect 4738 5807 4747 5827
rect 4767 5826 5323 5827
rect 4767 5807 5287 5826
rect 4738 5806 5287 5807
rect 5307 5806 5323 5826
rect 4738 5800 5323 5806
rect 5112 5776 5151 5780
rect 5357 5779 5391 5985
rect 5920 6000 5955 6006
rect 5920 5981 5925 6000
rect 5946 5981 5955 6000
rect 5920 5972 5955 5981
rect 6132 6002 6188 6007
rect 6132 5982 6139 6002
rect 6159 5982 6188 6002
rect 6132 5975 6188 5982
rect 6132 5974 6167 5975
rect 5924 5904 5953 5972
rect 5924 5870 6270 5904
rect 5112 5756 5120 5776
rect 5140 5756 5151 5776
rect 2463 5746 2498 5754
rect 2463 5726 2471 5746
rect 2491 5738 2498 5746
rect 2491 5726 2502 5738
rect 2463 5489 2502 5726
rect 3333 5703 3619 5704
rect 2818 5695 3621 5703
rect 2818 5678 2829 5695
rect 2819 5673 2829 5678
rect 2853 5678 3621 5695
rect 2853 5673 2858 5678
rect 2819 5660 2858 5673
rect 3363 5612 3398 5613
rect 3342 5605 3398 5612
rect 3342 5585 3371 5605
rect 3391 5585 3398 5605
rect 3342 5580 3398 5585
rect 3582 5603 3621 5678
rect 5112 5681 5151 5756
rect 5335 5774 5391 5779
rect 5335 5754 5342 5774
rect 5362 5754 5391 5774
rect 5335 5747 5391 5754
rect 5335 5746 5370 5747
rect 5875 5686 5914 5699
rect 5875 5681 5880 5686
rect 5112 5664 5880 5681
rect 5904 5681 5914 5686
rect 5904 5664 5915 5681
rect 5112 5656 5915 5664
rect 5114 5655 5400 5656
rect 6231 5633 6270 5870
rect 6231 5621 6242 5633
rect 6235 5613 6242 5621
rect 6262 5613 6270 5633
rect 6235 5605 6270 5613
rect 3582 5583 3593 5603
rect 3613 5583 3621 5603
rect 2463 5455 2809 5489
rect 2780 5387 2809 5455
rect 2566 5384 2601 5385
rect 2545 5377 2601 5384
rect 2545 5357 2574 5377
rect 2594 5357 2601 5377
rect 2545 5352 2601 5357
rect 2778 5378 2813 5387
rect 2778 5359 2787 5378
rect 2808 5359 2813 5378
rect 2778 5353 2813 5359
rect 3342 5374 3376 5580
rect 3582 5579 3621 5583
rect 3410 5553 3995 5559
rect 3410 5533 3426 5553
rect 3446 5552 3995 5553
rect 3446 5533 3966 5552
rect 3410 5532 3966 5533
rect 3986 5532 3995 5552
rect 3410 5524 3995 5532
rect 5617 5447 6202 5455
rect 5617 5427 5626 5447
rect 5646 5446 6202 5447
rect 5646 5427 6166 5446
rect 5617 5426 6166 5427
rect 6186 5426 6202 5446
rect 5617 5420 6202 5426
rect 5341 5412 5373 5413
rect 5338 5407 5373 5412
rect 5338 5387 5345 5407
rect 5365 5387 5373 5407
rect 6236 5399 6270 5605
rect 5338 5379 5373 5387
rect 3342 5366 3377 5374
rect 2545 5146 2579 5352
rect 3342 5346 3350 5366
rect 3370 5346 3377 5366
rect 3342 5341 3377 5346
rect 3342 5340 3374 5341
rect 2613 5325 3198 5331
rect 2613 5305 2629 5325
rect 2649 5324 3198 5325
rect 2649 5305 3169 5324
rect 2613 5304 3169 5305
rect 3189 5304 3198 5324
rect 2613 5296 3198 5304
rect 3278 5295 3308 5296
rect 3278 5268 3614 5295
rect 3278 5267 3313 5268
rect 2545 5138 2580 5146
rect 2545 5118 2553 5138
rect 2573 5118 2580 5138
rect 2545 5113 2580 5118
rect 2545 5092 2579 5113
rect 3278 5092 3308 5267
rect 3364 5200 3399 5201
rect 2545 5066 3308 5092
rect 2546 5065 2579 5066
rect 3278 5064 3308 5066
rect 3343 5193 3399 5200
rect 3343 5173 3372 5193
rect 3392 5173 3399 5193
rect 3343 5168 3399 5173
rect 3578 5195 3613 5268
rect 3578 5175 3585 5195
rect 3605 5175 3613 5195
rect 4720 5221 5305 5229
rect 4720 5201 4729 5221
rect 4749 5220 5305 5221
rect 4749 5201 5269 5220
rect 4720 5200 5269 5201
rect 5289 5200 5305 5220
rect 4720 5194 5305 5200
rect 3578 5168 3613 5175
rect 5339 5173 5373 5379
rect 6002 5387 6038 5396
rect 6002 5370 6011 5387
rect 6030 5370 6038 5387
rect 6002 5361 6038 5370
rect 6214 5394 6270 5399
rect 6214 5374 6221 5394
rect 6241 5374 6270 5394
rect 6214 5367 6270 5374
rect 6214 5366 6249 5367
rect 6008 5326 6034 5361
rect 6316 5326 6348 5327
rect 6008 5321 6348 5326
rect 6008 5303 6323 5321
rect 6345 5303 6348 5321
rect 6008 5298 6348 5303
rect 6316 5297 6348 5298
rect 2197 5045 2514 5048
rect 2197 5018 2200 5045
rect 2227 5018 2514 5045
rect 2197 5012 2514 5018
rect 2197 5009 2233 5012
rect 2478 4982 2514 5012
rect 2262 4978 2297 4979
rect 2241 4971 2297 4978
rect 2241 4951 2270 4971
rect 2290 4951 2297 4971
rect 2241 4946 2297 4951
rect 2476 4976 2514 4982
rect 2476 4950 2482 4976
rect 2508 4950 2514 4976
rect 2241 4747 2275 4946
rect 2476 4942 2514 4950
rect 3343 4962 3377 5168
rect 5103 5166 5138 5173
rect 3411 5141 3996 5147
rect 3411 5121 3427 5141
rect 3447 5140 3996 5141
rect 3447 5121 3967 5140
rect 3411 5120 3967 5121
rect 3987 5120 3996 5140
rect 3411 5112 3996 5120
rect 5103 5146 5111 5166
rect 5131 5146 5138 5166
rect 5103 5073 5138 5146
rect 5317 5168 5373 5173
rect 5317 5148 5324 5168
rect 5344 5148 5373 5168
rect 5317 5141 5373 5148
rect 5408 5275 5438 5277
rect 6137 5275 6170 5276
rect 5408 5249 6171 5275
rect 5317 5140 5352 5141
rect 5408 5074 5438 5249
rect 6137 5228 6171 5249
rect 6136 5223 6171 5228
rect 6136 5203 6143 5223
rect 6163 5203 6171 5223
rect 6136 5195 6171 5203
rect 5403 5073 5438 5074
rect 5102 5046 5438 5073
rect 5408 5045 5438 5046
rect 5518 5037 6103 5045
rect 5518 5017 5527 5037
rect 5547 5036 6103 5037
rect 5547 5017 6067 5036
rect 5518 5016 6067 5017
rect 6087 5016 6103 5036
rect 5518 5010 6103 5016
rect 5342 5000 5374 5001
rect 5339 4995 5374 5000
rect 5339 4975 5346 4995
rect 5366 4975 5374 4995
rect 6137 4989 6171 5195
rect 5339 4967 5374 4975
rect 3343 4954 3378 4962
rect 3343 4934 3351 4954
rect 3371 4934 3378 4954
rect 3343 4929 3378 4934
rect 3343 4928 3375 4929
rect 2309 4919 2894 4925
rect 2309 4899 2325 4919
rect 2345 4918 2894 4919
rect 2345 4899 2865 4918
rect 2309 4898 2865 4899
rect 2885 4898 2894 4918
rect 2309 4890 2894 4898
rect 4721 4809 5306 4817
rect 4721 4789 4730 4809
rect 4750 4808 5306 4809
rect 4750 4789 5270 4808
rect 4721 4788 5270 4789
rect 5290 4788 5306 4808
rect 4721 4782 5306 4788
rect 5095 4758 5134 4762
rect 5340 4761 5374 4967
rect 5904 4979 5938 4987
rect 5904 4961 5911 4979
rect 5930 4961 5938 4979
rect 5904 4954 5938 4961
rect 6115 4984 6171 4989
rect 6115 4964 6122 4984
rect 6142 4964 6171 4984
rect 6115 4957 6171 4964
rect 6115 4956 6150 4957
rect 5908 4924 5937 4954
rect 5908 4916 6290 4924
rect 5908 4897 6261 4916
rect 6282 4897 6290 4916
rect 5908 4892 6290 4897
rect 2241 4732 2278 4747
rect 2241 4712 2249 4732
rect 2269 4712 2278 4732
rect 2241 4709 2278 4712
rect 2055 4598 2092 4601
rect 2055 4578 2064 4598
rect 2084 4578 2092 4598
rect 2055 4563 2092 4578
rect 1439 4412 2024 4420
rect 1439 4392 1448 4412
rect 1468 4411 2024 4412
rect 1468 4392 1988 4411
rect 1439 4391 1988 4392
rect 2008 4391 2024 4411
rect 1439 4385 2024 4391
rect 958 4381 990 4382
rect 955 4376 990 4381
rect 955 4356 962 4376
rect 982 4356 990 4376
rect 2058 4364 2092 4563
rect 2036 4359 2092 4364
rect 955 4348 990 4356
rect 337 4190 922 4198
rect 337 4170 346 4190
rect 366 4189 922 4190
rect 366 4170 886 4189
rect 337 4169 886 4170
rect 906 4169 922 4189
rect 337 4163 922 4169
rect 956 4142 990 4348
rect 1818 4357 1853 4359
rect 1818 4351 1856 4357
rect 1818 4328 1826 4351
rect 1849 4328 1856 4351
rect 2036 4339 2043 4359
rect 2063 4339 2092 4359
rect 2036 4332 2092 4339
rect 2036 4331 2071 4332
rect 1818 4322 1856 4328
rect 1818 4309 1853 4322
rect 1816 4251 1853 4309
rect 720 4135 755 4142
rect 720 4115 728 4135
rect 748 4115 755 4135
rect 720 4042 755 4115
rect 934 4137 990 4142
rect 934 4117 941 4137
rect 961 4117 990 4137
rect 934 4110 990 4117
rect 1025 4244 1055 4246
rect 1754 4244 1787 4245
rect 1025 4218 1788 4244
rect 934 4109 969 4110
rect 1025 4043 1055 4218
rect 1754 4197 1788 4218
rect 1816 4234 1851 4251
rect 1816 4233 2110 4234
rect 1816 4232 2153 4233
rect 1816 4225 2158 4232
rect 1816 4199 2118 4225
rect 2149 4199 2158 4225
rect 1753 4192 1788 4197
rect 2109 4196 2158 4199
rect 1753 4172 1760 4192
rect 1780 4172 1788 4192
rect 2115 4191 2158 4196
rect 1753 4164 1788 4172
rect 1020 4042 1055 4043
rect 719 4015 1055 4042
rect 1025 4014 1055 4015
rect 1135 4006 1720 4014
rect 1135 3986 1144 4006
rect 1164 4005 1720 4006
rect 1164 3986 1684 4005
rect 1135 3985 1684 3986
rect 1704 3985 1720 4005
rect 1135 3979 1720 3985
rect 959 3969 991 3970
rect 956 3964 991 3969
rect 956 3944 963 3964
rect 983 3944 991 3964
rect 1754 3958 1788 4164
rect 956 3936 991 3944
rect 338 3778 923 3786
rect 338 3758 347 3778
rect 367 3777 923 3778
rect 367 3758 887 3777
rect 338 3757 887 3758
rect 907 3757 923 3777
rect 338 3751 923 3757
rect 712 3727 751 3731
rect 957 3730 991 3936
rect 1520 3951 1555 3957
rect 1520 3932 1525 3951
rect 1546 3932 1555 3951
rect 1520 3923 1555 3932
rect 1732 3953 1788 3958
rect 1732 3933 1739 3953
rect 1759 3933 1788 3953
rect 1732 3926 1788 3933
rect 1732 3925 1767 3926
rect 1524 3855 1553 3923
rect 1524 3821 1870 3855
rect 712 3707 720 3727
rect 740 3707 751 3727
rect 712 3632 751 3707
rect 935 3725 991 3730
rect 935 3705 942 3725
rect 962 3705 991 3725
rect 935 3698 991 3705
rect 935 3697 970 3698
rect 1475 3637 1514 3650
rect 1475 3632 1480 3637
rect 712 3615 1480 3632
rect 1504 3632 1514 3637
rect 1504 3615 1515 3632
rect 712 3607 1515 3615
rect 714 3606 1000 3607
rect 1831 3584 1870 3821
rect 1831 3572 1842 3584
rect 1835 3564 1842 3572
rect 1862 3564 1870 3584
rect 1835 3556 1870 3564
rect 1217 3398 1802 3406
rect 1217 3378 1226 3398
rect 1246 3397 1802 3398
rect 1246 3378 1766 3397
rect 1217 3377 1766 3378
rect 1786 3377 1802 3397
rect 1217 3371 1802 3377
rect 941 3363 973 3364
rect 938 3358 973 3363
rect 938 3338 945 3358
rect 965 3338 973 3358
rect 1836 3350 1870 3556
rect 938 3330 973 3338
rect 320 3172 905 3180
rect 320 3152 329 3172
rect 349 3171 905 3172
rect 349 3152 869 3171
rect 320 3151 869 3152
rect 889 3151 905 3171
rect 320 3145 905 3151
rect 939 3124 973 3330
rect 1604 3344 1635 3350
rect 1604 3325 1609 3344
rect 1630 3325 1635 3344
rect 1604 3283 1635 3325
rect 1814 3345 1870 3350
rect 1814 3325 1821 3345
rect 1841 3325 1870 3345
rect 1814 3318 1870 3325
rect 1814 3317 1849 3318
rect 1604 3255 1943 3283
rect 703 3117 738 3124
rect 703 3097 711 3117
rect 731 3097 738 3117
rect 703 3024 738 3097
rect 917 3119 973 3124
rect 917 3099 924 3119
rect 944 3099 973 3119
rect 917 3092 973 3099
rect 1008 3226 1038 3228
rect 1737 3226 1770 3227
rect 1008 3200 1771 3226
rect 917 3091 952 3092
rect 1008 3025 1038 3200
rect 1737 3179 1771 3200
rect 1736 3174 1771 3179
rect 1736 3154 1743 3174
rect 1763 3154 1771 3174
rect 1736 3146 1771 3154
rect 1003 3024 1038 3025
rect 702 2997 1038 3024
rect 1008 2996 1038 2997
rect 1118 2988 1703 2996
rect 1118 2968 1127 2988
rect 1147 2987 1703 2988
rect 1147 2968 1667 2987
rect 1118 2967 1667 2968
rect 1687 2967 1703 2987
rect 1118 2961 1703 2967
rect 942 2951 974 2952
rect 939 2946 974 2951
rect 939 2926 946 2946
rect 966 2926 974 2946
rect 1737 2940 1771 3146
rect 939 2918 974 2926
rect 321 2760 906 2768
rect 321 2740 330 2760
rect 350 2759 906 2760
rect 350 2740 870 2759
rect 321 2739 870 2740
rect 890 2739 906 2759
rect 321 2733 906 2739
rect 695 2709 734 2713
rect 940 2712 974 2918
rect 1504 2930 1538 2938
rect 1504 2912 1511 2930
rect 1530 2912 1538 2930
rect 1504 2905 1538 2912
rect 1715 2935 1771 2940
rect 1715 2915 1722 2935
rect 1742 2915 1771 2935
rect 1715 2908 1771 2915
rect 1715 2907 1750 2908
rect 1508 2875 1537 2905
rect 1508 2867 1890 2875
rect 1508 2848 1861 2867
rect 1882 2848 1890 2867
rect 1508 2843 1890 2848
rect 695 2689 703 2709
rect 723 2689 734 2709
rect 695 2614 734 2689
rect 918 2707 974 2712
rect 918 2687 925 2707
rect 945 2687 974 2707
rect 918 2680 974 2687
rect 918 2679 953 2680
rect 1458 2619 1497 2632
rect 1458 2614 1463 2619
rect 695 2597 1463 2614
rect 1487 2614 1497 2619
rect 1487 2597 1498 2614
rect 695 2589 1498 2597
rect 697 2588 983 2589
rect 1914 2570 1943 3255
rect 2251 3009 2278 4709
rect 5095 4738 5103 4758
rect 5123 4738 5134 4758
rect 3314 4685 3600 4686
rect 2799 4677 3602 4685
rect 2799 4660 2810 4677
rect 2800 4655 2810 4660
rect 2834 4660 3602 4677
rect 2834 4655 2839 4660
rect 2800 4642 2839 4655
rect 3344 4594 3379 4595
rect 3323 4587 3379 4594
rect 3323 4567 3352 4587
rect 3372 4567 3379 4587
rect 3323 4562 3379 4567
rect 3563 4585 3602 4660
rect 5095 4663 5134 4738
rect 5318 4756 5374 4761
rect 5318 4736 5325 4756
rect 5345 4736 5374 4756
rect 5318 4729 5374 4736
rect 5318 4728 5353 4729
rect 5858 4668 5897 4681
rect 5858 4663 5863 4668
rect 5095 4646 5863 4663
rect 5887 4663 5897 4668
rect 5887 4646 5898 4663
rect 5095 4638 5898 4646
rect 5097 4637 5383 4638
rect 3563 4565 3574 4585
rect 3594 4565 3602 4585
rect 6419 4614 6446 6314
rect 6754 6068 6783 6753
rect 7714 6734 8000 6735
rect 7199 6726 8002 6734
rect 7199 6709 7210 6726
rect 7200 6704 7210 6709
rect 7234 6709 8002 6726
rect 7234 6704 7239 6709
rect 7200 6691 7239 6704
rect 7744 6643 7779 6644
rect 7723 6636 7779 6643
rect 7723 6616 7752 6636
rect 7772 6616 7779 6636
rect 7723 6611 7779 6616
rect 7963 6634 8002 6709
rect 7963 6614 7974 6634
rect 7994 6614 8002 6634
rect 6807 6475 7189 6480
rect 6807 6456 6815 6475
rect 6836 6456 7189 6475
rect 6807 6448 7189 6456
rect 7160 6418 7189 6448
rect 6947 6415 6982 6416
rect 6926 6408 6982 6415
rect 6926 6388 6955 6408
rect 6975 6388 6982 6408
rect 6926 6383 6982 6388
rect 7159 6411 7193 6418
rect 7159 6393 7167 6411
rect 7186 6393 7193 6411
rect 7159 6385 7193 6393
rect 7723 6405 7757 6611
rect 7963 6610 8002 6614
rect 7791 6584 8376 6590
rect 7791 6564 7807 6584
rect 7827 6583 8376 6584
rect 7827 6564 8347 6583
rect 7791 6563 8347 6564
rect 8367 6563 8376 6583
rect 7791 6555 8376 6563
rect 7723 6397 7758 6405
rect 6926 6177 6960 6383
rect 7723 6377 7731 6397
rect 7751 6377 7758 6397
rect 7723 6372 7758 6377
rect 7723 6371 7755 6372
rect 6994 6356 7579 6362
rect 6994 6336 7010 6356
rect 7030 6355 7579 6356
rect 7030 6336 7550 6355
rect 6994 6335 7550 6336
rect 7570 6335 7579 6355
rect 6994 6327 7579 6335
rect 7659 6326 7689 6327
rect 7659 6299 7995 6326
rect 7659 6298 7694 6299
rect 6926 6169 6961 6177
rect 6926 6149 6934 6169
rect 6954 6149 6961 6169
rect 6926 6144 6961 6149
rect 6926 6123 6960 6144
rect 7659 6123 7689 6298
rect 7745 6231 7780 6232
rect 6926 6097 7689 6123
rect 6927 6096 6960 6097
rect 7659 6095 7689 6097
rect 7724 6224 7780 6231
rect 7724 6204 7753 6224
rect 7773 6204 7780 6224
rect 7724 6199 7780 6204
rect 7959 6226 7994 6299
rect 7959 6206 7966 6226
rect 7986 6206 7994 6226
rect 7959 6199 7994 6206
rect 6754 6040 7093 6068
rect 6848 6005 6883 6006
rect 6827 5998 6883 6005
rect 6827 5978 6856 5998
rect 6876 5978 6883 5998
rect 6827 5973 6883 5978
rect 7062 5998 7093 6040
rect 7062 5979 7067 5998
rect 7088 5979 7093 5998
rect 7062 5973 7093 5979
rect 7724 5993 7758 6199
rect 7792 6172 8377 6178
rect 7792 6152 7808 6172
rect 7828 6171 8377 6172
rect 7828 6152 8348 6171
rect 7792 6151 8348 6152
rect 8368 6151 8377 6171
rect 7792 6143 8377 6151
rect 7724 5985 7759 5993
rect 6827 5767 6861 5973
rect 7724 5965 7732 5985
rect 7752 5965 7759 5985
rect 7724 5960 7759 5965
rect 7724 5959 7756 5960
rect 6895 5946 7480 5952
rect 6895 5926 6911 5946
rect 6931 5945 7480 5946
rect 6931 5926 7451 5945
rect 6895 5925 7451 5926
rect 7471 5925 7480 5945
rect 6895 5917 7480 5925
rect 6827 5759 6862 5767
rect 6827 5739 6835 5759
rect 6855 5751 6862 5759
rect 6855 5739 6866 5751
rect 6827 5502 6866 5739
rect 7697 5716 7983 5717
rect 7182 5708 7985 5716
rect 7182 5691 7193 5708
rect 7183 5686 7193 5691
rect 7217 5691 7985 5708
rect 7217 5686 7222 5691
rect 7183 5673 7222 5686
rect 7727 5625 7762 5626
rect 7706 5618 7762 5625
rect 7706 5598 7735 5618
rect 7755 5598 7762 5618
rect 7706 5593 7762 5598
rect 7946 5616 7985 5691
rect 7946 5596 7957 5616
rect 7977 5596 7985 5616
rect 6827 5468 7173 5502
rect 7144 5400 7173 5468
rect 6930 5397 6965 5398
rect 6909 5390 6965 5397
rect 6909 5370 6938 5390
rect 6958 5370 6965 5390
rect 6909 5365 6965 5370
rect 7142 5391 7177 5400
rect 7142 5372 7151 5391
rect 7172 5372 7177 5391
rect 7142 5366 7177 5372
rect 7706 5387 7740 5593
rect 7946 5592 7985 5596
rect 7774 5566 8359 5572
rect 7774 5546 7790 5566
rect 7810 5565 8359 5566
rect 7810 5546 8330 5565
rect 7774 5545 8330 5546
rect 8350 5545 8359 5565
rect 7774 5537 8359 5545
rect 7706 5379 7741 5387
rect 6909 5159 6943 5365
rect 7706 5359 7714 5379
rect 7734 5359 7741 5379
rect 7706 5354 7741 5359
rect 7706 5353 7738 5354
rect 6977 5338 7562 5344
rect 6977 5318 6993 5338
rect 7013 5337 7562 5338
rect 7013 5318 7533 5337
rect 6977 5317 7533 5318
rect 7553 5317 7562 5337
rect 6977 5309 7562 5317
rect 7642 5308 7672 5309
rect 7642 5281 7978 5308
rect 7642 5280 7677 5281
rect 6909 5151 6944 5159
rect 6909 5131 6917 5151
rect 6937 5131 6944 5151
rect 6909 5126 6944 5131
rect 6909 5105 6943 5126
rect 7642 5105 7672 5280
rect 7728 5213 7763 5214
rect 6909 5079 7672 5105
rect 6910 5078 6943 5079
rect 7642 5077 7672 5079
rect 7707 5206 7763 5213
rect 7707 5186 7736 5206
rect 7756 5186 7763 5206
rect 7707 5181 7763 5186
rect 7942 5208 7977 5281
rect 7942 5188 7949 5208
rect 7969 5188 7977 5208
rect 7942 5181 7977 5188
rect 6561 5058 6878 5061
rect 6561 5031 6564 5058
rect 6591 5031 6878 5058
rect 6561 5025 6878 5031
rect 6561 5022 6597 5025
rect 6842 4995 6878 5025
rect 6626 4991 6661 4992
rect 6605 4984 6661 4991
rect 6605 4964 6634 4984
rect 6654 4964 6661 4984
rect 6605 4959 6661 4964
rect 6840 4989 6878 4995
rect 6840 4963 6846 4989
rect 6872 4963 6878 4989
rect 6605 4760 6639 4959
rect 6840 4955 6878 4963
rect 7707 4975 7741 5181
rect 7775 5154 8360 5160
rect 7775 5134 7791 5154
rect 7811 5153 8360 5154
rect 7811 5134 8331 5153
rect 7775 5133 8331 5134
rect 8351 5133 8360 5153
rect 7775 5125 8360 5133
rect 7707 4967 7742 4975
rect 7707 4947 7715 4967
rect 7735 4947 7742 4967
rect 7707 4942 7742 4947
rect 7707 4941 7739 4942
rect 6673 4932 7258 4938
rect 6673 4912 6689 4932
rect 6709 4931 7258 4932
rect 6709 4912 7229 4931
rect 6673 4911 7229 4912
rect 7249 4911 7258 4931
rect 6673 4903 7258 4911
rect 6605 4745 6642 4760
rect 6605 4725 6613 4745
rect 6633 4725 6642 4745
rect 6605 4722 6642 4725
rect 6419 4611 6456 4614
rect 6419 4591 6428 4611
rect 6448 4591 6456 4611
rect 6419 4576 6456 4591
rect 2407 4426 2789 4431
rect 2407 4407 2415 4426
rect 2436 4407 2789 4426
rect 2407 4399 2789 4407
rect 2760 4369 2789 4399
rect 2547 4366 2582 4367
rect 2526 4359 2582 4366
rect 2526 4339 2555 4359
rect 2575 4339 2582 4359
rect 2526 4334 2582 4339
rect 2759 4362 2793 4369
rect 2759 4344 2767 4362
rect 2786 4344 2793 4362
rect 2759 4336 2793 4344
rect 3323 4356 3357 4562
rect 3563 4561 3602 4565
rect 3391 4535 3976 4541
rect 3391 4515 3407 4535
rect 3427 4534 3976 4535
rect 3427 4515 3947 4534
rect 3391 4514 3947 4515
rect 3967 4514 3976 4534
rect 3391 4506 3976 4514
rect 5803 4425 6388 4433
rect 5803 4405 5812 4425
rect 5832 4424 6388 4425
rect 5832 4405 6352 4424
rect 5803 4404 6352 4405
rect 6372 4404 6388 4424
rect 5803 4398 6388 4404
rect 5322 4394 5354 4395
rect 5319 4389 5354 4394
rect 5319 4369 5326 4389
rect 5346 4369 5354 4389
rect 6422 4377 6456 4576
rect 6400 4372 6456 4377
rect 5319 4361 5354 4369
rect 3323 4348 3358 4356
rect 2526 4128 2560 4334
rect 3323 4328 3331 4348
rect 3351 4328 3358 4348
rect 3323 4323 3358 4328
rect 3323 4322 3355 4323
rect 2594 4307 3179 4313
rect 2594 4287 2610 4307
rect 2630 4306 3179 4307
rect 2630 4287 3150 4306
rect 2594 4286 3150 4287
rect 3170 4286 3179 4306
rect 2594 4278 3179 4286
rect 3259 4277 3289 4278
rect 3259 4250 3595 4277
rect 3259 4249 3294 4250
rect 2526 4120 2561 4128
rect 2526 4100 2534 4120
rect 2554 4100 2561 4120
rect 2526 4095 2561 4100
rect 2526 4074 2560 4095
rect 3259 4074 3289 4249
rect 3345 4182 3380 4183
rect 2526 4048 3289 4074
rect 2527 4047 2560 4048
rect 3259 4046 3289 4048
rect 3324 4175 3380 4182
rect 3324 4155 3353 4175
rect 3373 4155 3380 4175
rect 3324 4150 3380 4155
rect 3559 4177 3594 4250
rect 3559 4157 3566 4177
rect 3586 4157 3594 4177
rect 4701 4203 5286 4211
rect 4701 4183 4710 4203
rect 4730 4202 5286 4203
rect 4730 4183 5250 4202
rect 4701 4182 5250 4183
rect 5270 4182 5286 4202
rect 4701 4176 5286 4182
rect 3559 4150 3594 4157
rect 5320 4155 5354 4361
rect 6182 4370 6217 4372
rect 6182 4364 6220 4370
rect 6182 4341 6190 4364
rect 6213 4341 6220 4364
rect 6400 4352 6407 4372
rect 6427 4352 6456 4372
rect 6400 4345 6456 4352
rect 6400 4344 6435 4345
rect 6182 4335 6220 4341
rect 6182 4322 6217 4335
rect 6180 4264 6217 4322
rect 2349 4025 2381 4026
rect 2349 4020 2689 4025
rect 2349 4002 2352 4020
rect 2374 4002 2689 4020
rect 2349 3997 2689 4002
rect 2349 3996 2381 3997
rect 2663 3962 2689 3997
rect 2448 3956 2483 3957
rect 2427 3949 2483 3956
rect 2427 3929 2456 3949
rect 2476 3929 2483 3949
rect 2427 3924 2483 3929
rect 2659 3953 2695 3962
rect 2659 3936 2667 3953
rect 2686 3936 2695 3953
rect 2659 3927 2695 3936
rect 3324 3944 3358 4150
rect 5084 4148 5119 4155
rect 3392 4123 3977 4129
rect 3392 4103 3408 4123
rect 3428 4122 3977 4123
rect 3428 4103 3948 4122
rect 3392 4102 3948 4103
rect 3968 4102 3977 4122
rect 3392 4094 3977 4102
rect 5084 4128 5092 4148
rect 5112 4128 5119 4148
rect 5084 4055 5119 4128
rect 5298 4150 5354 4155
rect 5298 4130 5305 4150
rect 5325 4130 5354 4150
rect 5298 4123 5354 4130
rect 5389 4257 5419 4259
rect 6118 4257 6151 4258
rect 5389 4231 6152 4257
rect 5298 4122 5333 4123
rect 5389 4056 5419 4231
rect 6118 4210 6152 4231
rect 6180 4247 6215 4264
rect 6180 4246 6474 4247
rect 6180 4245 6517 4246
rect 6180 4238 6522 4245
rect 6180 4212 6482 4238
rect 6513 4212 6522 4238
rect 6117 4205 6152 4210
rect 6473 4209 6522 4212
rect 6117 4185 6124 4205
rect 6144 4185 6152 4205
rect 6479 4204 6522 4209
rect 6117 4177 6152 4185
rect 5384 4055 5419 4056
rect 5083 4028 5419 4055
rect 5389 4027 5419 4028
rect 5499 4019 6084 4027
rect 5499 3999 5508 4019
rect 5528 4018 6084 4019
rect 5528 3999 6048 4018
rect 5499 3998 6048 3999
rect 6068 3998 6084 4018
rect 5499 3992 6084 3998
rect 5323 3982 5355 3983
rect 5320 3977 5355 3982
rect 5320 3957 5327 3977
rect 5347 3957 5355 3977
rect 6118 3971 6152 4177
rect 5320 3949 5355 3957
rect 3324 3936 3359 3944
rect 2427 3718 2461 3924
rect 3324 3916 3332 3936
rect 3352 3916 3359 3936
rect 3324 3911 3359 3916
rect 3324 3910 3356 3911
rect 2495 3897 3080 3903
rect 2495 3877 2511 3897
rect 2531 3896 3080 3897
rect 2531 3877 3051 3896
rect 2495 3876 3051 3877
rect 3071 3876 3080 3896
rect 2495 3868 3080 3876
rect 4702 3791 5287 3799
rect 4702 3771 4711 3791
rect 4731 3790 5287 3791
rect 4731 3771 5251 3790
rect 4702 3770 5251 3771
rect 5271 3770 5287 3790
rect 4702 3764 5287 3770
rect 5076 3740 5115 3744
rect 5321 3743 5355 3949
rect 5884 3964 5919 3970
rect 5884 3945 5889 3964
rect 5910 3945 5919 3964
rect 5884 3936 5919 3945
rect 6096 3966 6152 3971
rect 6096 3946 6103 3966
rect 6123 3946 6152 3966
rect 6096 3939 6152 3946
rect 6096 3938 6131 3939
rect 5888 3868 5917 3936
rect 5888 3834 6234 3868
rect 5076 3720 5084 3740
rect 5104 3720 5115 3740
rect 2427 3710 2462 3718
rect 2427 3690 2435 3710
rect 2455 3702 2462 3710
rect 2455 3690 2466 3702
rect 2427 3453 2466 3690
rect 3297 3667 3583 3668
rect 2782 3659 3585 3667
rect 2782 3642 2793 3659
rect 2783 3637 2793 3642
rect 2817 3642 3585 3659
rect 2817 3637 2822 3642
rect 2783 3624 2822 3637
rect 3327 3576 3362 3577
rect 3306 3569 3362 3576
rect 3306 3549 3335 3569
rect 3355 3549 3362 3569
rect 3306 3544 3362 3549
rect 3546 3567 3585 3642
rect 5076 3645 5115 3720
rect 5299 3738 5355 3743
rect 5299 3718 5306 3738
rect 5326 3718 5355 3738
rect 5299 3711 5355 3718
rect 5299 3710 5334 3711
rect 5839 3650 5878 3663
rect 5839 3645 5844 3650
rect 5076 3628 5844 3645
rect 5868 3645 5878 3650
rect 5868 3628 5879 3645
rect 5076 3620 5879 3628
rect 5078 3619 5364 3620
rect 6195 3597 6234 3834
rect 6195 3585 6206 3597
rect 6199 3577 6206 3585
rect 6226 3577 6234 3597
rect 6199 3569 6234 3577
rect 3546 3547 3557 3567
rect 3577 3547 3585 3567
rect 2427 3419 2773 3453
rect 2744 3351 2773 3419
rect 2530 3348 2565 3349
rect 2509 3341 2565 3348
rect 2509 3321 2538 3341
rect 2558 3321 2565 3341
rect 2509 3316 2565 3321
rect 2742 3342 2777 3351
rect 2742 3323 2751 3342
rect 2772 3323 2777 3342
rect 2742 3317 2777 3323
rect 3306 3338 3340 3544
rect 3546 3543 3585 3547
rect 3374 3517 3959 3523
rect 3374 3497 3390 3517
rect 3410 3516 3959 3517
rect 3410 3497 3930 3516
rect 3374 3496 3930 3497
rect 3950 3496 3959 3516
rect 3374 3488 3959 3496
rect 5581 3411 6166 3419
rect 5581 3391 5590 3411
rect 5610 3410 6166 3411
rect 5610 3391 6130 3410
rect 5581 3390 6130 3391
rect 6150 3390 6166 3410
rect 5581 3384 6166 3390
rect 5305 3376 5337 3377
rect 5302 3371 5337 3376
rect 5302 3351 5309 3371
rect 5329 3351 5337 3371
rect 6200 3363 6234 3569
rect 5302 3343 5337 3351
rect 3306 3330 3341 3338
rect 2509 3110 2543 3316
rect 3306 3310 3314 3330
rect 3334 3310 3341 3330
rect 3306 3305 3341 3310
rect 3306 3304 3338 3305
rect 2577 3289 3162 3295
rect 2577 3269 2593 3289
rect 2613 3288 3162 3289
rect 2613 3269 3133 3288
rect 2577 3268 3133 3269
rect 3153 3268 3162 3288
rect 2577 3260 3162 3268
rect 3242 3259 3272 3260
rect 3242 3232 3578 3259
rect 3242 3231 3277 3232
rect 2509 3102 2544 3110
rect 2509 3082 2517 3102
rect 2537 3082 2544 3102
rect 2509 3077 2544 3082
rect 2509 3056 2543 3077
rect 3242 3056 3272 3231
rect 3328 3164 3363 3165
rect 2509 3030 3272 3056
rect 2510 3029 2543 3030
rect 3242 3028 3272 3030
rect 3307 3157 3363 3164
rect 3307 3137 3336 3157
rect 3356 3137 3363 3157
rect 3307 3132 3363 3137
rect 3542 3159 3577 3232
rect 3542 3139 3549 3159
rect 3569 3139 3577 3159
rect 4684 3185 5269 3193
rect 4684 3165 4693 3185
rect 4713 3184 5269 3185
rect 4713 3165 5233 3184
rect 4684 3164 5233 3165
rect 5253 3164 5269 3184
rect 4684 3158 5269 3164
rect 3542 3132 3577 3139
rect 5303 3137 5337 3343
rect 5968 3357 5999 3363
rect 5968 3338 5973 3357
rect 5994 3338 5999 3357
rect 5968 3296 5999 3338
rect 6178 3358 6234 3363
rect 6178 3338 6185 3358
rect 6205 3338 6234 3358
rect 6178 3331 6234 3338
rect 6178 3330 6213 3331
rect 5968 3268 6307 3296
rect 2251 2973 2605 3009
rect 2267 2972 2605 2973
rect 2579 2942 2605 2972
rect 2365 2940 2400 2941
rect 2344 2933 2400 2940
rect 2344 2913 2373 2933
rect 2393 2913 2400 2933
rect 2344 2908 2400 2913
rect 2573 2934 2614 2942
rect 2573 2916 2586 2934
rect 2604 2916 2614 2934
rect 2344 2702 2378 2908
rect 2573 2905 2614 2916
rect 3307 2926 3341 3132
rect 5067 3130 5102 3137
rect 3375 3105 3960 3111
rect 3375 3085 3391 3105
rect 3411 3104 3960 3105
rect 3411 3085 3931 3104
rect 3375 3084 3931 3085
rect 3951 3084 3960 3104
rect 3375 3076 3960 3084
rect 5067 3110 5075 3130
rect 5095 3110 5102 3130
rect 5067 3037 5102 3110
rect 5281 3132 5337 3137
rect 5281 3112 5288 3132
rect 5308 3112 5337 3132
rect 5281 3105 5337 3112
rect 5372 3239 5402 3241
rect 6101 3239 6134 3240
rect 5372 3213 6135 3239
rect 5281 3104 5316 3105
rect 5372 3038 5402 3213
rect 6101 3192 6135 3213
rect 6100 3187 6135 3192
rect 6100 3167 6107 3187
rect 6127 3167 6135 3187
rect 6100 3159 6135 3167
rect 5367 3037 5402 3038
rect 5066 3010 5402 3037
rect 5372 3009 5402 3010
rect 5482 3001 6067 3009
rect 5482 2981 5491 3001
rect 5511 3000 6067 3001
rect 5511 2981 6031 3000
rect 5482 2980 6031 2981
rect 6051 2980 6067 3000
rect 5482 2974 6067 2980
rect 5306 2964 5338 2965
rect 5303 2959 5338 2964
rect 5303 2939 5310 2959
rect 5330 2939 5338 2959
rect 6101 2953 6135 3159
rect 5303 2931 5338 2939
rect 3307 2918 3342 2926
rect 3307 2898 3315 2918
rect 3335 2898 3342 2918
rect 3307 2893 3342 2898
rect 3307 2892 3339 2893
rect 2412 2881 2997 2887
rect 2412 2861 2428 2881
rect 2448 2880 2997 2881
rect 2448 2861 2968 2880
rect 2412 2860 2968 2861
rect 2988 2860 2997 2880
rect 2412 2852 2997 2860
rect 4685 2773 5270 2781
rect 4685 2753 4694 2773
rect 4714 2772 5270 2773
rect 4714 2753 5234 2772
rect 4685 2752 5234 2753
rect 5254 2752 5270 2772
rect 4685 2746 5270 2752
rect 5059 2722 5098 2726
rect 5304 2725 5338 2931
rect 5868 2943 5902 2951
rect 5868 2925 5875 2943
rect 5894 2925 5902 2943
rect 5868 2918 5902 2925
rect 6079 2948 6135 2953
rect 6079 2928 6086 2948
rect 6106 2928 6135 2948
rect 6079 2921 6135 2928
rect 6079 2920 6114 2921
rect 5872 2888 5901 2918
rect 5872 2880 6254 2888
rect 5872 2861 6225 2880
rect 6246 2861 6254 2880
rect 5872 2856 6254 2861
rect 5059 2702 5067 2722
rect 5087 2702 5098 2722
rect 2344 2701 2379 2702
rect 2312 2694 2379 2701
rect 2312 2674 2352 2694
rect 2372 2674 2379 2694
rect 2312 2671 2379 2674
rect 2312 2668 2377 2671
rect 1883 2567 1948 2570
rect 1881 2564 1948 2567
rect 1881 2544 1888 2564
rect 1908 2544 1948 2564
rect 1881 2537 1948 2544
rect 1881 2536 1916 2537
rect 1263 2378 1848 2386
rect 1263 2358 1272 2378
rect 1292 2377 1848 2378
rect 1292 2358 1812 2377
rect 1263 2357 1812 2358
rect 1832 2357 1848 2377
rect 1263 2351 1848 2357
rect 921 2345 953 2346
rect 918 2340 953 2345
rect 918 2320 925 2340
rect 945 2320 953 2340
rect 918 2312 953 2320
rect 300 2154 885 2162
rect 300 2134 309 2154
rect 329 2153 885 2154
rect 329 2134 849 2153
rect 300 2133 849 2134
rect 869 2133 885 2153
rect 300 2127 885 2133
rect 919 2106 953 2312
rect 1648 2327 1681 2333
rect 1882 2330 1916 2536
rect 1648 2305 1653 2327
rect 1676 2305 1681 2327
rect 1648 2296 1681 2305
rect 1860 2325 1916 2330
rect 1860 2305 1867 2325
rect 1887 2305 1916 2325
rect 1860 2298 1916 2305
rect 1860 2297 1895 2298
rect 1650 2265 1677 2296
rect 2072 2265 2111 2277
rect 1650 2264 2113 2265
rect 1650 2242 2077 2264
rect 2101 2242 2113 2264
rect 1650 2234 2113 2242
rect 683 2099 718 2106
rect 683 2079 691 2099
rect 711 2079 718 2099
rect 683 2006 718 2079
rect 897 2101 953 2106
rect 897 2081 904 2101
rect 924 2081 953 2101
rect 897 2074 953 2081
rect 988 2208 1018 2210
rect 1717 2208 1750 2209
rect 988 2182 1751 2208
rect 897 2073 932 2074
rect 988 2007 1018 2182
rect 1717 2161 1751 2182
rect 1716 2156 1751 2161
rect 1716 2136 1723 2156
rect 1743 2136 1751 2156
rect 1716 2128 1751 2136
rect 983 2006 1018 2007
rect 682 1979 1018 2006
rect 988 1978 1018 1979
rect 1098 1970 1683 1978
rect 1098 1950 1107 1970
rect 1127 1969 1683 1970
rect 1127 1950 1647 1969
rect 1098 1949 1647 1950
rect 1667 1949 1683 1969
rect 1098 1943 1683 1949
rect 922 1933 954 1934
rect 919 1928 954 1933
rect 919 1908 926 1928
rect 946 1908 954 1928
rect 1717 1922 1751 2128
rect 919 1900 954 1908
rect 301 1742 886 1750
rect 301 1722 310 1742
rect 330 1741 886 1742
rect 330 1722 850 1741
rect 301 1721 850 1722
rect 870 1721 886 1741
rect 301 1715 886 1721
rect 675 1691 714 1695
rect 920 1694 954 1900
rect 1483 1915 1518 1921
rect 1483 1896 1488 1915
rect 1509 1896 1518 1915
rect 1483 1887 1518 1896
rect 1695 1917 1751 1922
rect 1695 1897 1702 1917
rect 1722 1897 1751 1917
rect 1695 1890 1751 1897
rect 1873 2068 1905 2080
rect 1873 2050 1880 2068
rect 1902 2050 1905 2068
rect 1695 1889 1730 1890
rect 1487 1819 1516 1887
rect 1487 1785 1833 1819
rect 675 1671 683 1691
rect 703 1671 714 1691
rect 675 1596 714 1671
rect 898 1689 954 1694
rect 898 1669 905 1689
rect 925 1669 954 1689
rect 898 1662 954 1669
rect 898 1661 933 1662
rect 1438 1601 1477 1614
rect 1438 1596 1443 1601
rect 675 1579 1443 1596
rect 1467 1596 1477 1601
rect 1467 1579 1478 1596
rect 675 1571 1478 1579
rect 677 1570 963 1571
rect 1794 1548 1833 1785
rect 1794 1536 1805 1548
rect 1798 1528 1805 1536
rect 1825 1528 1833 1548
rect 1798 1520 1833 1528
rect 1180 1362 1765 1370
rect 1180 1342 1189 1362
rect 1209 1361 1765 1362
rect 1209 1342 1729 1361
rect 1180 1341 1729 1342
rect 1749 1341 1765 1361
rect 1180 1335 1765 1341
rect 904 1327 936 1328
rect 901 1322 936 1327
rect 901 1302 908 1322
rect 928 1302 936 1322
rect 1799 1314 1833 1520
rect 901 1294 936 1302
rect 283 1136 868 1144
rect 283 1116 292 1136
rect 312 1135 868 1136
rect 312 1116 832 1135
rect 283 1115 832 1116
rect 852 1115 868 1135
rect 283 1109 868 1115
rect 902 1088 936 1294
rect 1565 1302 1601 1311
rect 1565 1285 1574 1302
rect 1593 1285 1601 1302
rect 1565 1276 1601 1285
rect 1777 1309 1833 1314
rect 1777 1289 1784 1309
rect 1804 1289 1833 1309
rect 1777 1282 1833 1289
rect 1777 1281 1812 1282
rect 1571 1241 1597 1276
rect 1873 1241 1905 2050
rect 2317 1983 2346 2668
rect 3277 2649 3563 2650
rect 2762 2641 3565 2649
rect 2762 2624 2773 2641
rect 2763 2619 2773 2624
rect 2797 2624 3565 2641
rect 2797 2619 2802 2624
rect 2763 2606 2802 2619
rect 3307 2558 3342 2559
rect 3286 2551 3342 2558
rect 3286 2531 3315 2551
rect 3335 2531 3342 2551
rect 3286 2526 3342 2531
rect 3526 2549 3565 2624
rect 5059 2627 5098 2702
rect 5282 2720 5338 2725
rect 5282 2700 5289 2720
rect 5309 2700 5338 2720
rect 5282 2693 5338 2700
rect 5282 2692 5317 2693
rect 5822 2632 5861 2645
rect 5822 2627 5827 2632
rect 5059 2610 5827 2627
rect 5851 2627 5861 2632
rect 5851 2610 5862 2627
rect 5059 2602 5862 2610
rect 5061 2601 5347 2602
rect 6278 2583 6307 3268
rect 6615 3022 6642 4722
rect 7678 4698 7964 4699
rect 7163 4690 7966 4698
rect 7163 4673 7174 4690
rect 7164 4668 7174 4673
rect 7198 4673 7966 4690
rect 7198 4668 7203 4673
rect 7164 4655 7203 4668
rect 7708 4607 7743 4608
rect 7687 4600 7743 4607
rect 7687 4580 7716 4600
rect 7736 4580 7743 4600
rect 7687 4575 7743 4580
rect 7927 4598 7966 4673
rect 7927 4578 7938 4598
rect 7958 4578 7966 4598
rect 6771 4439 7153 4444
rect 6771 4420 6779 4439
rect 6800 4420 7153 4439
rect 6771 4412 7153 4420
rect 7124 4382 7153 4412
rect 6911 4379 6946 4380
rect 6890 4372 6946 4379
rect 6890 4352 6919 4372
rect 6939 4352 6946 4372
rect 6890 4347 6946 4352
rect 7123 4375 7157 4382
rect 7123 4357 7131 4375
rect 7150 4357 7157 4375
rect 7123 4349 7157 4357
rect 7687 4369 7721 4575
rect 7927 4574 7966 4578
rect 7755 4548 8340 4554
rect 7755 4528 7771 4548
rect 7791 4547 8340 4548
rect 7791 4528 8311 4547
rect 7755 4527 8311 4528
rect 8331 4527 8340 4547
rect 7755 4519 8340 4527
rect 7687 4361 7722 4369
rect 6890 4141 6924 4347
rect 7687 4341 7695 4361
rect 7715 4341 7722 4361
rect 7687 4336 7722 4341
rect 7687 4335 7719 4336
rect 6958 4320 7543 4326
rect 6958 4300 6974 4320
rect 6994 4319 7543 4320
rect 6994 4300 7514 4319
rect 6958 4299 7514 4300
rect 7534 4299 7543 4319
rect 6958 4291 7543 4299
rect 7623 4290 7653 4291
rect 7623 4263 7959 4290
rect 7623 4262 7658 4263
rect 6890 4133 6925 4141
rect 6890 4113 6898 4133
rect 6918 4113 6925 4133
rect 6890 4108 6925 4113
rect 6890 4087 6924 4108
rect 7623 4087 7653 4262
rect 7709 4195 7744 4196
rect 6890 4061 7653 4087
rect 6891 4060 6924 4061
rect 7623 4059 7653 4061
rect 7688 4188 7744 4195
rect 7688 4168 7717 4188
rect 7737 4168 7744 4188
rect 7688 4163 7744 4168
rect 7923 4190 7958 4263
rect 7923 4170 7930 4190
rect 7950 4170 7958 4190
rect 7923 4163 7958 4170
rect 6713 4038 6745 4039
rect 6713 4033 7053 4038
rect 6713 4015 6716 4033
rect 6738 4015 7053 4033
rect 6713 4010 7053 4015
rect 6713 4009 6745 4010
rect 7027 3975 7053 4010
rect 6812 3969 6847 3970
rect 6791 3962 6847 3969
rect 6791 3942 6820 3962
rect 6840 3942 6847 3962
rect 6791 3937 6847 3942
rect 7023 3966 7059 3975
rect 7023 3949 7031 3966
rect 7050 3949 7059 3966
rect 7023 3940 7059 3949
rect 7688 3957 7722 4163
rect 7756 4136 8341 4142
rect 7756 4116 7772 4136
rect 7792 4135 8341 4136
rect 7792 4116 8312 4135
rect 7756 4115 8312 4116
rect 8332 4115 8341 4135
rect 7756 4107 8341 4115
rect 7688 3949 7723 3957
rect 6791 3731 6825 3937
rect 7688 3929 7696 3949
rect 7716 3929 7723 3949
rect 7688 3924 7723 3929
rect 7688 3923 7720 3924
rect 6859 3910 7444 3916
rect 6859 3890 6875 3910
rect 6895 3909 7444 3910
rect 6895 3890 7415 3909
rect 6859 3889 7415 3890
rect 7435 3889 7444 3909
rect 6859 3881 7444 3889
rect 6791 3723 6826 3731
rect 6791 3703 6799 3723
rect 6819 3715 6826 3723
rect 6819 3703 6830 3715
rect 6791 3466 6830 3703
rect 7661 3680 7947 3681
rect 7146 3672 7949 3680
rect 7146 3655 7157 3672
rect 7147 3650 7157 3655
rect 7181 3655 7949 3672
rect 7181 3650 7186 3655
rect 7147 3637 7186 3650
rect 7691 3589 7726 3590
rect 7670 3582 7726 3589
rect 7670 3562 7699 3582
rect 7719 3562 7726 3582
rect 7670 3557 7726 3562
rect 7910 3580 7949 3655
rect 7910 3560 7921 3580
rect 7941 3560 7949 3580
rect 6791 3432 7137 3466
rect 7108 3364 7137 3432
rect 6894 3361 6929 3362
rect 6873 3354 6929 3361
rect 6873 3334 6902 3354
rect 6922 3334 6929 3354
rect 6873 3329 6929 3334
rect 7106 3355 7141 3364
rect 7106 3336 7115 3355
rect 7136 3336 7141 3355
rect 7106 3330 7141 3336
rect 7670 3351 7704 3557
rect 7910 3556 7949 3560
rect 7738 3530 8323 3536
rect 7738 3510 7754 3530
rect 7774 3529 8323 3530
rect 7774 3510 8294 3529
rect 7738 3509 8294 3510
rect 8314 3509 8323 3529
rect 7738 3501 8323 3509
rect 7670 3343 7705 3351
rect 6873 3123 6907 3329
rect 7670 3323 7678 3343
rect 7698 3323 7705 3343
rect 7670 3318 7705 3323
rect 7670 3317 7702 3318
rect 6941 3302 7526 3308
rect 6941 3282 6957 3302
rect 6977 3301 7526 3302
rect 6977 3282 7497 3301
rect 6941 3281 7497 3282
rect 7517 3281 7526 3301
rect 6941 3273 7526 3281
rect 7606 3272 7636 3273
rect 7606 3245 7942 3272
rect 7606 3244 7641 3245
rect 6873 3115 6908 3123
rect 6873 3095 6881 3115
rect 6901 3095 6908 3115
rect 6873 3090 6908 3095
rect 6873 3069 6907 3090
rect 7606 3069 7636 3244
rect 7692 3177 7727 3178
rect 6873 3043 7636 3069
rect 6874 3042 6907 3043
rect 7606 3041 7636 3043
rect 7671 3170 7727 3177
rect 7671 3150 7700 3170
rect 7720 3150 7727 3170
rect 7671 3145 7727 3150
rect 7906 3172 7941 3245
rect 7906 3152 7913 3172
rect 7933 3152 7941 3172
rect 7906 3145 7941 3152
rect 6615 2986 6969 3022
rect 6631 2985 6969 2986
rect 6943 2955 6969 2985
rect 6729 2953 6764 2954
rect 6708 2946 6764 2953
rect 6708 2926 6737 2946
rect 6757 2926 6764 2946
rect 6708 2921 6764 2926
rect 6937 2947 6978 2955
rect 6937 2929 6950 2947
rect 6968 2929 6978 2947
rect 6708 2715 6742 2921
rect 6937 2918 6978 2929
rect 7671 2939 7705 3145
rect 7739 3118 8324 3124
rect 7739 3098 7755 3118
rect 7775 3117 8324 3118
rect 7775 3098 8295 3117
rect 7739 3097 8295 3098
rect 8315 3097 8324 3117
rect 7739 3089 8324 3097
rect 7671 2931 7706 2939
rect 7671 2911 7679 2931
rect 7699 2911 7706 2931
rect 7671 2906 7706 2911
rect 7671 2905 7703 2906
rect 6776 2894 7361 2900
rect 6776 2874 6792 2894
rect 6812 2893 7361 2894
rect 6812 2874 7332 2893
rect 6776 2873 7332 2874
rect 7352 2873 7361 2893
rect 6776 2865 7361 2873
rect 6708 2714 6743 2715
rect 6676 2707 6743 2714
rect 6676 2687 6716 2707
rect 6736 2687 6743 2707
rect 6676 2684 6743 2687
rect 6676 2681 6741 2684
rect 6247 2580 6312 2583
rect 6245 2577 6312 2580
rect 6245 2557 6252 2577
rect 6272 2557 6312 2577
rect 6245 2550 6312 2557
rect 6245 2549 6280 2550
rect 3526 2529 3537 2549
rect 3557 2529 3565 2549
rect 2370 2390 2752 2395
rect 2370 2371 2378 2390
rect 2399 2371 2752 2390
rect 2370 2363 2752 2371
rect 2723 2333 2752 2363
rect 2510 2330 2545 2331
rect 2489 2323 2545 2330
rect 2489 2303 2518 2323
rect 2538 2303 2545 2323
rect 2489 2298 2545 2303
rect 2722 2326 2756 2333
rect 2722 2308 2730 2326
rect 2749 2308 2756 2326
rect 2722 2300 2756 2308
rect 3286 2320 3320 2526
rect 3526 2525 3565 2529
rect 3354 2499 3939 2505
rect 3354 2479 3370 2499
rect 3390 2498 3939 2499
rect 3390 2479 3910 2498
rect 3354 2478 3910 2479
rect 3930 2478 3939 2498
rect 3354 2470 3939 2478
rect 5627 2391 6212 2399
rect 5627 2371 5636 2391
rect 5656 2390 6212 2391
rect 5656 2371 6176 2390
rect 5627 2370 6176 2371
rect 6196 2370 6212 2390
rect 5627 2364 6212 2370
rect 5285 2358 5317 2359
rect 5282 2353 5317 2358
rect 5282 2333 5289 2353
rect 5309 2333 5317 2353
rect 5282 2325 5317 2333
rect 3286 2312 3321 2320
rect 2489 2092 2523 2298
rect 3286 2292 3294 2312
rect 3314 2292 3321 2312
rect 3286 2287 3321 2292
rect 3286 2286 3318 2287
rect 2557 2271 3142 2277
rect 2557 2251 2573 2271
rect 2593 2270 3142 2271
rect 2593 2251 3113 2270
rect 2557 2250 3113 2251
rect 3133 2250 3142 2270
rect 2557 2242 3142 2250
rect 3222 2241 3252 2242
rect 3222 2214 3558 2241
rect 3222 2213 3257 2214
rect 2489 2084 2524 2092
rect 2489 2064 2497 2084
rect 2517 2064 2524 2084
rect 2489 2059 2524 2064
rect 2489 2038 2523 2059
rect 3222 2038 3252 2213
rect 3308 2146 3343 2147
rect 2489 2012 3252 2038
rect 2490 2011 2523 2012
rect 3222 2010 3252 2012
rect 3287 2139 3343 2146
rect 3287 2119 3316 2139
rect 3336 2119 3343 2139
rect 3287 2114 3343 2119
rect 3522 2141 3557 2214
rect 3522 2121 3529 2141
rect 3549 2121 3557 2141
rect 4664 2167 5249 2175
rect 4664 2147 4673 2167
rect 4693 2166 5249 2167
rect 4693 2147 5213 2166
rect 4664 2146 5213 2147
rect 5233 2146 5249 2166
rect 4664 2140 5249 2146
rect 3522 2114 3557 2121
rect 5283 2119 5317 2325
rect 6012 2340 6045 2346
rect 6246 2343 6280 2549
rect 6012 2318 6017 2340
rect 6040 2318 6045 2340
rect 6012 2309 6045 2318
rect 6224 2338 6280 2343
rect 6224 2318 6231 2338
rect 6251 2318 6280 2338
rect 6224 2311 6280 2318
rect 6224 2310 6259 2311
rect 6014 2278 6041 2309
rect 6436 2278 6475 2290
rect 6014 2277 6477 2278
rect 6014 2255 6441 2277
rect 6465 2255 6477 2277
rect 6014 2247 6477 2255
rect 2317 1955 2656 1983
rect 2411 1920 2446 1921
rect 2390 1913 2446 1920
rect 2390 1893 2419 1913
rect 2439 1893 2446 1913
rect 2390 1888 2446 1893
rect 2625 1913 2656 1955
rect 2625 1894 2630 1913
rect 2651 1894 2656 1913
rect 2625 1888 2656 1894
rect 3287 1908 3321 2114
rect 5047 2112 5082 2119
rect 3355 2087 3940 2093
rect 3355 2067 3371 2087
rect 3391 2086 3940 2087
rect 3391 2067 3911 2086
rect 3355 2066 3911 2067
rect 3931 2066 3940 2086
rect 3355 2058 3940 2066
rect 5047 2092 5055 2112
rect 5075 2092 5082 2112
rect 5047 2019 5082 2092
rect 5261 2114 5317 2119
rect 5261 2094 5268 2114
rect 5288 2094 5317 2114
rect 5261 2087 5317 2094
rect 5352 2221 5382 2223
rect 6081 2221 6114 2222
rect 5352 2195 6115 2221
rect 5261 2086 5296 2087
rect 5352 2020 5382 2195
rect 6081 2174 6115 2195
rect 6080 2169 6115 2174
rect 6080 2149 6087 2169
rect 6107 2149 6115 2169
rect 6080 2141 6115 2149
rect 5347 2019 5382 2020
rect 5046 1992 5382 2019
rect 5352 1991 5382 1992
rect 5462 1983 6047 1991
rect 5462 1963 5471 1983
rect 5491 1982 6047 1983
rect 5491 1963 6011 1982
rect 5462 1962 6011 1963
rect 6031 1962 6047 1982
rect 5462 1956 6047 1962
rect 5286 1946 5318 1947
rect 5283 1941 5318 1946
rect 5283 1921 5290 1941
rect 5310 1921 5318 1941
rect 6081 1935 6115 2141
rect 5283 1913 5318 1921
rect 3287 1900 3322 1908
rect 2390 1682 2424 1888
rect 3287 1880 3295 1900
rect 3315 1880 3322 1900
rect 3287 1875 3322 1880
rect 3287 1874 3319 1875
rect 2458 1861 3043 1867
rect 2458 1841 2474 1861
rect 2494 1860 3043 1861
rect 2494 1841 3014 1860
rect 2458 1840 3014 1841
rect 3034 1840 3043 1860
rect 2458 1832 3043 1840
rect 4665 1755 5250 1763
rect 4665 1735 4674 1755
rect 4694 1754 5250 1755
rect 4694 1735 5214 1754
rect 4665 1734 5214 1735
rect 5234 1734 5250 1754
rect 4665 1728 5250 1734
rect 5039 1704 5078 1708
rect 5284 1707 5318 1913
rect 5847 1928 5882 1934
rect 5847 1909 5852 1928
rect 5873 1909 5882 1928
rect 5847 1900 5882 1909
rect 6059 1930 6115 1935
rect 6059 1910 6066 1930
rect 6086 1910 6115 1930
rect 6059 1903 6115 1910
rect 6237 2081 6269 2093
rect 6237 2063 6244 2081
rect 6266 2063 6269 2081
rect 6059 1902 6094 1903
rect 5851 1832 5880 1900
rect 5851 1798 6197 1832
rect 5039 1684 5047 1704
rect 5067 1684 5078 1704
rect 2390 1674 2425 1682
rect 2390 1654 2398 1674
rect 2418 1666 2425 1674
rect 2418 1654 2429 1666
rect 2390 1417 2429 1654
rect 3260 1631 3546 1632
rect 2745 1623 3548 1631
rect 2745 1606 2756 1623
rect 2746 1601 2756 1606
rect 2780 1606 3548 1623
rect 2780 1601 2785 1606
rect 2746 1588 2785 1601
rect 3290 1540 3325 1541
rect 3269 1533 3325 1540
rect 3269 1513 3298 1533
rect 3318 1513 3325 1533
rect 3269 1508 3325 1513
rect 3509 1531 3548 1606
rect 5039 1609 5078 1684
rect 5262 1702 5318 1707
rect 5262 1682 5269 1702
rect 5289 1682 5318 1702
rect 5262 1675 5318 1682
rect 5262 1674 5297 1675
rect 5802 1614 5841 1627
rect 5802 1609 5807 1614
rect 5039 1592 5807 1609
rect 5831 1609 5841 1614
rect 5831 1592 5842 1609
rect 5039 1584 5842 1592
rect 5041 1583 5327 1584
rect 6158 1561 6197 1798
rect 6158 1549 6169 1561
rect 6162 1541 6169 1549
rect 6189 1541 6197 1561
rect 6162 1533 6197 1541
rect 3509 1511 3520 1531
rect 3540 1511 3548 1531
rect 2390 1383 2736 1417
rect 2707 1315 2736 1383
rect 2493 1312 2528 1313
rect 1571 1213 1905 1241
rect 2472 1305 2528 1312
rect 2472 1285 2501 1305
rect 2521 1285 2528 1305
rect 2472 1280 2528 1285
rect 2705 1306 2740 1315
rect 2705 1287 2714 1306
rect 2735 1287 2740 1306
rect 2705 1281 2740 1287
rect 3269 1302 3303 1508
rect 3509 1507 3548 1511
rect 3337 1481 3922 1487
rect 3337 1461 3353 1481
rect 3373 1480 3922 1481
rect 3373 1461 3893 1480
rect 3337 1460 3893 1461
rect 3913 1460 3922 1480
rect 3337 1452 3922 1460
rect 5544 1375 6129 1383
rect 5544 1355 5553 1375
rect 5573 1374 6129 1375
rect 5573 1355 6093 1374
rect 5544 1354 6093 1355
rect 6113 1354 6129 1374
rect 5544 1348 6129 1354
rect 5268 1340 5300 1341
rect 5265 1335 5300 1340
rect 5265 1315 5272 1335
rect 5292 1315 5300 1335
rect 6163 1327 6197 1533
rect 5265 1307 5300 1315
rect 3269 1294 3304 1302
rect 666 1081 701 1088
rect 666 1061 674 1081
rect 694 1061 701 1081
rect 666 988 701 1061
rect 880 1083 936 1088
rect 880 1063 887 1083
rect 907 1063 936 1083
rect 880 1056 936 1063
rect 971 1190 1001 1192
rect 1700 1190 1733 1191
rect 971 1164 1734 1190
rect 880 1055 915 1056
rect 971 989 1001 1164
rect 1700 1143 1734 1164
rect 1699 1138 1734 1143
rect 1699 1118 1706 1138
rect 1726 1118 1734 1138
rect 1699 1110 1734 1118
rect 966 988 1001 989
rect 665 961 1001 988
rect 971 960 1001 961
rect 1081 952 1666 960
rect 1081 932 1090 952
rect 1110 951 1666 952
rect 1110 932 1630 951
rect 1081 931 1630 932
rect 1650 931 1666 951
rect 1081 925 1666 931
rect 905 915 937 916
rect 902 910 937 915
rect 902 890 909 910
rect 929 890 937 910
rect 1700 904 1734 1110
rect 2472 1074 2506 1280
rect 3269 1274 3277 1294
rect 3297 1274 3304 1294
rect 3269 1269 3304 1274
rect 3269 1268 3301 1269
rect 2540 1253 3125 1259
rect 2540 1233 2556 1253
rect 2576 1252 3125 1253
rect 2576 1233 3096 1252
rect 2540 1232 3096 1233
rect 3116 1232 3125 1252
rect 2540 1224 3125 1232
rect 3205 1223 3235 1224
rect 3205 1196 3541 1223
rect 3205 1195 3240 1196
rect 2472 1066 2507 1074
rect 2472 1046 2480 1066
rect 2500 1046 2507 1066
rect 2472 1041 2507 1046
rect 2472 1020 2506 1041
rect 3205 1020 3235 1195
rect 3291 1128 3326 1129
rect 2472 994 3235 1020
rect 2473 993 2506 994
rect 3205 992 3235 994
rect 3270 1121 3326 1128
rect 3270 1101 3299 1121
rect 3319 1101 3326 1121
rect 3270 1096 3326 1101
rect 3505 1123 3540 1196
rect 3505 1103 3512 1123
rect 3532 1103 3540 1123
rect 4647 1149 5232 1157
rect 4647 1129 4656 1149
rect 4676 1148 5232 1149
rect 4676 1129 5196 1148
rect 4647 1128 5196 1129
rect 5216 1128 5232 1148
rect 4647 1122 5232 1128
rect 3505 1096 3540 1103
rect 5266 1101 5300 1307
rect 5929 1315 5965 1324
rect 5929 1298 5938 1315
rect 5957 1298 5965 1315
rect 5929 1289 5965 1298
rect 6141 1322 6197 1327
rect 6141 1302 6148 1322
rect 6168 1302 6197 1322
rect 6141 1295 6197 1302
rect 6141 1294 6176 1295
rect 5935 1254 5961 1289
rect 6237 1254 6269 2063
rect 6681 1996 6710 2681
rect 7641 2662 7927 2663
rect 7126 2654 7929 2662
rect 7126 2637 7137 2654
rect 7127 2632 7137 2637
rect 7161 2637 7929 2654
rect 7161 2632 7166 2637
rect 7127 2619 7166 2632
rect 7671 2571 7706 2572
rect 7650 2564 7706 2571
rect 7650 2544 7679 2564
rect 7699 2544 7706 2564
rect 7650 2539 7706 2544
rect 7890 2562 7929 2637
rect 7890 2542 7901 2562
rect 7921 2542 7929 2562
rect 6734 2403 7116 2408
rect 6734 2384 6742 2403
rect 6763 2384 7116 2403
rect 6734 2376 7116 2384
rect 7087 2346 7116 2376
rect 6874 2343 6909 2344
rect 6853 2336 6909 2343
rect 6853 2316 6882 2336
rect 6902 2316 6909 2336
rect 6853 2311 6909 2316
rect 7086 2339 7120 2346
rect 7086 2321 7094 2339
rect 7113 2321 7120 2339
rect 7086 2313 7120 2321
rect 7650 2333 7684 2539
rect 7890 2538 7929 2542
rect 7718 2512 8303 2518
rect 7718 2492 7734 2512
rect 7754 2511 8303 2512
rect 7754 2492 8274 2511
rect 7718 2491 8274 2492
rect 8294 2491 8303 2511
rect 7718 2483 8303 2491
rect 7650 2325 7685 2333
rect 6853 2105 6887 2311
rect 7650 2305 7658 2325
rect 7678 2305 7685 2325
rect 7650 2300 7685 2305
rect 7650 2299 7682 2300
rect 6921 2284 7506 2290
rect 6921 2264 6937 2284
rect 6957 2283 7506 2284
rect 6957 2264 7477 2283
rect 6921 2263 7477 2264
rect 7497 2263 7506 2283
rect 6921 2255 7506 2263
rect 7586 2254 7616 2255
rect 7586 2227 7922 2254
rect 7586 2226 7621 2227
rect 6853 2097 6888 2105
rect 6853 2077 6861 2097
rect 6881 2077 6888 2097
rect 6853 2072 6888 2077
rect 6853 2051 6887 2072
rect 7586 2051 7616 2226
rect 7672 2159 7707 2160
rect 6853 2025 7616 2051
rect 6854 2024 6887 2025
rect 7586 2023 7616 2025
rect 7651 2152 7707 2159
rect 7651 2132 7680 2152
rect 7700 2132 7707 2152
rect 7651 2127 7707 2132
rect 7886 2154 7921 2227
rect 7886 2134 7893 2154
rect 7913 2134 7921 2154
rect 7886 2127 7921 2134
rect 6681 1968 7020 1996
rect 6775 1933 6810 1934
rect 6754 1926 6810 1933
rect 6754 1906 6783 1926
rect 6803 1906 6810 1926
rect 6754 1901 6810 1906
rect 6989 1926 7020 1968
rect 6989 1907 6994 1926
rect 7015 1907 7020 1926
rect 6989 1901 7020 1907
rect 7651 1921 7685 2127
rect 7719 2100 8304 2106
rect 7719 2080 7735 2100
rect 7755 2099 8304 2100
rect 7755 2080 8275 2099
rect 7719 2079 8275 2080
rect 8295 2079 8304 2099
rect 7719 2071 8304 2079
rect 7651 1913 7686 1921
rect 6754 1695 6788 1901
rect 7651 1893 7659 1913
rect 7679 1893 7686 1913
rect 7651 1888 7686 1893
rect 7651 1887 7683 1888
rect 6822 1874 7407 1880
rect 6822 1854 6838 1874
rect 6858 1873 7407 1874
rect 6858 1854 7378 1873
rect 6822 1853 7378 1854
rect 7398 1853 7407 1873
rect 6822 1845 7407 1853
rect 6754 1687 6789 1695
rect 6754 1667 6762 1687
rect 6782 1679 6789 1687
rect 6782 1667 6793 1679
rect 6754 1430 6793 1667
rect 7624 1644 7910 1645
rect 7109 1636 7912 1644
rect 7109 1619 7120 1636
rect 7110 1614 7120 1619
rect 7144 1619 7912 1636
rect 7144 1614 7149 1619
rect 7110 1601 7149 1614
rect 7654 1553 7689 1554
rect 7633 1546 7689 1553
rect 7633 1526 7662 1546
rect 7682 1526 7689 1546
rect 7633 1521 7689 1526
rect 7873 1544 7912 1619
rect 7873 1524 7884 1544
rect 7904 1524 7912 1544
rect 6754 1396 7100 1430
rect 7071 1328 7100 1396
rect 6857 1325 6892 1326
rect 5935 1226 6269 1254
rect 6836 1318 6892 1325
rect 6836 1298 6865 1318
rect 6885 1298 6892 1318
rect 6836 1293 6892 1298
rect 7069 1319 7104 1328
rect 7069 1300 7078 1319
rect 7099 1300 7104 1319
rect 7069 1294 7104 1300
rect 7633 1315 7667 1521
rect 7873 1520 7912 1524
rect 7701 1494 8286 1500
rect 7701 1474 7717 1494
rect 7737 1493 8286 1494
rect 7737 1474 8257 1493
rect 7701 1473 8257 1474
rect 8277 1473 8286 1493
rect 7701 1465 8286 1473
rect 7633 1307 7668 1315
rect 902 882 937 890
rect 284 724 869 732
rect 284 704 293 724
rect 313 723 869 724
rect 313 704 833 723
rect 284 703 833 704
rect 853 703 869 723
rect 284 697 869 703
rect 658 673 697 677
rect 903 676 937 882
rect 1467 894 1501 902
rect 1467 876 1474 894
rect 1493 876 1501 894
rect 1467 869 1501 876
rect 1678 899 1734 904
rect 1678 879 1685 899
rect 1705 879 1734 899
rect 1678 872 1734 879
rect 3270 890 3304 1096
rect 5030 1094 5065 1101
rect 3338 1069 3923 1075
rect 3338 1049 3354 1069
rect 3374 1068 3923 1069
rect 3374 1049 3894 1068
rect 3338 1048 3894 1049
rect 3914 1048 3923 1068
rect 3338 1040 3923 1048
rect 5030 1074 5038 1094
rect 5058 1074 5065 1094
rect 5030 1001 5065 1074
rect 5244 1096 5300 1101
rect 5244 1076 5251 1096
rect 5271 1076 5300 1096
rect 5244 1069 5300 1076
rect 5335 1203 5365 1205
rect 6064 1203 6097 1204
rect 5335 1177 6098 1203
rect 5244 1068 5279 1069
rect 5335 1002 5365 1177
rect 6064 1156 6098 1177
rect 6063 1151 6098 1156
rect 6063 1131 6070 1151
rect 6090 1131 6098 1151
rect 6063 1123 6098 1131
rect 5330 1001 5365 1002
rect 5029 974 5365 1001
rect 5335 973 5365 974
rect 5445 965 6030 973
rect 5445 945 5454 965
rect 5474 964 6030 965
rect 5474 945 5994 964
rect 5445 944 5994 945
rect 6014 944 6030 964
rect 5445 938 6030 944
rect 5269 928 5301 929
rect 5266 923 5301 928
rect 5266 903 5273 923
rect 5293 903 5301 923
rect 6064 917 6098 1123
rect 6836 1087 6870 1293
rect 7633 1287 7641 1307
rect 7661 1287 7668 1307
rect 7633 1282 7668 1287
rect 7633 1281 7665 1282
rect 6904 1266 7489 1272
rect 6904 1246 6920 1266
rect 6940 1265 7489 1266
rect 6940 1246 7460 1265
rect 6904 1245 7460 1246
rect 7480 1245 7489 1265
rect 6904 1237 7489 1245
rect 7569 1236 7599 1237
rect 7569 1209 7905 1236
rect 7569 1208 7604 1209
rect 6836 1079 6871 1087
rect 6836 1059 6844 1079
rect 6864 1059 6871 1079
rect 6836 1054 6871 1059
rect 6836 1033 6870 1054
rect 7569 1033 7599 1208
rect 7655 1141 7690 1142
rect 6836 1007 7599 1033
rect 6837 1006 6870 1007
rect 7569 1005 7599 1007
rect 7634 1134 7690 1141
rect 7634 1114 7663 1134
rect 7683 1114 7690 1134
rect 7634 1109 7690 1114
rect 7869 1136 7904 1209
rect 7869 1116 7876 1136
rect 7896 1116 7904 1136
rect 7869 1109 7904 1116
rect 5266 895 5301 903
rect 3270 882 3305 890
rect 1678 871 1713 872
rect 1471 839 1500 869
rect 3270 862 3278 882
rect 3298 862 3305 882
rect 3270 857 3305 862
rect 3270 856 3302 857
rect 1471 831 1853 839
rect 1471 812 1824 831
rect 1845 812 1853 831
rect 1471 807 1853 812
rect 4648 737 5233 745
rect 4648 717 4657 737
rect 4677 736 5233 737
rect 4677 717 5197 736
rect 4648 716 5197 717
rect 5217 716 5233 736
rect 4648 710 5233 716
rect 658 653 666 673
rect 686 653 697 673
rect 658 578 697 653
rect 881 671 937 676
rect 881 651 888 671
rect 908 651 937 671
rect 881 644 937 651
rect 5022 686 5061 690
rect 5267 689 5301 895
rect 5831 907 5865 915
rect 5831 889 5838 907
rect 5857 889 5865 907
rect 5831 882 5865 889
rect 6042 912 6098 917
rect 6042 892 6049 912
rect 6069 892 6098 912
rect 6042 885 6098 892
rect 7634 903 7668 1109
rect 7702 1082 8287 1088
rect 7702 1062 7718 1082
rect 7738 1081 8287 1082
rect 7738 1062 8258 1081
rect 7702 1061 8258 1062
rect 8278 1061 8287 1081
rect 7702 1053 8287 1061
rect 7634 895 7669 903
rect 6042 884 6077 885
rect 5835 852 5864 882
rect 7634 875 7642 895
rect 7662 875 7669 895
rect 7634 870 7669 875
rect 7634 869 7666 870
rect 5835 844 6217 852
rect 5835 825 6188 844
rect 6209 825 6217 844
rect 5835 820 6217 825
rect 5022 666 5030 686
rect 5050 666 5061 686
rect 881 643 916 644
rect 2116 596 2167 627
rect 1421 583 1460 596
rect 1421 578 1426 583
rect 658 561 1426 578
rect 1450 578 1460 583
rect 1450 561 1461 578
rect 658 553 1461 561
rect 2116 570 2133 596
rect 2161 570 2167 596
rect 660 552 946 553
rect 2116 547 2167 570
rect 2196 602 2242 633
rect 4040 631 4083 639
rect 2196 571 2210 602
rect 2238 571 2242 602
rect 2196 564 2242 571
rect 4034 624 4089 631
rect 4034 599 4047 624
rect 4079 599 4089 624
rect 498 536 559 545
rect 498 509 506 536
rect 542 530 559 536
rect 600 530 675 534
rect 542 528 675 530
rect 542 509 606 528
rect 498 492 606 509
rect 651 492 675 528
rect 498 490 675 492
rect 600 460 675 490
rect 2129 355 2160 547
rect 2115 334 2161 355
rect 2115 313 2122 334
rect 2143 313 2161 334
rect 2115 309 2161 313
rect 2115 306 2150 309
rect 1497 148 2082 156
rect 1497 128 1506 148
rect 1526 147 2082 148
rect 1526 128 2046 147
rect 1497 127 2046 128
rect 2066 127 2082 147
rect 1497 121 2082 127
rect 2116 100 2150 306
rect 2198 240 2232 564
rect 4034 507 4089 599
rect 5022 591 5061 666
rect 5245 684 5301 689
rect 5245 664 5252 684
rect 5272 664 5301 684
rect 5245 657 5301 664
rect 5245 656 5280 657
rect 6480 609 6531 640
rect 5785 596 5824 609
rect 5785 591 5790 596
rect 5022 574 5790 591
rect 5814 591 5824 596
rect 5814 574 5825 591
rect 5022 566 5825 574
rect 6480 583 6497 609
rect 6525 583 6531 609
rect 5024 565 5310 566
rect 6480 560 6531 583
rect 6560 615 6606 646
rect 8404 644 8447 652
rect 6560 584 6574 615
rect 6602 584 6606 615
rect 6560 577 6606 584
rect 8398 637 8453 644
rect 8398 612 8411 637
rect 8443 612 8453 637
rect 4034 475 4045 507
rect 4085 475 4089 507
rect 4862 549 4923 558
rect 4862 522 4870 549
rect 4906 543 4923 549
rect 4964 543 5039 547
rect 4906 541 5039 543
rect 4906 522 4970 541
rect 4862 505 4970 522
rect 5015 505 5039 541
rect 4862 503 5039 505
rect 4034 462 4089 475
rect 4964 473 5039 503
rect 6493 368 6524 560
rect 6479 347 6525 368
rect 6479 326 6486 347
rect 6507 326 6525 347
rect 6479 322 6525 326
rect 6479 319 6514 322
rect 4618 282 4649 287
rect 2198 220 2204 240
rect 2224 220 2232 240
rect 2198 214 2232 220
rect 3820 262 4654 282
rect 1877 94 1920 98
rect 1877 70 1888 94
rect 1911 70 1920 94
rect 1877 66 1920 70
rect 2094 95 2150 100
rect 2094 75 2101 95
rect 2121 75 2150 95
rect 2094 68 2150 75
rect 2094 67 2129 68
rect 1884 2 1915 66
rect 3820 2 3846 262
rect 4604 260 4650 262
rect 4604 239 4611 260
rect 4632 239 4650 260
rect 4684 252 5777 285
rect 4604 235 4650 239
rect 4604 232 4639 235
rect 3986 74 4571 82
rect 3986 54 3995 74
rect 4015 73 4571 74
rect 4015 54 4535 73
rect 3986 53 4535 54
rect 4555 53 4571 73
rect 3986 47 4571 53
rect 4605 26 4639 232
rect 4686 166 4729 252
rect 4686 146 4693 166
rect 4713 146 4729 166
rect 4686 135 4729 146
rect 4583 21 4639 26
rect 1884 -21 3847 2
rect 4583 1 4590 21
rect 4610 1 4639 21
rect 4583 -6 4639 1
rect 5746 9 5775 252
rect 5861 161 6446 169
rect 5861 141 5870 161
rect 5890 160 6446 161
rect 5890 141 6410 160
rect 5861 140 6410 141
rect 6430 140 6446 160
rect 5861 134 6446 140
rect 6243 114 6286 116
rect 6239 108 6290 114
rect 6480 113 6514 319
rect 6562 253 6596 577
rect 8398 520 8453 612
rect 8398 488 8409 520
rect 8449 488 8453 520
rect 8398 475 8453 488
rect 6562 233 6568 253
rect 6588 233 6596 253
rect 6562 227 6596 233
rect 6239 84 6255 108
rect 6278 84 6290 108
rect 6239 75 6290 84
rect 6458 108 6514 113
rect 6458 88 6465 108
rect 6485 88 6514 108
rect 6458 81 6514 88
rect 6458 80 6493 81
rect 6243 9 6286 75
rect 4583 -7 4618 -6
rect 5746 -19 6286 9
rect 5749 -21 6286 -19
rect 1892 -23 3847 -21
rect 6243 -23 6286 -21
<< via1 >>
rect 2200 5018 2227 5045
rect 2118 4199 2149 4225
rect 6564 5031 6591 5058
rect 6482 4212 6513 4238
rect 2133 570 2161 596
rect 2210 571 2238 602
rect 606 492 651 528
rect 6497 583 6525 609
rect 6574 584 6602 615
rect 4045 475 4085 507
rect 4970 505 5015 541
rect 8409 488 8449 520
<< metal2 >>
rect 6559 5058 6596 5062
rect 2195 5045 2232 5049
rect 2195 5018 2200 5045
rect 2227 5018 2232 5045
rect 6559 5031 6564 5058
rect 6591 5031 6596 5058
rect 6559 5021 6596 5031
rect 2195 5008 2232 5018
rect 2110 4225 2158 4243
rect 2110 4199 2118 4225
rect 2149 4199 2158 4225
rect 2110 4167 2158 4199
rect 2118 621 2158 4167
rect 2199 2271 2225 5008
rect 6474 4238 6522 4256
rect 6474 4212 6482 4238
rect 6513 4212 6522 4238
rect 6474 4180 6522 4212
rect 2197 633 2225 2271
rect 6482 634 6522 4180
rect 6563 2284 6589 5021
rect 6561 646 6589 2284
rect 2118 596 2164 621
rect 2118 570 2133 596
rect 2161 570 2164 596
rect 2118 551 2164 570
rect 2196 602 2242 633
rect 2196 571 2210 602
rect 2238 571 2242 602
rect 2196 564 2242 571
rect 6482 609 6528 634
rect 6482 583 6497 609
rect 6525 583 6528 609
rect 6482 564 6528 583
rect 6560 615 6606 646
rect 6560 584 6574 615
rect 6602 584 6606 615
rect 6560 577 6606 584
rect 6486 560 6528 564
rect 2122 547 2164 551
rect 4956 541 5031 553
rect 592 528 667 540
rect 592 492 606 528
rect 651 515 667 528
rect 2109 515 2203 520
rect 651 507 4089 515
rect 651 492 4045 507
rect 592 475 4045 492
rect 4085 475 4089 507
rect 4956 505 4970 541
rect 5015 528 5031 541
rect 6473 528 6567 533
rect 5015 520 8453 528
rect 5015 505 8409 520
rect 4956 488 8409 505
rect 8449 488 8453 520
rect 4956 479 8453 488
rect 6473 476 6567 479
rect 592 466 4089 475
rect 2109 463 2203 466
<< labels >>
rlabel locali 373 8244 395 8259 1 d0
rlabel locali 427 8432 456 8438 1 vdd
rlabel locali 424 8133 453 8139 1 gnd
rlabel space 530 8151 559 8160 1 gnd
rlabel nwell 562 8409 585 8412 1 vdd
rlabel locali 374 7832 396 7847 1 d0
rlabel locali 428 8020 457 8026 1 vdd
rlabel locali 425 7721 454 7727 1 gnd
rlabel space 531 7739 560 7748 1 gnd
rlabel nwell 563 7997 586 8000 1 vdd
rlabel locali 264 8677 288 8707 1 vref
rlabel locali 356 7226 378 7241 1 d0
rlabel locali 410 7414 439 7420 1 vdd
rlabel locali 407 7115 436 7121 1 gnd
rlabel space 513 7133 542 7142 1 gnd
rlabel nwell 545 7391 568 7394 1 vdd
rlabel locali 357 6814 379 6829 1 d0
rlabel locali 411 7002 440 7008 1 vdd
rlabel locali 408 6703 437 6709 1 gnd
rlabel space 514 6721 543 6730 1 gnd
rlabel nwell 546 6979 569 6982 1 vdd
rlabel locali 1225 8248 1254 8254 1 vdd
rlabel locali 1222 7949 1251 7955 1 gnd
rlabel space 1328 7967 1357 7976 1 gnd
rlabel nwell 1360 8225 1383 8228 1 vdd
rlabel locali 1165 8056 1187 8073 1 d1
rlabel locali 1208 7230 1237 7236 1 vdd
rlabel locali 1205 6931 1234 6937 1 gnd
rlabel space 1311 6949 1340 6958 1 gnd
rlabel nwell 1343 7207 1366 7210 1 vdd
rlabel locali 1148 7038 1170 7055 1 d1
rlabel locali 1307 7640 1336 7646 1 vdd
rlabel locali 1304 7341 1333 7347 1 gnd
rlabel space 1410 7359 1439 7368 1 gnd
rlabel nwell 1442 7617 1465 7620 1 vdd
rlabel locali 1249 7448 1269 7472 1 d2
rlabel locali 336 6208 358 6223 1 d0
rlabel locali 390 6396 419 6402 1 vdd
rlabel locali 387 6097 416 6103 1 gnd
rlabel space 493 6115 522 6124 1 gnd
rlabel nwell 525 6373 548 6376 1 vdd
rlabel locali 337 5796 359 5811 1 d0
rlabel locali 391 5984 420 5990 1 vdd
rlabel locali 388 5685 417 5691 1 gnd
rlabel space 494 5703 523 5712 1 gnd
rlabel nwell 526 5961 549 5964 1 vdd
rlabel locali 319 5190 341 5205 1 d0
rlabel locali 373 5378 402 5384 1 vdd
rlabel locali 370 5079 399 5085 1 gnd
rlabel space 476 5097 505 5106 1 gnd
rlabel nwell 508 5355 531 5358 1 vdd
rlabel locali 320 4778 342 4793 1 d0
rlabel locali 374 4966 403 4972 1 vdd
rlabel locali 371 4667 400 4673 1 gnd
rlabel space 477 4685 506 4694 1 gnd
rlabel nwell 509 4943 532 4946 1 vdd
rlabel locali 1188 6212 1217 6218 1 vdd
rlabel locali 1185 5913 1214 5919 1 gnd
rlabel space 1291 5931 1320 5940 1 gnd
rlabel nwell 1323 6189 1346 6192 1 vdd
rlabel locali 1128 6020 1150 6037 1 d1
rlabel locali 1171 5194 1200 5200 1 vdd
rlabel locali 1168 4895 1197 4901 1 gnd
rlabel space 1274 4913 1303 4922 1 gnd
rlabel nwell 1306 5171 1329 5174 1 vdd
rlabel locali 1111 5002 1133 5019 1 d1
rlabel locali 1270 5604 1299 5610 1 vdd
rlabel locali 1267 5305 1296 5311 1 gnd
rlabel space 1373 5323 1402 5332 1 gnd
rlabel nwell 1405 5581 1428 5584 1 vdd
rlabel locali 1212 5412 1232 5436 1 d2
rlabel locali 1353 6620 1382 6626 1 vdd
rlabel locali 1350 6321 1379 6327 1 gnd
rlabel space 1456 6339 1485 6348 1 gnd
rlabel nwell 1488 6597 1511 6600 1 vdd
rlabel locali 1297 6434 1317 6447 1 d3
rlabel locali 300 4172 322 4187 1 d0
rlabel locali 354 4360 383 4366 1 vdd
rlabel locali 351 4061 380 4067 1 gnd
rlabel space 457 4079 486 4088 1 gnd
rlabel nwell 489 4337 512 4340 1 vdd
rlabel locali 301 3760 323 3775 1 d0
rlabel locali 355 3948 384 3954 1 vdd
rlabel locali 352 3649 381 3655 1 gnd
rlabel space 458 3667 487 3676 1 gnd
rlabel nwell 490 3925 513 3928 1 vdd
rlabel locali 283 3154 305 3169 1 d0
rlabel locali 337 3342 366 3348 1 vdd
rlabel locali 334 3043 363 3049 1 gnd
rlabel space 440 3061 469 3070 1 gnd
rlabel nwell 472 3319 495 3322 1 vdd
rlabel locali 284 2742 306 2757 1 d0
rlabel locali 338 2930 367 2936 1 vdd
rlabel locali 335 2631 364 2637 1 gnd
rlabel space 441 2649 470 2658 1 gnd
rlabel nwell 473 2907 496 2910 1 vdd
rlabel locali 1152 4176 1181 4182 1 vdd
rlabel locali 1149 3877 1178 3883 1 gnd
rlabel space 1255 3895 1284 3904 1 gnd
rlabel nwell 1287 4153 1310 4156 1 vdd
rlabel locali 1092 3984 1114 4001 1 d1
rlabel locali 1135 3158 1164 3164 1 vdd
rlabel locali 1132 2859 1161 2865 1 gnd
rlabel space 1238 2877 1267 2886 1 gnd
rlabel nwell 1270 3135 1293 3138 1 vdd
rlabel locali 1075 2966 1097 2983 1 d1
rlabel locali 1234 3568 1263 3574 1 vdd
rlabel locali 1231 3269 1260 3275 1 gnd
rlabel space 1337 3287 1366 3296 1 gnd
rlabel nwell 1369 3545 1392 3548 1 vdd
rlabel locali 1176 3376 1196 3400 1 d2
rlabel locali 263 2136 285 2151 1 d0
rlabel locali 317 2324 346 2330 1 vdd
rlabel locali 314 2025 343 2031 1 gnd
rlabel space 420 2043 449 2052 1 gnd
rlabel nwell 452 2301 475 2304 1 vdd
rlabel locali 264 1724 286 1739 1 d0
rlabel locali 318 1912 347 1918 1 vdd
rlabel locali 315 1613 344 1619 1 gnd
rlabel space 421 1631 450 1640 1 gnd
rlabel nwell 453 1889 476 1892 1 vdd
rlabel locali 246 1118 268 1133 1 d0
rlabel locali 300 1306 329 1312 1 vdd
rlabel locali 297 1007 326 1013 1 gnd
rlabel space 403 1025 432 1034 1 gnd
rlabel nwell 435 1283 458 1286 1 vdd
rlabel locali 247 706 269 721 1 d0
rlabel locali 301 894 330 900 1 vdd
rlabel locali 298 595 327 601 1 gnd
rlabel space 404 613 433 622 1 gnd
rlabel nwell 436 871 459 874 1 vdd
rlabel locali 1115 2140 1144 2146 1 vdd
rlabel locali 1112 1841 1141 1847 1 gnd
rlabel space 1218 1859 1247 1868 1 gnd
rlabel nwell 1250 2117 1273 2120 1 vdd
rlabel locali 1055 1948 1077 1965 1 d1
rlabel locali 1098 1122 1127 1128 1 vdd
rlabel locali 1095 823 1124 829 1 gnd
rlabel space 1201 841 1230 850 1 gnd
rlabel nwell 1233 1099 1256 1102 1 vdd
rlabel locali 1038 930 1060 947 1 d1
rlabel locali 1197 1532 1226 1538 1 vdd
rlabel locali 1194 1233 1223 1239 1 gnd
rlabel space 1300 1251 1329 1260 1 gnd
rlabel nwell 1332 1509 1355 1512 1 vdd
rlabel locali 1139 1340 1159 1364 1 d2
rlabel locali 1280 2548 1309 2554 1 vdd
rlabel locali 1277 2249 1306 2255 1 gnd
rlabel space 1383 2267 1412 2276 1 gnd
rlabel nwell 1415 2525 1438 2528 1 vdd
rlabel locali 1224 2362 1244 2375 1 d3
rlabel locali 1456 4582 1485 4588 1 vdd
rlabel locali 1453 4283 1482 4289 1 gnd
rlabel space 1559 4301 1588 4310 1 gnd
rlabel nwell 1591 4559 1614 4562 1 vdd
rlabel locali 1402 4392 1421 4409 1 d4
rlabel locali 2912 4901 2931 4918 5 d4
rlabel nwell 2719 4748 2742 4751 5 vdd
rlabel space 2745 5000 2774 5009 5 gnd
rlabel locali 2851 5021 2880 5027 5 gnd
rlabel locali 2848 4722 2877 4728 5 vdd
rlabel locali 3089 6935 3109 6948 5 d3
rlabel nwell 2895 6782 2918 6785 5 vdd
rlabel space 2921 7034 2950 7043 5 gnd
rlabel locali 3027 7055 3056 7061 5 gnd
rlabel locali 3024 6756 3053 6762 5 vdd
rlabel locali 3174 7946 3194 7970 5 d2
rlabel nwell 2978 7798 3001 7801 5 vdd
rlabel space 3004 8050 3033 8059 5 gnd
rlabel locali 3110 8071 3139 8077 5 gnd
rlabel locali 3107 7772 3136 7778 5 vdd
rlabel locali 3273 8363 3295 8380 5 d1
rlabel nwell 3077 8208 3100 8211 5 vdd
rlabel space 3103 8460 3132 8469 5 gnd
rlabel locali 3209 8481 3238 8487 5 gnd
rlabel locali 3206 8182 3235 8188 5 vdd
rlabel locali 3256 7345 3278 7362 5 d1
rlabel nwell 3060 7190 3083 7193 5 vdd
rlabel space 3086 7442 3115 7451 5 gnd
rlabel locali 3192 7463 3221 7469 5 gnd
rlabel locali 3189 7164 3218 7170 5 vdd
rlabel nwell 3874 8436 3897 8439 5 vdd
rlabel space 3900 8688 3929 8697 5 gnd
rlabel locali 4006 8709 4035 8715 5 gnd
rlabel locali 4003 8410 4032 8416 5 vdd
rlabel locali 4064 8589 4086 8604 5 d0
rlabel nwell 3875 8024 3898 8027 5 vdd
rlabel space 3901 8276 3930 8285 5 gnd
rlabel locali 4007 8297 4036 8303 5 gnd
rlabel locali 4004 7998 4033 8004 5 vdd
rlabel locali 4065 8177 4087 8192 5 d0
rlabel nwell 3857 7418 3880 7421 5 vdd
rlabel space 3883 7670 3912 7679 5 gnd
rlabel locali 3989 7691 4018 7697 5 gnd
rlabel locali 3986 7392 4015 7398 5 vdd
rlabel locali 4047 7571 4069 7586 5 d0
rlabel nwell 3858 7006 3881 7009 5 vdd
rlabel space 3884 7258 3913 7267 5 gnd
rlabel locali 3990 7279 4019 7285 5 gnd
rlabel locali 3987 6980 4016 6986 5 vdd
rlabel locali 4048 7159 4070 7174 5 d0
rlabel locali 3137 5910 3157 5934 5 d2
rlabel nwell 2941 5762 2964 5765 5 vdd
rlabel space 2967 6014 2996 6023 5 gnd
rlabel locali 3073 6035 3102 6041 5 gnd
rlabel locali 3070 5736 3099 5742 5 vdd
rlabel locali 3236 6327 3258 6344 5 d1
rlabel nwell 3040 6172 3063 6175 5 vdd
rlabel space 3066 6424 3095 6433 5 gnd
rlabel locali 3172 6445 3201 6451 5 gnd
rlabel locali 3169 6146 3198 6152 5 vdd
rlabel locali 3219 5309 3241 5326 5 d1
rlabel nwell 3023 5154 3046 5157 5 vdd
rlabel space 3049 5406 3078 5415 5 gnd
rlabel locali 3155 5427 3184 5433 5 gnd
rlabel locali 3152 5128 3181 5134 5 vdd
rlabel nwell 3837 6400 3860 6403 5 vdd
rlabel space 3863 6652 3892 6661 5 gnd
rlabel locali 3969 6673 3998 6679 5 gnd
rlabel locali 3966 6374 3995 6380 5 vdd
rlabel locali 4027 6553 4049 6568 5 d0
rlabel nwell 3838 5988 3861 5991 5 vdd
rlabel space 3864 6240 3893 6249 5 gnd
rlabel locali 3970 6261 3999 6267 5 gnd
rlabel locali 3967 5962 3996 5968 5 vdd
rlabel locali 4028 6141 4050 6156 5 d0
rlabel nwell 3820 5382 3843 5385 5 vdd
rlabel space 3846 5634 3875 5643 5 gnd
rlabel locali 3952 5655 3981 5661 5 gnd
rlabel locali 3949 5356 3978 5362 5 vdd
rlabel locali 4010 5535 4032 5550 5 d0
rlabel nwell 3821 4970 3844 4973 5 vdd
rlabel space 3847 5222 3876 5231 5 gnd
rlabel locali 3953 5243 3982 5249 5 gnd
rlabel locali 3950 4944 3979 4950 5 vdd
rlabel locali 4011 5123 4033 5138 5 d0
rlabel locali 3016 2863 3036 2876 5 d3
rlabel nwell 2822 2710 2845 2713 5 vdd
rlabel space 2848 2962 2877 2971 5 gnd
rlabel locali 2954 2983 2983 2989 5 gnd
rlabel locali 2951 2684 2980 2690 5 vdd
rlabel locali 3101 3874 3121 3898 5 d2
rlabel nwell 2905 3726 2928 3729 5 vdd
rlabel space 2931 3978 2960 3987 5 gnd
rlabel locali 3037 3999 3066 4005 5 gnd
rlabel locali 3034 3700 3063 3706 5 vdd
rlabel locali 3200 4291 3222 4308 5 d1
rlabel nwell 3004 4136 3027 4139 5 vdd
rlabel space 3030 4388 3059 4397 5 gnd
rlabel locali 3136 4409 3165 4415 5 gnd
rlabel locali 3133 4110 3162 4116 5 vdd
rlabel locali 3183 3273 3205 3290 5 d1
rlabel nwell 2987 3118 3010 3121 5 vdd
rlabel space 3013 3370 3042 3379 5 gnd
rlabel locali 3119 3391 3148 3397 5 gnd
rlabel locali 3116 3092 3145 3098 5 vdd
rlabel nwell 3801 4364 3824 4367 5 vdd
rlabel space 3827 4616 3856 4625 5 gnd
rlabel locali 3933 4637 3962 4643 5 gnd
rlabel locali 3930 4338 3959 4344 5 vdd
rlabel locali 3991 4517 4013 4532 5 d0
rlabel nwell 3802 3952 3825 3955 5 vdd
rlabel space 3828 4204 3857 4213 5 gnd
rlabel locali 3934 4225 3963 4231 5 gnd
rlabel locali 3931 3926 3960 3932 5 vdd
rlabel locali 3992 4105 4014 4120 5 d0
rlabel nwell 3784 3346 3807 3349 5 vdd
rlabel space 3810 3598 3839 3607 5 gnd
rlabel locali 3916 3619 3945 3625 5 gnd
rlabel locali 3913 3320 3942 3326 5 vdd
rlabel locali 3974 3499 3996 3514 5 d0
rlabel nwell 3785 2934 3808 2937 5 vdd
rlabel space 3811 3186 3840 3195 5 gnd
rlabel locali 3917 3207 3946 3213 5 gnd
rlabel locali 3914 2908 3943 2914 5 vdd
rlabel locali 3975 3087 3997 3102 5 d0
rlabel locali 3064 1838 3084 1862 5 d2
rlabel nwell 2868 1690 2891 1693 5 vdd
rlabel space 2894 1942 2923 1951 5 gnd
rlabel locali 3000 1963 3029 1969 5 gnd
rlabel locali 2997 1664 3026 1670 5 vdd
rlabel locali 3163 2255 3185 2272 5 d1
rlabel nwell 2967 2100 2990 2103 5 vdd
rlabel space 2993 2352 3022 2361 5 gnd
rlabel locali 3099 2373 3128 2379 5 gnd
rlabel locali 3096 2074 3125 2080 5 vdd
rlabel locali 3146 1237 3168 1254 5 d1
rlabel nwell 2950 1082 2973 1085 5 vdd
rlabel space 2976 1334 3005 1343 5 gnd
rlabel locali 3082 1355 3111 1361 5 gnd
rlabel locali 3079 1056 3108 1062 5 vdd
rlabel nwell 3764 2328 3787 2331 5 vdd
rlabel space 3790 2580 3819 2589 5 gnd
rlabel locali 3896 2601 3925 2607 5 gnd
rlabel locali 3893 2302 3922 2308 5 vdd
rlabel locali 3954 2481 3976 2496 5 d0
rlabel nwell 3765 1916 3788 1919 5 vdd
rlabel space 3791 2168 3820 2177 5 gnd
rlabel locali 3897 2189 3926 2195 5 gnd
rlabel locali 3894 1890 3923 1896 5 vdd
rlabel locali 3955 2069 3977 2084 5 d0
rlabel nwell 3747 1310 3770 1313 5 vdd
rlabel space 3773 1562 3802 1571 5 gnd
rlabel locali 3879 1583 3908 1589 5 gnd
rlabel locali 3876 1284 3905 1290 5 vdd
rlabel locali 3937 1463 3959 1478 5 d0
rlabel nwell 3748 898 3771 901 5 vdd
rlabel space 3774 1150 3803 1159 5 gnd
rlabel locali 3880 1171 3909 1177 5 gnd
rlabel locali 3877 872 3906 878 5 vdd
rlabel locali 3938 1051 3960 1066 5 d0
rlabel nwell 1649 295 1672 298 1 vdd
rlabel space 1617 37 1646 46 1 gnd
rlabel locali 1511 19 1540 25 1 gnd
rlabel locali 1514 318 1543 324 1 vdd
rlabel locali 1456 131 1471 144 1 d5
rlabel locali 4737 8257 4759 8272 1 d0
rlabel locali 4791 8445 4820 8451 1 vdd
rlabel locali 4788 8146 4817 8152 1 gnd
rlabel space 4894 8164 4923 8173 1 gnd
rlabel nwell 4926 8422 4949 8425 1 vdd
rlabel locali 4738 7845 4760 7860 1 d0
rlabel locali 4792 8033 4821 8039 1 vdd
rlabel locali 4789 7734 4818 7740 1 gnd
rlabel space 4895 7752 4924 7761 1 gnd
rlabel nwell 4927 8010 4950 8013 1 vdd
rlabel locali 4720 7239 4742 7254 1 d0
rlabel locali 4774 7427 4803 7433 1 vdd
rlabel locali 4771 7128 4800 7134 1 gnd
rlabel space 4877 7146 4906 7155 1 gnd
rlabel nwell 4909 7404 4932 7407 1 vdd
rlabel locali 4721 6827 4743 6842 1 d0
rlabel locali 4775 7015 4804 7021 1 vdd
rlabel locali 4772 6716 4801 6722 1 gnd
rlabel space 4878 6734 4907 6743 1 gnd
rlabel nwell 4910 6992 4933 6995 1 vdd
rlabel locali 5589 8261 5618 8267 1 vdd
rlabel locali 5586 7962 5615 7968 1 gnd
rlabel space 5692 7980 5721 7989 1 gnd
rlabel nwell 5724 8238 5747 8241 1 vdd
rlabel locali 5529 8069 5551 8086 1 d1
rlabel locali 5572 7243 5601 7249 1 vdd
rlabel locali 5569 6944 5598 6950 1 gnd
rlabel space 5675 6962 5704 6971 1 gnd
rlabel nwell 5707 7220 5730 7223 1 vdd
rlabel locali 5512 7051 5534 7068 1 d1
rlabel locali 5671 7653 5700 7659 1 vdd
rlabel locali 5668 7354 5697 7360 1 gnd
rlabel space 5774 7372 5803 7381 1 gnd
rlabel nwell 5806 7630 5829 7633 1 vdd
rlabel locali 5613 7461 5633 7485 1 d2
rlabel locali 4700 6221 4722 6236 1 d0
rlabel locali 4754 6409 4783 6415 1 vdd
rlabel locali 4751 6110 4780 6116 1 gnd
rlabel space 4857 6128 4886 6137 1 gnd
rlabel nwell 4889 6386 4912 6389 1 vdd
rlabel locali 4701 5809 4723 5824 1 d0
rlabel locali 4755 5997 4784 6003 1 vdd
rlabel locali 4752 5698 4781 5704 1 gnd
rlabel space 4858 5716 4887 5725 1 gnd
rlabel nwell 4890 5974 4913 5977 1 vdd
rlabel locali 4683 5203 4705 5218 1 d0
rlabel locali 4737 5391 4766 5397 1 vdd
rlabel locali 4734 5092 4763 5098 1 gnd
rlabel space 4840 5110 4869 5119 1 gnd
rlabel nwell 4872 5368 4895 5371 1 vdd
rlabel locali 4684 4791 4706 4806 1 d0
rlabel locali 4738 4979 4767 4985 1 vdd
rlabel locali 4735 4680 4764 4686 1 gnd
rlabel space 4841 4698 4870 4707 1 gnd
rlabel nwell 4873 4956 4896 4959 1 vdd
rlabel locali 5552 6225 5581 6231 1 vdd
rlabel locali 5549 5926 5578 5932 1 gnd
rlabel space 5655 5944 5684 5953 1 gnd
rlabel nwell 5687 6202 5710 6205 1 vdd
rlabel locali 5492 6033 5514 6050 1 d1
rlabel locali 5535 5207 5564 5213 1 vdd
rlabel locali 5532 4908 5561 4914 1 gnd
rlabel space 5638 4926 5667 4935 1 gnd
rlabel nwell 5670 5184 5693 5187 1 vdd
rlabel locali 5475 5015 5497 5032 1 d1
rlabel locali 5634 5617 5663 5623 1 vdd
rlabel locali 5631 5318 5660 5324 1 gnd
rlabel space 5737 5336 5766 5345 1 gnd
rlabel nwell 5769 5594 5792 5597 1 vdd
rlabel locali 5576 5425 5596 5449 1 d2
rlabel locali 5717 6633 5746 6639 1 vdd
rlabel locali 5714 6334 5743 6340 1 gnd
rlabel space 5820 6352 5849 6361 1 gnd
rlabel nwell 5852 6610 5875 6613 1 vdd
rlabel locali 5661 6447 5681 6460 1 d3
rlabel locali 4664 4185 4686 4200 1 d0
rlabel locali 4718 4373 4747 4379 1 vdd
rlabel locali 4715 4074 4744 4080 1 gnd
rlabel space 4821 4092 4850 4101 1 gnd
rlabel nwell 4853 4350 4876 4353 1 vdd
rlabel locali 4665 3773 4687 3788 1 d0
rlabel locali 4719 3961 4748 3967 1 vdd
rlabel locali 4716 3662 4745 3668 1 gnd
rlabel space 4822 3680 4851 3689 1 gnd
rlabel nwell 4854 3938 4877 3941 1 vdd
rlabel locali 4647 3167 4669 3182 1 d0
rlabel locali 4701 3355 4730 3361 1 vdd
rlabel locali 4698 3056 4727 3062 1 gnd
rlabel space 4804 3074 4833 3083 1 gnd
rlabel nwell 4836 3332 4859 3335 1 vdd
rlabel locali 4648 2755 4670 2770 1 d0
rlabel locali 4702 2943 4731 2949 1 vdd
rlabel locali 4699 2644 4728 2650 1 gnd
rlabel space 4805 2662 4834 2671 1 gnd
rlabel nwell 4837 2920 4860 2923 1 vdd
rlabel locali 5516 4189 5545 4195 1 vdd
rlabel locali 5513 3890 5542 3896 1 gnd
rlabel space 5619 3908 5648 3917 1 gnd
rlabel nwell 5651 4166 5674 4169 1 vdd
rlabel locali 5456 3997 5478 4014 1 d1
rlabel locali 5499 3171 5528 3177 1 vdd
rlabel locali 5496 2872 5525 2878 1 gnd
rlabel space 5602 2890 5631 2899 1 gnd
rlabel nwell 5634 3148 5657 3151 1 vdd
rlabel locali 5439 2979 5461 2996 1 d1
rlabel locali 5598 3581 5627 3587 1 vdd
rlabel locali 5595 3282 5624 3288 1 gnd
rlabel space 5701 3300 5730 3309 1 gnd
rlabel nwell 5733 3558 5756 3561 1 vdd
rlabel locali 5540 3389 5560 3413 1 d2
rlabel locali 4627 2149 4649 2164 1 d0
rlabel locali 4681 2337 4710 2343 1 vdd
rlabel locali 4678 2038 4707 2044 1 gnd
rlabel space 4784 2056 4813 2065 1 gnd
rlabel nwell 4816 2314 4839 2317 1 vdd
rlabel locali 4628 1737 4650 1752 1 d0
rlabel locali 4682 1925 4711 1931 1 vdd
rlabel locali 4679 1626 4708 1632 1 gnd
rlabel space 4785 1644 4814 1653 1 gnd
rlabel nwell 4817 1902 4840 1905 1 vdd
rlabel locali 4610 1131 4632 1146 1 d0
rlabel locali 4664 1319 4693 1325 1 vdd
rlabel locali 4661 1020 4690 1026 1 gnd
rlabel space 4767 1038 4796 1047 1 gnd
rlabel nwell 4799 1296 4822 1299 1 vdd
rlabel locali 4611 719 4633 734 1 d0
rlabel locali 4665 907 4694 913 1 vdd
rlabel locali 4662 608 4691 614 1 gnd
rlabel space 4768 626 4797 635 1 gnd
rlabel nwell 4800 884 4823 887 1 vdd
rlabel locali 5479 2153 5508 2159 1 vdd
rlabel locali 5476 1854 5505 1860 1 gnd
rlabel space 5582 1872 5611 1881 1 gnd
rlabel nwell 5614 2130 5637 2133 1 vdd
rlabel locali 5419 1961 5441 1978 1 d1
rlabel locali 5462 1135 5491 1141 1 vdd
rlabel locali 5459 836 5488 842 1 gnd
rlabel space 5565 854 5594 863 1 gnd
rlabel nwell 5597 1112 5620 1115 1 vdd
rlabel locali 5402 943 5424 960 1 d1
rlabel locali 5561 1545 5590 1551 1 vdd
rlabel locali 5558 1246 5587 1252 1 gnd
rlabel space 5664 1264 5693 1273 1 gnd
rlabel nwell 5696 1522 5719 1525 1 vdd
rlabel locali 5503 1353 5523 1377 1 d2
rlabel locali 5644 2561 5673 2567 1 vdd
rlabel locali 5641 2262 5670 2268 1 gnd
rlabel space 5747 2280 5776 2289 1 gnd
rlabel nwell 5779 2538 5802 2541 1 vdd
rlabel locali 5588 2375 5608 2388 1 d3
rlabel locali 5820 4595 5849 4601 1 vdd
rlabel locali 5817 4296 5846 4302 1 gnd
rlabel space 5923 4314 5952 4323 1 gnd
rlabel nwell 5955 4572 5978 4575 1 vdd
rlabel locali 5766 4405 5785 4422 1 d4
rlabel locali 7276 4914 7295 4931 5 d4
rlabel nwell 7083 4761 7106 4764 5 vdd
rlabel space 7109 5013 7138 5022 5 gnd
rlabel locali 7215 5034 7244 5040 5 gnd
rlabel locali 7212 4735 7241 4741 5 vdd
rlabel locali 7453 6948 7473 6961 5 d3
rlabel nwell 7259 6795 7282 6798 5 vdd
rlabel space 7285 7047 7314 7056 5 gnd
rlabel locali 7391 7068 7420 7074 5 gnd
rlabel locali 7388 6769 7417 6775 5 vdd
rlabel locali 7538 7959 7558 7983 5 d2
rlabel nwell 7342 7811 7365 7814 5 vdd
rlabel space 7368 8063 7397 8072 5 gnd
rlabel locali 7474 8084 7503 8090 5 gnd
rlabel locali 7471 7785 7500 7791 5 vdd
rlabel locali 7637 8376 7659 8393 5 d1
rlabel nwell 7441 8221 7464 8224 5 vdd
rlabel space 7467 8473 7496 8482 5 gnd
rlabel locali 7573 8494 7602 8500 5 gnd
rlabel locali 7570 8195 7599 8201 5 vdd
rlabel locali 7620 7358 7642 7375 5 d1
rlabel nwell 7424 7203 7447 7206 5 vdd
rlabel space 7450 7455 7479 7464 5 gnd
rlabel locali 7556 7476 7585 7482 5 gnd
rlabel locali 7553 7177 7582 7183 5 vdd
rlabel locali 8556 8711 8584 8729 5 gnd
rlabel nwell 8238 8449 8261 8452 5 vdd
rlabel space 8264 8701 8293 8710 5 gnd
rlabel locali 8370 8722 8399 8728 5 gnd
rlabel locali 8367 8423 8396 8429 5 vdd
rlabel locali 8428 8602 8450 8617 5 d0
rlabel nwell 8239 8037 8262 8040 5 vdd
rlabel space 8265 8289 8294 8298 5 gnd
rlabel locali 8371 8310 8400 8316 5 gnd
rlabel locali 8368 8011 8397 8017 5 vdd
rlabel locali 8429 8190 8451 8205 5 d0
rlabel nwell 8221 7431 8244 7434 5 vdd
rlabel space 8247 7683 8276 7692 5 gnd
rlabel locali 8353 7704 8382 7710 5 gnd
rlabel locali 8350 7405 8379 7411 5 vdd
rlabel locali 8411 7584 8433 7599 5 d0
rlabel nwell 8222 7019 8245 7022 5 vdd
rlabel space 8248 7271 8277 7280 5 gnd
rlabel locali 8354 7292 8383 7298 5 gnd
rlabel locali 8351 6993 8380 6999 5 vdd
rlabel locali 8412 7172 8434 7187 5 d0
rlabel locali 7501 5923 7521 5947 5 d2
rlabel nwell 7305 5775 7328 5778 5 vdd
rlabel space 7331 6027 7360 6036 5 gnd
rlabel locali 7437 6048 7466 6054 5 gnd
rlabel locali 7434 5749 7463 5755 5 vdd
rlabel locali 7600 6340 7622 6357 5 d1
rlabel nwell 7404 6185 7427 6188 5 vdd
rlabel space 7430 6437 7459 6446 5 gnd
rlabel locali 7536 6458 7565 6464 5 gnd
rlabel locali 7533 6159 7562 6165 5 vdd
rlabel locali 7583 5322 7605 5339 5 d1
rlabel nwell 7387 5167 7410 5170 5 vdd
rlabel space 7413 5419 7442 5428 5 gnd
rlabel locali 7519 5440 7548 5446 5 gnd
rlabel locali 7516 5141 7545 5147 5 vdd
rlabel nwell 8201 6413 8224 6416 5 vdd
rlabel space 8227 6665 8256 6674 5 gnd
rlabel locali 8333 6686 8362 6692 5 gnd
rlabel locali 8330 6387 8359 6393 5 vdd
rlabel locali 8391 6566 8413 6581 5 d0
rlabel nwell 8202 6001 8225 6004 5 vdd
rlabel space 8228 6253 8257 6262 5 gnd
rlabel locali 8334 6274 8363 6280 5 gnd
rlabel locali 8331 5975 8360 5981 5 vdd
rlabel locali 8392 6154 8414 6169 5 d0
rlabel nwell 8184 5395 8207 5398 5 vdd
rlabel space 8210 5647 8239 5656 5 gnd
rlabel locali 8316 5668 8345 5674 5 gnd
rlabel locali 8313 5369 8342 5375 5 vdd
rlabel locali 8374 5548 8396 5563 5 d0
rlabel nwell 8185 4983 8208 4986 5 vdd
rlabel space 8211 5235 8240 5244 5 gnd
rlabel locali 8317 5256 8346 5262 5 gnd
rlabel locali 8314 4957 8343 4963 5 vdd
rlabel locali 8375 5136 8397 5151 5 d0
rlabel locali 7380 2876 7400 2889 5 d3
rlabel nwell 7186 2723 7209 2726 5 vdd
rlabel space 7212 2975 7241 2984 5 gnd
rlabel locali 7318 2996 7347 3002 5 gnd
rlabel locali 7315 2697 7344 2703 5 vdd
rlabel locali 7465 3887 7485 3911 5 d2
rlabel nwell 7269 3739 7292 3742 5 vdd
rlabel space 7295 3991 7324 4000 5 gnd
rlabel locali 7401 4012 7430 4018 5 gnd
rlabel locali 7398 3713 7427 3719 5 vdd
rlabel locali 7564 4304 7586 4321 5 d1
rlabel nwell 7368 4149 7391 4152 5 vdd
rlabel space 7394 4401 7423 4410 5 gnd
rlabel locali 7500 4422 7529 4428 5 gnd
rlabel locali 7497 4123 7526 4129 5 vdd
rlabel locali 7547 3286 7569 3303 5 d1
rlabel nwell 7351 3131 7374 3134 5 vdd
rlabel space 7377 3383 7406 3392 5 gnd
rlabel locali 7483 3404 7512 3410 5 gnd
rlabel locali 7480 3105 7509 3111 5 vdd
rlabel nwell 8165 4377 8188 4380 5 vdd
rlabel space 8191 4629 8220 4638 5 gnd
rlabel locali 8297 4650 8326 4656 5 gnd
rlabel locali 8294 4351 8323 4357 5 vdd
rlabel locali 8355 4530 8377 4545 5 d0
rlabel nwell 8166 3965 8189 3968 5 vdd
rlabel space 8192 4217 8221 4226 5 gnd
rlabel locali 8298 4238 8327 4244 5 gnd
rlabel locali 8295 3939 8324 3945 5 vdd
rlabel locali 8356 4118 8378 4133 5 d0
rlabel nwell 8148 3359 8171 3362 5 vdd
rlabel space 8174 3611 8203 3620 5 gnd
rlabel locali 8280 3632 8309 3638 5 gnd
rlabel locali 8277 3333 8306 3339 5 vdd
rlabel locali 8338 3512 8360 3527 5 d0
rlabel nwell 8149 2947 8172 2950 5 vdd
rlabel space 8175 3199 8204 3208 5 gnd
rlabel locali 8281 3220 8310 3226 5 gnd
rlabel locali 8278 2921 8307 2927 5 vdd
rlabel locali 8339 3100 8361 3115 5 d0
rlabel locali 7428 1851 7448 1875 5 d2
rlabel nwell 7232 1703 7255 1706 5 vdd
rlabel space 7258 1955 7287 1964 5 gnd
rlabel locali 7364 1976 7393 1982 5 gnd
rlabel locali 7361 1677 7390 1683 5 vdd
rlabel locali 7527 2268 7549 2285 5 d1
rlabel nwell 7331 2113 7354 2116 5 vdd
rlabel space 7357 2365 7386 2374 5 gnd
rlabel locali 7463 2386 7492 2392 5 gnd
rlabel locali 7460 2087 7489 2093 5 vdd
rlabel locali 7510 1250 7532 1267 5 d1
rlabel nwell 7314 1095 7337 1098 5 vdd
rlabel space 7340 1347 7369 1356 5 gnd
rlabel locali 7446 1368 7475 1374 5 gnd
rlabel locali 7443 1069 7472 1075 5 vdd
rlabel nwell 8128 2341 8151 2344 5 vdd
rlabel space 8154 2593 8183 2602 5 gnd
rlabel locali 8260 2614 8289 2620 5 gnd
rlabel locali 8257 2315 8286 2321 5 vdd
rlabel locali 8318 2494 8340 2509 5 d0
rlabel nwell 8129 1929 8152 1932 5 vdd
rlabel space 8155 2181 8184 2190 5 gnd
rlabel locali 8261 2202 8290 2208 5 gnd
rlabel locali 8258 1903 8287 1909 5 vdd
rlabel locali 8319 2082 8341 2097 5 d0
rlabel nwell 8111 1323 8134 1326 5 vdd
rlabel space 8137 1575 8166 1584 5 gnd
rlabel locali 8243 1596 8272 1602 5 gnd
rlabel locali 8240 1297 8269 1303 5 vdd
rlabel locali 8301 1476 8323 1491 5 d0
rlabel nwell 8112 911 8135 914 5 vdd
rlabel space 8138 1163 8167 1172 5 gnd
rlabel locali 8244 1184 8273 1190 5 gnd
rlabel locali 8241 885 8270 891 5 vdd
rlabel locali 8302 1064 8324 1079 5 d0
rlabel nwell 6013 308 6036 311 1 vdd
rlabel space 5981 50 6010 59 1 gnd
rlabel locali 5875 32 5904 38 1 gnd
rlabel locali 5878 331 5907 337 1 vdd
rlabel locali 5820 144 5835 157 1 d5
rlabel locali 4376 91 4398 106 1 vout
rlabel nwell 4138 221 4161 224 1 vdd
rlabel space 4106 -37 4135 -28 1 gnd
rlabel locali 4000 -55 4029 -49 1 gnd
rlabel locali 4003 244 4032 250 1 vdd
rlabel locali 3939 54 3962 70 1 d6
<< end >>

* SPICE3 file created from 10bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_10002_n7915# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1 a_26555_3913# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_14463_5570# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3 a_5497_n9531# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_30648_4032# d0 a_31137_3926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5 a_9220_5937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6 a_3180_n3469# a_3437_n3485# a_2382_n3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7 vdd d0 a_21008_3144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8 a_4769_2265# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9 vdd d2 a_11534_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 vdd d0 a_34185_7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X11 a_30704_7086# d0 a_31193_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X12 a_9202_5331# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X13 a_23057_3521# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X14 a_9402_3901# a_9184_3901# a_8913_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X15 a_11998_n7378# a_12251_n7582# a_11196_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X16 vdd d3 a_11308_n8376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X17 gnd d3 a_28679_n8388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X18 a_28531_n5726# a_28788_n5742# a_28436_n5128# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X19 gnd d0 a_16722_2152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X20 vdd d4 a_33047_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X21 a_6986_5378# d0 a_7783_5606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X22 a_30711_7304# d0 a_31192_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X23 a_31119_3320# d1 a_31917_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X24 a_1514_7158# d2 a_1565_6667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X25 a_16358_n7579# a_16362_n7391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X26 a_29401_n10026# a_26195_n9957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X27 a_26284_4019# a_26291_4237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X28 a_33062_3379# d0 a_33859_3607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X29 a_4790_n2589# d1 a_5588_n2638# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_13095_n5062# d0 a_13586_n5256# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X31 a_2545_1470# d0 a_3347_1109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X32 a_12101_2329# a_12358_2139# a_11303_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X33 a_2438_n6707# d0 a_3236_n6523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X34 a_17496_1158# d0 a_17977_1246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X35 gnd d3 a_15599_n4317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X36 a_32796_n5329# a_33053_n5345# a_32717_n4125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X37 gnd d0 a_29712_1133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X38 a_19838_1913# a_20091_1900# a_19788_3110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X39 gnd d0 a_29784_5617# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X40 a_17597_6755# a_17599_7048# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X41 a_17449_n9608# a_17454_n9932# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X42 a_4609_8067# a_4616_8285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X43 a_4987_2265# a_4769_2265# a_4512_2360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X44 a_3253_n7541# a_3257_n7353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X45 a_11327_3354# a_11580_3341# a_11241_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X46 a_10182_6573# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X47 a_17870_n6660# a_17652_n6660# a_17395_n6554# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X48 a_1482_5651# a_1276_6140# a_696_6324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X49 a_14551_3653# a_14345_4142# a_13765_4326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X50 a_31013_n8322# d1 a_31810_n8783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X51 a_4828_n4213# a_4610_n4213# a_4339_n4118# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X52 a_2138_n6113# d3 a_2314_n8147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X53 a_12174_6401# a_12431_6211# a_11376_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X54 a_26358_n4237# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X55 vdd d0 a_29728_2563# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X56 a_4988_1853# d1 a_5773_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X57 a_28399_n3092# a_28652_n3296# a_28349_n4300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X58 gnd d1 a_20103_n8771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X59 a_10875_n6326# d3 a_10978_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X60 a_11158_3123# d2 a_11204_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X61 a_26087_n4142# d0 a_26576_n4237# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X62 a_26538_n2613# a_26320_n2613# a_26063_n2507# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X63 a_3379_3734# a_3636_3544# a_2586_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X64 a_4864_n6249# d1 a_5661_n6710# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X65 a_3456_7629# a_3470_8412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X66 a_28784_8633# d0 a_29586_8272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X67 a_6023_6561# a_5805_6561# a_5924_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X68 a_27553_3123# a_27335_3123# a_26755_3307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X69 a_26065_n3025# d0 a_26556_n3219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X70 a_28657_1507# a_28914_1317# a_28575_2115# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X71 a_30487_n6191# d0 a_30976_n6286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 a_20554_n3705# a_20571_n4499# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X73 a_33753_n8421# a_34006_n8625# a_32951_n8793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X74 vdd d0 a_12197_n4940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X75 gnd d0 a_29568_n4952# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X76 a_30684_6068# a_30691_6286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X77 a_25191_7654# a_25205_8437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X78 a_21926_5025# a_21933_5243# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X79 a_26265_2708# a_26267_3001# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X80 a_24156_2946# d2 a_24239_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X81 a_20647_n8795# a_20900_n8999# a_19850_n8567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X82 a_1229_n2802# a_1023_n3410# a_443_n3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X83 vdd d1 a_11400_n4712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X84 gnd d0 a_16741_3582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X85 a_13331_6781# a_13333_7074# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X86 a_15568_2116# d1 a_15654_1331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X87 a_3253_n7541# a_3510_n7557# a_2455_n7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X88 a_23042_n3666# d3 a_23141_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X89 a_26649_n8309# d1 a_27446_n8770# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X90 a_26735_2289# a_26517_2289# a_26254_2201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X91 gnd d1 a_33171_n6773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X92 a_25615_n10665# a_25872_n10681# a_17125_n10728# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X93 a_15491_n3503# a_15744_n3707# a_15392_n3093# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 gnd d1 a_15837_n8797# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X95 a_6678_n8160# d2 a_6757_n9364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X96 a_2603_4347# d0 a_3396_4752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X97 a_15641_6188# a_15898_5998# a_15595_7208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X98 a_24202_1926# a_24455_1913# a_24152_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X99 a_6684_n5292# a_6941_n5308# a_6605_n4088# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X100 gnd d0 a_20791_n2479# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X101 a_29531_5630# a_29545_6413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X102 a_26735_2289# d1 a_27521_1616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X103 a_15641_6188# d1 a_15727_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X104 a_22124_847# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X105 a_7563_n4912# a_7567_n4724# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X106 a_26809_5949# a_26591_5949# a_26318_5956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X107 a_1334_n8733# a_1116_n8500# a_536_n8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X108 a_33715_n6797# a_33968_n7001# a_32918_n6569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X109 a_30795_n8322# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X110 a_20730_2728# a_20734_2551# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X111 a_25078_1311# a_25082_1134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X112 a_16309_n4337# a_16304_n4937# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X113 a_2365_n2635# d0 a_3163_n2451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X114 a_14291_1088# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X115 a_24100_n2660# d0 a_24898_n2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X116 a_26195_n9957# a_29658_n10042# a_28608_n9610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 vdd d0 a_16722_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X118 a_14587_5689# a_14381_6178# a_13802_5950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X119 a_33748_n9021# a_34005_n9037# a_32955_n8605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X120 a_28533_2958# a_28786_2945# a_28426_5173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X121 a_20754_3569# a_21007_3556# a_19957_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X122 a_4917_n9715# a_4699_n9715# a_4436_n9426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X123 gnd d0 a_8090_8647# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X124 a_22938_2093# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X125 a_27388_6177# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X126 gnd d1 a_28807_n6760# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X127 a_18957_2488# a_18739_2488# a_18863_2607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X128 a_32951_n8793# a_33208_n8809# a_32869_n9401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X129 gnd d0 a_29641_n9024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 gnd d0 a_20845_n5533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X131 a_11134_n9376# d1 a_11216_n8768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X132 vdd d0 a_29712_1133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X133 a_24132_n9188# a_24385_n9392# a_24049_n8172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X134 a_27589_5159# a_27371_5159# a_26792_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 gnd d1 a_7076_n7754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X136 a_7711_1122# a_7706_1711# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X137 a_4506_2177# a_4512_2360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X138 a_1307_n3641# a_1105_n2802# a_1224_n2625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_4645_n6661# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X140 a_23011_6165# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X141 a_29351_n6784# a_29604_n6988# a_28554_n6556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X142 a_12141_4600# a_12157_5383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X143 a_21798_n9121# d0 a_22289_n9315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X144 a_11323_3531# a_11580_3341# a_11241_4139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X145 vdd d0 a_3473_n5933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X146 gnd d1 a_11453_n7766# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X147 a_245_n4612# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X148 a_14831_403# a_14649_4548# a_14764_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X149 a_25204_8849# a_25208_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X150 a_5579_n8923# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X151 a_21993_8480# a_20844_8659# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X152 a_31783_n3691# d3 a_31882_n3868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X153 a_17850_5924# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X154 a_7620_n7778# a_7873_n7982# a_6823_n7550# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X155 a_4700_n9303# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X156 gnd d0 a_33895_n2929# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X157 a_32918_n6569# d0 a_33715_n6797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X158 a_23254_7712# a_23048_8201# a_22469_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X159 a_5759_7581# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X160 a_21941_5944# d0 a_22432_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X161 a_5703_n8923# d2 a_5749_n7903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X162 a_24022_n3080# d1 a_24121_n3490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X163 a_7711_1122# a_7964_1109# a_6909_1483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X164 a_185_4383# d0 a_660_4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X165 a_26430_n8721# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X166 a_17395_n6554# d0 a_17870_n6660# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X167 a_2494_6993# d2 a_2573_8186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X168 a_31735_5172# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X169 gnd d1 a_33098_n2701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X170 a_26410_n7703# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X171 a_1380_n7713# a_1178_n6874# a_1302_n6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X172 a_6090_378# a_5908_4523# a_6023_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X173 a_13785_4932# a_13567_4932# a_13296_5038# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X174 a_4845_n5231# d1 a_5630_n4851# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X175 a_6856_n9774# a_7113_n9790# a_6761_n9176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X176 a_7784_5194# a_7779_5783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X177 gnd d0 a_8001_3145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X178 a_18678_n3653# a_18476_n2814# a_18595_n2637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X179 a_10150_1604# a_9944_2093# a_9364_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X180 vdd d0 a_16741_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X181 a_24214_n8580# d0 a_25011_n8808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X182 gnd d1 a_15961_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X183 a_18450_n6476# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X184 a_26094_n4360# a_26100_n4543# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X185 a_27932_283# d6 a_26029_208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X186 a_55_n8395# d0 a_536_n8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X187 a_18812_3098# d2 a_18863_2607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X188 a_28608_n9610# a_28861_n9814# a_28509_n9200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X189 a_228_7036# d0 a_717_6930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X190 vdd d0 a_21061_6198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X191 a_32058_n5902# a_31840_n5902# a_31882_n3868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X192 vdd d1 a_20047_n5717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X193 a_2603_4347# d0 a_3400_4575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X194 vdd d0 a_25244_n7994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X195 gnd d1 a_20300_8418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X196 a_17449_n9608# d0 a_17924_n9714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X197 a_22358_2277# a_22140_2277# a_21883_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X198 a_515_8360# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X199 a_17487_841# a_17489_940# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 gnd d1 a_28951_3353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X201 gnd d1 a_33152_n5755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X202 a_27118_n2429# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X203 a_78_n9596# d0 a_553_n9702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X204 gnd d1 a_16034_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X205 a_2393_n9351# d1 a_2479_n8555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X206 a_14826_284# d5 a_12951_197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X207 a_30721_n4662# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X208 a_30701_n3644# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X209 a_18751_n7725# a_18549_n6886# a_18673_n6886# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X210 gnd d1 a_7003_n3682# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X211 a_22359_1865# d1 a_23144_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X212 vdd d1 a_2712_n7741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X213 gnd d0 a_12340_1533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 a_16525_5219# a_16778_5206# a_15723_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_17869_7354# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X216 a_25024_n10014# a_21818_n9945# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X217 a_20750_3746# a_21007_3556# a_19957_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X218 a_2536_6150# d1 a_2618_5542# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X219 gnd d1 a_29024_7425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X220 a_13133_n7197# a_13140_n7415# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X221 a_23394_6573# a_23176_6573# a_23295_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 a_4609_8067# d0 a_5098_7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X223 vdd d0 a_8073_7629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X224 a_10323_n5877# a_10105_n5877# a_10220_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X225 a_9183_4313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X226 a_7547_n3706# a_7800_n3910# a_6750_n3478# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X227 a_26610_7379# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X228 gnd d0 a_7893_n9000# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X229 a_6678_5149# d3 a_6785_2934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X230 a_9241_n6261# a_9023_n6261# a_8750_n6067# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X231 a_1240_4104# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X232 a_8733_n5148# a_8740_n5366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X233 a_10223_5676# d2 a_10301_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X234 a_28602_7207# d2 a_28652_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X235 a_11994_n7566# a_11998_n7378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X236 a_3379_3734# a_3383_3557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X237 a_20717_1533# a_20970_1520# a_19920_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X238 a_16468_2577# a_16721_2564# a_15671_2349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X239 a_21740_n5549# d0 a_22215_n5655# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 vdd d0 a_12215_n5546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X241 a_11417_8444# d0 a_12214_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X242 a_15580_n8781# d0 a_16382_n8409# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X243 a_28287_n10602# d5 a_27694_n5889# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X244 vdd d0 a_34149_5218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X245 a_5080_7355# d1 a_5878_7171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X246 a_3432_6788# a_3689_6598# a_2639_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X247 vdd d0 a_16615_n7595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X248 a_32135_6598# a_31917_6598# a_32041_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X249 a_4682_n8697# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X250 a_29458_1558# a_29711_1545# a_28661_1330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X251 gnd d1 a_33388_7438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X252 a_30711_7304# a_30717_7487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X253 a_33679_n4761# a_33693_n5555# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X254 a_9965_n2650# a_9747_n2417# a_9167_n2601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X255 a_27245_n9555# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X256 a_29454_1735# a_29458_1558# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X257 gnd d1 a_2802_1280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X258 a_13151_n8116# a_13153_n8215# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X259 a_15654_1331# d0 a_16447_1736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 a_28494_n3690# d0 a_29296_n3318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X261 a_13258_2709# d0 a_13749_2896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X262 a_31958_5701# a_31752_6190# a_31173_5962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X263 a_33733_n7403# a_33986_n7607# a_32931_n7775# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X264 a_28468_n7352# a_28725_n7368# a_28422_n8372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X265 vdd d0 a_8001_3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X266 a_17353_n4335# d0 a_17834_n4624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X267 gnd d2 a_15645_n3297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X268 vdd d1 a_15961_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X269 a_23811_n10590# d4 a_23873_n6138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X270 a_18885_7170# a_18667_7170# a_18087_7354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X271 a_10121_n7738# a_9919_n6899# a_10038_n6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_11065_n5116# a_11318_n5320# a_10982_n4100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X273 a_1358_5532# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 a_13585_n5668# d1 a_14371_n4876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X275 a_11233_n9786# d0 a_12031_n9602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X276 a_13368_n5256# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X277 a_26160_n8214# a_26167_n8432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X278 vdd d1 a_28951_3353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X279 vdd d2 a_7121_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X280 vdd d1 a_16034_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X281 a_9219_6349# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X282 a_13097_n5161# d0 a_13586_n5256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X283 a_13548_n3632# a_13330_n3632# a_13073_n3526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X284 a_20537_n2687# a_20790_n2891# a_19740_n2459# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 a_24334_4549# a_24591_4359# a_24239_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X286 a_29401_n10026# a_29658_n10042# a_28608_n9610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X287 a_31536_n5496# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X288 a_26539_n2201# d1 a_27336_n2662# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X289 gnd d0 a_16578_n5971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 vdd d0 a_12340_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X291 a_6601_n4276# d2 a_6647_n3256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X292 a_6831_1914# a_7084_1901# a_6781_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X293 vdd d0 a_3547_n9593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X294 a_30957_n5268# a_30739_n5268# a_30466_n5074# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X295 a_2586_3329# a_2839_3316# a_2500_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_2536_6150# d1 a_2622_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X297 vdd d1 a_29024_7425# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X298 a_463_n4612# d1 a_1261_n4661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X299 a_11396_7603# d0 a_12198_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X300 a_4828_n4213# a_4610_n4213# a_4337_n4019# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X301 a_17382_n6153# a_17389_n6371# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X302 a_18031_4300# a_17813_4300# a_17550_4212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X303 a_19773_n4683# a_20030_n4699# a_19691_n5291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X304 a_1186_1050# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X305 a_13659_n9328# d1 a_14444_n8948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X306 a_26358_n4237# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X307 a_17148_133# a_25910_208# a_21680_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X308 a_29278_n2712# a_29292_n3506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X309 gnd d1 a_20083_n7753# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X310 a_26538_n2613# a_26320_n2613# a_26057_n2324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X311 a_4863_n6661# d1 a_5661_n6710# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X312 vdd d0 a_12413_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X313 gnd d4 a_2571_4946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X314 a_20713_1710# a_20970_1520# a_19920_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X315 a_19937_2323# a_20190_2310# a_19838_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X316 a_1560_6548# a_1358_5532# a_1482_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X317 a_28353_n4112# d2 a_28432_n5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 a_16464_2754# a_16721_2564# a_15671_2349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X319 a_4752_1247# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X320 a_5698_n8746# a_5480_n8513# a_4900_n8697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X321 a_15491_n3503# d0 a_16288_n3731# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X322 a_228_7036# a_235_7254# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X323 a_27172_n5483# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X324 a_13658_n9740# a_13440_n9740# a_13177_n9451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X325 a_9437_6349# a_9219_6349# a_8962_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X326 a_8802_n8603# d0 a_9277_n8709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X327 gnd d0 a_29548_n3934# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X328 a_21868_1872# a_21870_1971# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X329 a_2314_5136# a_2571_4946# a_1721_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X330 a_4579_6249# a_4585_6432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X331 a_24227_n9786# d0 a_25029_n9414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X332 a_33692_n5967# a_33949_n5983# a_32899_n5551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X333 a_25188_7419# a_25445_7229# a_24390_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X334 vdd d5 a_15438_n10619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X335 a_23047_n3843# d3 a_23141_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_32841_n2685# a_33098_n2701# a_32759_n3293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X337 a_26648_n8721# d1 a_27446_n8770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X338 gnd d1 a_28751_n3706# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X339 a_29454_1735# a_29711_1545# a_28661_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X340 a_7531_n2276# a_7784_n2480# a_6729_n2648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X341 a_5851_2489# a_5649_1473# a_5768_1063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X342 a_21956_6444# a_21961_6768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X343 a_28730_5579# d0 a_29528_5395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X344 a_20768_4352# a_20772_4175# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X345 gnd d1 a_15817_n7779# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X346 a_25607_n2057# a_24898_n2476# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X347 a_26321_n2201# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X348 vdd d2 a_7014_n9380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X349 vdd d1 a_28788_n5742# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X350 a_16268_n2489# a_16272_n2301# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X351 a_17759_1246# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X352 vdd d1 a_2802_1280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X353 a_15654_1331# d0 a_16451_1559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X354 a_33895_5643# a_34148_5630# a_33098_5415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_19907_6162# d1 a_19989_5554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X356 gnd d0 a_25351_2551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X357 a_21866_1354# d0 a_22341_1259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X358 a_6601_n4276# a_6858_n4292# a_6498_n6314# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X359 a_30795_n8322# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X360 a_33873_4390# a_33877_4213# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X361 a_10220_n7915# a_10002_n7915# a_10126_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X362 gnd d2 a_28762_n9404# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X363 a_25115_3347# a_25119_3170# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X364 a_30775_n7304# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X365 a_16361_n7803# a_16614_n8007# a_15564_n7575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X366 a_28678_2348# d0 a_29471_2753# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X367 a_18105_7960# a_17887_7960# a_17616_8066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X368 a_26333_6456# d0 a_26808_6361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X369 a_24049_5161# d3 a_24156_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X370 a_31716_4154# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X371 a_15419_n8185# a_15672_n8389# a_15243_n6151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 vdd d1 a_11363_n2676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X373 vdd d0 a_25155_n2492# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X374 gnd d0 a_25424_6623# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 gnd d2 a_15682_n5333# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X376 a_13566_5344# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X377 a_13766_3914# a_13548_3914# a_13277_4020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X378 a_13440_n9740# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X379 a_n25_n4105# d0 a_464_n4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X380 a_162_3182# a_168_3365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X381 a_30502_n7110# a_30504_n7209# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X382 a_22178_3901# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X383 a_26121_n6079# d0 a_26612_n6273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X384 a_31917_3136# a_31699_3136# a_31120_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X385 a_11101_n7152# d1 a_11196_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X386 a_2423_n5501# d0 a_3220_n5729# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X387 a_11123_n3678# a_11380_n3694# a_11028_n3080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X388 a_13729_1878# a_13511_1878# a_13240_1984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X389 a_21800_n9220# d0 a_22289_n9315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X390 a_17977_1246# a_17759_1246# a_17502_1341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X391 a_245_n4612# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_2582_3506# a_2839_3316# a_2500_4114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X393 gnd d1 a_2929_8406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X394 a_27599_2513# d3 a_27698_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X395 a_8930_4926# a_8932_5025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X396 a_1820_246# a_1602_246# a_1721_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 a_26756_2895# a_26538_2895# a_26267_3001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X398 a_25188_7419# a_25192_7242# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X399 a_18574_2080# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X400 a_5579_n8923# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 a_16361_n7803# a_16378_n8597# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X402 a_4700_n9303# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X403 a_9421_4919# a_9203_4919# a_8932_5025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X404 a_31990_7208# a_31772_7208# a_31193_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X405 a_3396_4752# a_3400_4575# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X406 a_n10_n5024# a_n8_n5123# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X407 a_19757_n3477# d0 a_20550_n3893# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X408 a_12013_n8996# a_12270_n9012# a_11220_n8580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X409 a_17417_n8090# d0 a_17908_n8284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X410 a_30438_n3355# a_30444_n3538# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X411 gnd d0 a_20918_n9605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X412 a_26410_n7703# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X413 a_19933_2500# a_20190_2310# a_19838_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X414 a_13313_n2614# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X415 gnd d0 a_12451_7229# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X416 a_643_3270# d1 a_1441_3086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_1380_n7713# a_1178_n6874# a_1297_n6697# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X418 a_14128_n3448# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X419 a_20610_n6759# a_20624_n7553# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X420 a_16506_4201# a_16759_4188# a_15704_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X421 a_8686_n2312# a_8692_n2495# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X422 a_2504_3937# d1 a_2599_4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X423 gnd d2 a_24528_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 a_318_n8684# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X425 a_30728_8322# a_30734_8505# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X426 a_7821_7230# a_7816_7819# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X427 a_16308_n4749# a_16561_n4953# a_15511_n4521# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 a_4532_3378# a_4534_3896# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X429 gnd d0 a_25335_1121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X430 a_3273_n8559# a_3530_n8575# a_2475_n8743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X431 a_27714_283# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X432 a_24952_n5530# a_24956_n5342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X433 a_24194_n7562# d0 a_24991_n7790# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X434 a_15243_n6151# a_15496_n6355# a_15181_n10603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X435 a_8976_7279# d0 a_9457_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X436 a_716_7342# d1 a_1514_7158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X437 a_35_n7377# d0 a_516_n7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X438 a_30427_n2520# a_30429_n3038# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X439 a_29496_3182# a_29749_3169# a_28694_3543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X440 a_14582_5160# a_14364_5160# a_13784_5344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X441 a_22199_n4225# d1 a_22996_n4686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X442 a_22921_1075# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X443 a_15522_3136# d2 a_15572_1939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X444 a_31834_5582# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X445 vdd d4 a_15676_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X446 a_32552_n10615# d4 a_32610_n6351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X447 a_10260_7712# d2 a_10306_6692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X448 a_19654_n3255# d1 a_19740_n2459# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X449 a_33891_5820# a_34148_5630# a_33098_5415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X450 a_19907_6162# d1 a_19993_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X451 vdd d0 a_25351_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X452 a_20611_n6347# a_20864_n6551# a_19809_n6719# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X453 a_26592_n5667# a_26374_n5667# a_26117_n5561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X454 a_2360_n7127# d1 a_2459_n7537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X455 a_13123_n6397# d0 a_13604_n6686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X456 a_30701_n3644# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X457 vdd d0 a_34130_4200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X458 a_33877_4213# a_33872_4802# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X459 a_24407_8621# d0 a_25209_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X460 vdd d0 a_20917_n10017# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X461 a_31737_n4711# d2 a_31788_n3868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X462 a_23176_3111# a_22958_3111# a_22378_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X463 vdd d6 a_12949_n10693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X464 a_18067_6336# d1 a_18853_5663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X465 a_28678_2348# d0 a_29475_2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X466 a_7816_7819# a_7820_7642# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X467 a_7838_8248# a_8091_8235# a_7036_8609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_4605_7450# a_4607_7968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X469 a_8926_4408# a_8930_4926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X470 vdd d0 a_25424_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X471 a_23976_n4100# a_24229_n4304# a_23869_n6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X472 a_5686_3509# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X473 gnd d0 a_25208_n5958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X474 a_10323_n5877# a_10105_n5877# a_10147_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X475 a_2318_4959# d3 a_2494_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X476 a_16381_n8821# a_16634_n9025# a_15584_n8593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X477 a_11160_n5714# d0 a_11962_n5342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X478 a_28531_n5726# d0 a_29329_n5542# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X479 a_16345_n6373# a_16598_n6577# a_15543_n6745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 a_162_3182# d0 a_643_3270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X481 vdd d2 a_2757_3924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X482 a_15691_3367# d0 a_16484_3772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X483 a_13346_7475# d0 a_13821_7380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X484 a_29312_n4524# a_29569_n4540# a_28514_n4708# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X485 a_30691_6286# d0 a_31172_6374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X486 gnd d2 a_11498_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X487 a_33872_4802# a_33876_4625# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X488 a_15560_n7763# d0 a_16362_n7391# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X489 a_27373_n4698# d2 a_27424_n3855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X490 a_13146_n7598# a_13151_n8116# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X491 a_7710_1534# a_7963_1521# a_6913_1306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X492 a_30938_4944# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X493 a_31773_n6747# d2 a_31856_n7763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X494 a_19826_n7737# a_20083_n7753# a_19731_n7139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X495 a_30882_1890# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 a_22431_6349# a_22213_6349# a_21950_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X497 a_6085_259# d4 a_6682_4972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X498 a_26501_859# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X499 a_13247_2202# a_13253_2385# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X500 a_3347_1109# a_3600_1096# a_2545_1470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X501 a_8746_n5549# a_8750_n6067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X502 a_17797_2870# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X503 a_26629_n7291# a_26411_n7291# a_26140_n7196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X504 vdd d0 a_7911_n9606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X505 a_n38_n3305# d0 a_443_n3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X506 a_17389_n6371# d0 a_17870_n6660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X507 a_9965_n2650# a_9747_n2417# a_9168_n2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X508 a_9256_8385# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X509 a_27245_n9555# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X510 a_14148_n4466# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X511 a_30881_2302# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X512 gnd d0 a_34022_n10055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X513 a_17616_n4624# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X514 vdd d0 a_12288_n9618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X515 a_23869_n6326# d3 a_23976_n4100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X516 a_15342_n4301# d2 a_15388_n3281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X517 a_2504_3937# d1 a_2603_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X518 a_19794_n5513# d0 a_20587_n5929# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 a_4517_2684# d0 a_5008_2871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X520 a_13569_n4238# a_13351_n4238# a_13078_n4044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_17359_n4518# d0 a_17834_n4624# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X522 vdd d0 a_25335_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X523 a_17333_n3317# d0 a_17814_n3606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X524 a_8876_1971# a_8883_2189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X525 a_31173_5962# d1 a_31958_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X526 a_15543_n6745# d0 a_16345_n6373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X527 a_14165_n5484# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X528 a_11237_n9598# d0 a_8824_n9945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X529 a_33697_n5367# a_33692_n5967# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X530 a_13043_n2107# a_13050_n2325# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X531 a_2577_8009# d1 a_2676_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X532 a_13368_n5256# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X533 a_21710_n4130# a_21717_n4348# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X534 a_8658_196# d7 a_8757_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X535 a_24214_n8580# a_24467_n8784# a_24128_n9376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X536 a_20731_2316# a_20735_2139# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X537 a_13548_n3632# a_13330_n3632# a_13067_n3343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 a_33152_8469# d0 a_33945_8874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X539 a_27118_n2429# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X540 a_17539_3377# d0 a_18014_3282# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X541 a_12105_2152# a_12358_2139# a_11303_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 gnd d0 a_20863_n6963# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X543 a_2492_n9761# d0 a_3294_n9389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X544 vdd d1 a_7276_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X545 a_28612_4151# a_28869_3961# a_28533_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X546 a_23115_n7738# a_22913_n6899# a_23037_n6899# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X547 a_12161_5206# a_12414_5193# a_11359_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X548 a_1519_7687# a_1313_8176# a_734_7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X549 a_7834_8425# a_8091_8235# a_7036_8609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X550 vdd d2 a_28689_n5332# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X551 a_28711_4561# d0 a_29509_4377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X552 a_20043_8608# d0 a_20841_8424# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X553 a_27518_n3855# a_27300_n3855# a_27424_n3855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X554 a_4572_n2589# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X555 a_17579_6030# a_17586_6248# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X556 a_17599_7048# d0 a_18088_6942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 vdd d2 a_33089_n7381# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X558 a_15671_2349# a_15924_2336# a_15572_1939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 a_9384_3295# d1 a_10182_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X560 a_13658_n9740# d1 a_14444_n8948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_4808_n3195# a_4590_n3195# a_4317_n3001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X562 a_12832_197# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_19753_n3665# a_20010_n3681# a_19658_n3067# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X564 vdd d3 a_32970_n4329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X565 vdd d0 a_12160_n2904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X566 a_33876_4625# a_34129_4612# a_33079_4397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X567 a_7820_7642# a_7834_8425# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X568 a_19875_3949# d1 a_19970_4536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X569 a_8759_n6384# d0 a_9240_n6673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X570 a_8796_n8420# a_8802_n8603# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X571 a_15691_3367# d0 a_16488_3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X572 a_28784_8633# d0 a_29582_8449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X573 a_8872_1354# d0 a_9347_1259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X574 a_9059_n8709# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X575 a_28661_1330# a_28914_1317# a_28575_2115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X576 a_125_1146# a_131_1329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X577 a_12101_2329# a_12105_2152# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X578 a_5630_n4851# a_5424_n5459# a_4845_n5231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X579 a_14334_n2840# d2 a_14412_n3679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X580 a_21903_3390# d0 a_22378_3295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X581 a_5698_n8746# a_5480_n8513# a_4901_n8285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X582 a_7706_1711# a_7963_1521# a_6913_1306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X583 a_4210_172# a_5966_259# a_6090_378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X584 a_6930_2324# a_7183_2311# a_6831_1914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X585 a_17395_n6554# a_17397_n7072# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X586 a_8782_n7585# d0 a_9257_n7691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_11059_4984# d3 a_11235_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X588 a_9820_n6489# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X589 a_20786_5782# a_20790_5605# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X590 a_29296_n3318# a_29291_n3918# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X591 a_15568_2116# d1 a_15650_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X592 a_9129_1259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X593 gnd d0 a_33986_n7607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X594 a_258_8455# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X595 gnd d0 a_7857_n6552# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X596 a_5878_7171# a_5660_7171# a_5081_6943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X597 a_3437_6199# a_3432_6788# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X598 a_26321_n2201# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X599 gnd d0 a_12234_n6564# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X600 a_28426_n8184# d2 a_28505_n9388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X601 a_11290_1318# d0 a_12083_1723# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X602 a_23873_n6138# a_24126_n6342# a_23811_n10590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X603 a_32062_2526# a_31844_2526# a_31963_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X604 a_21727_n5148# a_21734_n5366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X605 a_6787_n5514# d0 a_7584_n5742# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X606 a_11143_n4696# d0 a_11941_n4512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X607 a_30638_3232# d0 a_31119_3320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X608 a_13131_n7098# d0 a_13622_n7292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X609 a_10220_n7915# a_10002_n7915# a_10121_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X610 gnd d0 a_29621_n8006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X611 a_26666_n9327# a_26448_n9327# a_26177_n9232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X612 a_22233_7367# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X613 a_30775_n7304# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X614 vdd d3 a_6931_n8364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X615 a_24225_7195# a_24482_7005# a_24053_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X616 a_11024_n3268# d1 a_11110_n2472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X617 a_8883_2189# a_8889_2372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X618 a_27191_n6501# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X619 gnd d0 a_427_n2164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X620 vdd d2 a_20128_3936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X621 a_23300_6692# a_23130_7593# a_23249_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X622 a_24902_n2288# a_24897_n2888# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X623 a_32976_4164# d1 a_33058_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X624 a_23141_n3843# d4 a_23317_n5877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X625 a_4826_4907# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 a_1385_n7890# d3 a_1479_n7890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X627 a_26394_n6273# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X628 a_16465_2342# a_16469_2165# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X629 vdd d2 a_15862_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X630 a_16520_5808# a_16777_5618# a_15727_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X631 a_33053_8059# a_33306_8046# a_32970_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X632 a_33152_8469# d0 a_33949_8697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X633 a_25081_1546# a_25334_1533# a_24284_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 a_30902_2908# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X635 a_n45_n3087# d0 a_444_n3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X636 a_26123_n6178# d0 a_26612_n6273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X637 vdd d0 a_16759_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X638 a_15580_n8781# a_15837_n8797# a_15498_n9389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X639 a_29389_n8408# a_29642_n8612# a_28587_n8780# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X640 gnd d5 a_24068_n10606# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X641 a_32893_3148# a_33150_2958# a_32790_5186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X642 vdd d0 a_12233_n6976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X643 a_33840_2177# a_33835_2766# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X644 a_20043_8608# d0 a_20845_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X645 a_225_n3594# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X646 a_4971_835# d1 a_5768_1063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X647 gnd d3 a_33223_7030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X648 gnd d1 a_20263_6382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X649 a_30957_n5268# a_30739_n5268# a_30468_n5173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X650 a_464_n4200# d1 a_1261_n4661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X651 a_15667_2526# a_15924_2336# a_15572_1939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X652 gnd d0 a_33933_n4553# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_9438_5937# d1 a_10223_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X654 a_4568_5414# a_4570_5932# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X655 a_29568_7666# a_29582_8449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X656 a_215_6236# d0 a_696_6324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X657 a_6781_3111# d2 a_6827_2091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X658 a_3380_3322# a_3384_3145# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X659 a_33872_4802# a_34129_4612# a_33079_4397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X660 a_18777_n3830# d4 a_18953_n5864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X661 a_3183_n3693# a_3200_n4487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X662 a_23048_8201# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X663 a_26247_1983# d0 a_26736_1877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_19875_3949# d1 a_19974_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X665 a_27327_n8947# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X666 a_29295_n3730# a_29312_n4524# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X667 a_31482_n2442# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X668 a_24137_n4696# d0 a_24939_n4324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X669 a_11993_n7978# a_12250_n7994# a_11200_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X670 a_28472_n7164# d1 a_28567_n7762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X671 gnd d0 a_16524_n2917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X672 a_17397_n7072# d0 a_17888_n7266# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X673 gnd d0 a_7784_n2480# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X674 a_28494_n3690# a_28751_n3706# a_28399_n3092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X675 a_13313_n2614# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X676 vdd d1 a_28844_n8796# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X677 vdd d0 a_3493_n6539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X678 a_26237_1183# d0 a_26718_1271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X679 a_20570_n4911# a_20574_n4723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X680 a_10343_271# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X681 gnd d1 a_29004_6407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X682 a_28550_n6744# a_28807_n6760# a_28468_n7352# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X683 a_26230_965# a_26237_1183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X684 a_18656_1472# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X685 gnd d1 a_15727_n2689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X686 a_33912_6661# a_33929_7444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X687 a_18637_n4850# d2 a_18683_n3830# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X688 a_6926_2501# a_7183_2311# a_6831_1914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X689 a_19731_n7139# a_19984_n7343# a_19681_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X690 a_13658_n9740# a_13440_n9740# a_13183_n9634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X691 a_8796_n8420# d0 a_9277_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X692 a_26254_2201# d0 a_26735_2289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X693 a_18105_7960# a_17887_7960# a_17614_7967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X694 a_30702_6793# a_30704_7086# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X695 a_298_n7666# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X696 a_23037_n6899# d2 a_23115_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X697 a_4427_n9109# a_4429_n9208# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X698 a_2442_n6519# d0 a_3239_n6747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X699 a_16288_n3731# a_16541_n3935# a_15491_n3503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X700 a_27677_6704# d3 a_27771_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X701 a_41_n7560# d0 a_516_n7666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X702 a_25029_n9414# a_25282_n9618# a_24227_n9786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X703 a_2356_n7315# d1 a_2442_n6519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X704 a_26718_1271# d1 a_27516_1087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X705 a_19689_4971# a_19942_4958# a_19092_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X706 a_22198_n4637# d1 a_22996_n4686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X707 a_9364_2277# a_9146_2277# a_8883_2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 gnd d3 a_28606_n4316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X709 a_10048_n3666# a_9846_n2827# a_9970_n2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X710 a_32862_n3515# d0 a_33655_n3931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X711 a_22179_n3207# d1 a_22964_n2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X712 a_7543_n3894# a_7547_n3706# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X713 a_28579_1938# d1 a_28674_2525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 a_14687_n5890# a_14469_n5890# a_14511_n3856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X715 a_20628_n7365# a_20623_n7965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X716 a_13386_n6686# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X717 a_11290_1318# d0 a_12087_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X718 a_12177_6636# a_12194_7419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X719 a_46_n8078# a_48_n8177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X720 a_31618_n4888# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X721 a_14592_2514# a_14390_1498# a_14514_1617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X722 a_6930_2324# d0 a_7727_2552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X723 a_30919_3926# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X724 a_26592_n5667# a_26374_n5667# a_26111_n5378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 vdd d4 a_32867_n6367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X726 a_30475_n5391# a_30481_n5574# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X727 a_32610_n6351# d3 a_32713_n4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X728 a_3166_n2675# a_3419_n2879# a_2369_n2447# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X729 a_6647_n3256# d1 a_6729_n2648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 a_16322_n5543# a_16579_n5559# a_15524_n5727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X731 a_17212_n839# d8 a_17125_n10728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X732 a_2287_n3055# a_2540_n3259# a_2237_n4263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X733 a_26303_5037# a_26310_5255# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X734 a_10109_2501# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X735 a_22469_7973# a_22251_7973# a_21978_7980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X736 a_13641_n8722# a_13423_n8722# a_13166_n8616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X737 a_22178_n3619# a_21960_n3619# a_21697_n3330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X738 a_4590_n3195# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X739 a_1721_246# d4 a_2314_5136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X740 a_32976_4164# d1 a_33062_3379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X741 a_30992_7998# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X742 gnd d5 a_32809_n10631# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X743 a_23020_1485# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X744 a_1477_5122# a_1259_5122# a_680_4894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X745 vdd d0 a_12178_n3510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X746 a_1602_246# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X747 gnd d0 a_8073_7629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X748 a_33049_8236# a_33306_8046# a_32970_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X749 a_5567_2081# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X750 a_28432_n5316# d1 a_28514_n4708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_25077_1723# a_25334_1533# a_24284_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X752 a_31210_7998# a_30992_7998# a_30719_8005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X753 a_19727_n7327# d1 a_19813_n6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X754 a_31136_4338# a_30918_4338# a_30661_4433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X755 a_33748_n9021# a_33752_n8833# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X756 a_21851_854# d0 a_22342_847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X757 a_13440_n9740# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X758 a_5676_n3831# a_5506_n4851# a_5630_n4851# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X759 a_17504_1859# d0 a_17995_1852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X760 gnd d1 a_2659_n4687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X761 a_22468_8385# a_22250_8385# a_21993_8480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X762 a_27254_n4875# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X763 a_21421_n10664# d6 a_21322_n10664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X764 a_3220_n5729# a_3473_n5933# a_2423_n5501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X765 a_27378_n4875# d2 a_27424_n3855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X766 vdd d0 a_20790_n2891# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X767 a_11417_8444# d0 a_12210_8849# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X768 a_10879_n6138# d3 a_11051_n8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X769 vdd d3 a_33223_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X770 a_7584_n5742# a_7600_n6536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X771 vdd d1 a_20263_6382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X772 a_7568_n4312# a_7563_n4912# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X773 a_8696_n3112# a_8703_n3330# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X774 a_31778_n6924# d2 a_31856_n7763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X775 gnd d0 a_34149_5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_30717_7487# a_30719_8005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X777 a_27414_n6911# a_27208_n7519# a_26629_n7291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X778 a_2423_n5501# a_2676_n5705# a_2324_n5091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X779 a_19658_n3067# a_19911_n3271# a_19608_n4275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X780 a_26029_208# a_30203_209# a_30322_209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X781 gnd d2 a_20091_1900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 vdd d6 a_30320_n10705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X783 a_17212_n839# d9 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X784 a_2369_n2447# d0 a_3166_n2675# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X785 a_24301_2336# d0 a_25094_2741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 vdd d1 a_7096_n8772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X787 a_22123_1259# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X788 a_10327_2501# a_10109_2501# a_10233_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X789 a_24104_n2472# d0 a_24901_n2700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X790 a_2566_2311# a_2819_2298# a_2467_1901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X791 a_14148_n4466# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X792 a_26590_6361# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X793 gnd d0 a_3727_8222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X794 a_17616_n4624# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X795 a_23115_n7738# d3 a_23214_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X796 a_14128_n3448# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X797 a_21868_1872# d0 a_22359_1865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X798 a_19030_6560# d4 a_19097_377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X799 a_28734_5402# d0 a_29531_5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X800 a_12193_7831# a_12197_7654# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X801 a_26074_n3342# a_26080_n3525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X802 a_17596_n3606# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X803 a_10467_390# a_10285_4535# a_10327_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X804 a_22197_4919# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X805 a_8679_n2094# d0 a_9168_n2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X806 vdd d0 a_20844_n5945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X807 a_12174_6401# a_12178_6224# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X808 a_17339_n3500# d0 a_17814_n3606# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X809 gnd d1 a_24430_n6748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X810 a_31958_5701# d2 a_32036_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X811 a_19794_n5513# a_20047_n5717# a_19695_n5103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X812 gnd d2 a_28832_1925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 a_30902_n2626# a_30684_n2626# a_30427_n2520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X814 a_23222_2501# d3 a_23321_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X815 a_22379_2883# a_22161_2883# a_21890_2989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X816 a_31705_n2852# a_31499_n3460# a_30920_n3232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X817 a_9130_847# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X818 vdd d4 a_11312_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X819 a_28579_1938# d1 a_28678_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X820 vdd d1 a_24610_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X821 a_11997_n7790# a_12014_n8584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X822 a_9222_n5243# d1 a_10007_n4863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X823 a_12014_n8584# a_12018_n8396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X824 a_24194_n7562# a_24447_n7766# a_24095_n7152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X825 a_14691_2514# a_14473_2514# a_14592_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X826 a_8714_n4031# a_8716_n4130# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X827 vdd d0 a_20987_2538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X828 a_27480_2513# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X829 a_13333_7074# d0 a_13822_6968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X830 a_17689_n8696# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X831 a_22341_1259# a_22123_1259# a_21866_1354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X832 a_24338_4372# a_24591_4359# a_24239_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X833 vdd d1 a_24627_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X834 a_30954_6374# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X835 a_31120_2908# a_30902_2908# a_30631_3014# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X836 a_23394_6573# d4 a_23461_390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X837 a_21680_n2312# a_21686_n2495# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X838 a_31761_1510# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X839 a_13056_n2508# a_13058_n3026# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X840 a_22198_n4637# a_21980_n4637# a_21723_n4531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X841 a_27518_n3855# a_27300_n3855# a_27419_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X842 a_21890_2989# a_21897_3207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X843 a_25135_4600# a_25151_5383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X844 a_32841_n2685# d0 a_33639_n2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 a_15605_4152# d1 a_15687_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X846 a_18853_5663# a_18647_6152# a_18068_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X847 a_11396_7603# d0 a_12194_7419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X848 a_10978_n4288# d2 a_11028_n3080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X849 a_1223_3086# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X850 gnd d4 a_28683_4983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 a_13258_2709# a_13260_3002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X852 a_7036_8609# d0 a_7834_8425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X853 gnd d2 a_33196_1938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X854 a_15682_8047# a_15935_8034# a_15599_7031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X855 a_4599_7267# d0 a_5080_7355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X856 a_607_822# a_389_822# a_116_829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 a_24225_7195# d2 a_24271_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_8765_n6567# d0 a_9240_n6673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X859 a_13236_1367# a_13238_1885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X860 a_7640_n8796# a_7654_n9590# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X861 a_7654_n9590# a_7658_n9402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X862 a_13331_n3220# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X863 vdd d0 a_20881_n7569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X864 a_27626_7195# d2 a_27677_6704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X865 vdd d1 a_15781_n5743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X866 gnd d4 a_28503_n6354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_19850_n8567# d0 a_20643_n8983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X868 a_15498_n9389# a_15755_n9405# a_15419_n8185# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X869 a_5666_n6887# a_5460_n7495# a_4881_n7267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X870 a_8804_n9121# d0 a_9295_n9315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X871 a_27446_n8770# a_27228_n8537# a_26648_n8721# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X872 a_25192_7242# a_25445_7229# a_24390_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X873 a_14221_n8538# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X874 vdd d0 a_29531_n2916# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X875 a_16501_4790# a_16758_4600# a_15708_4385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X876 vdd d2 a_28652_n3296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X877 a_24301_2336# d0 a_25098_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X878 a_4789_3283# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X879 a_4863_6943# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X880 a_32790_n8197# d2 a_32873_n9213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X881 a_11179_n6732# d0 a_11977_n6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X882 a_7637_n8572# a_7641_n8384# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X883 a_17760_834# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X884 a_7581_n5518# a_7838_n5534# a_6783_n5702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X885 a_11904_n2476# a_12161_n2492# a_11106_n2660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X886 a_19792_2933# a_20045_2920# a_19685_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 a_13404_n7292# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X888 a_30719_8005# a_30721_8104# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X889 a_4900_n8697# a_4682_n8697# a_4425_n8591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X890 vdd d0 a_3727_8222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X891 a_29291_n3918# a_29548_n3934# a_28498_n3502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X892 a_26666_n9327# a_26448_n9327# a_26175_n9133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X893 a_498_7342# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X894 a_13569_n4238# a_13351_n4238# a_13080_n4143# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X895 a_209_n2164# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X896 a_8757_196# a_8539_196# a_8658_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X897 a_23099_n5877# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X898 a_13547_4326# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X899 a_30665_4951# a_30667_5050# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X900 a_5008_2871# a_4790_2871# a_4519_2977# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X901 a_8920_4225# a_8926_4408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X902 a_26140_n7196# a_26147_n7414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X903 a_27191_n6501# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X904 a_33766_n9627# a_34023_n9643# a_32968_n9811# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X905 a_12197_7654# a_12211_8437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X906 a_26338_6780# d0 a_26829_6967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X907 a_23214_n7915# d4 a_23317_n5877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 a_31082_1284# a_30864_1284# a_30601_1196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X909 a_31737_n4711# a_31519_n4478# a_30939_n4662# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X910 a_13603_7380# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X911 a_24952_n5530# a_25209_n5546# a_24154_n5714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X912 a_3342_1698# a_3346_1521# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X913 a_6839_n8756# d0 a_7637_n8572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X914 a_26394_n6273# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X915 a_21740_n5549# a_21744_n6067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X916 a_26537_3307# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X917 a_3179_n3881# a_3183_n3693# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X918 a_30721_8104# a_30728_8322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X919 a_7817_7407# a_7821_7230# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X920 a_11183_n6544# d0 a_11980_n6772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X921 vdd d1 a_2912_7388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X922 a_28554_n6556# d0 a_29347_n6972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X923 a_15560_n7763# a_15817_n7779# a_15465_n7165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X924 a_31742_n4888# a_31536_n5496# a_30957_n5268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X925 a_29369_n7390# a_29622_n7594# a_28567_n7762# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X926 a_31156_4944# a_30938_4944# a_30665_4951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X927 a_6963_4537# a_7220_4347# a_6868_3950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X928 a_18014_3282# a_17796_3282# a_17533_3194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X929 a_26123_n6178# a_26130_n6396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X930 vdd d0 a_20808_n3497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X931 a_734_7948# a_516_7948# a_243_7955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X932 a_26230_965# d0 a_26719_859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X933 a_26291_4237# d0 a_26772_4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X934 a_27492_n7750# a_27290_n6911# a_27414_n6911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X935 a_65_n9195# a_72_n9413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X936 a_15605_4152# d1 a_15691_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X937 a_22070_n9727# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X938 a_14293_n3856# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X939 a_33728_n8003# a_33985_n8019# a_32935_n7587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X940 a_716_7342# a_498_7342# a_241_7437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X941 gnd d0 a_21098_8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X942 gnd d0 a_33913_n3535# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X943 a_15474_n2485# d0 a_16267_n2901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X944 a_8993_8297# a_8999_8480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X945 a_7036_8609# d0 a_7838_8248# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X946 a_5805_3099# a_5587_3099# a_5007_3283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X947 a_18850_n7902# d4 a_18953_n5864# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X948 a_19920_1305# a_20173_1292# a_19834_2090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X949 a_15678_8224# a_15935_8034# a_15599_7031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X950 a_27373_n4698# a_27155_n4465# a_26575_n4649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X951 gnd d1 a_7256_6383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_27327_n8947# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X953 a_31482_n2442# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X954 a_499_n6648# a_281_n6648# a_18_n6359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X955 gnd d0 a_16832_8260# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X956 a_17399_n7171# d0 a_17888_n7266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X957 a_24117_n3678# d0 a_24919_n3306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X958 a_15388_n3281# d1 a_15470_n2673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X959 a_4573_n2177# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X960 gnd d1 a_33332_4384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X961 a_16575_8450# a_16579_8273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X962 vdd d1 a_28824_n7778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X963 a_9059_n8709# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X964 a_17634_n5230# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X965 a_5630_n4851# a_5424_n5459# a_4844_n5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X966 a_20845_8247# a_20840_8836# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X967 a_14329_n2663# d2 a_14412_n3679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X968 a_12142_4188# a_12137_4777# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X969 a_29582_8449# a_29839_8259# a_28784_8633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X970 gnd d2 a_2577_n5295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X971 a_9402_3901# a_9184_3901# a_8911_3908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X972 a_31882_n3868# a_31664_n3868# a_31783_n3691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X973 a_7654_n9590# a_7911_n9606# a_6856_n9774# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X974 a_298_n7666# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_11138_n9188# d1 a_11237_n9598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X976 a_1446_3615# a_1240_4104# a_661_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X977 a_6937_8199# a_7194_8009# a_6858_7006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X978 a_26260_2384# a_26265_2708# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X979 a_29332_n5766# a_29348_n6560# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X980 a_29316_n4336# a_29311_n4936# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X981 a_30940_n4250# a_30722_n4250# a_30449_n4056# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_31783_n3691# a_31581_n2852# a_31705_n2852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X983 a_6831_1914# d1 a_6926_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X984 a_30661_4433# a_30665_4951# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X985 a_5097_8373# a_4879_8373# a_4622_8468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X986 a_29364_n7990# a_29621_n8006# a_28571_n7574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X987 a_18684_8188# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X988 a_30920_n3232# a_30702_n3232# a_30431_n3137# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X989 gnd d0 a_16597_n6989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X990 a_10048_n3666# a_9846_n2827# a_9965_n2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X991 a_17380_n6054# a_17382_n6153# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X992 a_22178_n3619# d1 a_22964_n2827# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X993 a_11961_n5754# a_12214_n5958# a_11164_n5526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 a_17924_n9714# d1 a_18710_n8922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_15429_n5129# d1 a_15524_n5727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X996 a_133_1847# d0 a_624_1840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X997 a_2492_n9761# a_2749_n9777# a_2397_n9163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X998 a_28606_7030# d2 a_28685_8223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X999 vdd d0 a_33912_n3947# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1000 a_21790_n8420# a_21796_n8603# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1001 a_30548_n9463# d0 a_31029_n9752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1002 a_14619_7196# a_14401_7196# a_13821_7380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1003 a_20661_n9589# a_20918_n9605# a_19863_n9773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1004 vdd d1 a_33115_n3719# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1005 a_24407_8621# d0 a_25205_8437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1006 a_26340_7073# a_26347_7291# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1007 a_4495_1342# d0 a_4970_1247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1008 gnd d0 a_25407_5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1009 a_13641_n8722# a_13423_n8722# a_13160_n8433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1010 a_22216_n5243# a_21998_n5243# a_21727_n5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1011 gnd d0 a_34186_7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1012 a_17487_841# d0 a_17978_834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1013 a_13621_n7704# a_13403_n7704# a_13146_n7598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1014 gnd d8 a_17382_n10744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 a_3473_8647# a_3726_8634# a_2676_8419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 gnd d2 a_24348_n7356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1017 a_32796_n5329# d1 a_32882_n4533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1018 a_17316_n2299# a_17322_n2482# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1019 a_17322_n2482# a_17324_n3000# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1020 a_22160_3295# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1021 a_6750_n3478# d0 a_7543_n3894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1022 a_17575_5413# a_17577_5931# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1023 a_28715_4384# d0 a_29512_4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1024 a_6806_n6532# d0 a_7599_n6948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1025 a_25172_6224# a_25167_6813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1026 a_23031_7183# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1027 a_5676_n3831# a_5506_n4851# a_5625_n4674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1028 a_4568_5414# d0 a_5043_5319# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1029 a_22795_n5471# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1030 a_7526_n2876# a_7783_n2892# a_6733_n2460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1031 a_17798_n2176# d1 a_18595_n2637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1032 a_27254_n4875# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_4901_n8285# a_4683_n8285# a_4410_n8091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1034 gnd d1 a_2639_n3669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1035 a_32614_n6163# d3 a_32786_n8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1036 a_5460_n7495# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1037 a_32713_n4313# a_32970_n4329# a_32610_n6351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1038 a_20665_n9401# a_20660_n10001# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1039 a_16977_n2070# d0 a_17798_n2176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1040 a_1586_2476# a_1368_2476# a_1487_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1041 a_21581_184# a_23337_271# a_23461_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1042 a_26611_n6685# a_26393_n6685# a_26130_n6396# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 a_18812_6560# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1044 a_32790_5186# d3 a_32897_2971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1045 vdd d1 a_24591_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1046 a_25081_1546# a_25095_2329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1047 a_12692_n10677# d5 a_15181_n10603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1048 a_14329_n2663# a_14111_n2430# a_13532_n2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1049 a_1659_6548# d4 a_1726_365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1050 vdd d0 a_21098_8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1051 a_4429_n9208# a_4436_n9426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1052 a_16395_n9615# a_16399_n9427# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1053 a_17797_n2588# a_17579_n2588# a_17316_n2299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1054 vdd d1 a_7256_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1055 gnd d0 a_3529_n8987# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1056 a_n25_n4105# a_n18_n4323# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1057 a_28505_n9388# d1 a_28587_n8780# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1058 vdd d0 a_16832_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1059 a_5924_6561# d3 a_6023_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1060 a_28514_n4708# a_28771_n4724# a_28432_n5316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1061 a_25167_6813# a_25171_6636# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1062 a_5081_6943# a_4863_6943# a_4592_7049# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1063 a_29275_n2488# a_29279_n2300# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1064 vdd d1 a_33332_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1065 a_32914_n6757# a_33171_n6773# a_32832_n7365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1066 a_23120_n7915# d3 a_23214_n7915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1067 a_9364_2277# d1 a_10150_1604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1068 a_11993_n7978# a_11997_n7790# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1069 gnd d0 a_29729_2151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1070 a_4770_1853# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1071 a_16579_8273# a_16574_8862# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1072 gnd d0 a_29801_6635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1073 a_17596_n3606# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1074 a_480_n5630# a_262_n5630# a_n1_n5341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1075 a_83_n9920# a_3546_n10005# a_2496_n9573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1076 a_8709_n3513# a_8714_n4031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1077 a_18632_n4673# d2 a_18683_n3830# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1078 a_15181_n10603# a_15438_n10619# a_12692_n10677# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1079 a_24100_n2660# a_24357_n2676# a_24018_n3268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1080 a_3384_3145# a_3637_3132# a_2582_3506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1081 a_2618_5542# d0 a_3420_5181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1082 vdd d0 a_16778_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1083 a_31209_8410# d1 a_31995_7737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1084 a_11204_2103# d1 a_11290_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1085 a_19777_n4495# d0 a_20574_n4723# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1086 a_2573_8186# d1 a_2655_7578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1087 a_8244_n10653# d6 a_10916_n10590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1088 gnd d1 a_20190_2310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1089 a_11924_n3718# a_11941_n4512# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1090 a_6831_1914# d1 a_6930_2324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1091 a_31691_n8960# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1092 a_30902_n2626# a_30684_n2626# a_30421_n2337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1093 a_405_2252# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1094 a_15704_4562# d0 a_16506_4201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1095 a_17586_6248# d0 a_18067_6336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1096 gnd d3 a_2747_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1097 a_18936_6679# d3 a_19030_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_6674_n8348# a_6931_n8364# a_6502_n6126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1099 a_26355_7992# d0 a_26846_7985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1100 a_3289_n9989# a_83_n9920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1101 a_32882_n4533# d0 a_33675_n4949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1102 a_2442_n6519# a_2695_n6723# a_2356_n7315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1103 a_9221_n5655# d1 a_10007_n4863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 a_17777_1852# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1105 a_11417_8444# a_11670_8431# a_11318_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1106 a_28606_7030# d2 a_28689_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1107 a_5550_1063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1108 a_10145_1075# a_9927_1075# a_9348_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_17669_n7678# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1110 a_606_1234# a_388_1234# a_125_1146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1111 a_24280_1495# a_24537_1305# a_24198_2103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1112 gnd d7 a_8501_n10669# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1113 a_22198_n4637# a_21980_n4637# a_21717_n4348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 a_26347_7291# a_26353_7474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1115 vdd d0 a_34186_7254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1116 a_22178_n3619# a_21960_n3619# a_21703_n3513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1117 a_17850_5924# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1118 a_3469_8824# a_3726_8634# a_2676_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1119 a_3272_n8971# a_3276_n8783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1120 a_13711_1272# a_13493_1272# a_13230_1184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1121 a_30975_n6698# a_30757_n6698# a_30500_n6592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1122 a_26500_1271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1123 a_17924_n9714# a_17706_n9714# a_17449_n9608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1124 a_11945_n4324# a_12198_n4528# a_11143_n4696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1125 a_12018_n8396# a_12013_n8996# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1126 a_21943_6043# d0 a_22432_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1127 a_22033_n7691# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1128 vdd d2 a_15718_n7369# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1129 a_18557_1062# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1130 a_13104_n5379# a_13110_n5562# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1131 a_30203_209# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1132 a_21933_5243# d0 a_22414_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1133 a_22342_847# a_22124_847# a_21853_953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1134 a_22341_1259# d1 a_23139_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1135 a_9077_n9315# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1136 a_27553_6585# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1137 a_15645_6011# d1 a_15744_6421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1138 a_13785_4932# a_13567_4932# a_13294_4939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1139 a_24202_1926# d1 a_24297_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1140 a_17995_1852# a_17777_1852# a_17506_1958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1141 a_32041_6717# d3 a_32135_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1142 a_8806_n9220# d0 a_9295_n9315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 a_19830_n7549# d0 a_20623_n7965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1144 a_14308_2106# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1145 a_28349_n4300# d2 a_28399_n3092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1146 a_27446_n8770# a_27228_n8537# a_26649_n8309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1147 a_24901_n2700# a_25154_n2904# a_24104_n2472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1148 a_20606_n6947# a_20863_n6963# a_19813_n6531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1149 a_27414_n6911# a_27208_n7519# a_26628_n7703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1150 a_33639_n2501# a_33896_n2517# a_32841_n2685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1151 a_21860_1171# a_21866_1354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1152 a_22414_5331# d1 a_23212_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1153 a_28648_6187# d1 a_28734_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1154 a_14201_n7520# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1155 a_27694_n5889# a_27476_n5889# a_27591_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1156 a_22959_n2650# d2 a_23042_n3666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1157 a_5060_6337# a_4842_6337# a_4579_6249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1158 vdd d0 a_16651_n10043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1159 a_18705_n8745# d2 a_18756_n7902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1160 a_27298_1087# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1161 a_17125_n10728# d7 a_21421_n10664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1162 a_6674_n8348# d2 a_6724_n7140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1163 a_11127_n3490# d0 a_11924_n3718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1164 vdd d0 a_29586_n5558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1165 a_4880_n7679# a_4662_n7679# a_4405_n7573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1166 vdd d0 a_29729_2151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1167 vdd d0 a_29801_6635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1168 a_31844_2526# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1169 a_9039_n7691# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1170 a_2369_n2447# a_2622_n2651# a_2283_n3243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1171 a_24955_n5754# a_24971_n6548# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1172 a_6785_2934# a_7038_2921# a_6678_5149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1173 a_18775_1062# a_18557_1062# a_17977_1246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1174 a_3380_3322# a_3637_3132# a_2582_3506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1175 a_11340_4549# a_11597_4359# a_11245_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1176 a_14490_n7928# a_14320_n8948# a_14439_n8771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1177 a_28535_n5538# d0 a_29332_n5766# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1178 a_16340_n6973# a_16597_n6989# a_15547_n6557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1179 a_23099_n5877# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1180 a_26245_1884# a_26247_1983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1181 vdd d1 a_20190_2310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1182 a_24059_n5116# d1 a_24154_n5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1183 a_21690_n3112# a_21697_n3330# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1184 a_1721_246# d5 a_1820_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1185 a_21781_n8103# d0 a_22272_n8297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1186 a_3220_n5729# a_3236_n6523# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1187 gnd d2 a_6941_n5308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1188 vdd d2 a_2650_n9367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1189 a_31705_n2852# a_31499_n3460# a_30919_n3644# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1190 a_3453_7394# a_3710_7204# a_2655_7578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1191 a_14371_n4876# a_14165_n5484# a_13585_n5668# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1192 a_17851_n5642# a_17633_n5642# a_17376_n5536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1193 a_14707_284# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1194 a_6819_n7738# d0 a_7617_n7554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1195 a_1492_2595# a_1322_3496# a_1446_3615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1196 a_11413_8621# a_11670_8431# a_11318_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1197 a_16524_5631# a_16777_5618# a_15727_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1198 a_21960_n3619# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1199 a_22271_n8709# a_22053_n8709# a_21790_n8420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1200 vdd d2 a_24455_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1201 a_2599_4524# d0 a_3397_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1202 a_7600_n6536# a_7857_n6552# a_6802_n6720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1203 vdd d1 a_28914_1317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1204 a_24049_n8172# a_24302_n8376# a_23873_n6138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1205 a_389_822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1206 vdd d1 a_19993_n2663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1207 a_17093_n839# d9 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1208 a_30624_2397# d0 a_31099_2302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1209 a_16272_n2301# a_16525_n2505# a_15470_n2673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1210 a_4309_172# a_4091_172# a_4210_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1211 a_27492_n7750# a_27290_n6911# a_27409_n6734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1212 a_1043_n4428# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1213 gnd d0 a_3616_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1214 a_22070_n9727# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 a_13532_n2202# a_13314_n2202# a_13043_n2107# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1216 a_1133_n9518# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1217 a_28604_n9798# d0 a_29402_n9614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1218 a_14293_n3856# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1219 a_426_2858# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1220 a_258_8455# d0 a_733_8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1221 gnd d1 a_24484_n9802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1222 a_5024_4301# d1 a_5810_3628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1223 a_27373_n4698# a_27155_n4465# a_26576_n4237# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1224 a_32717_n4125# d2 a_32800_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1225 a_537_n8272# a_319_n8272# a_48_n8177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1226 a_27341_n2839# a_27135_n3447# a_26555_n3631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1227 gnd d0 a_16562_n4541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1228 a_20755_3157# a_21008_3144# a_19953_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1229 gnd d0 a_8091_8235# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1230 a_2241_n4075# d2 a_2320_n5279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1231 a_13331_n3220# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1232 a_6913_1306# a_7166_1293# a_6827_2091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1233 a_13531_2896# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1234 a_24202_1926# d1 a_24301_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1235 gnd d0 a_25388_4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1236 a_9964_3111# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1237 a_554_n9290# a_336_n9290# a_63_n9096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1238 a_13170_n9233# a_13177_n9451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1239 gnd d3 a_20118_6992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1240 a_336_n9290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1241 a_23103_2501# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1242 vdd d0 a_29785_5205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1243 a_24271_6175# d1 a_24357_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1244 gnd d1 a_29041_8443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1245 a_14221_n8538# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1246 a_26050_n2106# a_26057_n2324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1247 a_31783_n3691# a_31581_n2852# a_31700_n2675# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_27558_3652# d2 a_27604_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 a_5966_259# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1250 a_13530_3308# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1251 a_15415_n8373# d2 a_15461_n7353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1252 a_30920_n3232# a_30702_n3232# a_30429_n3038# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1253 a_16267_n2901# a_16524_n2917# a_15474_n2485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1254 a_10002_n4686# d2 a_10053_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1255 a_18504_n9530# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1256 a_30976_n6286# a_30758_n6286# a_30485_n6092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1257 a_426_n2576# d1 a_1224_n2625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1258 a_32895_n5739# d0 a_33693_n5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1259 a_30559_n9970# a_34022_n10055# a_32972_n9623# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1260 a_11055_5161# d3 a_11162_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1261 a_13838_8398# a_13620_8398# a_13357_8310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1262 a_644_2858# a_426_2858# a_155_2964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1263 gnd d4 a_24306_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1264 a_33676_n4537# a_33933_n4553# a_32878_n4721# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1265 gnd d2 a_2720_1888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1266 gnd d0 a_12430_6623# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1267 a_14597_2633# a_14427_3534# a_14546_3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1268 a_27434_3533# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1269 a_6930_2324# d0 a_7723_2729# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1270 a_30554_n9646# d0 a_31029_n9752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1271 a_3204_n4299# a_3457_n4503# a_2402_n4671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1272 a_16542_6237# a_16537_6826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1273 a_31810_n8783# a_31592_n8550# a_31013_n8322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1274 a_13838_8398# d1 a_14624_7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 a_20823_7818# a_21080_7628# a_20030_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1276 a_31778_n6924# a_31572_n7532# a_30992_n7716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1277 a_21943_6043# a_21950_6261# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1278 a_26828_7379# a_26610_7379# a_26347_7291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1279 a_21322_n10664# d5 a_23811_n10590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_22216_n5243# a_21998_n5243# a_21725_n5049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1281 a_24018_n3268# a_24275_n3284# a_23972_n4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1282 a_13621_n7704# a_13403_n7704# a_13140_n7415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1283 a_78_n9596# a_83_n9920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1284 a_29475_2576# a_29728_2563# a_28678_2348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1285 a_6854_7183# a_7111_6993# a_6682_4972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1286 a_500_n6236# d1 a_1297_n6697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1287 a_18377_n2404# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1288 a_24152_3123# a_24409_2933# a_24049_5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1289 gnd d3 a_33150_2958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1290 a_15502_n9201# d1 a_15597_n9799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1291 a_21980_n4637# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1292 a_29368_n7802# a_29385_n8596# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1293 a_24053_4984# d3 a_24225_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1294 vdd d0 a_33985_n8019# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1295 a_22795_n5471# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1296 a_19792_2933# d2 a_19871_4126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1297 gnd d0 a_16651_n10043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1298 a_17797_n2588# d1 a_18595_n2637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1299 gnd d0 a_7964_1109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1300 a_27591_n7927# a_27373_n7927# a_27497_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1301 a_2599_4524# d0 a_3401_4163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1302 a_23074_n8935# a_22868_n9543# a_22288_n9727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1303 vdd d0 a_7856_n6964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1304 gnd d2 a_20021_n9379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1305 a_17370_n5353# a_17376_n5536# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1306 vdd d0 a_20828_n4515# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1307 a_31798_3546# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1308 a_29548_6648# a_29801_6635# a_28751_6420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1309 a_516_7948# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1310 vdd d3 a_33043_n8401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1311 a_31880_1100# a_31662_1100# a_31083_872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1312 vdd d0 a_3616_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1313 a_13223_966# d0 a_13712_860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1314 a_14283_n6912# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1315 a_24919_n3306# a_25172_n3510# a_24117_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 vdd d1 a_28734_n2688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1317 a_4315_n2483# a_4317_n3001# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1318 a_20624_n7553# a_20881_n7569# a_19826_n7737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1319 a_2314_n8147# d2 a_2393_n9351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1320 a_24975_n6360# a_25228_n6564# a_24173_n6732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1321 a_11183_n6544# a_11436_n6748# a_11097_n7340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1322 a_17835_n4212# a_17617_n4212# a_17346_n4117# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1323 a_21944_n2189# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1324 gnd d1 a_2892_6370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1325 a_15744_6421# d0 a_16537_6826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1326 a_20550_n3893# a_20554_n3705# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1327 gnd d0 a_12341_1121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1328 a_21905_3908# a_21907_4007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1329 gnd d0 a_3509_n7969# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1330 a_443_n3594# a_225_n3594# a_n32_n3488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1331 a_31871_7618# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1332 a_20751_3334# a_21008_3144# a_19953_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1333 a_499_n6648# a_281_n6648# a_24_n6542# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1334 a_8930_4926# d0 a_9421_4919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1335 vdd d0 a_8091_8235# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1336 a_17871_n6248# d1 a_18668_n6709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1337 a_11277_6175# a_11534_5985# a_11231_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1338 a_8876_1971# d0 a_9365_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1339 vdd d0 a_8074_7217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1340 a_16362_n7391# a_16357_n7991# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1341 gnd d3 a_2567_n8351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1342 a_17634_n5230# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1343 a_9184_3901# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1344 a_28734_5402# d0 a_29527_5807# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1345 a_26611_6967# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1346 a_31882_n3868# a_31664_n3868# a_31788_n3868# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1347 a_19736_n2647# d0 a_20534_n2463# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1348 a_606_1234# d1 a_1404_1050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1349 a_4442_n9609# a_4447_n9933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1350 a_16469_2165# a_16722_2152# a_15667_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1351 vdd d1 a_29041_8443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1352 a_20533_n2875# a_20537_n2687# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1353 a_9147_1865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1354 a_5768_1063# d2 a_5851_2489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1355 a_32790_5186# a_33047_4996# a_32197_296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1356 a_29384_n9008# a_29641_n9024# a_28591_n8592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1357 a_22017_n6261# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1358 a_18087_7354# a_17869_7354# a_17612_7449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1359 a_30940_n4250# a_30722_n4250# a_30451_n4155# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1360 a_21914_4225# d0 a_22395_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1361 a_6858_7006# d2 a_6941_8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1362 a_19685_n8159# d2 a_19764_n9363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1363 a_5542_n6887# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1364 a_28652_6010# a_28905_5997# a_28602_7207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1365 a_13766_3914# a_13548_3914# a_13275_3921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1366 a_30063_n10689# d5 a_32552_n10615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1367 gnd d1 a_24610_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1368 a_17326_n3099# a_17333_n3317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1369 a_12141_4600# a_12394_4587# a_11344_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 vdd d0 a_12430_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1371 a_24970_n6960# a_25227_n6976# a_24177_n6544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1372 a_29459_1146# a_29712_1133# a_28657_1507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1373 a_6761_n9176# d1 a_6860_n9586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1374 vdd d0 a_33932_n4965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1375 a_4519_2977# a_4526_3195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1376 a_17925_n9302# d1 a_18710_n8922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1377 a_24173_n6732# d0 a_24975_n6360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1378 a_4791_n2177# a_4573_n2177# a_4302_n2082# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1379 a_20730_2728# a_20987_2538# a_19937_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1380 gnd d0 a_20987_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1381 a_16484_3772# a_16488_3595# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1382 a_21783_n8202# a_21790_n8420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1383 a_10255_7183# a_10037_7183# a_9457_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1384 a_32882_n4533# a_33135_n4737# a_32796_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1385 a_4769_2265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1386 a_7723_2729# a_7727_2552# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1387 a_1276_6140# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1388 a_11945_n4324# a_11940_n4924# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1389 a_22395_4313# d1 a_23181_3640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1390 vdd d0 a_7783_n2892# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1391 a_30975_6980# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1392 a_15650_1508# d0 a_16448_1324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1393 a_4419_n8408# d0 a_4900_n8697# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1394 a_9421_4919# a_9203_4919# a_8930_4926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1395 a_1339_n8910# d2 a_1385_n7890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1396 a_29471_2753# a_29728_2563# a_28678_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1397 a_32552_n10615# a_32809_n10631# a_30063_n10689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1398 a_33728_n8003# a_33732_n7815# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1399 a_17924_n9714# a_17706_n9714# a_17443_n9425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1400 a_16305_n4525# a_16309_n4337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1401 a_5805_6561# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1402 a_n12_n4506# a_n10_n5024# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1403 a_18853_5663# d2 a_18931_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1404 a_23317_n5877# a_24068_n10606# a_21322_n10664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1405 a_31120_2908# d1 a_31917_3136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1406 a_135_1946# a_142_2164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1407 a_9077_n9315# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1408 a_16524_5631# a_16538_6414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1409 a_22452_6955# d1 a_23249_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1410 a_4592_7049# a_4599_7267# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1411 a_9240_n6673# d1 a_10038_n6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1412 a_29544_6825# a_29801_6635# a_28751_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1413 a_8913_4007# a_8920_4225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1414 a_24227_n9786# a_24484_n9802# a_24132_n9188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1415 a_32759_n3293# d1 a_32841_n2685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1416 gnd d0 a_25192_n4528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1417 gnd d3 a_2494_n4279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1418 a_24229_7018# d2 a_24308_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1419 a_17344_n4018# a_17346_n4117# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1420 a_26517_2289# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1421 a_27631_7724# a_27425_8213# a_26846_7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1422 a_18586_n8922# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1423 a_14329_n2663# a_14111_n2430# a_13531_n2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1424 vdd d1 a_2892_6370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1425 a_6787_n5514# a_7040_n5718# a_6688_n5104# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 a_15744_6421# d0 a_16541_6649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1427 a_22964_n2827# d2 a_23042_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1428 vout a_17093_n839# a_17212_n839# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1429 vdd d0 a_12341_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1430 vdd d0 a_33969_n6589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1431 gnd d0 a_3710_7204# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1432 a_21956_6444# d0 a_22431_6349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1433 a_18710_n8922# d2 a_18756_n7902# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1434 vdd d4 a_6755_n6330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1435 a_16561_7667# a_16814_7654# a_15764_7439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1436 a_3436_6611# a_3453_7394# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1437 vdd d2 a_24492_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1438 a_24055_n5304# d1 a_24137_n4696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1439 a_480_n5630# a_262_n5630# a_5_n5524# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1440 a_6023_6561# a_5805_6561# a_5929_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1441 a_33753_n8421# a_33748_n9021# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1442 a_7600_n6536# a_7604_n6348# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1443 a_17994_2264# d1 a_18780_1591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1444 vdd d0 a_12414_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1445 a_20714_1298# a_20971_1108# a_19916_1482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1446 gnd d1 a_24374_n3694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1447 a_22054_n8297# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1448 a_16465_2342# a_16722_2152# a_15667_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1449 a_2467_1901# d1 a_2566_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1450 a_19834_2090# d1 a_19920_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1451 a_22234_n6673# a_22016_n6673# a_21759_n6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1452 gnd d1 a_2839_3316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1453 a_31691_n8960# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1454 a_20574_n4723# a_20827_n4927# a_19777_n4495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1455 vdd d2 a_20201_8008# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1456 a_9438_5937# a_9220_5937# a_8949_6043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1457 a_31995_7737# a_31789_8226# a_31210_7998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1458 a_21761_n7085# d0 a_22252_n7279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1459 a_8694_n3013# a_8696_n3112# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1460 a_6720_n7328# d1 a_6802_n6720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1461 a_22877_n4863# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1462 a_17851_n5642# a_17633_n5642# a_17370_n5353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1463 a_29455_1323# a_29712_1133# a_28657_1507# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1464 a_24975_n6360# a_24970_n6960# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1465 gnd d0 a_25264_n9012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1466 a_444_n3182# a_226_n3182# a_n47_n2988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1467 a_2672_8596# a_2929_8406# a_2577_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1468 a_7526_n2876# a_7530_n2688# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1469 a_11216_n8768# d0 a_12018_n8396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1470 a_22251_n7691# a_22033_n7691# a_21770_n7402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1471 a_30429_n3038# a_30431_n3137# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1472 vdd d0 a_7874_n7570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1473 a_30451_n4155# d0 a_30940_n4250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1474 a_20713_1710# a_20717_1533# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1475 a_30429_n3038# d0 a_30920_n3232# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1476 a_26736_1877# d1 a_27521_1616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1477 a_31119_3320# a_30901_3320# a_30638_3232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_30938_4944# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1479 a_27932_283# a_27714_283# a_27838_402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1480 a_6967_4360# a_7220_4347# a_6868_3950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1481 a_15650_1508# d0 a_16452_1147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1482 a_33839_2589# a_33856_3372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1483 a_3240_n6335# a_3235_n6935# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1484 a_8236_n2045# a_8679_n2094# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1485 a_8987_n4225# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1486 a_1023_n3410# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1487 a_13532_n2202# a_13314_n2202# a_12613_n2057# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1488 a_24154_n5714# a_24411_n5730# a_24059_n5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1489 a_9184_n3619# a_8966_n3619# a_8703_n3330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1490 gnd d1 a_2732_n8759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1491 a_15507_n4709# d0 a_16305_n4525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1492 a_733_8360# d1 a_1519_7687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1493 a_20644_n8571# a_20648_n8383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1494 a_189_4901# a_191_5000# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1495 a_28674_2525# d0 a_29472_2341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1496 gnd d3 a_15779_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1497 a_33928_7856# a_33932_7679# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1498 a_537_n8272# a_319_n8272# a_46_n8078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1499 a_14587_5689# a_14381_6178# a_13801_6362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1500 a_27341_n2839# a_27135_n3447# a_26556_n3219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1501 a_517_n7254# a_299_n7254# a_28_n7159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1502 gnd d0 a_16542_n3523# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1503 vdd d0 a_33896_n2517# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1504 a_15723_5580# d0 a_16525_5219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1505 a_1565_6667# a_1395_7568# a_1514_7158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1506 a_28468_n7352# d1 a_28554_n6556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1507 a_21462_184# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1508 gnd d0 a_25425_6211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1509 a_13567_4932# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1510 a_14402_n6735# a_14184_n6502# a_13604_n6686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1511 a_29586_8272# a_29839_8259# a_28784_8633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1512 a_27589_5159# a_27371_5159# a_26791_5343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1513 a_24229_7018# d2 a_24312_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1514 a_13605_n6274# a_13387_n6274# a_13116_n6179# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1515 a_7617_n7554# a_7621_n7366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1516 a_23011_6165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1517 a_9257_n7691# a_9039_n7691# a_8782_n7585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1518 gnd d3 a_7111_6993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1519 a_25168_6401# a_25172_6224# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1520 a_4412_n8190# d0 a_4901_n8285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1521 a_14201_n7520# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1522 a_10007_n4863# d2 a_10053_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1523 a_22141_1865# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1524 a_11101_n7152# a_11354_n7356# a_11051_n8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1525 gnd d0 a_3420_n2467# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1526 a_18050_5318# a_17832_5318# a_17569_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1527 a_11231_7195# a_11488_7005# a_11059_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1528 gnd d0 a_16635_n8613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1529 a_13221_867# a_13223_966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1530 a_33038_2538# a_33295_2348# a_32943_1951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1531 a_16557_7844# a_16814_7654# a_15764_7439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1532 a_15781_8457# a_16034_8444# a_15682_8047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1533 a_23254_7712# a_23048_8201# a_22468_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1534 a_1406_n3818# a_1188_n3818# a_1307_n3641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1535 a_4482_941# d0 a_4971_835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1536 a_3184_n3281# a_3437_n3485# a_2382_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1537 a_31778_n6924# a_31572_n7532# a_30993_n7304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1538 a_14490_n7928# a_14320_n8948# a_14444_n8948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1539 a_28771_7438# a_29024_7425# a_28685_8223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_30601_1196# d0 a_31082_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1541 a_23176_6573# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1542 a_9295_n9315# d1 a_10080_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1543 a_1079_n6464# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1544 vdd d1 a_2839_3316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1545 vdd d1 a_15744_n3707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1546 a_7816_7819# a_8073_7629# a_7023_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1547 a_1404_1050# d2 a_1487_2476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1548 a_30322_209# d6 a_26029_208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1549 a_15781_8457# d0 a_16574_8862# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1550 a_499_n6648# d1 a_1297_n6697# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1551 gnd d0 a_29605_n6576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1552 a_18377_n2404# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1553 gnd d0 a_3474_n5521# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 a_28535_n5538# a_28788_n5742# a_28436_n5128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1555 a_8967_6768# d0 a_9458_6955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1556 a_21980_n4637# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1557 a_21960_n3619# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1558 a_22271_n8709# a_22053_n8709# a_21796_n8603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1559 a_27591_n7927# a_27373_n7927# a_27492_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1560 a_7710_1534# a_7724_2317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1561 a_26338_6780# a_26340_7073# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1562 a_23074_n8935# a_22868_n9543# a_22289_n9315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1563 vdd d1 a_15854_n9815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1564 a_16447_1736# a_16451_1559# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1565 a_28771_7438# d0 a_29564_7843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1566 a_18777_n3830# a_18559_n3830# a_18678_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1567 a_28395_n3280# d1 a_28481_n2484# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1568 a_13080_n4143# a_13087_n4361# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1569 a_33892_5408# a_34149_5218# a_33094_5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1570 a_32800_n5141# a_33053_n5345# a_32717_n4125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 a_26147_n7414# d0 a_26628_n7703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1572 a_1043_n4428# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1573 a_14283_n6912# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1574 a_9204_n4637# a_8986_n4637# a_8729_n4531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1575 a_1133_n9518# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1576 a_17835_n4212# a_17617_n4212# a_17344_n4018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1577 gnd d1 a_24591_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1578 a_3179_n3881# a_3436_n3897# a_2386_n3465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1579 a_6651_n3068# d1 a_6750_n3478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1580 a_28674_2525# d0 a_29476_2164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1581 a_24918_n3718# a_24935_n4512# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1582 gnd d1 a_24574_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1583 a_23394_6573# a_23176_6573# a_23300_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1584 a_2138_n6113# d3 a_2310_n8335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1585 a_17870_n6660# d1 a_18668_n6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 a_9385_2883# a_9167_2883# a_8894_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 a_2237_n4263# a_2494_n4279# a_2134_n6301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1588 vdd d0 a_25425_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1589 a_4363_n5354# a_4369_n5537# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1590 a_31752_6190# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1591 a_13821_7380# a_13603_7380# a_13346_7475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1592 vdd d0 a_29604_n6988# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1593 a_1240_4104# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1594 gnd d0 a_7820_n4928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_10218_5147# d2 a_10301_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1596 a_6843_n8568# d0 a_7640_n8796# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1597 a_18705_n8745# a_18487_n8512# a_17907_n8696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1598 a_28436_n5128# d1 a_28535_n5538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1599 a_6827_2091# d1 a_6909_1483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1600 a_4555_5013# a_4562_5231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1601 a_22814_n6489# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1602 a_18667_7170# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1603 a_2618_5542# d0 a_3416_5358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1604 a_15687_3544# d0 a_16485_3360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1605 gnd d0 a_12197_n4940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_17908_n8284# a_17690_n8284# a_17419_n8189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1607 a_9384_3295# a_9166_3295# a_8909_3390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1608 a_22017_n6261# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1609 a_30682_5969# d0 a_31173_5962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1610 a_17629_8467# d0 a_18104_8372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1611 a_35_n7377# a_41_n7560# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1612 a_14417_n3856# a_14247_n4876# a_14371_n4876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1613 gnd d1 a_11400_n4712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1614 a_32202_415# a_32020_4560# a_32135_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1615 a_5081_6943# d1 a_5878_7171# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1616 a_20026_7590# a_20283_7400# a_19944_8198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1617 a_18504_n9530# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1618 a_3257_n7353# a_3510_n7557# a_2455_n7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1619 a_14514_1617# d2 a_14592_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1620 gnd d0 a_16704_1546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1621 a_4375_n6154# a_4382_n6372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1622 a_15777_8634# a_16034_8444# a_15682_8047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1623 a_25012_n8396# a_25007_n8996# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1624 a_282_n6236# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1625 a_21421_n10664# a_25872_n10681# a_17125_n10728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1626 a_19685_5148# d3 a_19792_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1627 a_10233_2620# a_10063_3521# a_10182_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1628 a_3383_3557# a_3397_4340# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1629 a_5098_7961# d1 a_5883_7700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1630 a_6766_n4684# d0 a_7564_n4500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1631 a_6688_n5104# a_6941_n5308# a_6605_n4088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1632 a_9474_8385# d1 a_10260_7712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1633 a_19608_n4275# a_19865_n4291# a_19505_n6313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1634 a_8787_n8103# a_8789_n8202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1635 a_32862_n3515# a_33115_n3719# a_32763_n3105# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1636 a_31810_n8783# a_31592_n8550# a_31012_n8734# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1637 a_28767_7615# a_29024_7425# a_28685_8223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1638 a_1215_n8910# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1639 a_252_8272# a_258_8455# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1640 a_3469_8824# a_3473_8647# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1641 a_28481_n2484# d0 a_29274_n2900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1642 a_4549_4396# a_4553_4914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1643 a_17813_4300# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1644 a_22996_n4686# a_22778_n4453# a_22198_n4637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1645 gnd d0 a_7963_1521# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1646 a_4399_n7390# d0 a_4880_n7679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1647 a_20030_7413# d0 a_20827_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1648 a_26100_n4543# d0 a_26575_n4649# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1649 a_17653_n6248# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1650 a_31100_1890# a_30882_1890# a_30609_1897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1651 a_15781_8457# d0 a_16578_8685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1652 a_9258_n7279# a_9040_n7279# a_8767_n7085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1653 a_4447_n9933# a_7910_n10018# a_6860_n9586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1654 a_5661_n6710# a_5443_n6477# a_4863_n6661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1655 a_26074_n3342# d0 a_26555_n3631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1656 a_30500_n6592# d0 a_30975_n6698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 a_4626_n5643# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1658 a_26280_3402# a_26282_3920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1659 a_21993_8480# d0 a_22468_8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1660 a_1060_n5446# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1661 a_12156_5795# a_12413_5605# a_11363_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1662 vdd d1 a_24447_n7766# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1663 a_21796_n8603# a_21798_n9121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1664 a_1358_5532# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1665 a_23181_3640# d2 a_23227_2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1666 a_6682_4972# d3 a_6858_7006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1667 a_29458_1558# a_29472_2341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1668 a_22162_n2189# a_21944_n2189# a_21243_n2044# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1669 a_11307_2336# d0 a_12100_2741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1670 a_8723_n4348# a_8729_n4531# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1671 a_32955_n8605# a_33208_n8809# a_32869_n9401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1672 a_16272_n2301# a_16267_n2901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1673 a_28771_7438# d0 a_29568_7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1674 a_30721_8104# d0 a_31210_7998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1675 a_9219_6349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1676 vdd d2 a_24312_n5320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1677 a_17363_n5135# a_17370_n5353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1678 a_23141_n3843# a_22923_n3843# a_23047_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1679 a_14345_4142# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1680 a_33148_8646# d0 a_33946_8462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1681 a_29544_6825# a_29548_6648# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1682 a_30624_2397# a_30629_2721# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1683 a_17370_n5353# d0 a_17851_n5642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1684 a_25136_4188# a_25131_4777# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1685 a_6770_n4496# d0 a_7567_n4724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1686 a_18586_n8922# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1687 vdd d0 a_29549_n3522# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1688 a_2417_3098# d2 a_2463_2078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1689 a_11380_6408# d0 a_12173_6813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1690 a_12161_5206# a_12156_5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1691 a_9475_7973# a_9257_7973# a_8986_8079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1692 a_6440_n10578# d4 a_6502_n6126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1693 vdd d1 a_24574_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1694 a_30728_8322# d0 a_31209_8410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1695 a_4842_6337# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1696 a_27335_3123# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_32918_n6569# d0 a_33711_n6985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1698 a_22235_n6261# d1 a_23032_n6722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1699 a_30919_3926# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1700 a_30680_5451# a_30682_5969# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1701 a_23130_7593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1702 a_25192_7242# a_25187_7831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1703 a_1544_4510# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1704 a_24022_n3080# d1 a_24117_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1705 a_31856_n7763# a_31654_n6924# a_31778_n6924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1706 a_17526_2976# a_17533_3194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1707 a_30975_6980# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1708 a_15687_3544# d0 a_16489_3183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1709 vdd d2 a_28869_3961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1710 a_11344_4372# a_11597_4359# a_11245_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_30475_n5391# d0 a_30956_n5680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1712 a_33839_2589# a_34092_2576# a_33042_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1713 a_11940_n4924# a_11944_n4736# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1714 a_6860_n9586# a_7113_n9790# a_6761_n9176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_25171_6636# a_25424_6623# a_24374_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1716 a_32869_n9401# d1 a_32955_n8605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1717 a_22234_n6673# a_22016_n6673# a_21753_n6384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1718 a_7707_1299# a_7964_1109# a_6909_1483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1719 a_24214_n8580# d0 a_25007_n8996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1720 vdd d0 a_16704_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1721 gnd d1 a_15924_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1722 a_5732_2489# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1723 a_22877_n4863# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1724 a_5851_2489# a_5649_1473# a_5773_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1725 a_32197_296# d4 a_32794_5009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1726 a_30974_7392# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1727 a_23120_n7915# a_22950_n8935# a_23074_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1728 a_31699_3136# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1729 a_n55_n2287# a_n49_n2470# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1730 a_2490_7170# d2 a_2540_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1731 gnd d0 a_25244_n7994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_11196_n7750# d0 a_11998_n7378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1733 a_32078_296# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1734 a_21813_n9621# a_21818_n9945# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1735 a_30431_n3137# d0 a_30920_n3232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1736 a_17759_1246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1737 a_11231_7195# d2 a_11277_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1738 a_14597_2633# d3 a_14691_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1739 a_3252_n7953# a_3256_n7765# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1740 gnd d1 a_28914_1317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1741 a_20571_n4499# a_20575_n4311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1742 a_4499_1959# d0 a_4988_1853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1743 a_2393_n9351# d1 a_2475_n8743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 a_21860_1171# d0 a_22341_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1745 a_11286_1495# d0 a_12084_1311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1746 a_15346_n4113# d2 a_15429_n5129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1747 a_8987_n4225# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1748 vdd d0 a_7963_1521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1749 a_30629_2721# d0 a_31120_2908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1750 a_9203_4919# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1751 a_9222_n5243# a_9004_n5243# a_8733_n5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1752 a_19948_8021# d1 a_20047_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1753 a_31772_7208# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1754 a_8967_n3207# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1755 a_22234_6955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1756 a_1334_n8733# d2 a_1385_n7890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1757 a_7580_n5930# a_7584_n5742# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1758 a_26327_6273# d0 a_26808_6361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1759 gnd d1 a_2712_n7741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1760 vdd d0 a_16541_n3935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1761 a_15487_n3691# d0 a_16285_n3507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1762 a_26593_n5255# d1 a_27378_n4875# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1763 a_517_n7254# a_299_n7254# a_26_n7060# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1764 a_24198_2103# d1 a_24280_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1765 a_8343_n10653# d7 a_4050_n10652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1766 a_15346_n4113# a_15599_n4317# a_15239_n6339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_11307_2336# d0 a_12104_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1768 a_9801_n5471# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1769 a_27599_2513# a_27397_1497# a_27516_1087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1770 a_9857_n8525# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1771 a_14402_n6735# a_14184_n6502# a_13605_n6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1772 a_24275_5998# a_24528_5985# a_24225_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1773 a_14649_4548# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1774 a_33148_8646# d0 a_33950_8285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1775 a_31917_3136# a_31699_3136# a_31119_3320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1776 a_25082_1134# a_25335_1121# a_24280_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1777 a_26808_6361# d1 a_27594_5688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1778 a_14546_6586# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1779 a_25607_n2057# d0 a_26539_n2201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1780 a_13605_n6274# a_13387_n6274# a_13114_n6080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1781 a_30466_n5074# a_30468_n5173# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1782 a_24271_6175# d1 a_24353_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1783 a_15580_n8781# d0 a_16378_n8597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1784 a_11380_6408# d0 a_12177_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1785 a_14364_5160# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1786 a_1820_246# a_1602_246# a_1726_365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1787 a_15419_5174# a_15676_4984# a_14826_284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1788 a_13333_7074# a_13340_7292# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1789 a_3277_n8371# a_3272_n8971# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1790 gnd d0 a_16615_n7595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1791 a_31990_7208# a_31772_7208# a_31192_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1792 a_24173_n6732# a_24430_n6748# a_24091_n7340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1793 a_206_5919# d0 a_697_5912# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1794 a_11940_n4924# a_12197_n4940# a_11147_n4508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1795 a_31120_2908# a_30902_2908# a_30629_2721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1796 a_33749_n8609# a_33753_n8421# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1797 a_15392_n3093# d1 a_15491_n3503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1798 a_20827_7641# a_21080_7628# a_20030_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1799 a_33835_2766# a_34092_2576# a_33042_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1800 a_33049_8236# d1 a_33135_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1801 a_9294_n9727# d1 a_10080_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1802 a_1079_n6464# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1803 a_25167_6813# a_25424_6623# a_24374_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1804 a_28472_n7164# a_28725_n7368# a_28422_n8372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1805 a_2419_n5689# d0 a_3217_n5505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1806 a_29275_n2488# a_29532_n2504# a_28477_n2672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1807 vdd d1 a_20173_1292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1808 a_26160_n8214# d0 a_26649_n8309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1809 vdd d1 a_15924_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1810 a_23811_n10590# d4 a_23869_n6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1811 a_717_6930# d1 a_1514_7158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1812 a_26111_n5378# a_26117_n5561# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1813 a_2500_4114# a_2757_3924# a_2421_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1814 a_32786_n8385# d2 a_32836_n7177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1815 a_26301_4938# d0 a_26792_4931# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1816 a_24914_n3906# a_24918_n3718# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1817 a_1334_n8733# a_1116_n8500# a_537_n8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1818 a_4480_842# a_4482_941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1819 a_624_1840# a_406_1840# a_133_1847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1820 a_30449_n4056# d0 a_30940_n4250# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1821 gnd d0 a_3599_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1822 a_1582_n5852# a_1364_n5852# a_1479_n7890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1823 vdd d0 a_16614_n8007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1824 vdd d2 a_7084_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1825 a_11286_1495# d0 a_12088_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1826 a_4534_3896# a_4536_3995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1827 a_23037_n6899# a_22831_n7507# a_22251_n7691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1828 a_2655_7578# d0 a_3453_7394# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1829 a_26153_n7597# d0 a_26628_n7703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1830 a_22213_6349# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1831 a_6926_2501# d0 a_7728_2140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1832 a_5007_3283# d1 a_5805_3099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1833 a_13050_n2325# d0 a_13531_n2614# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1834 a_9204_n4637# a_8986_n4637# a_8723_n4348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1835 vdd d3 a_2674_2908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1836 a_9168_n2189# d1 a_9965_n2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1837 a_8236_n2045# a_7527_n2464# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1838 a_24357_5390# d0 a_25154_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1839 a_1023_n3410# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1840 a_30680_5451# d0 a_31155_5356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1841 a_18068_5924# d1 a_18853_5663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1842 a_9184_n3619# a_8966_n3619# a_8709_n3513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1843 vdd d3 a_15672_n8389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1844 a_4622_8468# a_3473_8647# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1845 a_17815_n3194# a_17597_n3194# a_17324_n3000# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1846 gnd d3 a_11415_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1847 gnd d0 a_3547_n9593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1848 a_24049_n8172# d2 a_24132_n9188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1849 a_2639_6383# a_2892_6370# a_2540_5973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1850 a_19777_n4495# a_20030_n4699# a_19691_n5291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1851 a_13350_8092# d0 a_13839_7986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1852 gnd d0 a_8074_7217# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1853 a_25078_1311# a_25335_1121# a_24280_1495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1854 a_18705_n8745# a_18487_n8512# a_17908_n8284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1855 a_31137_3926# a_30919_3926# a_30648_4032# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1856 a_6823_n7550# d0 a_7620_n7778# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1857 a_10982_n4100# d2 a_11061_n5304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1858 a_18953_n5864# a_18735_n5864# a_18850_n7902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1859 a_19790_n5701# d0 a_20592_n5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1860 a_4302_n2082# a_4309_n2300# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1861 a_27698_2513# a_27480_2513# a_27599_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1862 a_24939_n4324# a_24934_n4924# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1863 a_26340_7073# d0 a_26829_6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1864 a_21243_n2044# a_21673_n2094# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1865 a_17888_n7266# a_17670_n7266# a_17399_n7171# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1866 a_4828_n4213# d1 a_5625_n4674# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1867 a_13357_8310# d0 a_13838_8398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1868 a_13110_n5562# d0 a_13585_n5668# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1869 a_14417_n3856# a_14247_n4876# a_14366_n4699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1870 a_16394_n10027# a_13188_n9958# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1871 a_33696_n5779# a_33949_n5983# a_32899_n5551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1872 a_22431_6349# a_22213_6349# a_21956_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1873 a_3397_4340# a_3401_4163# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1874 a_26501_859# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1875 a_32845_n2497# a_33098_n2701# a_32759_n3293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1876 a_20827_7641# a_20841_8424# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1877 a_31210_7998# a_30992_7998# a_30721_8104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1878 a_25008_n8584# a_25265_n8600# a_24210_n8768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1879 a_282_n6236# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1880 a_28608_n9610# d0 a_26195_n9957# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1881 a_13821_7380# d1 a_14619_7196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1882 a_1406_n3818# a_1188_n3818# a_1312_n3818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1883 a_7019_7591# a_7276_7401# a_6937_8199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1884 a_20734_2551# a_20987_2538# a_19937_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1885 a_15682_8047# d1 a_15777_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1886 a_4050_n10652# d6 a_2175_n10565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1887 gnd d1 a_28788_n5742# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1888 a_26247_1983# a_26254_2201# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1889 gnd d2 a_7014_n9380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1890 a_28509_n9200# d1 a_28608_n9610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1891 a_29455_1323# a_29459_1146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1892 a_1313_8176# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1893 a_1261_n4661# a_1043_n4428# a_464_n4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1894 a_30648_4032# a_30655_4250# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1895 a_26357_n4649# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1896 a_15419_5174# d3 a_15522_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1897 a_19695_n5103# d1 a_19794_n5513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1898 a_6605_n4088# a_6858_n4292# a_6498_n6314# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1899 a_22996_n4686# a_22778_n4453# a_22199_n4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1900 a_21961_6768# a_21963_7061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1901 vdd d1 a_15764_n4725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1902 gnd d1 a_11543_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1903 a_22964_n2827# a_22758_n3435# a_22178_n3619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1904 a_24095_n7152# d1 a_24194_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1905 a_9457_7367# a_9239_7367# a_8976_7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1906 a_29351_n6784# a_29365_n7578# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1907 a_4388_n6555# a_4390_n7073# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1908 a_5878_7171# d2 a_5929_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1909 a_5661_n6710# a_5443_n6477# a_4864_n6249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 a_26080_n3525# d0 a_26555_n3631# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1911 a_28685_8223# d1 a_28767_7615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1912 a_30522_n8128# d0 a_31013_n8322# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1913 a_4626_n5643# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1914 a_1060_n5446# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1915 a_21581_184# d6 a_21680_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1916 a_32020_4560# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1917 a_7023_7414# d0 a_7820_7642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1918 a_23976_n4100# d2 a_24059_n5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1919 gnd d0 a_25155_n2492# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 a_17543_3994# d0 a_18032_3888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1921 a_27833_283# d4 a_28430_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1922 a_464_n4200# a_246_n4200# a_n25_n4105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1923 gnd d1 a_2819_2298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1924 a_18549_n6886# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1925 a_32899_n5551# d0 a_33696_n5779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1926 a_18777_n3830# a_18559_n3830# a_18683_n3830# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1927 a_23141_n3843# a_22923_n3843# a_23042_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1928 a_6806_n6532# a_7059_n6736# a_6720_n7328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1929 vdd d5 a_2333_n10581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1930 a_17376_n5536# d0 a_17851_n5642# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1931 a_33929_7444# a_33933_7267# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1932 a_11127_n3490# a_11380_n3694# a_11028_n3080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1933 a_17562_5012# a_17569_5230# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1934 a_3199_n4899# a_3456_n4915# a_2406_n4483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1935 vdd d3 a_24229_n4304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1936 a_1519_7687# a_1313_8176# a_733_8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1937 a_2635_6560# a_2892_6370# a_2540_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1938 gnd d1 a_33225_n9827# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1939 a_9385_2883# d1 a_10182_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1940 a_8759_n6384# a_8765_n6567# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1941 a_6498_n6314# d3 a_6605_n4088# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1942 a_17399_n7171# a_17406_n7389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1943 a_17376_n5536# a_17380_n6054# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1944 a_12017_n8808# a_12270_n9012# a_11220_n8580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1945 a_8909_3390# a_8911_3908# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1946 a_1565_6667# d3 a_1659_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1947 a_31856_n7763# a_31654_n6924# a_31773_n6747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 a_4590_6756# d0 a_5081_6943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1949 a_3180_n3469# a_3184_n3281# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1950 a_8866_1171# d0 a_9347_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1951 a_10075_n8758# d2 a_10126_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1952 a_31172_6374# a_30954_6374# a_30691_6286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1953 a_19871_4126# a_20128_3936# a_19792_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1954 a_24394_7426# d0 a_25187_7831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1955 a_17556_4395# a_17560_4913# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1956 a_3277_n8371# a_3530_n8575# a_2475_n8743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1957 a_10150_1604# d2 a_10228_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1958 a_24194_n7562# d0 a_24987_n7978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1959 a_21763_n7184# a_21770_n7402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1960 a_16561_7667# a_16575_8450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1961 a_30524_n8227# a_30531_n8445# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1962 a_9747_n2417# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1963 a_24914_n3906# a_25171_n3922# a_24121_n3490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1964 a_32931_n7775# d0 a_33733_n7403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1965 a_23120_n7915# a_22950_n8935# a_23069_n8758# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1966 a_4309_n2300# d0 a_4790_n2589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1967 a_16502_4378# a_16759_4188# a_15704_4562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1968 gnd d2 a_15935_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1969 a_24297_2513# d0 a_25099_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1970 a_5878_7171# a_5660_7171# a_5080_7355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1971 a_31995_7737# d2 a_32041_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1972 a_11925_n3306# a_11920_n3906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1973 vdd d3 a_20045_2920# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1974 a_15682_8047# d1 a_15781_8457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1975 a_23873_n6138# d3 a_24045_n8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1976 a_17612_7449# a_17614_7967# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1977 a_19654_n3255# d1 a_19736_n2647# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1978 a_26254_2201# a_26260_2384# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1979 a_32062_2526# a_31844_2526# a_31968_2645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1980 a_32970_7043# a_33223_7030# a_32794_5009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1981 a_7748_3158# a_7743_3747# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1982 a_30655_4250# a_30661_4433# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1983 a_5883_7700# a_5677_8189# a_5097_8373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1984 a_26846_7985# a_26628_7985# a_26355_7992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1985 a_20010_6395# a_20263_6382# a_19911_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1986 a_1215_n8910# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1987 a_16285_n3507# a_16289_n3319# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1988 a_2360_n7127# d1 a_2455_n7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1989 a_9222_n5243# a_9004_n5243# a_8731_n5049# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1990 a_20790_5605# a_20804_6388# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1991 a_8967_n3207# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1992 a_9278_n8297# a_9060_n8297# a_8787_n8103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1993 gnd d6 a_12949_n10693# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 a_26094_n4360# d0 a_26575_n4649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1995 a_28685_8223# d1 a_28771_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1996 a_17653_n6248# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1997 vdd d3 a_28786_2945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1998 a_19740_n2459# d0 a_20537_n2687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1999 a_9944_2093# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 vdd d1 a_24467_n8784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2001 a_18850_n7902# a_18632_n7902# a_18756_n7902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2002 a_16448_1324# a_16452_1147# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2003 a_6941_8022# d1 a_7040_8432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2004 a_13236_1367# d0 a_13711_1272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2005 a_5081_6943# a_4863_6943# a_4590_6756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2006 a_28751_6420# a_29004_6407# a_28652_6010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2007 a_26845_8397# a_26627_8397# a_26370_8492# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2008 a_9420_5331# d1 a_10218_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2009 a_21680_n2312# d0 a_22161_n2601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2010 a_204_5401# d0 a_679_5306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2011 a_9801_n5471# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2012 vdd d3 a_24302_n8376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2013 a_9857_n8525# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2014 a_17324_n3000# a_17326_n3099# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2015 a_27626_7195# a_27408_7195# a_26829_6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2016 a_30739_n5268# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2017 a_21781_n8103# a_21783_n8202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2018 a_26050_n2106# d0 a_26539_n2201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2019 vdd d2 a_11391_n9392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2020 a_14390_1498# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2021 a_5924_6561# a_5722_5545# a_5841_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2022 a_13309_5439# d0 a_13784_5344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2023 a_29316_n4336# a_29569_n4540# a_28514_n4708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2024 a_15560_n7763# d0 a_16358_n7579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2025 a_7567_n4724# a_7820_n4928# a_6770_n4496# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2026 a_26282_3920# d0 a_26773_3913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2027 a_16285_n3507# a_16542_n3523# a_15487_n3691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2028 a_19830_n7549# a_20083_n7753# a_19731_n7139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2029 a_13170_n9233# d0 a_13659_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2030 a_17832_5318# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2031 a_6502_n6126# a_6755_n6330# a_6440_n10578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2032 a_33042_2361# a_33295_2348# a_32943_1951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2033 a_23048_8201# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2034 a_26245_1884# d0 a_26736_1877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2035 a_4585_6432# d0 a_5060_6337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2036 a_26612_n6273# d1 a_27409_n6734# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2037 a_13363_8493# a_12214_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2038 a_21717_n4348# a_21723_n4531# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2039 a_33098_5415# a_33351_5402# a_33012_6200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2040 a_31029_n9752# d1 a_31815_n8960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2041 a_6729_n2648# d0 a_7531_n2276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2042 a_10343_271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2043 vdd d2 a_11461_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2044 a_22250_8385# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2045 a_23869_n6326# d3 a_23972_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2046 gnd d5 a_28445_n10618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2047 a_24394_7426# d0 a_25191_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2048 a_11106_n2660# d0 a_11908_n2288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2049 a_1259_5122# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2050 a_9023_n6261# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2051 a_7820_7642# a_8073_7629# a_7023_7414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2052 a_33042_2361# d0 a_33835_2766# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2053 a_15543_n6745# d0 a_16341_n6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2054 vdd d2 a_15935_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2055 a_28514_n4708# d0 a_29316_n4336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2056 vdd d1 a_7166_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2057 vdd d4 a_24126_n6342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2058 a_5851_2489# d3 a_5950_2489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2059 a_5098_7961# a_4880_7961# a_4609_8067# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2060 a_15564_n7575# d0 a_16361_n7803# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2061 vdd d1 a_24394_n4712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2062 a_9364_2277# a_9146_2277# a_8889_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2063 a_3470_8412# a_3474_8235# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2064 a_11134_n9376# a_11391_n9392# a_11055_n8172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2065 a_1302_n6874# a_1096_n7482# a_517_n7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2066 a_1409_1579# a_1203_2068# a_624_1840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2067 a_1582_n5852# a_1364_n5852# a_1406_n3818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2068 a_19933_2500# d0 a_20731_2316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2069 a_1441_3086# d2 a_1492_2595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2070 a_30903_n2214# d1 a_31700_n2675# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2071 a_32966_7220# a_33223_7030# a_32794_5009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2072 a_20006_6572# a_20263_6382# a_19911_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2073 a_23037_n6899# a_22831_n7507# a_22252_n7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2074 a_32968_n9811# d0 a_33770_n9439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2075 a_19861_7182# d2 a_19907_6162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2076 a_20624_n7553# a_20628_n7365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2077 a_15243_n6151# d3 a_15419_n8185# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2078 a_33896_5231# a_34149_5218# a_33094_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2079 a_13056_n2508# d0 a_13531_n2614# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2080 a_2492_n9761# d0 a_3290_n9577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2081 a_9167_n2601# d1 a_9965_n2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2082 a_26320_6055# a_26327_6273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2083 a_3217_n5505# a_3474_n5521# a_2419_n5689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2084 a_28575_2115# a_28832_1925# a_28529_3135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2085 a_4988_1853# a_4770_1853# a_4497_1860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2086 a_15429_n5129# a_15682_n5333# a_15346_n4113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2087 a_10109_2501# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2088 gnd d0 a_7910_n10018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2089 a_8932_5025# a_8939_5243# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2090 a_2314_5136# d3 a_2417_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2091 a_11277_6175# d1 a_11363_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2092 gnd d0 a_25408_5193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2093 a_4480_842# a_7707_1299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2094 gnd d2 a_33089_n7381# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2095 a_3474_8235# a_3727_8222# a_2672_8596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2096 a_1477_5122# a_1259_5122# a_679_5306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2097 a_3290_n9577# a_3294_n9389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2098 a_19757_n3477# a_20010_n3681# a_19658_n3067# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2099 a_11281_5998# d1 a_11380_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2100 gnd d0 a_12160_n2904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2101 vdd d0 a_29642_n8612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2102 a_10285_4535# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2103 a_28711_4561# d0 a_29513_4200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2104 a_7531_n2276# a_7526_n2876# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2105 a_18673_n6886# a_18467_n7494# a_17888_n7266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2106 a_5407_n4441# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2107 a_18953_n5864# a_18735_n5864# a_18777_n3830# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2108 a_13367_n5668# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2109 a_5768_1063# a_5550_1063# a_4971_835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2110 vdd d1 a_15980_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2111 a_17888_n7266# a_17670_n7266# a_17397_n7072# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2112 a_4827_n4625# d1 a_5625_n4674# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2113 a_13728_2290# a_13510_2290# a_13247_2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2114 a_11055_5161# a_11312_4971# a_10462_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2115 a_4808_n3195# d1 a_5593_n2815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2116 a_10223_5676# a_10017_6165# a_9438_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2117 a_696_6324# a_478_6324# a_215_6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2118 a_26029_208# a_30203_209# a_27932_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2119 a_14473_2514# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2120 a_3216_n5917# a_3220_n5729# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2121 a_1224_n2625# a_1006_n2392# a_426_n2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2122 a_11196_n7750# a_11453_n7766# a_11101_n7152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2123 a_24988_n7566# a_25245_n7582# a_24190_n7750# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2124 a_4317_n3001# d0 a_4808_n3195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2125 a_22123_1259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2126 a_15511_n4521# d0 a_16308_n4749# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2127 a_24370_6585# a_24627_6395# a_24275_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2128 vdd d6 a_21579_n10680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2129 a_19957_3341# d0 a_20750_3746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2130 a_26718_1271# a_26500_1271# a_26237_1183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2131 a_32897_2971# d2 a_32980_3987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2132 a_15181_n10603# d4 a_15243_n6151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2133 a_13801_6362# a_13583_6362# a_13320_6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2134 a_15425_n5317# d1 a_15511_n4521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2135 a_8872_1354# a_8874_1872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2136 a_26590_6361# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2137 a_31861_n7940# d3 a_31955_n7940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2138 gnd d1 a_28771_n4724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2139 a_18957_2488# d4 a_19097_377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2140 a_22950_n8935# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2141 a_23222_2501# a_23020_1485# a_23139_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2142 a_9060_n8297# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2143 a_17541_3895# a_17543_3994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2144 a_10467_390# a_10285_4535# a_10400_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2145 gnd d3 a_6931_n8364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2146 a_22964_n2827# a_22758_n3435# a_22179_n3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2147 a_26102_n5061# d0 a_26593_n5255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2148 a_20030_7413# d0 a_20823_7818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2149 a_9240_n6673# a_9022_n6673# a_8765_n6567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2150 a_33042_2361# d0 a_33839_2589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2151 a_22431_6349# d1 a_23217_5676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2152 a_26158_n8115# d0 a_26649_n8309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2153 a_30524_n8227# d0 a_31013_n8322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2154 a_26791_5343# a_26573_5343# a_26310_5255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2155 a_30502_n7110# d0 a_30993_n7304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2156 a_19809_n6719# d0 a_20611_n6347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2157 gnd d3 a_11308_n8376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2158 a_24991_n7790# a_25008_n8584# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2159 a_31029_n9752# a_30811_n9752# a_30554_n9646# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2160 a_9883_n4863# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2161 a_14624_7725# d2 a_14670_6705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2162 a_26104_n5160# a_26111_n5378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2163 a_1479_n7890# a_1261_n7890# a_1385_n7890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2164 a_14826_284# d4 a_15419_5174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2165 a_23295_6573# a_23093_5557# a_23212_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2166 a_13060_n3125# a_13067_n3343# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2167 a_17577_5931# d0 a_18068_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2168 a_4375_n6154# d0 a_4864_n6249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2169 a_13311_5957# a_13313_6056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2170 a_19933_2500# d0 a_20735_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2171 a_31742_n4888# d2 a_31788_n3868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2172 vdd d0 a_3419_n2879# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2173 a_31083_872# a_30865_872# a_30592_879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2174 vdd d0 a_16634_n9025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2175 a_14691_2514# a_14473_2514# a_14597_2633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2176 gnd d2 a_2830_7996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2177 a_15584_n8593# a_15837_n8797# a_15498_n9389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2178 a_30954_6374# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2179 a_29369_n7390# a_29364_n7990# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2180 a_23321_2501# d4 a_23461_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2181 a_32873_n9213# d1 a_32968_n9811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2182 vdd d0 a_12377_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2183 a_12951_197# a_14707_284# a_14826_284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2184 a_18853_5663# a_18647_6152# a_18067_6336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2185 a_3470_8412# a_3727_8222# a_2672_8596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2186 a_17580_n2176# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2187 a_607_822# a_389_822# a_118_928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2188 a_11997_n7790# a_12250_n7994# a_11200_n7562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2189 a_2421_2921# d2 a_2500_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2190 a_10080_n8935# d2 a_10126_n7915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2191 gnd d0 a_3493_n6539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2192 a_28554_n6556# a_28807_n6760# a_28468_n7352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2193 vdd d1 a_2676_n5705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2194 a_33732_n7815# a_33985_n8019# a_32935_n7587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2195 a_20592_n5329# a_20845_n5533# a_19790_n5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2196 a_9401_4313# d1 a_10187_3640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2197 a_19546_n10577# d5 a_18953_n5864# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2198 a_2442_n6519# d0 a_3235_n6935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 a_13104_n5379# d0 a_13585_n5668# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2200 a_442_4288# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2201 a_32832_n7365# d1 a_32918_n6569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2202 a_21980_8079# a_21987_8297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2203 a_9747_n2417# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2204 a_17487_841# a_20714_1298# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2205 vdd d1 a_29004_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2206 a_9457_7367# d1 a_10255_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2207 a_17760_834# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2208 a_12031_n9602# a_12288_n9618# a_11233_n9786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2209 a_19957_3341# d0 a_20754_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2210 a_21851_854# a_21853_953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2211 vdd d2 a_11281_n3284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2212 a_15727_5403# a_15980_5390# a_15641_6188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2213 a_13290_4421# d0 a_13765_4326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2214 a_17796_3282# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2215 a_22359_1865# a_22141_1865# a_21868_1872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2216 a_516_7948# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2217 a_4827_n4625# a_4609_n4625# a_4352_n4519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2218 a_13326_6457# a_13331_6781# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2219 a_1261_n4661# a_1043_n4428# a_463_n4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2220 a_19944_8198# d1 a_20026_7590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2221 a_26357_n4649# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2222 vdd d3 a_7038_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2223 a_30882_1890# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2224 gnd d4 a_32867_n6367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2225 a_498_7342# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2226 a_24128_n9376# d1 a_24214_n8580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2227 a_16326_n5355# a_16579_n5559# a_15524_n5727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2228 a_26538_2895# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2229 a_5587_3099# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2230 a_19948_8021# d1 a_20043_8608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2231 a_21776_n7585# a_21781_n8103# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2232 a_19764_n9363# a_20021_n9379# a_19685_n8159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2233 a_30537_n8628# a_30539_n9146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2234 a_7003_6396# a_7256_6383# a_6904_5986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2235 a_26280_3402# d0 a_26755_3307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2236 a_13621_7986# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2237 a_10916_n10590# d5 a_10323_n5877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2238 a_13547_4326# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2239 a_18850_n7902# a_18632_n7902# a_18751_n7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2240 a_8932_5025# d0 a_9421_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2241 a_4549_4396# d0 a_5024_4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2242 a_33079_4397# a_33332_4384# a_32980_3987# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2243 a_5929_6680# a_5759_7581# a_5883_7700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2244 a_18683_n3830# a_18513_n4850# a_18632_n4673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2245 a_21686_n2495# d0 a_22161_n2601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_13641_n8722# d1 a_14439_n8771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2247 a_4373_n6055# a_4375_n6154# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2248 gnd d0 a_12178_n3510# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2249 a_13748_3308# a_13530_3308# a_13267_3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2250 a_9184_3901# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2251 a_15595_7208# a_15852_7018# a_15423_4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2252 a_23115_n7738# a_22913_n6899# a_23032_n6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2253 a_24059_n5116# a_24312_n5320# a_23976_n4100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2254 a_26611_6967# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2255 a_26537_3307# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2256 a_13620_8398# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2257 a_18032_3888# a_17814_3888# a_17541_3895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2258 a_28432_n5316# a_28689_n5332# a_28353_n4112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2259 a_4572_n2589# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2260 vdd d2 a_11498_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2261 a_11363_5390# d0 a_12156_5795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2262 a_11980_n6772# a_11994_n7566# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2263 a_32832_n7365# a_33089_n7381# a_32786_n8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2264 a_29569_7254# a_29564_7843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2265 a_29296_n3318# a_29549_n3522# a_28494_n3690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_26228_866# d0 a_26719_859# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2267 gnd d0 a_20790_n2891# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2268 a_14401_7196# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 gnd d0 a_3617_2114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2270 a_18031_4300# a_17813_4300# a_17556_4395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2271 a_30794_n8734# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2272 gnd d0 a_34005_n9037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2273 gnd d6 a_30320_n10705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2274 a_17217_n720# d9 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2275 vdd d1 a_7203_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2276 a_2369_n2447# d0 a_3162_n2863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2277 a_31609_n9568# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2278 a_26611_n6685# d1 a_27409_n6734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2279 a_15524_n5727# d0 a_16326_n5355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2280 a_21680_184# d7 a_17148_133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2281 a_24308_8211# d1 a_24390_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2282 gnd d1 a_7096_n8772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2283 a_3432_6788# a_3436_6611# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2284 a_24104_n2472# d0 a_24897_n2888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2285 a_12125_3170# a_12120_3759# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2286 a_27677_6704# a_27507_7605# a_27626_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2287 a_18812_3098# a_18594_3098# a_18015_2870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2288 a_29315_n4748# a_29329_n5542# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2289 a_5728_n5865# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2290 a_25154_5618# a_25407_5605# a_24357_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2291 a_23456_271# d4 a_24053_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2292 a_9820_n6489# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2293 a_9168_n2189# a_8950_n2189# a_8679_n2094# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2294 a_33049_8236# d1 a_33131_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2295 a_7800_6624# a_7817_7407# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2296 gnd d0 a_25389_4175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2297 a_17361_n5036# a_17363_n5135# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2298 a_26243_1366# a_26245_1884# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2299 a_30644_3415# a_30646_3933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2300 vdd d2 a_11354_n7356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2301 a_9023_n6261# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2302 gnd d0 a_20844_n5945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2303 a_n18_n4323# d0 a_463_n4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2304 a_7760_4765# a_7764_4588# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2305 a_2494_6993# d2 a_2577_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2306 gnd d0 a_8054_6199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2307 a_1446_3615# a_1240_4104# a_660_4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2308 a_2562_2488# a_2819_2298# a_2467_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2309 a_32951_n8793# d0 a_33753_n8421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2310 a_21807_n9438# d0 a_22288_n9727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2311 a_20537_n2687# a_20551_n3481# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2312 a_13531_2896# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2313 a_20551_n3481# a_20555_n3293# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2314 a_29312_n4524# a_29316_n4336# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2315 a_14412_n3679# d3 a_14511_n3856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2316 a_15526_2959# d2 a_15609_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2317 a_26448_n9327# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2318 vdd d0 a_16652_n9631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2319 a_1368_2476# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2320 a_30902_n2626# d1 a_31700_n2675# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2321 gnd d0 a_12431_6211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2322 a_4302_n2082# d0 a_4791_n2177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2323 a_8740_n5366# d0 a_9221_n5655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2324 a_6926_2501# d0 a_7724_2317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2325 a_15572_1939# a_15825_1926# a_15522_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2326 a_10002_n4686# a_9784_n4453# a_9204_n4637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2327 a_6999_6573# a_7256_6383# a_6904_5986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2328 a_17454_n9932# a_20917_n10017# a_19867_n9585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2329 a_4489_1159# d0 a_4970_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2330 a_33835_2766# a_33839_2589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2331 a_1487_2476# a_1285_1460# a_1404_1050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2332 a_32759_n3293# a_33016_n3309# a_32713_n4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2333 a_23337_271# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2334 a_27516_1087# d2 a_27599_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2335 a_25155_5206# a_25150_5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2336 a_28587_n8780# d0 a_29389_n8408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2337 a_33075_4574# a_33332_4384# a_32980_3987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2338 a_10978_n4288# d2 a_11024_n3268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2339 a_696_6324# d1 a_1482_5651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2340 a_29476_2164# a_29729_2151# a_28674_2525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2341 a_22840_n2827# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2342 vdd d0 a_29622_n7594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2343 a_4562_5231# d0 a_5043_5319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2344 gnd d0 a_7838_n5534# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2345 a_16521_5396# a_16778_5206# a_15723_5580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2346 gnd d0 a_3709_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2347 gnd d0 a_20881_n7569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2348 a_30739_n5268# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2349 a_5407_n4441# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2350 gnd d1 a_15781_n5743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2351 a_5387_n3423# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2352 a_26772_4325# a_26554_4325# a_26291_4237# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2353 gnd d0 a_12215_n5546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2354 a_3257_n7353# a_3252_n7953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2355 a_15502_n9201# a_15755_n9405# a_15419_n8185# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2356 a_1586_2476# a_1368_2476# a_1492_2595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2357 a_2494_6993# a_2747_6980# a_2318_4959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2358 a_9438_5937# a_9220_5937# a_8947_5944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2359 a_30704_7086# a_30711_7304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2360 a_29549_6236# a_29802_6223# a_28747_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2361 a_4807_n3607# d1 a_5593_n2815# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2362 a_10075_n8758# a_9857_n8525# a_9277_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2363 vdd d0 a_3617_2114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2364 a_13168_n9134# d0 a_13659_n9328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2365 a_33729_n7591# a_33733_n7403# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2366 a_3236_n6523# a_3493_n6539# a_2438_n6707# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2367 a_24308_8211# d1 a_24394_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2368 a_19681_n8347# d2 a_19731_n7139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2369 a_17575_5413# d0 a_18050_5318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2370 a_388_1234# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2371 a_15740_6598# d0 a_16538_6414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2372 a_11908_n2288# a_12161_n2492# a_11106_n2660# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2373 a_24987_n7978# a_24991_n7790# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2374 a_31030_n9340# d1 a_31815_n8960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2375 a_4845_n5231# a_4627_n5231# a_4356_n5136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2376 a_26375_n5255# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2377 a_22950_n8935# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2378 vdd d0 a_25389_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2379 a_28430_4996# d3 a_28606_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2380 a_13493_1272# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2381 a_13311_5957# d0 a_13802_5950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2382 vdd d0 a_25372_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2383 a_26104_n5160# d0 a_26593_n5255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2384 a_461_5306# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2385 a_23249_7183# a_23031_7183# a_22452_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2386 a_4881_n7267# d1 a_5666_n6887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2387 vdd d0 a_7837_n5946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2388 vdd d2 a_19911_n3271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2389 a_20750_3746# a_20754_3569# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2390 a_31210_7998# d1 a_31995_7737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2391 a_9240_n6673# a_9022_n6673# a_8759_n6384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2392 a_10978_n4288# a_11235_n4304# a_10875_n6326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2393 a_5640_6153# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2394 a_5950_2489# a_5732_2489# a_5851_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2395 a_30504_n7209# d0 a_30993_n7304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2396 a_31029_n9752# a_30811_n9752# a_30548_n9463# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 vdd d0 a_12214_n5958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2398 a_9883_n4863# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2399 a_33770_n9439# a_34023_n9643# a_32968_n9811# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2400 vdd d1 a_7040_n5718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2401 a_31618_n4888# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2402 a_15584_n8593# d0 a_16381_n8821# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2403 a_7023_7414# d0 a_7816_7819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2404 a_2237_n4263# d2 a_2287_n3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2405 a_18088_6942# a_17870_6942# a_17599_7048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2406 a_30646_3933# a_30648_4032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2407 a_21905_3908# d0 a_22396_3901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2408 a_13567_4932# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2409 gnd d1 a_11580_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2410 vdd d1 a_11417_n5730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2411 a_17777_1852# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2412 a_26666_n9327# d1 a_27451_n8947# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2413 a_10145_1075# a_9927_1075# a_9347_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2414 a_12142_4188# a_12395_4175# a_11340_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2415 vdd d0 a_12431_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2416 a_606_1234# a_388_1234# a_131_1329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2417 a_680_4894# a_462_4894# a_189_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2418 gnd d0 a_20988_2126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2419 gnd d2 a_20164_5972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2420 a_15564_n7575# a_15817_n7779# a_15465_n7165# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2421 a_6783_n5702# d0 a_7585_n5330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2422 gnd d0 a_20808_n3497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2423 gnd d1 a_11653_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2424 a_5625_n7903# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2425 a_13711_1272# a_13493_1272# a_13236_1367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2426 a_15708_4385# a_15961_4372# a_15609_3975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2427 a_28498_n3502# d0 a_29295_n3730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2428 a_25095_2329# a_25099_2152# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2429 a_26665_n9739# a_26447_n9739# a_26184_n9450# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2430 a_10038_n6722# d2 a_10121_n7738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2431 a_29472_2341# a_29729_2151# a_28674_2525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2432 a_11158_3123# d2 a_11208_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2433 gnd d2 a_28905_5997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2434 gnd d0 a_29765_4599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2435 a_18557_1062# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2436 vdd d2 a_2613_n7331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2437 a_3163_n2451# a_3420_n2467# a_2365_n2635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2438 a_24117_n3678# d0 a_24915_n3494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2439 vdd d0 a_3709_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2440 a_2324_n5091# d1 a_2423_n5501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2441 a_19608_n4275# d2 a_19658_n3067# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2442 a_22342_847# d1 a_23139_1075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2443 a_24919_n3306# a_24914_n3906# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2444 a_8909_3390# d0 a_9384_3295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2445 a_14764_6586# a_14546_6586# a_14665_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2446 a_18915_4522# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2447 a_28698_3366# a_28951_3353# a_28612_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2448 a_18751_n7725# d3 a_18850_n7902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2449 a_13340_7292# d0 a_13821_7380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2450 gnd d1 a_28824_n7778# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2451 a_13367_n5668# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2452 a_30957_n5268# d1 a_31742_n4888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2453 a_31193_6980# a_30975_6980# a_30704_7086# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2454 a_32968_n9811# a_33225_n9827# a_32873_n9213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2455 a_24154_n5714# d0 a_24956_n5342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2456 a_29545_6413# a_29802_6223# a_28747_6597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2457 a_6839_n8756# a_7096_n8772# a_6757_n9364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2458 a_11138_n9188# d1 a_11233_n9786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 a_19685_5148# a_19942_4958# a_19092_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2460 a_1322_3496# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2461 a_8969_7061# d0 a_9458_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2462 a_28529_3135# d2 a_28575_2115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2463 a_22415_4919# d1 a_23212_5147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2464 a_31209_8410# a_30991_8410# a_30728_8322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2465 a_11216_n8768# a_11473_n8784# a_11134_n9376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2466 a_24198_2103# a_24455_1913# a_24152_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2467 vdd d5 a_19704_n10593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2468 a_5060_6337# a_4842_6337# a_4585_6432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2469 a_21680_184# a_21462_184# a_19191_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2470 a_15740_6598# d0 a_16542_6237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2471 a_14509_1088# a_14291_1088# a_13711_1272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2472 a_3419_5593# a_3433_6376# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2473 a_24297_2513# d0 a_25095_2329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2474 vdd d0 a_3546_n10005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2475 a_4827_n4625# a_4609_n4625# a_4346_n4336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2476 a_10187_3640# d2 a_10233_2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2477 a_16562_7255# a_16815_7242# a_15760_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2478 a_30487_n6191# a_30494_n6409# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2479 a_2496_n9573# a_2749_n9777# a_2397_n9163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2480 a_3203_n4711# a_3217_n5505# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2481 gnd d0 a_33912_n3947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2482 a_4807_n3607# a_4589_n3607# a_4332_n3501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2483 a_31844_2526# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2484 a_3363_2539# a_3616_2526# a_2566_2311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2485 a_31856_n7763# d3 a_31955_n7940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2486 a_24353_5567# d0 a_25151_5383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2487 a_61_n8578# d0 a_536_n8684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2488 a_15511_n4521# a_15764_n4725# a_15425_n5317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2489 a_28730_5579# d0 a_29532_5218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2490 a_20665_n9401# a_20918_n9605# a_19863_n9773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2491 a_6937_8199# d1 a_7019_7591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2492 a_28529_3135# a_28786_2945# a_28426_5173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2493 vdd d0 a_25282_n9618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2494 a_4553_4914# a_4555_5013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2495 a_18067_6336# a_17849_6336# a_17586_6248# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2496 a_26316_5438# a_26318_5956# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2497 a_7653_n10002# a_4447_n9933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2498 a_32796_n5329# d1 a_32878_n4721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2499 a_4512_2360# a_4517_2684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2500 a_10462_271# d4 a_11055_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2501 a_6941_8022# d1 a_7036_8609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2502 a_21708_n4031# d0 a_22199_n4225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2503 a_5552_n3831# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2504 a_30611_1996# d0 a_31100_1890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2505 gnd d1 a_11363_n2676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2506 a_21950_6261# a_21956_6444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2507 a_3343_1286# a_3347_1109# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2508 vdd d1 a_11580_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2509 vdd d0 a_34075_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2510 a_4373_n6055# d0 a_4864_n6249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2511 gnd d0 a_16814_7654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2512 a_13621_n7704# d1 a_14407_n6912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2513 a_24231_n9598# d0 a_21818_n9945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2514 a_18751_n7725# a_18549_n6886# a_18668_n6709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2515 a_19865_7005# a_20118_6992# a_19689_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2516 a_12138_4365# a_12395_4175# a_11340_4549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2517 a_4610_n4213# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2518 a_7530_n2688# a_7783_n2892# a_6733_n2460# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2519 a_155_2964# d0 a_644_2858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2520 vdd d0 a_20988_2126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2521 a_10136_7593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2522 vdd d1 a_20120_n9789# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2523 a_5588_n2638# d2 a_5671_n3654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2524 a_30618_2214# d0 a_31099_2302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2525 a_30684_6068# d0 a_31173_5962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2526 a_4309_172# a_4091_172# a_1820_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2527 vdd d1 a_11653_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2528 a_26320_n2613# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2529 a_15704_4562# a_15961_4372# a_15609_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2530 a_26117_n5561# a_26121_n6079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2531 a_2397_n9163# d1 a_2496_n9573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2532 a_426_2858# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2533 a_24053_4984# a_24306_4971# a_23456_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2534 a_30794_n8734# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2535 a_8984_7980# a_8986_8079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2536 a_6766_n4684# a_7023_n4700# a_6684_n5292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2537 a_25099_2152# a_25094_2741# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2538 a_14427_3534# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2539 a_5025_3889# d1 a_5810_3628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2540 a_30774_n7716# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2541 gnd d0 a_33985_n8019# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2542 a_20660_n10001# a_20917_n10017# a_19867_n9585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2543 gnd d1 a_24411_n5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2544 a_19863_n9773# d0 a_20665_n9401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2545 a_22414_5331# a_22196_5331# a_21933_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2546 a_10875_n6326# a_11132_n6342# a_10817_n10590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2547 a_11162_2946# d2 a_11241_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 a_31099_2302# d1 a_31885_1629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2549 a_11998_n7378# a_11993_n7978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2550 a_11143_n4696# a_11400_n4712# a_11061_n5304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2551 vdd d1 a_2929_8406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2552 a_28694_3543# a_28951_3353# a_28612_4151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2553 a_5728_n5865# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2554 a_6688_n5104# d1 a_6783_n5702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2555 a_32918_n6569# a_33171_n6773# a_32832_n7365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2556 vdd d0 a_25154_n2904# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2557 a_11051_n8360# d2 a_11101_n7152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2558 a_31155_5356# d1 a_31953_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2559 a_8806_n9220# a_8813_n9438# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2560 a_6963_4537# d0 a_7761_4353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2561 a_14500_7606# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2562 a_26649_n8309# a_26431_n8309# a_26158_n8115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2563 a_n12_n4506# d0 a_463_n4612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2564 a_6090_378# d5 a_4210_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2565 a_30667_5050# a_30674_5268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2566 a_11307_2336# a_11560_2323# a_11208_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2567 a_25171_6636# a_25188_7419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2568 a_18031_4300# d1 a_18817_3627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2569 a_208_6018# a_215_6236# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2570 a_8244_n10653# d6 a_12692_n10677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2571 a_27553_3123# d2 a_27604_2632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2572 a_21813_n9621# d0 a_22288_n9727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2573 a_15597_n9799# d0 a_16399_n9427# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2574 gnd d0 a_29659_n9630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2575 a_19768_n9175# d1 a_19867_n9585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2576 a_6678_n8160# a_6931_n8364# a_6502_n6126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2577 a_29333_n5354# a_29328_n5954# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2578 a_14417_n3856# d3 a_14511_n3856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2579 vdd d1 a_2622_n2651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2580 a_24239_3962# a_24492_3949# a_24156_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2581 a_28616_3974# d1 a_28711_4561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2582 a_26448_n9327# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2583 a_18863_2607# a_18693_3508# a_18812_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2584 a_16558_7432# a_16815_7242# a_15760_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2585 a_21818_n9945# a_25281_n10030# a_24231_n9598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2586 a_31662_1100# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2587 a_3359_2716# a_3616_2526# a_2566_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2588 a_2573_8186# d1 a_2659_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2589 a_14597_2633# a_14427_3534# a_14551_3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2590 a_13548_n3632# d1 a_14334_n2840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2591 gnd d1 a_24664_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2592 a_8746_n5549# d0 a_9221_n5655# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2593 a_29495_3594# a_29509_4377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2594 a_17426_n8407# d0 a_17907_n8696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2595 a_13839_7986# d1 a_14624_7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2596 a_10002_n4686# a_9784_n4453# a_9205_n4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2597 a_29388_n8820# a_29641_n9024# a_28591_n8592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2598 a_31737_n4711# a_31519_n4478# a_30940_n4250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2599 a_9475_7973# a_9257_7973# a_8984_7980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2600 a_26828_7379# a_26610_7379# a_26353_7474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2601 a_9970_n2827# a_9764_n3435# a_9184_n3619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2602 gnd d3 a_24482_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2603 a_11277_6175# d1 a_11359_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2604 gnd d0 a_16721_2564# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2605 vdd d2 a_33196_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2606 a_28567_n7762# d0 a_29369_n7390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2607 a_7817_7407# a_8074_7217# a_7019_7591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2608 a_26167_n8432# a_26173_n8615# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2609 a_18683_n3830# a_18513_n4850# a_18637_n4850# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2610 a_26829_6967# d1 a_27626_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2611 a_13642_n8310# d1 a_14439_n8771# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2612 a_15777_8634# d0 a_16575_8450# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2613 vdd d0 a_16814_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2614 a_31536_n5496# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2615 a_22840_n2827# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2616 gnd d2 a_15718_n7369# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2617 a_25114_3759# a_25371_3569# a_24321_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2618 a_4543_4213# a_4549_4396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2619 a_2076_n10565# a_2333_n10581# a_2175_n10565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2620 a_4319_n3100# a_4326_n3318# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2621 a_9474_8385# a_9256_8385# a_8999_8480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2622 a_5024_4301# a_4806_4301# a_4543_4213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2623 vdd d0 a_16525_n2505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2624 a_28422_n8372# a_28679_n8388# a_28250_n6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2625 gnd d1 a_20066_n6735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2626 a_11160_n5714# d0 a_11958_n5530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2627 gnd d0 a_29711_1545# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2628 a_5387_n3423# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2629 a_12137_4777# a_12141_4600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2630 a_32202_415# d5 a_30322_209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2631 a_28767_7615# d0 a_29565_7431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2632 a_21888_2696# a_21890_2989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2633 a_10075_n8758# a_9857_n8525# a_9278_n8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2634 a_20610_n6759# a_20863_n6963# a_19813_n6531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2635 a_10043_n6899# a_9837_n7507# a_9257_n7691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2636 a_33675_n4949# a_33679_n4761# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2637 a_27594_5688# d2 a_27672_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2638 vdd d4 a_19762_n6329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2639 a_717_6930# a_499_6930# a_228_7036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2640 a_22913_n6899# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2641 a_31609_n9568# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2642 a_21976_7462# a_21978_7980# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2643 a_27172_n5483# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2644 a_661_3876# a_443_3876# a_170_3883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2645 gnd d0 a_8053_6611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2646 a_17125_n10728# d7 a_25615_n10665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2647 gnd d0 a_7911_n9606# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2648 a_32858_n3703# d0 a_33660_n3331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2649 a_6674_n8348# d2 a_6720_n7328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2650 vdd d2 a_33126_n9417# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2651 a_8874_1872# d0 a_9365_1865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2652 a_4845_n5231# a_4627_n5231# a_4354_n5037# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2653 gnd d0 a_29586_n5558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2654 a_26375_n5255# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2655 a_30631_3014# d0 a_31120_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2656 a_13822_6968# a_13604_6968# a_13333_7074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2657 a_19846_n8755# a_20103_n8771# a_19764_n9363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2658 a_6963_4537# d0 a_7765_4176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2659 a_9203_4919# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2660 a_22234_6955# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2661 a_3343_1286# a_3600_1096# a_2545_1470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2662 a_14490_n7928# d3 a_14584_n7928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2663 a_11164_n5526# d0 a_11961_n5754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2664 a_33131_7628# a_33388_7438# a_33049_8236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2665 a_28535_n5538# d0 a_29328_n5954# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2666 a_11303_2513# a_11560_2323# a_11208_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2667 a_660_4288# a_442_4288# a_185_4383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2668 a_16344_n6785# a_16597_n6989# a_15547_n6557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2669 a_29311_n4936# a_29568_n4952# a_28518_n4520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2670 a_6860_n9586# d0 a_7653_n10002# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2671 a_19916_1482# d0 a_20714_1298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2672 a_9385_2883# a_9167_2883# a_8896_2989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2673 a_11065_n5116# d1 a_11164_n5526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2674 a_14402_n6735# d2 a_14485_n7751# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2675 a_5703_n8923# a_5497_n9531# a_4917_n9715# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2676 gnd d2 a_2650_n9367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2677 a_11944_n4736# a_11958_n5530# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2678 a_28616_3974# d1 a_28715_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2679 vdd d0 a_3457_n4503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2680 gnd d0 a_16705_1134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2681 a_2463_2078# a_2720_1888# a_2417_3098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2682 a_26665_n9739# d1 a_27451_n8947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2683 a_13569_n4238# d1 a_14366_n4699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2684 vdd d1 a_24664_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2685 a_7604_n6348# a_7857_n6552# a_6802_n6720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2686 a_148_2347# d0 a_623_2252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2687 a_27425_8213# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 a_17851_n5642# d1 a_18637_n4850# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2689 a_28349_n4300# a_28606_n4316# a_28246_n6338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2690 gnd d1 a_19993_n2663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2691 a_17093_n839# d9 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2692 vdd d0 a_7910_n10018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2693 a_22396_3901# d1 a_23181_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2694 gnd d0 a_12377_3569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_5625_n7903# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2696 gnd d2 a_7157_5973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2697 a_27341_n2839# d2 a_27419_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2698 a_11941_n4512# a_11945_n4324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2699 vdd d0 a_16721_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2700 vdd d0 a_12287_n10030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2701 a_29274_n2900# a_29278_n2712# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2702 a_2310_n8335# d2 a_2360_n7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2703 a_30812_n9340# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2704 a_8244_n10653# a_8501_n10669# a_8343_n10653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2705 a_13568_n4650# a_13350_n4650# a_13087_n4361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2706 a_33949_8697# a_33639_n2501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2707 a_208_6018# d0 a_697_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2708 gnd d2 a_33233_3974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2709 a_15777_8634# d0 a_16579_8273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2710 a_30322_209# a_32078_296# a_32202_415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2711 a_16488_3595# a_16502_4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2712 a_8686_n2312# d0 a_9167_n2601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2713 a_13260_3002# a_13267_3220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2714 a_5805_6561# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2715 a_15650_1508# a_15907_1318# a_15568_2116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2716 vdd d4 a_2571_4946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2717 a_32717_n4125# d2 a_32796_n5329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2718 a_12157_5383# a_12414_5193# a_11359_5567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2719 a_18848_5134# d2 a_18931_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2720 vdd d1 a_7059_n6736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2721 a_10228_2501# a_10026_1485# a_10150_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2722 vdd d0 a_29711_1545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2723 gnd d1 a_28931_2335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2724 a_18756_n7902# d3 a_18850_n7902# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2725 vdd d0 a_25172_n3510# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2726 a_13313_6056# d0 a_13802_5950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2727 a_16574_8862# a_16578_8685# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2728 vdd d1 a_11436_n6748# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2729 vdd d0 a_25228_n6564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2730 vdd d0 a_7980_2539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2731 a_28767_7615# d0 a_29569_7254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2732 a_31789_8226# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2733 a_4753_835# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2734 a_17419_n8189# d0 a_17908_n8284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2735 a_6819_n7738# a_7076_n7754# a_6724_n7140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2736 a_27631_7724# a_27425_8213# a_26845_8397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2737 a_10561_271# d6 a_8658_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2738 a_7581_n5518# a_7585_n5330# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2739 a_2496_n9573# d0 a_83_n9920# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2740 a_26303_5037# d0 a_26792_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2741 a_8950_n2189# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2742 vdd d0 a_25388_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2743 a_30685_n2214# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2744 a_11376_6585# d0 a_12174_6401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2745 a_21950_6261# d0 a_22431_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2746 a_13728_2290# d1 a_14514_1617# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2747 vdd d0 a_8053_6611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2748 a_30719_8005# d0 a_31210_7998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2749 a_318_n8684# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2750 a_13110_n5562# a_13114_n6080# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2751 a_27694_n5889# a_28445_n10618# a_28287_n10602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2752 a_23139_1075# d2 a_23222_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2753 a_33680_n4349# a_33933_n4553# a_32878_n4721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2754 a_2586_3329# d0 a_3379_3734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2755 a_4807_n3607# a_4589_n3607# a_4326_n3318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2756 a_7761_4353# a_7765_4176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2757 a_13784_5344# d1 a_14582_5160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2758 a_6787_n5514# d0 a_7580_n5930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2759 a_24275_5998# d1 a_24370_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 gnd d1 a_33278_1330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2761 a_24974_n6772# a_24988_n7566# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2762 a_24956_n5342# a_24951_n5942# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2763 a_15526_2959# a_15779_2946# a_15419_5174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2764 a_18630_5134# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2765 a_13330_n3632# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2766 a_28587_n8780# a_28844_n8796# a_28505_n9388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2767 a_11024_n3268# d1 a_11106_n2660# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2768 a_24022_n3080# a_24275_n3284# a_23972_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2769 a_33840_2177# a_34093_2164# a_33038_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2770 a_22395_4313# a_22177_4313# a_21914_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2771 a_30976_n6286# d1 a_31773_n6747# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2772 a_2659_7401# d0 a_3452_7806# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2773 a_1395_7568# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 a_5060_6337# d1 a_5846_5664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2775 a_31995_7737# a_31789_8226# a_31209_8410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2776 a_21710_n4130# d0 a_22199_n4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2777 a_5552_n3831# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2778 a_17669_n7678# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2779 a_25172_6224# a_25425_6211# a_24370_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2780 a_13129_n6580# d0 a_13604_n6686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2781 a_32763_n3105# d1 a_32858_n3703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2782 a_21688_n3013# d0 a_22179_n3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2783 vdd d0 a_16705_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2784 a_3221_n5317# a_3216_n5917# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2785 vdd d1 a_33135_n4737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2786 a_31137_3926# a_30919_3926# a_30646_3933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2787 a_15599_7031# a_15852_7018# a_15423_4997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2788 a_4610_n4213# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2789 a_5469_n2815# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2790 a_33836_2354# a_33840_2177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2791 gnd d0 a_7856_n6964# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2792 a_20844_8659# a_21097_8646# a_20047_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2793 a_16325_n5767# a_16341_n6561# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2794 a_31917_6598# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2795 a_31193_6980# a_30975_6980# a_30702_6793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2796 a_30975_n6698# a_30757_n6698# a_30494_n6409# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2797 a_10053_n3843# a_9883_n4863# a_10007_n4863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2798 a_30865_872# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2799 a_22216_n5243# d1 a_23001_n4863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2800 a_5593_n2815# d2 a_5671_n3654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2801 gnd d0 a_20828_n4515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2802 a_31761_1510# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2803 a_22272_n8297# d1 a_23069_n8758# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2804 a_26320_n2613# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2805 gnd d0 a_12233_n6976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2806 gnd d3 a_33043_n8401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2807 a_32895_n5739# a_33152_n5755# a_32800_n5141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2808 a_17426_n8407# a_17432_n8590# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2809 a_4412_n8190# a_4419_n8408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2810 a_17432_n8590# a_17434_n9108# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2811 a_22994_5147# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2812 gnd d1 a_28734_n2688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2813 a_20628_n7365# a_20881_n7569# a_19826_n7737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2814 vdd d0 a_7964_1109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2815 a_32610_n6351# a_32867_n6367# a_32552_n10615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2816 a_734_7948# d1 a_1519_7687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2817 a_3204_n4299# a_3199_n4899# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2818 a_26665_n9739# a_26447_n9739# a_26190_n9633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2819 a_5480_n8513# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2820 a_30774_n7716# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2821 a_6746_n3666# a_7003_n3682# a_6651_n3068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2822 gnd d1 a_7203_3329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2823 a_31192_7392# a_30974_7392# a_30717_7487# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2824 a_19788_3110# d2 a_19838_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2825 a_13267_3220# a_13273_3403# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2826 a_26102_n5061# a_26104_n5160# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2827 a_20606_n6947# a_20610_n6759# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2828 a_4683_n8285# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2829 a_1565_6667# a_1395_7568# a_1519_7687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2830 vdd d1 a_28931_2335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2831 a_n55_n2287# d0 a_426_n2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2832 a_28498_n3502# a_28751_n3706# a_28399_n3092# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2833 gnd d1 a_28844_n8796# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2834 a_21924_4926# d0 a_22415_4919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2835 a_12124_3582# a_12138_4365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2836 vdd d2 a_24528_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2837 a_5661_n6710# d2 a_5744_n7726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2838 vdd d0 a_12271_n8600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2839 a_27694_n5889# a_27476_n5889# a_27518_n3855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2840 a_26393_n6685# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2841 a_12100_2741# a_12104_2564# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2842 a_26629_n7291# a_26411_n7291# a_26138_n7097# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2843 a_23032_n6722# a_22814_n6489# a_22234_n6673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2844 a_11241_4139# d1 a_11323_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2845 a_n32_n3488# d0 a_443_n3594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2846 a_21322_n10664# a_21579_n10680# a_21421_n10664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2847 a_31885_1629# d2 a_31963_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2848 gnd d0 a_3689_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2849 a_2283_n3243# d1 a_2369_n2447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2850 a_8896_2989# a_8903_3207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2851 a_29329_n5542# a_29586_n5558# a_28531_n5726# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2852 a_4880_n7679# a_4662_n7679# a_4399_n7390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2853 a_8776_n7402# a_8782_n7585# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2854 a_17560_4913# a_17562_5012# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2855 a_11376_6585# d0 a_12178_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2856 a_11318_8034# a_11571_8021# a_11235_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 vdd d0 a_20827_n4927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2858 a_22141_1865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2859 a_27771_6585# d4 a_27838_402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2860 gnd d0 a_3672_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2861 a_18050_5318# a_17832_5318# a_17575_5413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2862 a_5773_1592# a_5567_2081# a_4987_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2863 a_27446_n8770# d2 a_27497_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2864 a_30956_n5680# a_30738_n5680# a_30481_n5574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2865 a_21939_5426# a_21941_5944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2866 a_2586_3329# d0 a_3383_3557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2867 a_33932_7679# a_34185_7666# a_33135_7451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2868 a_6761_n9176# d1 a_6856_n9774# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2869 gnd d0 a_33932_n4965# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2870 a_20751_3334# a_20755_3157# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2871 a_24173_n6732# d0 a_24971_n6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2872 a_30517_n7610# a_30522_n8128# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2873 a_28575_2115# d1 a_28661_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2874 a_4480_842# d0 a_4971_835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2875 a_2076_n10565# d4 a_2138_n6113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2876 vdd d1 a_33278_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2877 gnd d1 a_16017_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2878 a_17406_n7389# d0 a_17887_n7678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2879 a_4532_3378# d0 a_5007_3283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2880 a_28648_6187# a_28905_5997# a_28602_7207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2881 a_9970_n2827# a_9764_n3435# a_9185_n3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2882 a_24321_3354# a_24574_3341# a_24235_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2883 gnd d0 a_7783_n2892# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2884 a_23176_6573# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2885 a_20828_7229# a_21081_7216# a_20026_7590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2886 vdd d0 a_3492_n6951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2887 a_16977_n2070# a_17309_n2081# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2888 a_33836_2354# a_34093_2164# a_33038_2538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2889 a_12137_4777# a_12394_4587# a_11344_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2890 a_17633_n5642# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2891 a_2659_7401# d0 a_3456_7629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2892 a_9167_2883# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2893 a_25168_6401# a_25425_6211# a_24370_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2894 a_17599_7048# a_17606_7266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2895 a_13603_7380# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2896 vdd d1 a_2695_n6723# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2897 a_15388_n3281# a_15645_n3297# a_15342_n4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2898 a_15470_n2673# d0 a_16272_n2301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2899 a_20587_n5929# a_20844_n5945# a_19794_n5513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2900 a_4592_7049# d0 a_5081_6943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2901 a_13622_n7292# d1 a_14407_n6912# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2902 a_24152_3123# d2 a_24198_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2903 a_14511_n3856# d4 a_14687_n5890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2904 a_27521_1616# a_27315_2105# a_26736_1877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2905 a_20840_8836# a_21097_8646# a_20047_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2906 a_10026_1485# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2907 a_9166_3295# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2908 vdd d0 a_7821_n4516# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2909 gnd d0 a_3600_1096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2910 a_7604_n6348# a_7599_n6948# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2911 a_24231_n9598# a_24484_n9802# a_24132_n9188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2912 a_16451_1559# a_16704_1546# a_15654_1331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2913 a_19447_n10577# d4 a_19509_n6125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2914 a_27135_n3447# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2915 vdd d0 a_12198_n4528# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2916 a_10043_n6899# a_9837_n7507# a_9258_n7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2917 a_10063_3521# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2918 a_26556_n3219# a_26338_n3219# a_26065_n3025# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2919 a_28426_5173# d3 a_28529_3135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2920 a_16321_n5955# a_16578_n5971# a_15528_n5539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2921 a_18015_2870# d1 a_18812_3098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2922 gnd d0 a_33969_n6589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2923 a_16451_1559# a_16465_2342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2924 a_336_n9290# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2925 gnd d1 a_11633_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2926 a_3457_7217# a_3452_7806# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2927 gnd d0 a_29838_8671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_14366_n7928# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 vdd d2 a_6977_n7344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2930 a_31885_1629# a_31679_2118# a_31100_1890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2931 a_4356_n5136# a_4363_n5354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2932 vdd d0 a_12177_n3922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2933 a_28430_4996# d3 a_28602_7207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2934 a_16537_6826# a_16541_6649# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2935 a_26649_n8309# a_26431_n8309# a_26160_n8214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2936 gnd d0 a_25372_3157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2937 a_11241_4139# d1 a_11327_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2938 a_13424_n8310# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2939 a_31953_5172# a_31735_5172# a_31156_4944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2940 a_11147_n4508# d0 a_11944_n4736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2941 a_2402_n4671# d0 a_3204_n4299# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2942 a_1441_3086# a_1223_3086# a_643_3270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2943 a_11314_8211# a_11571_8021# a_11235_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2944 vdd d0 a_3672_5580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2945 a_17623_8284# d0 a_18104_8372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2946 a_5703_n8923# a_5497_n9531# a_4918_n9303# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2947 a_14407_n6912# d2 a_14485_n7751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2948 a_13348_7993# d0 a_13839_7986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2949 a_13133_n7197# d0 a_13622_n7292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2950 a_22432_5937# a_22214_5937# a_21943_6043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2951 a_16399_n9427# a_16652_n9631# a_15597_n9799# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2952 vdd d0 a_3437_n3485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2953 a_33928_7856# a_34185_7666# a_33135_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2954 a_6909_1483# d0 a_7707_1299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2955 a_10233_2620# a_10063_3521# a_10187_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2956 a_13568_n4650# d1 a_14366_n4699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2957 a_11216_n8768# d0 a_12014_n8584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2958 a_3452_7806# a_3456_7629# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2959 a_643_3270# a_425_3270# a_162_3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2960 a_13549_n3220# d1 a_14334_n2840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2961 a_623_2252# d1 a_1409_1579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2962 gnd d0 a_7874_n7570# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2963 a_7724_2317# a_7728_2140# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2964 a_9475_7973# d1 a_10260_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2965 a_20735_2139# a_20988_2126# a_19933_2500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2966 vdd d1 a_16017_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2967 a_27217_n2839# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2968 a_9257_7973# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2969 a_18104_8372# d1 a_18890_7699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2970 a_21800_n9220# a_21807_n9438# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2971 a_24317_3531# a_24574_3341# a_24235_4139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2972 a_26284_4019# d0 a_26773_3913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2973 a_21941_5944# a_21943_6043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2974 a_20824_7406# a_21081_7216# a_20026_7590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2975 vdd d7 a_25872_n10681# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2976 a_33860_3195# a_33855_3784# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2977 a_17496_1158# a_17502_1341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2978 a_28505_n9388# a_28762_n9404# a_28426_n8184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2979 a_131_1329# a_133_1847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2980 a_717_6930# a_499_6930# a_226_6743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2981 a_5588_n2638# a_5370_n2405# a_4790_n2589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2982 a_8692_n2495# d0 a_9167_n2601# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2983 a_13765_4326# d1 a_14551_3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2984 a_19691_n5291# a_19948_n5307# a_19612_n4087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2985 a_23176_3111# d2 a_23227_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2986 a_11097_n7340# d1 a_11183_n6544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2987 a_7019_7591# d0 a_7821_7230# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2988 a_n27_n4006# a_n25_n4105# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2989 a_28468_n7352# d1 a_28550_n6744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2990 a_24091_n7340# a_24348_n7356# a_24045_n8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2991 vdd d2 a_33053_n5345# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2992 a_9_n6042# d0 a_500_n6236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2993 a_18611_4116# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2994 a_263_n5218# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2995 a_26411_n7291# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2996 a_26755_3307# d1 a_27553_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2997 gnd d0 a_21043_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2998 a_14345_4142# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2999 a_16447_1736# a_16704_1546# a_15654_1331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3000 a_23461_390# d5 a_21581_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 gnd d0 a_29822_7241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3002 vdd d2 a_6904_n3272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3003 a_23144_1604# a_22938_2093# a_22358_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3004 a_33877_4213# a_34130_4200# a_33075_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3005 a_1586_2476# d4 a_1726_365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3006 gnd d0 a_29531_n2916# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3007 a_26576_n4237# a_26358_n4237# a_26087_n4142# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3008 a_17541_3895# d0 a_18032_3888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3009 a_5098_7961# a_4880_7961# a_4607_7968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3010 a_30685_n2214# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3011 a_13351_n4238# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3012 gnd d2 a_28652_n3296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3013 a_14546_3124# a_14328_3124# a_13749_2896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3014 a_4842_6337# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3015 a_24_n6542# a_26_n7060# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3016 a_20551_n3481# a_20808_n3497# a_19753_n3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3017 vdd d0 a_20901_n8587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3018 a_27335_3123# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3019 a_7779_5783# a_7783_5606# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3020 a_204_5401# a_206_5919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3021 a_13230_1184# a_13236_1367# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3022 a_481_n5218# d1 a_1266_n4838# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3023 a_32845_n2497# d0 a_33638_n2913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3024 a_6682_4972# a_6935_4959# a_6085_259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3025 a_33659_n3743# a_33676_n4537# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3026 vdd d0 a_29838_8671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3027 a_10301_6573# a_10099_5557# a_10218_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3028 a_33660_n3331# a_33913_n3535# a_32858_n3703# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3029 gnd d0 a_34006_n8625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3030 a_19920_1305# d0 a_20713_1710# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3031 a_15671_2349# d0 a_16464_2754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3032 a_5043_5319# a_4825_5319# a_4562_5231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3033 a_22975_4129# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3034 a_13326_6457# d0 a_13801_6362# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3035 a_31555_n6514# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3036 a_14485_n7751# d3 a_14584_n7928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3037 a_13330_n3632# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3038 vdd d0 a_20880_n7981# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3039 a_28567_n7762# a_28824_n7778# a_28472_n7164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3040 a_13386_n6686# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3041 a_30975_n6698# d1 a_31773_n6747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3042 a_17849_6336# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3043 a_30758_n6286# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3044 gnd d1 a_15744_n3707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3045 a_17707_n9302# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3046 a_8859_953# a_8866_1171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3047 a_18931_6560# d3 a_19030_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3048 a_27397_1497# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3049 a_28661_1330# d0 a_29454_1735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3050 vdd d3 a_33150_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3051 a_21690_n3112# d0 a_22179_n3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3052 a_26316_5438# d0 a_26791_5343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3053 a_8813_n9438# d0 a_9294_n9727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3054 a_24956_n5342# a_25209_n5546# a_24154_n5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3055 a_11164_n5526# a_11417_n5730# a_11065_n5116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3056 gnd d0 a_34075_1558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3057 a_31699_3136# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3058 a_27300_n3855# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3059 a_5469_n2815# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3060 a_23217_5676# d2 a_23295_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3061 a_21961_6768# d0 a_22452_6955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3062 gnd d0 a_25171_n3922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3063 a_17353_n4335# a_17359_n4518# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3064 a_4590_n3195# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3065 a_11183_n6544# d0 a_11976_n6960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3066 a_24992_n7378# a_24987_n7978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3067 a_20714_1298# a_20718_1121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3068 a_20731_2316# a_20988_2126# a_19933_2500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3069 a_13303_5256# a_13309_5439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3070 a_31013_n8322# a_30795_n8322# a_30524_n8227# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3071 gnd d1 a_15854_n9815# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3072 a_14592_2514# d3 a_14691_2514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3073 a_10053_n3843# a_9883_n4863# a_10002_n4686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3074 a_22215_n5655# d1 a_23001_n4863# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3075 a_17852_n5230# d1 a_18637_n4850# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3076 a_11903_n2888# a_12160_n2904# a_11110_n2472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3077 a_28395_n3280# d1 a_28477_n2672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3078 a_3872_n2032# a_3163_n2451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3079 a_4497_1860# d0 a_4988_1853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3080 a_27470_5569# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3081 a_17616_8066# a_17623_8284# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3082 a_22271_n8709# d1 a_23069_n8758# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3083 gnd d2 a_2793_5960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3084 a_22252_n7279# d1 a_23037_n6899# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3085 gnd d0 a_3653_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3086 a_31772_7208# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3087 a_33655_n3931# a_33912_n3947# a_32862_n3515# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3088 vdd d0 a_34005_n9037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3089 a_27336_n2662# d2 a_27419_n3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3090 a_18739_2488# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3091 a_30812_n9340# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3092 a_3183_n3693# a_3436_n3897# a_2386_n3465# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3093 a_5480_n8513# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3094 a_13568_n4650# a_13350_n4650# a_13093_n4544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3095 a_6651_n3068# d1 a_6746_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3096 a_16381_n8821# a_16395_n9615# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3097 a_208_n2576# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3098 a_14665_6586# d3 a_14764_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3099 vdd d1 a_33208_n8809# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3100 a_1266_n4838# d2 a_1312_n3818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3101 a_2360_n7127# a_2613_n7331# a_2310_n8335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3102 a_21998_n5243# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3103 a_6729_n2648# a_6986_n2664# a_6647_n3256# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3104 a_12138_4365# a_12142_4188# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3105 a_24939_n4324# a_25192_n4528# a_24137_n4696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3106 a_2241_n4075# a_2494_n4279# a_2134_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3107 a_n49_n2470# d0 a_426_n2576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3108 a_26846_7985# a_26628_7985# a_26357_8091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3109 a_4663_n7267# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3110 a_33765_n10039# a_34022_n10055# a_32972_n9623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3111 a_24239_3962# d1 a_24338_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3112 a_17519_2359# d0 a_17994_2264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3113 gnd d0 a_29604_n6988# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3114 a_3276_n8783# a_3290_n9577# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3115 a_14649_4548# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3116 a_24951_n5942# a_25208_n5958# a_24158_n5526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3117 a_19916_1482# a_20173_1292# a_19834_2090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3118 a_6843_n8568# d0 a_7636_n8984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3119 a_26809_5949# d1 a_27594_5688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3120 vdd d0 a_12251_n7582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3121 a_8703_n3330# a_8709_n3513# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3122 vdd d0 a_29822_7241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3123 a_28436_n5128# d1 a_28531_n5726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3124 a_7658_n9402# a_7911_n9606# a_6856_n9774# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3125 a_6023_6561# d4 a_6090_378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3126 a_5749_n7903# a_5579_n8923# a_5703_n8923# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3127 a_20660_n10001# a_17454_n9932# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3128 a_29368_n7802# a_29621_n8006# a_28571_n7574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3129 a_17579_6030# d0 a_18068_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3130 a_406_1840# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3131 vdd d0 a_20807_n3909# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3132 a_27451_n8947# d2 a_27497_n7927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3133 a_21744_n6067# d0 a_22235_n6261# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3134 a_241_7437# a_243_7955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3135 vdd d2 a_19984_n7343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3136 a_19920_1305# d0 a_20717_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3137 a_27558_3652# a_27352_4141# a_26773_3913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3138 a_2417_3098# a_2674_2908# a_2314_5136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3139 vdd d3 a_19865_n4291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3140 a_3401_4163# a_3396_4752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3141 a_15671_2349# d0 a_16468_2577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3142 vdd d1 a_7113_n9790# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3143 a_19612_n4087# a_19865_n4291# a_19505_n6313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3144 a_21883_2372# d0 a_22358_2277# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3145 a_20643_n8983# a_20647_n8795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3146 a_21763_n7184# d0 a_22252_n7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3147 a_24121_n3490# d0 a_24918_n3718# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3148 a_11162_2946# a_11415_2933# a_11055_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3149 a_41_n7560# a_46_n8078# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3150 a_27833_283# d5 a_27932_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3151 a_1721_246# d4 a_2318_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3152 a_4309_n2300# a_4315_n2483# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3153 a_17633_n5642# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3154 a_29402_n9614# a_29659_n9630# a_28604_n9798# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3155 a_24390_7603# d0 a_25192_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3156 a_17689_n8696# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3157 a_18050_5318# d1 a_18848_5134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3158 a_28661_1330# d0 a_29458_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3159 a_553_n9702# a_335_n9702# a_78_n9596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3160 a_14469_n5890# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3161 a_8866_1171# a_8872_1354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3162 a_7821_7230# a_8074_7217# a_7019_7591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3163 a_7653_n10002# a_7910_n10018# a_6860_n9586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3164 a_33038_2538# d0 a_33836_2354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3165 a_3217_n5505# a_3221_n5317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3166 a_5846_5664# a_5640_6153# a_5061_5925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3167 a_27336_n2662# a_27118_n2429# a_26539_n2201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3168 a_25118_3582# a_25371_3569# a_24321_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3169 vdd d0 a_25407_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3170 vdd d0 a_33950_n5571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3171 a_4517_2684# a_4519_2977# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3172 a_29476_2164# a_29471_2753# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3173 a_17513_2176# a_17519_2359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3174 a_10037_7183# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3175 vdd d0 a_7801_n3498# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3176 vdd d0 a_3653_4562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3177 a_22213_6349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3178 a_27135_n3447# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3179 a_20047_8431# d0 a_20840_8836# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3180 a_26808_6361# a_26590_6361# a_26327_6273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3181 a_30674_5268# d0 a_31155_5356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3182 a_33823_1159# a_33818_1748# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3183 a_252_8272# d0 a_733_8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3184 gnd d4 a_2391_n6317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3185 a_19809_n6719# a_20066_n6735# a_19727_n7327# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3186 a_22215_n5655# a_21997_n5655# a_21740_n5549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3187 a_29548_6648# a_29565_7431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3188 a_32939_2128# d1 a_33021_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3189 a_13275_3921# a_13277_4020# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3190 a_30421_n2337# a_30427_n2520# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3191 a_11290_1318# a_11543_1305# a_11204_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3192 a_24104_n2472# a_24357_n2676# a_24018_n3268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3193 a_30864_1284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3194 a_3437_6199# a_3690_6186# a_2635_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3195 a_12088_1134# a_12083_1723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3196 a_19447_n10577# a_19704_n10593# a_19546_n10577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3197 a_n62_n2069# d0 a_427_n2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3198 a_33135_7451# a_33388_7438# a_33049_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3199 vdd d2 a_28832_1925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3200 a_27698_2513# a_27480_2513# a_27604_2632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3201 a_13404_n7292# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3202 a_4900_n8697# a_4682_n8697# a_4419_n8408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3203 a_32869_n9401# d1 a_32951_n8793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3204 a_2382_n3653# d0 a_3184_n3281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3205 a_17316_n2299# d0 a_17797_n2588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3206 a_24935_n4512# a_24939_n4324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3207 a_31963_2526# a_31761_1510# a_31880_1100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3208 vdd d0 a_12467_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3209 a_27838_402# a_27656_4547# a_27698_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3210 a_4369_n5537# a_4373_n6055# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3211 a_6868_3950# a_7121_3937# a_6785_2934# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3212 gnd d0 a_21024_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3213 a_27771_6585# a_27553_6585# a_27677_6704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3214 a_22996_n4686# d2 a_23047_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3215 a_21943_n2601# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3216 a_11196_n7750# d0 a_11994_n7566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3217 vdd d2 a_28725_n7368# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3218 a_1313_8176# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3219 a_33135_7451# d0 a_33928_7856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3220 a_243_7955# a_245_8054# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3221 a_11977_n6548# a_12234_n6564# a_11179_n6732# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3222 a_2138_n6113# a_2391_n6317# a_2076_n10565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3223 a_8804_n9121# a_8806_n9220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3224 vdd d4 a_28683_4983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3225 gnd d2 a_11318_n5320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3226 a_9457_7367# a_9239_7367# a_8982_7462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3227 a_5007_3283# a_4789_3283# a_4526_3195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3228 a_n49_n2470# a_n47_n2988# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3229 a_5588_n2638# a_5370_n2405# a_4791_n2177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3230 a_1514_7158# a_1296_7158# a_717_6930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3231 a_13586_n5256# a_13368_n5256# a_13097_n5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3232 a_8714_n4031# d0 a_9205_n4225# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3233 a_24225_7195# d2 a_24275_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3234 a_20026_7590# d0 a_20824_7406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3235 a_33038_2538# d0 a_33840_2177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3236 a_21770_n7402# a_21776_n7585# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3237 a_226_n3182# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3238 a_13140_n7415# a_13146_n7598# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3239 a_15654_1331# a_15907_1318# a_15568_2116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3240 a_18890_7699# d2 a_18936_6679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3241 a_8343_n10653# d7 a_8244_n10653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3242 a_11904_n2476# a_11908_n2288# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3243 a_10306_6692# a_10136_7593# a_10255_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3244 a_11_n6141# d0 a_500_n6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3245 a_7743_3747# a_8000_3557# a_6950_3342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3246 vdd d0 a_29658_n10042# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3247 a_8740_n5366# a_8746_n5549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3248 a_33655_n3931# a_33659_n3743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3249 gnd d0 a_7980_2539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3250 a_1482_5651# d2 a_1560_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3251 a_29545_6413# a_29549_6236# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3252 a_31880_1100# a_31662_1100# a_31082_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3253 a_20047_8431# d0 a_20844_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3254 a_13221_867# d0 a_13712_860# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3255 a_7637_n8572# a_7894_n8588# a_6839_n8756# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3256 a_28349_n4300# d2 a_28395_n3280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3257 a_30955_5962# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3258 a_26173_n8615# a_26175_n9133# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3259 a_17886_8372# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3260 a_13123_n6397# a_13129_n6580# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3261 a_26576_n4237# a_26358_n4237# a_26085_n4043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3262 gnd d0 a_8036_5593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3263 a_8962_6444# d0 a_9437_6349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3264 a_13129_n6580# a_13131_n7098# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3265 a_8859_953# d0 a_9348_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3266 a_19509_n6125# a_19762_n6329# a_19447_n10577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3267 vdd d0 a_12378_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3268 a_19788_3110# a_20045_2920# a_19685_5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3269 a_26556_n3219# a_26338_n3219# a_26067_n3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3270 a_24338_4372# d0 a_25131_4777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3271 gnd d0 a_34112_3594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3272 a_32939_2128# d1 a_33025_1343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3273 a_24177_n6544# a_24430_n6748# a_24091_n7340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3274 a_32873_n9213# a_33126_n9417# a_32790_n8197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3275 a_5677_8189# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3276 a_26628_7985# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3277 a_480_n5630# d1 a_1266_n4838# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3278 a_23254_7712# d2 a_23300_6692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3279 a_8729_n4531# a_8731_n5049# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3280 a_11944_n4736# a_12197_n4940# a_11147_n4508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3281 a_14366_n7928# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3282 a_1560_6548# d3 a_1659_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3283 a_27378_n4875# a_27172_n5483# a_26592_n5667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3284 a_2455_n7725# d0 a_3257_n7353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3285 a_14247_n4876# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3286 a_3433_6376# a_3690_6186# a_2635_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3287 a_607_822# d1 a_1404_1050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3288 a_31172_6374# a_30954_6374# a_30697_6469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3289 a_31555_n6514# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3290 a_15392_n3093# d1 a_15487_n3691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3291 a_28602_7207# a_28859_7017# a_28430_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3292 a_5649_1473# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3293 a_6913_1306# d0 a_7706_1711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3294 a_13424_n8310# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3295 a_15239_n6339# d3 a_15342_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3296 a_9076_n9727# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3297 a_6605_n4088# d2 a_6688_n5104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3298 a_26627_8397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3299 a_15470_n2673# a_15727_n2689# a_15388_n3281# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3300 a_17707_n9302# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3301 a_29279_n2300# a_29532_n2504# a_28477_n2672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3302 vdd d1 a_7220_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3303 a_8819_n9621# d0 a_9294_n9727# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3304 a_31955_n7940# a_31737_n7940# a_31856_n7763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3305 a_33680_n4349# a_33675_n4949# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3306 a_8911_3908# a_8913_4007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3307 a_27408_7195# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3308 a_27300_n3855# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3309 vdd d0 a_21024_4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3310 a_32786_n8385# d2 a_32832_n7365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3311 a_31990_7208# d2 a_32041_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3312 a_33638_n2913# a_33895_n2929# a_32845_n2497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3313 a_5722_5545# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3314 a_4405_n7573# d0 a_4880_n7679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3315 a_31013_n8322# a_30795_n8322# a_30522_n8128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3316 a_11907_n2700# a_11921_n3494# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3317 a_33135_7451# d0 a_33932_7679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3318 a_30993_n7304# a_30775_n7304# a_30504_n7209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3319 a_11921_n3494# a_11925_n3306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3320 a_8999_8480# a_7837_8660# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3321 a_33053_8059# d1 a_33148_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3322 a_19953_3518# a_20210_3328# a_19871_4126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3323 gnd d0 a_16614_n8007# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3324 a_5443_n6477# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3325 a_27217_n2839# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3326 vdd d1 a_7293_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3327 a_4562_5231# a_4568_5414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3328 a_26228_866# a_26230_965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3329 a_22251_n7691# d1 a_23037_n6899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3330 a_191_5000# d0 a_680_4894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3331 vdd d0 a_29585_n5970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3332 a_4864_n6249# a_4646_n6249# a_4373_n6055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3333 a_13240_1984# d0 a_13729_1878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3334 a_18890_7699# a_18684_8188# a_18105_7960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3335 gnd d3 a_15672_n8389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3336 a_15524_n5727# a_15781_n5743# a_15429_n5129# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3337 a_12156_5795# a_12160_5618# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3338 a_20026_7590# d0 a_20828_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3339 a_8658_196# a_12832_197# a_12951_197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3340 vdd d0 a_3599_1508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3341 a_7564_n4500# a_7821_n4516# a_6766_n4684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3342 a_5460_n7495# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3343 a_24049_n8172# d2 a_24128_n9376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3344 a_208_n2576# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3345 a_13548_3914# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3346 gnd d1 a_20246_5364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3347 a_11061_n5304# d1 a_11147_n4508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3348 a_13230_1184# d0 a_13711_1272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3349 gnd d1 a_15997_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3350 vdd d1 a_33188_n7791# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3351 a_21998_n5243# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3352 a_9421_4919# d1 a_10218_5147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3353 a_198_5218# d0 a_679_5306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3354 a_20808_6211# a_21061_6198# a_20006_6572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3355 a_22289_n9315# a_22071_n9315# a_21800_n9220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3356 a_4663_n7267# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3357 a_29274_n2900# a_29531_n2916# a_28481_n2484# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3358 a_13247_2202# d0 a_13728_2290# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3359 a_263_n5218# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3360 a_26538_2895# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3361 a_6823_n7550# d0 a_7616_n7966# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3362 a_31100_1890# a_30882_1890# a_30611_1996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3363 gnd d1 a_28987_5389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3364 a_13621_7986# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3365 a_17834_n4624# d1 a_18632_n4673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3366 a_5924_6561# a_5722_5545# a_5846_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3367 a_2402_n4671# a_2659_n4687# a_2320_n5279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3368 a_13303_5256# d0 a_13784_5344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3369 a_7838_8248# a_7833_8837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3370 a_11359_5567# d0 a_12157_5383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3371 a_17815_n3194# d1 a_18600_n2814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3372 a_13711_1272# d1 a_14509_1088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3373 a_5749_n7903# a_5579_n8923# a_5698_n8746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3374 a_22868_n9543# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3375 a_16399_n9427# a_16394_n10027# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3376 a_7599_n6948# a_7856_n6964# a_6806_n6532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3377 a_22234_n6673# d1 a_23032_n6722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3378 a_6909_1483# a_7166_1293# a_6827_2091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3379 a_30458_n4373# d0 a_30939_n4662# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3380 a_8757_196# d8 a_17217_n720# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3381 a_18088_6942# a_17870_6942# a_17597_6755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3382 a_15572_1939# d1 a_15667_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3383 a_20571_n4499# a_20828_n4515# a_19773_n4683# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3384 a_10182_3111# a_9964_3111# a_9385_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3385 a_21907_4007# d0 a_22396_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3386 a_13351_n4238# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3387 a_17324_n3000# d0 a_17815_n3194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3388 a_1203_2068# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3389 a_17832_5318# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3390 a_33075_4574# d0 a_33873_4390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3391 vdd d3 a_20118_6992# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3392 a_21746_n6166# d0 a_22235_n6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3393 a_16538_6414# a_16542_6237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3394 a_25012_n8396# a_25265_n8600# a_24210_n8768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3395 a_13531_n2614# a_13313_n2614# a_13056_n2508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3396 a_18032_3888# a_17814_3888# a_17543_3994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3397 a_4579_6249# d0 a_5060_6337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3398 a_30481_n5574# d0 a_30956_n5680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3399 a_14334_n2840# a_14128_n3448# a_13549_n3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3400 a_12105_2152# a_12100_2741# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3401 a_29406_n9426# a_29401_n10026# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3402 vdd d3 a_15852_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3403 a_28575_2115# d1 a_28657_1507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3404 a_18931_6560# a_18729_5544# a_18848_5134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3405 a_4050_n10652# d6 a_3951_n10652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3406 a_17995_1852# d1 a_18780_1591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3407 a_22378_3295# a_22160_3295# a_21897_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3408 a_536_n8684# a_318_n8684# a_61_n8578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3409 a_28509_n9200# d1 a_28604_n9798# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3410 a_63_n9096# d0 a_554_n9290# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3411 a_6913_1306# d0 a_7710_1534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3412 a_25155_5206# a_25408_5193# a_24353_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3413 a_19867_n9585# d0 a_20660_n10001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3414 a_1259_5122# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3415 a_20804_6388# a_20808_6211# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3416 a_22378_3295# d1 a_23176_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3417 a_553_n9702# a_335_n9702# a_72_n9413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3418 a_16288_n3731# a_16305_n4525# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3419 a_22451_7367# a_22233_7367# a_21970_7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3420 a_12197_7654# a_12450_7641# a_11400_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3421 a_27290_n6911# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3422 a_1409_1579# a_1203_2068# a_623_2252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3423 a_24988_n7566# a_24992_n7378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3424 a_16340_n6973# a_16344_n6785# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3425 a_29513_4200# a_29508_4789# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3426 a_33053_8059# d1 a_33152_8469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3427 a_18863_2607# d3 a_18957_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3428 a_31119_3320# a_30901_3320# a_30644_3415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3429 a_32899_n5551# d0 a_33692_n5967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3430 vdd d1 a_6986_n2664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3431 a_281_n6648# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3432 a_4499_1959# a_4506_2177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3433 a_478_6324# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3434 gnd d5 a_2333_n10581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3435 a_33675_n4949# a_33932_n4965# a_32882_n4533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3436 a_24053_4984# d3 a_24229_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3437 gnd d3 a_24229_n4304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3438 a_3203_n4711# a_3456_n4915# a_2406_n4483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3439 a_4988_1853# a_4770_1853# a_4499_1959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3440 vdd d1 a_2819_2298# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3441 vdd d1 a_20246_5364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3442 a_26318_5956# d0 a_26809_5949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3443 a_198_5218# a_204_5401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3444 a_1261_n4661# d2 a_1312_n3818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3445 a_13583_6362# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3446 a_22215_n5655# a_21997_n5655# a_21734_n5366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3447 gnd d0 a_16634_n9025# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3448 vdd d0 a_25462_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3449 a_6498_n6314# d3 a_6601_n4276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3450 a_15727_5403# d0 a_16524_5631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3451 a_24284_1318# d0 a_25077_1723# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3452 a_31581_n2852# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3453 a_3346_1521# a_3360_2304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3454 a_11245_3962# a_11498_3949# a_11162_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3455 vdd d0 a_29569_n4540# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3456 a_10285_4535# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3457 a_209_n2164# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3458 a_20644_n8571# a_20901_n8587# a_19846_n8755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3459 a_4553_4914# d0 a_5044_4907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3460 a_26573_5343# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3461 a_215_6236# a_221_6419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3462 a_17994_2264# a_17776_2264# a_17513_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3463 gnd d1 a_11670_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3464 gnd d2 a_15825_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3465 a_17579_n2588# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3466 a_7780_5371# a_7784_5194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3467 a_5768_1063# a_5550_1063# a_4970_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3468 vdd d3 a_2747_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3469 a_28246_n6338# a_28503_n6354# a_28188_n10602# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3470 a_15572_1939# d1 a_15671_2349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3471 a_23093_5557# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3472 a_10223_5676# a_10017_6165# a_9437_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3473 a_9039_n7691# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3474 a_696_6324# a_478_6324# a_221_6419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3475 gnd d3 a_11488_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3476 a_14473_2514# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3477 a_26736_1877# a_26518_1877# a_26245_1884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3478 a_32931_n7775# d0 a_33729_n7591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3479 a_28422_n8372# d2 a_28472_n7164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3480 a_20623_n7965# a_20880_n7981# a_19830_n7549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3481 a_24974_n6772# a_25227_n6976# a_24177_n6544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3482 a_12017_n8808# a_12031_n9602# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3483 a_17834_n4624# a_17616_n4624# a_17359_n4518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3484 a_23001_n4863# d2 a_23047_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3485 a_21943_n2601# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3486 a_28715_4384# a_28968_4371# a_28616_3974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3487 a_33712_n6573# a_33969_n6589# a_32914_n6757# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3488 a_26718_1271# a_26500_1271# a_26243_1366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3489 a_18637_n4850# a_18431_n5458# a_17852_n5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3490 a_28246_n6338# d3 a_28353_n4112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3491 a_9_n6042# a_11_n6141# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3492 a_12120_3759# a_12377_3569# a_11327_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3493 a_13801_6362# a_13583_6362# a_13326_6457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3494 a_20611_n6347# a_20606_n6947# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3495 a_21783_n8202# d0 a_22272_n8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3496 gnd d0 a_8017_4575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3497 a_26735_2289# a_26517_2289# a_26260_2384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3498 a_14371_n4876# a_14165_n5484# a_13586_n5256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3499 a_21697_n3330# a_21703_n3513# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3500 a_30458_n4373# a_30464_n4556# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3501 a_22432_5937# d1 a_23217_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3502 a_8999_8480# d0 a_9474_8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3503 a_13586_n5256# a_13368_n5256# a_13095_n5062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3504 a_26791_5343# a_26573_5343# a_26316_5438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3505 a_8716_n4130# d0 a_9205_n4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3506 a_19740_n2459# d0 a_20533_n2875# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3507 a_27516_1087# a_27298_1087# a_26719_859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3508 a_12193_7831# a_12450_7641# a_11400_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3509 a_19092_258# d4 a_19685_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3510 a_8694_n3013# d0 a_9185_n3207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3511 gnd d1 a_24467_n8784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3512 a_14619_7196# d2 a_14670_6705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3513 a_27336_n2662# a_27118_n2429# a_26538_n2613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3514 a_8874_1872# a_8876_1971# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3515 a_23295_6573# a_23093_5557# a_23217_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3516 a_22016_n6673# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3517 a_14111_n2430# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3518 a_7019_7591# d0 a_7817_7407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3519 a_31083_872# a_30865_872# a_30594_978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3520 a_29348_n6560# a_29605_n6576# a_28550_n6744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3521 vdd d0 a_16561_n4953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3522 a_32713_n4313# d2 a_32763_n3105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3523 a_25910_208# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3524 a_n18_n4323# a_n12_n4506# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3525 a_25118_3582# a_25132_4365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3526 a_8962_6444# a_8967_6768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3527 a_14444_n8948# a_14238_n9556# a_13658_n9740# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3528 gnd d2 a_11391_n9392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3529 a_4790_n2589# a_4572_n2589# a_4315_n2483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3530 a_22938_2093# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3531 a_28747_6597# a_29004_6407# a_28652_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3532 a_7617_n7554# a_7874_n7570# a_6819_n7738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3533 a_25094_2741# a_25098_2564# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3534 a_8787_n8103# d0 a_9278_n8297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3535 a_21883_2372# a_21888_2696# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3536 a_8679_n2094# a_8686_n2312# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3537 vdd d3 a_15599_n4317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3538 gnd d0 a_16831_8672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3539 a_24284_1318# d0 a_25081_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3540 a_8966_n3619# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3541 a_6781_3111# a_7038_2921# a_6678_5149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3542 a_9277_n8709# a_9059_n8709# a_8796_n8420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3543 a_680_4894# a_462_4894# a_191_5000# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3544 a_18735_n5864# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3545 gnd d0 a_29766_4187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3546 a_172_3982# d0 a_661_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3547 a_30414_n2119# a_30421_n2337# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3548 a_13177_n9451# a_13183_n9634# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3549 a_11924_n3718# a_12177_n3922# a_11127_n3490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3550 a_14247_n4876# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3551 vdd d0 a_3710_7204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3552 a_6729_n2648# d0 a_7527_n2464# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3553 vdd d1 a_11670_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3554 a_16562_7255# a_16557_7844# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3555 vdd d0 a_34165_6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3556 gnd d2 a_7194_8009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3557 a_22161_n2601# a_21943_n2601# a_21686_n2495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3558 gnd d1 a_20227_4346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3559 a_21963_7061# a_21970_7279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3560 a_9076_n9727# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3561 a_11106_n2660# d0 a_11904_n2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3562 a_5759_7581# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3563 a_2320_n5279# a_2577_n5295# a_2241_n4075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3564 a_9402_3901# d1 a_10187_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3565 vdd d1 a_15800_n6761# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3566 a_179_4200# d0 a_660_4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3567 gnd d1 a_20283_7400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3568 a_8539_196# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3569 a_13050_n2325# a_13056_n2508# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3570 a_17814_3888# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3571 a_33749_n8609# a_34006_n8625# a_32951_n8793# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3572 a_28514_n4708# d0 a_29312_n4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3573 gnd d4 a_24126_n6342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3574 a_15564_n7575# d0 a_16357_n7991# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3575 a_28711_4561# a_28968_4371# a_28616_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3576 gnd d1 a_24394_n4712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3577 a_26267_3001# d0 a_26756_2895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3578 a_5061_5925# a_4843_5925# a_4572_6031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3579 a_4427_n9109# d0 a_4918_n9303# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3580 vdd d0 a_33968_n7001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3581 a_11138_n9188# a_11391_n9392# a_11055_n8172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3582 a_13284_4238# d0 a_13765_4326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3583 a_2463_2078# d1 a_2545_1470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3584 a_22359_1865# a_22141_1865# a_21870_1971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3585 a_17309_n2081# d0 a_17798_n2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3586 a_19097_377# a_18915_4522# a_18957_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3587 a_30993_n7304# a_30775_n7304# a_30502_n7110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3588 a_31172_6374# d1 a_31958_5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3589 vdd d0 a_8017_4575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3590 a_5443_n6477# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3591 a_6785_2934# d2 a_6864_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3592 a_32968_n9811# d0 a_33766_n9627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3593 a_15243_n6151# d3 a_15415_n8373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3594 a_33693_n5555# a_33950_n5571# a_32895_n5739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3595 a_3364_2127# a_3617_2114# a_2562_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3596 a_2540_5973# a_2793_5960# a_2490_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3597 a_9240_6955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3598 a_17813_4300# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3599 a_4354_n5037# a_4356_n5136# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3600 a_13749_2896# a_13531_2896# a_13258_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3601 a_28608_n9610# d0 a_29401_n10026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3602 a_6946_3519# a_7203_3329# a_6864_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3603 a_32036_6598# a_31834_5582# a_31953_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3604 a_26274_3219# d0 a_26755_3307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3605 a_464_n4200# a_246_n4200# a_n27_n4006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3606 a_246_n4200# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3607 a_8857_854# a_8859_953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3608 a_26612_n6273# a_26394_n6273# a_26123_n6178# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3609 a_7544_n3482# a_7801_n3498# a_6746_n3666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3610 a_18594_3098# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3611 a_27507_7605# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3612 vdd d0 a_7894_n8588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3613 a_4543_4213# d0 a_5024_4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3614 a_11028_n3080# d1 a_11127_n3490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3615 a_22289_n9315# a_22071_n9315# a_21798_n9121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3616 gnd d1 a_7239_5365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3617 a_13748_3308# a_13530_3308# a_13273_3403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3618 a_13822_6968# a_13604_6968# a_13331_6781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3619 gnd d0 a_29642_n8612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3620 a_18414_n4440# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3621 a_18936_6679# a_18766_7580# a_18885_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3622 a_517_n7254# d1 a_1302_n6874# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3623 a_24239_3962# d1 a_24334_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3624 gnd d0 a_16815_7242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3625 a_18394_n3422# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3626 a_7620_n7778# a_7637_n8572# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3627 a_7801_6212# a_8054_6199# a_6999_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3628 a_16394_n10027# a_16651_n10043# a_15601_n9611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3629 a_23461_390# a_23279_4535# a_23321_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3630 gnd d1 a_33315_3366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3631 a_443_n3594# a_225_n3594# a_n38_n3305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3632 a_17814_n3606# d1 a_18600_n2814# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3633 a_11220_n8580# d0 a_12017_n8808# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3634 a_17597_n3194# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3635 a_22868_n9543# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3636 a_2382_n3653# a_2639_n3669# a_2287_n3055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3637 vdd d0 a_7873_n7982# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3638 a_15597_n9799# a_15854_n9815# a_15502_n9201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3639 a_30464_n4556# d0 a_30939_n4662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3640 a_30438_n3355# d0 a_30919_n3644# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3641 a_9348_847# a_9130_847# a_8857_854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3642 a_17556_4395# d0 a_18031_4300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3643 vdd d0 a_20845_n5533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3644 vdd d0 a_21080_7628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3645 a_27497_n7927# a_27327_n8947# a_27451_n8947# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3646 a_31700_n2675# a_31482_n2442# a_30902_n2626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3647 a_30601_1196# a_30607_1379# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3648 vdd d4 a_24306_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3649 vdd d0 a_16831_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3650 a_14320_n8948# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3651 a_15599_7031# d2 a_15678_8224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3652 a_n1_n5341# a_5_n5524# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3653 a_8986_n4637# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3654 a_13531_n2614# a_13313_n2614# a_13050_n2325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3655 a_26029_208# d7 a_17148_133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3656 a_26158_n8115# a_26160_n8214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3657 a_24992_n7378# a_25245_n7582# a_24190_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3658 a_15511_n4521# d0 a_16304_n4937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3659 a_16284_n3919# a_16288_n3731# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3660 gnd d6 a_21579_n10680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3661 a_3272_n8971# a_3529_n8987# a_2479_n8555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3662 a_6757_n9364# d1 a_6843_n8568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3663 vdd d3 a_7111_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3664 a_2475_n8743# d0 a_3277_n8371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3665 a_27677_6704# a_27507_7605# a_27631_7724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3666 a_2393_n9351# a_2650_n9367# a_2314_n8147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3667 a_24231_n9598# d0 a_25024_n10014# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3668 a_15181_n10603# d4 a_15239_n6339# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3669 a_26370_8492# d0 a_26845_8397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3670 a_516_n7666# a_298_n7666# a_41_n7560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3671 a_4354_n5037# d0 a_4845_n5231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3672 a_1285_1460# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3673 a_7743_3747# a_7747_3570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3674 a_17888_n7266# d1 a_18673_n6886# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3675 vdd d0 a_33895_n2929# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3676 vdd d1 a_20227_4346# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3677 a_25204_8849# a_25461_8659# a_24411_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3678 a_4315_n2483# d0 a_4790_n2589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3679 a_24390_7603# d0 a_25188_7419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3680 a_9146_2277# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3681 a_31955_n7940# a_31737_n7940# a_31861_n7940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3682 a_33676_n4537# a_33680_n4349# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3683 a_17333_n3317# a_17339_n3500# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3684 a_27290_n6911# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3685 a_19809_n6719# d0 a_20607_n6535# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3686 a_19792_2933# d2 a_19875_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3687 a_13604_n6686# a_13386_n6686# a_13129_n6580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3688 a_3456_7629# a_3709_7616# a_2659_7401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3689 a_33733_n7403# a_33728_n8003# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3690 a_20534_n2463# a_20791_n2479# a_19736_n2647# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3691 a_31788_n3868# a_31618_n4888# a_31742_n4888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3692 a_4425_n8591# d0 a_4900_n8697# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3693 a_26554_4325# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3694 a_2175_n10565# d5 a_1582_n5852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3695 a_2463_2078# d1 a_2549_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3696 gnd d0 a_3419_n2879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3697 a_1368_2476# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3698 vdd d0 a_16579_n5559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3699 a_155_2964# a_162_3182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3700 a_30661_4433# d0 a_31136_4338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3701 a_12215_8260# a_12210_8849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3702 a_11323_3531# d0 a_12125_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3703 a_3360_2304# a_3617_2114# a_2562_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3704 a_20807_6623# a_21060_6610# a_20010_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3705 a_18632_n7902# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3706 a_30717_7487# d0 a_31192_7392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3707 a_4864_n6249# a_4646_n6249# a_4375_n6154# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3708 a_26333_6456# a_26338_6780# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3709 a_15584_n8593# d0 a_16377_n9009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3710 a_30734_8505# a_29585_8684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3711 a_26829_6967# a_26611_6967# a_26340_7073# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3712 vdd d0 a_25191_n4940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3713 a_23337_271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3714 vdd d1 a_7239_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3715 a_27424_n3855# a_27254_n4875# a_27378_n4875# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3716 a_31581_n2852# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3717 a_10233_2620# d3 a_10327_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3718 vdd d0 a_16815_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3719 a_26167_n8432# d0 a_26648_n8721# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3720 gnd d0 a_3473_n5933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3721 a_25115_3347# a_25372_3157# a_24317_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3722 vdd d1 a_33315_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3723 a_20006_6572# d0 a_20804_6388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3724 a_30901_3320# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3725 a_6868_3950# d1 a_6967_4360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3726 a_6684_n5292# d1 a_6770_n4496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3727 a_17835_n4212# d1 a_18632_n4673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3728 a_9347_1259# d1 a_10145_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3729 a_26772_4325# a_26554_4325# a_26297_4420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3730 gnd d1 a_2676_n5705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3731 a_10817_n10590# d4 a_10879_n6138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3732 a_4987_2265# d1 a_5773_1592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3733 a_17217_n720# a_17029_133# a_17148_133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3734 a_19546_n10577# d5 a_19447_n10577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3735 a_22923_n3843# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3736 a_31192_7392# d1 a_31990_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3737 a_15599_7031# d2 a_15682_8047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3738 a_32832_n7365# d1 a_32914_n6757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3739 a_6827_2091# d1 a_6913_1306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3740 a_388_1234# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3741 a_17569_5230# d0 a_18050_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3742 gnd d0 a_12467_8659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3743 a_20623_n7965# a_20627_n7777# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3744 a_22054_n8297# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3745 a_462_4894# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3746 a_17834_n4624# a_17616_n4624# a_17353_n4335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3747 a_19911_5985# a_20164_5972# a_19861_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3748 a_14334_n2840# a_14128_n3448# a_13548_n3632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3749 a_1224_n2625# d2 a_1307_n3641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3750 a_17814_n3606# a_17596_n3606# a_17339_n3500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3751 gnd d2 a_11281_n3284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3752 a_13511_1878# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3753 a_4971_835# a_4753_835# a_4480_842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3754 a_11400_7426# a_11653_7413# a_11314_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3755 a_24934_n4924# a_25191_n4940# a_24141_n4508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3756 a_13493_1272# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3757 gnd d1 a_20047_n5717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3758 a_17506_1958# a_17513_2176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3759 a_24128_n9376# d1 a_24210_n8768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3760 a_461_5306# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3761 a_21907_4007# a_21914_4225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3762 a_5640_6153# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3763 a_19768_n9175# a_20021_n9379# a_19685_n8159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3764 a_29512_4612# a_29765_4599# a_28715_4384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3765 a_24137_n4696# a_24394_n4712# a_24055_n5304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3766 a_13510_2290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3767 a_12035_n9414# a_12030_n10014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3768 a_8696_n3112# d0 a_9185_n3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3769 a_3452_7806# a_3709_7616# a_2659_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3770 gnd d1 a_24447_n7766# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3771 a_17907_n8696# a_17689_n8696# a_17432_n8590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3772 a_21926_5025# d0 a_22415_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3773 a_22016_n6673# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3774 a_624_1840# a_406_1840# a_135_1946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3775 a_14291_1088# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3776 a_5841_5135# a_5623_5135# a_5044_4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3777 a_7747_3570# a_8000_3557# a_6950_3342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3778 a_11061_n5304# a_11318_n5320# a_10982_n4100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3779 a_18595_n2637# d2 a_18678_n3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3780 a_12157_5383# a_12161_5206# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3781 a_14444_n8948# a_14238_n9556# a_13659_n9328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3782 a_281_n6648# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3783 a_20754_3569# a_20768_4352# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3784 a_20803_6800# a_21060_6610# a_20010_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3785 a_14665_6586# a_14463_5570# a_14582_5160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3786 a_18647_6152# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3787 a_18957_2488# a_18739_2488# a_18858_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3788 a_28430_4996# a_28683_4983# a_27833_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3789 a_32836_n7177# a_33089_n7381# a_32786_n8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3790 a_11233_n9786# d0 a_12035_n9414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3791 a_20648_n8383# a_20643_n8983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3792 a_31882_n3868# d4 a_32058_n5902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3793 a_32943_1951# a_33196_1938# a_32893_3148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3794 a_2676_8419# d0 a_3469_8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3795 gnd d0 a_12378_3157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3796 a_20840_8836# a_20844_8659# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3797 a_8767_n7085# d0 a_9258_n7279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3798 a_14412_n3679# a_14210_n2840# a_14329_n2663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3799 a_3364_2127# a_3359_2716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3800 a_13240_1984# a_13247_2202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3801 a_17434_n9108# a_17436_n9207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3802 a_9004_n5243# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3803 gnd d1 a_33368_6420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3804 a_17652_n6660# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3805 a_15524_n5727# d0 a_16322_n5543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3806 a_18735_n5864# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3807 a_9257_n7691# a_9039_n7691# a_8776_n7402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3808 a_21243_n2044# d0 a_22162_n2189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3809 a_28287_n10602# d5 a_28188_n10602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3810 vdd d2 a_2540_n3259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3811 vdd d2 a_15755_n9405# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3812 a_16305_n4525# a_16562_n4541# a_15507_n4709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3813 a_18915_4522# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3814 a_30618_2214# a_30624_2397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3815 a_24901_n2700# a_24915_n3494# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3816 a_24915_n3494# a_24919_n3306# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3817 a_22161_n2601# a_21943_n2601# a_21680_n2312# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3818 a_8692_n2495# a_8694_n3013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3819 a_28606_7030# a_28859_7017# a_28430_4996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3820 vdd d0 a_7981_2127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3821 a_1726_365# a_1544_4510# a_1586_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3822 a_33818_1748# a_34075_1558# a_33025_1343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3823 a_17417_n8090# a_17419_n8189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3824 a_13221_867# a_16448_1324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3825 a_28353_n4112# d2 a_28436_n5128# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3826 gnd d1 a_7220_4347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3827 a_644_2858# d1 a_1441_3086# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3828 a_13622_n7292# a_13404_n7292# a_13133_n7197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3829 a_61_n8578# a_63_n9096# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3830 vdd d1 a_15907_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3831 vdd d0 a_29548_n3934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3832 a_28494_n3690# d0 a_29292_n3506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3833 a_4429_n9208# d0 a_4918_n9303# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3834 a_18637_n4850# a_18431_n5458# a_17851_n5642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3835 a_10150_1604# a_9944_2093# a_9365_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3836 a_20607_n6535# a_20611_n6347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3837 vdd d0 a_8054_6199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3838 a_10182_3111# d2 a_10233_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3839 a_11396_7603# a_11653_7413# a_11314_8211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3840 a_7727_2552# a_7744_3335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3841 a_427_n2164# a_209_n2164# a_n62_n2069# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3842 a_19957_3341# a_20210_3328# a_19871_4126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3843 gnd d1 a_7293_8419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3844 a_2582_3506# d0 a_3380_3322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3845 a_26591_5949# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3846 a_23317_n5877# a_23099_n5877# a_23214_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3847 a_30451_n4155# a_30458_n4373# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3848 a_7706_1711# a_7710_1534# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3849 a_7616_n7966# a_7620_n7778# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3850 a_1479_n7890# a_1261_n7890# a_1380_n7713# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3851 vdd d0 a_34023_n9643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3852 vdd d3 a_15779_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3853 a_4495_1342# a_4497_1860# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3854 a_22196_5331# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3855 a_21933_5243# a_21939_5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3856 a_2549_1293# d0 a_3342_1698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3857 vdd d0 a_25209_n5546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3858 a_18067_6336# a_17849_6336# a_17592_6431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3859 a_26612_n6273# a_26394_n6273# a_26121_n6079# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3860 a_32763_n3105# a_33016_n3309# a_32713_n4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3861 a_15498_n9389# d1 a_15584_n8593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3862 a_10255_7183# d2 a_10306_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3863 a_1006_n2392# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3864 a_32020_4560# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3865 gnd d4 a_19942_4958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3866 a_15744_6421# a_15997_6408# a_15645_6011# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3867 a_28587_n8780# d0 a_29385_n8596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3868 a_14831_403# d5 a_12951_197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3869 a_7547_n3706# a_7564_n4500# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3870 a_8767_n7085# a_8769_n7184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3871 a_1096_n7482# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3872 a_241_7437# d0 a_716_7342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3873 a_19097_377# d5 a_19191_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3874 a_14111_n2430# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3875 a_11318_8034# d1 a_11413_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3876 a_22358_2277# d1 a_23144_1604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3877 gnd d0 a_29622_n7594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3878 a_13087_n4361# a_13093_n4544# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3879 a_18394_n3422# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3880 a_26153_n7597# a_26158_n8115# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3881 a_153_2671# d0 a_644_2858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3882 a_28734_5402# a_28987_5389# a_28648_6187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3883 a_14551_3653# d2 a_14597_2633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3884 a_24198_2103# d1 a_24284_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3885 a_26355_7992# a_26357_8091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3886 vdd d2 a_15682_n5333# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3887 a_20845_8247# a_21098_8234# a_20043_8608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3888 a_14511_n3856# a_14293_n3856# a_14417_n3856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3889 a_11200_n7562# d0 a_11997_n7790# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3890 a_2676_8419# d0 a_3473_8647# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3891 a_8967_6768# a_8969_7061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3892 a_30444_n3538# d0 a_30919_n3644# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3893 a_28399_n3092# d1 a_28498_n3502# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3894 a_27497_n7927# a_27327_n8947# a_27446_n8770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3895 a_31700_n2675# a_31482_n2442# a_30903_n2214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3896 a_18693_3508# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3897 a_22432_5937# a_22214_5937# a_21941_5944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3898 a_9205_n4225# d1 a_10002_n4686# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3899 a_8986_n4637# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3900 a_4791_n2177# a_4573_n2177# a_3872_n2032# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3901 a_14427_3534# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3902 vdd d1 a_33368_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3903 a_3240_n6335# a_3493_n6539# a_2438_n6707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3904 a_9221_n5655# a_9003_n5655# a_8746_n5549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3905 a_4622_8468# d0 a_5097_8373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3906 a_19681_n8347# d2 a_19727_n7327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3907 a_21708_n4031# a_21710_n4130# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3908 a_8966_n3619# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3909 a_9277_n8709# a_9059_n8709# a_8802_n8603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3910 a_32135_6598# d4 a_32202_415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3911 a_24411_8444# a_24664_8431# a_24312_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3912 a_7641_n8384# a_7636_n8984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3913 a_22414_5331# a_22196_5331# a_21939_5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3914 a_23139_1075# a_22921_1075# a_22342_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3915 a_3433_6376# a_3437_6199# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3916 a_17908_n8284# a_17690_n8284# a_17417_n8090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3917 a_15491_n3503# d0 a_16284_n3919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3918 a_5671_n3654# d3 a_5770_n3831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3919 a_31100_1890# d1 a_31885_1629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3920 gnd d3 a_15852_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3921 a_3252_n7953# a_3509_n7969# a_2459_n7537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3922 a_18467_n7494# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3923 a_30063_n10689# a_30320_n10705# a_25615_n10665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3924 a_6724_n7140# d1 a_6823_n7550# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3925 a_9257_7973# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3926 a_516_n7666# a_298_n7666# a_35_n7377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3927 vdd d0 a_25281_n10030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3928 a_24227_n9786# d0 a_25025_n9602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3929 a_4356_n5136# d0 a_4845_n5231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3930 a_32135_6598# a_31917_6598# a_32036_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3931 gnd d5 a_15438_n10619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3932 a_31156_4944# d1 a_31953_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3933 a_4337_n4019# d0 a_4828_n4213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3934 a_14500_7606# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3935 a_2310_n8335# a_2567_n8351# a_2138_n6113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3936 a_33660_n3331# a_33655_n3931# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3937 a_6085_259# d5 a_4210_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3938 gnd d2 a_19911_n3271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3939 a_23212_5147# a_22994_5147# a_22415_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3940 a_10982_n4100# a_11235_n4304# a_10875_n6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3941 a_4382_n6372# a_4388_n6555# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3942 a_18032_3888# d1 a_18817_3627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3943 a_6440_n10578# a_6697_n10594# a_3951_n10652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3944 a_9256_8385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3945 a_26057_n2324# d0 a_26538_n2613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3946 a_4806_4301# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3947 gnd d0 a_3690_6186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3948 gnd d0 a_12214_n5958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3949 vdd d1 a_2749_n9777# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3950 a_2237_n4263# d2 a_2283_n3243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3951 a_29388_n8820# a_29402_n9614# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3952 vdd d0 a_20864_n6551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3953 a_18051_4906# a_17833_4906# a_17562_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3954 a_18863_2607# a_18693_3508# a_18817_3627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3955 a_29475_2576# a_29492_3359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3956 a_55_n8395# a_61_n8578# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3957 a_30592_879# a_33819_1336# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3958 a_17526_2976# d0 a_18015_2870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3959 a_2582_3506# d0 a_3384_3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3960 a_33933_7267# a_34186_7254# a_33131_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3961 a_11245_3962# d1 a_11344_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3962 a_18632_n7902# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3963 a_29564_7843# a_29568_7666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3964 a_499_6930# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3965 a_185_4383# a_189_4901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3966 a_26130_n6396# a_26136_n6579# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3967 a_19681_n8347# a_19938_n8363# a_19509_n6125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3968 a_7800_6624# a_8053_6611# a_7003_6396# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3969 a_17533_3194# d0 a_18014_3282# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3970 a_2655_7578# d0 a_3457_7217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3971 a_23001_n4863# a_22795_n5471# a_22215_n5655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3972 a_2423_n5501# d0 a_3216_n5917# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3973 a_27424_n3855# a_27254_n4875# a_27373_n4698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3974 a_11318_8034# d1 a_11417_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3975 a_15727_5403# d0 a_16520_5808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3976 gnd d0 a_25462_8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3977 a_13604_6968# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3978 a_32800_n5141# d1 a_32899_n5551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3979 a_537_n8272# d1 a_1334_n8733# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3980 a_26173_n8615# d0 a_26648_n8721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3981 a_18414_n4440# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3982 a_5024_4301# a_4806_4301# a_4549_4396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3983 a_3167_n2263# a_3420_n2467# a_2365_n2635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3984 a_25011_n8808# a_25025_n9602# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3985 a_19608_n4275# d2 a_19654_n3255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3986 a_2324_n5091# d1 a_2419_n5689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3987 a_4699_n9715# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3988 a_31099_2302# a_30881_2302# a_30618_2214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3989 a_21890_2989# d0 a_22379_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3990 a_20841_8424# a_21098_8234# a_20043_8608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3991 a_9167_2883# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3992 vdd d2 a_28905_5997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3993 a_12832_197# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3994 vdd d0 a_29765_4599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3995 a_6999_6573# d0 a_7797_6389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3996 a_6843_n8568# a_7096_n8772# a_6757_n9364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3997 a_22923_n3843# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3998 a_733_8360# a_515_8360# a_252_8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3999 a_1441_6548# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4000 vdd d2 a_24385_n9392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4001 a_16452_1147# a_16705_1134# a_15650_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4002 a_23214_n7915# a_22996_n7915# a_23120_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4003 a_5810_3628# a_5604_4117# a_5025_3889# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4004 a_1105_n2802# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4005 a_14320_n8948# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4006 a_13284_4238# a_13290_4421# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4007 a_27589_5159# d2 a_27672_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4008 a_11220_n8580# a_11473_n8784# a_11134_n9376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4009 gnd d5 a_19704_n10593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4010 a_24407_8621# a_24664_8431# a_24312_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4011 a_21897_3207# d0 a_22378_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4012 a_21963_7061# d0 a_22452_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4013 a_25008_n8584# a_25012_n8396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4014 a_1229_n2802# d2 a_1307_n3641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4015 a_9168_n2189# a_8950_n2189# a_8236_n2045# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4016 a_661_3876# a_443_3876# a_172_3982# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4017 a_17814_n3606# a_17596_n3606# a_17333_n3317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4018 a_15543_n6745# a_15800_n6761# a_15461_n7353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4019 gnd d0 a_3546_n10005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4020 a_28652_6010# d1 a_28747_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4021 a_12124_3582# a_12377_3569# a_11327_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4022 vdd d1 a_24357_n2676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4023 a_26772_4325# d1 a_27558_3652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4024 a_6904_5986# a_7157_5973# a_6854_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4025 a_16271_n2713# a_16285_n3507# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4026 a_32980_3987# a_33233_3974# a_32897_2971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4027 a_24095_n7152# d1 a_24190_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4028 a_27604_2632# a_27434_3533# a_27553_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4029 a_6900_6163# d1 a_6982_5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4030 a_24117_n3678# a_24374_n3694# a_24022_n3080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4031 vdd d0 a_3690_6186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4032 a_13494_860# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4033 a_26845_8397# d1 a_27631_7724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4034 vdd d0 a_3673_5168# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4035 a_1297_n6697# d2 a_1380_n7713# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4036 a_17887_n7678# a_17669_n7678# a_17412_n7572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4037 a_18476_n2814# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4038 vdd d1 a_11543_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4039 a_20591_n5741# a_20607_n6535# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4040 a_20575_n4311# a_20570_n4911# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4041 a_33929_7444# a_34186_7254# a_33131_7628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4042 a_26592_n5667# d1 a_27378_n4875# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4043 a_18600_n2814# d2 a_18678_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4044 a_25007_n8996# a_25264_n9012# a_24214_n8580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4045 a_142_2164# d0 a_623_2252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4046 a_14624_7725# a_14418_8214# a_13839_7986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4047 a_27425_8213# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4048 gnd d1 a_20120_n9789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4049 a_23300_6692# a_23130_7593# a_23254_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4050 a_8813_n9438# a_8819_n9621# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4051 a_31955_n7940# d4 a_32058_n5902# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4052 a_7796_6801# a_8053_6611# a_7003_6396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4053 a_20010_6395# d0 a_20803_6800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4054 a_2397_n9163# d1 a_2492_n9761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4055 a_9004_n5243# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4056 a_6770_n4496# a_7023_n4700# a_6684_n5292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4057 a_15419_n8185# d2 a_15502_n9201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4058 a_2475_n8743# a_2732_n8759# a_2393_n9351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4059 a_17690_n8284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4060 a_9295_n9315# a_9077_n9315# a_8806_n9220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4061 a_19863_n9773# d0 a_20661_n9589# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4062 a_11903_n2888# a_11907_n2700# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4063 a_21978_7980# d0 a_22469_7973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4064 a_10879_n6138# a_11132_n6342# a_10817_n10590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4065 a_30531_n8445# d0 a_31012_n8734# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4066 a_11147_n4508# a_11400_n4712# a_11061_n5304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4067 a_33025_1343# a_33278_1330# a_32939_2128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4068 a_18668_n6709# d2 a_18751_n7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4069 vdd d5 a_11074_n10606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4070 a_22177_4313# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4071 gnd d0 a_25154_n2904# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4072 gnd d0 a_34165_6648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4073 a_4382_n6372# d0 a_4863_n6661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4074 a_17977_1246# d1 a_18775_1062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4075 a_31789_8226# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4076 a_9874_n9543# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4077 a_4753_835# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4078 gnd d0 a_21044_5180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4079 a_4419_n8408# a_4425_n8591# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4080 a_16448_1324# a_16705_1134# a_15650_1508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4081 a_10147_n3843# d4 a_10323_n5877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4082 a_4091_172# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4083 gnd d1 a_24554_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4084 a_12030_n10014# a_8824_n9945# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4085 gnd d0 a_12288_n9618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4086 a_13729_1878# d1 a_14514_1617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4087 a_11231_7195# d2 a_11281_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4088 a_19768_n9175# d1 a_19863_n9773# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4089 a_9365_1865# a_9147_1865# a_8874_1872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4090 gnd d1 a_2622_n2651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4091 a_4843_5925# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4092 a_13350_8092# a_13357_8310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4093 a_16378_n8597# a_16635_n8613# a_15580_n8781# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4094 a_27714_283# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4095 a_3363_2539# a_3380_3322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4096 a_27672_6585# d3 a_27771_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4097 vdd d0 a_29839_8259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4098 a_23317_n5877# a_23099_n5877# a_23141_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4099 a_1404_1050# a_1186_1050# a_607_822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4100 a_30481_n5574# a_30485_n6092# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4101 a_26719_859# d1 a_27516_1087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4102 a_15667_2526# d0 a_16465_2342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4103 a_29532_5218# a_29527_5807# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4104 a_31834_5582# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4105 a_33098_5415# d0 a_33891_5820# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4106 a_235_7254# a_241_7437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4107 a_6950_3342# a_7203_3329# a_6864_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4108 a_17550_4212# a_17556_4395# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4109 a_18630_5134# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4110 a_6900_6163# d1 a_6986_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4111 a_20647_n8795# a_20661_n9589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4112 a_22395_4313# a_22177_4313# a_21920_4408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4113 a_20661_n9589# a_20665_n9401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4114 a_16308_n4749# a_16322_n5543# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4115 a_5061_5925# d1 a_5846_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4116 a_1395_7568# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4117 a_15465_n7165# d1 a_15564_n7575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4118 a_11143_n4696# d0 a_11945_n4324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4119 a_28567_n7762# d0 a_29365_n7578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4120 a_24271_6175# a_24528_5985# a_24225_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4121 a_11344_4372# d0 a_12137_4777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4122 a_28657_1507# d0 a_29455_1323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4123 a_16502_4378# a_16506_4201# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4124 a_19937_2323# d0 a_20734_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4125 gnd d3 a_24302_n8376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4126 a_1582_n5852# a_2333_n10581# a_2175_n10565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4127 gnd d4 a_6935_4959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4128 a_11051_n8360# a_11308_n8376# a_10879_n6138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4129 a_21703_n3513# a_21708_n4031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4130 gnd d0 a_34076_1146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4131 a_28426_n8184# a_28679_n8388# a_28250_n6150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4132 a_30464_n4556# a_30466_n5074# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4133 gnd d0 a_16525_n2505# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4134 a_32935_n7587# d0 a_33732_n7815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4135 gnd d2 a_28689_n5332# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4136 a_23181_3640# a_22975_4129# a_22396_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4137 a_30865_872# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4138 a_30629_2721# a_30631_3014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4139 a_10043_n6899# d2 a_10121_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4140 a_14511_n3856# a_14293_n3856# a_14412_n3679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4141 a_170_3883# a_172_3982# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4142 a_26447_n9739# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4143 a_3419_5593# a_3672_5580# a_2622_5365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4144 a_29527_5807# a_29531_5630# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4145 gnd d3 a_32970_n4329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4146 a_25119_3170# a_25114_3759# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4147 a_20010_6395# d0 a_20807_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4148 a_3872_n2032# a_4302_n2082# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4149 a_5567_2081# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4150 a_148_2347# a_153_2671# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4151 a_22994_5147# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4152 gnd d0 a_3654_4150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4153 gnd d0 a_21080_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4154 a_9204_n4637# d1 a_10002_n4686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4155 a_14412_n3679# a_14210_n2840# a_14334_n2840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4156 a_32893_3148# d2 a_32939_2128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4157 a_9221_n5655# a_9003_n5655# a_8740_n5366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4158 a_9185_n3207# d1 a_9970_n2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4159 a_18_n6359# a_24_n6542# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4160 a_25135_4600# a_25388_4587# a_24338_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4161 a_6856_n9774# d0 a_7658_n9402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4162 a_17652_n6660# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4163 a_12104_2564# a_12121_3347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4164 a_5676_n3831# d3 a_5770_n3831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4165 a_33021_1520# a_33278_1330# a_32939_2128# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4166 a_118_928# d0 a_607_822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4167 a_15764_7439# a_16017_7426# a_15678_8224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4168 a_28571_n7574# d0 a_29368_n7802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4169 a_26267_3001# a_26274_3219# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4170 a_19850_n8567# a_20103_n8771# a_19764_n9363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4171 a_4339_n4118# d0 a_4828_n4213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4172 a_25208_8672# a_25461_8659# a_24411_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4173 vdd d0 a_21044_5180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4174 vdd d0 a_16524_n2917# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4175 a_11164_n5526# d0 a_11957_n5942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4176 a_18710_n8922# a_18504_n9530# a_17925_n9302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4177 a_28250_n6150# d3 a_28426_n8184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4178 a_33094_5592# a_33351_5402# a_33012_6200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4179 a_26063_n2507# d0 a_26538_n2613# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4180 vdd d1 a_24554_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4181 a_29315_n4748# a_29568_n4952# a_28518_n4520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4182 a_27315_2105# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4183 a_27698_2513# d4 a_27838_402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4184 a_13183_n9634# a_13188_n9958# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4185 a_33025_1343# d0 a_33822_1571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4186 a_15764_7439# d0 a_16557_7844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4187 a_221_6419# a_226_6743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4188 gnd d0 a_3457_n4503# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4189 a_4901_n8285# d1 a_5698_n8746# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4190 a_16284_n3919# a_16541_n3935# a_15491_n3503# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4191 a_13357_8310# a_13363_8493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4192 a_13183_n9634# d0 a_13658_n9740# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4193 a_26063_n2507# a_26065_n3025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4194 a_18780_1591# a_18574_2080# a_17995_1852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4195 a_4536_3995# d0 a_5025_3889# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4196 a_11323_3531# d0 a_12121_3347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4197 a_31953_5172# d2 a_32036_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4198 a_25025_n9602# a_25282_n9618# a_24227_n9786# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4199 a_19916_1482# d0 a_20718_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4200 a_30955_5962# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4201 vdd d2 a_24275_n3284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4202 a_15667_2526# d0 a_16469_2165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4203 a_15609_3975# a_15862_3962# a_15526_2959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4204 vdd d3 a_11415_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4205 a_33098_5415# d0 a_33895_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4206 a_33016_6023# d1 a_33111_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4207 a_4309_172# d7 a_8757_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4208 a_6733_n2460# d0 a_7530_n2688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4209 a_26130_n6396# d0 a_26611_n6685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4210 a_18595_n2637# a_18377_n2404# a_17797_n2588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4211 a_11380_6408# a_11633_6395# a_11281_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4212 a_18549_n6886# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4213 a_1116_n8500# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4214 a_8986_8079# a_8993_8297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4215 a_23001_n4863# a_22795_n5471# a_22216_n5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4216 a_32610_n6351# d3 a_32717_n4125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4217 a_7603_n6760# a_7617_n7554# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4218 a_4050_n10652# a_8501_n10669# a_8343_n10653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4219 a_11110_n2472# d0 a_11907_n2700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4220 a_28657_1507# d0 a_29459_1146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4221 a_17798_n2176# a_17580_n2176# a_17309_n2081# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4222 a_31679_2118# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4223 a_9022_n6673# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4224 vdd d0 a_34076_1146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4225 a_19846_n8755# d0 a_20648_n8383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4226 a_16525_5219# a_16520_5808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4227 a_4699_n9715# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4228 a_25119_3170# a_25372_3157# a_24317_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4229 a_27521_1616# a_27315_2105# a_26735_2289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4230 vdd d0 a_25408_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4231 a_28518_n4520# d0 a_29315_n4748# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4232 a_20841_8424# a_20845_8247# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4233 vdd d5 a_32809_n10631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4234 a_4790_2871# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4235 a_6868_3950# d1 a_6963_4537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4236 a_14485_n7751# a_14283_n6912# a_14407_n6912# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4237 gnd d0 a_25172_n3510# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4238 a_1223_3086# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4239 a_19689_4971# d3 a_19861_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4240 gnd d0 a_25228_n6564# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4241 gnd d1 a_11436_n6748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4242 a_3415_5770# a_3672_5580# a_2622_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4243 a_28188_n10602# d4 a_28250_n6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4244 a_30609_1897# d0 a_31100_1890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4245 a_28432_n5316# d1 a_28518_n4520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4246 vdd d0 a_3654_4150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4247 a_22214_5937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4248 a_32972_n9623# d0 a_30559_n9970# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4249 a_24137_n4696# d0 a_24935_n4512# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4250 a_6823_n7550# a_7076_n7754# a_6724_n7140# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4251 a_23214_n7915# a_22996_n7915# a_23115_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4252 a_1105_n2802# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4253 a_10063_3521# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4254 a_30665_4951# d0 a_31156_4944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4255 a_2496_n9573# d0 a_3289_n9989# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4256 a_17406_n7389# a_17412_n7572# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4257 a_17612_7449# d0 a_18087_7354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4258 a_425_3270# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4259 a_243_7955# d0 a_734_7948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4260 a_11200_n7562# a_11453_n7766# a_11101_n7152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4261 a_25029_n9414# a_25024_n10014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4262 a_3216_n5917# a_3473_n5933# a_2423_n5501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4263 a_24018_n3268# d1 a_24104_n2472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4264 a_21761_n7085# a_21763_n7184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4265 a_13131_n7098# a_13133_n7197# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4266 a_3184_n3281# a_3179_n3881# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4267 a_15760_7616# a_16017_7426# a_15678_8224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4268 a_15419_5174# d3 a_15526_2959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4269 a_4607_7968# a_4609_8067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4270 a_31885_1629# a_31679_2118# a_31099_2302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4271 a_26274_3219# a_26280_3402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4272 a_29347_n6972# a_29351_n6784# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4273 a_6502_n6126# d3 a_6678_n8160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4274 a_33656_n3519# a_33660_n3331# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4275 a_499_6930# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4276 a_8731_n5049# a_8733_n5148# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4277 a_2356_n7315# d1 a_2438_n6707# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4278 a_31953_5172# a_31735_5172# a_31155_5356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4279 a_13548_3914# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4280 a_1178_n6874# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4281 a_22831_n7507# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4282 a_8911_3908# d0 a_9402_3901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4283 vdd d0 a_25227_n6976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4284 a_32943_1951# d1 a_33042_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4285 a_15764_7439# d0 a_16561_7667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4286 a_1302_n6874# d2 a_1380_n7713# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4287 a_31958_5701# a_31752_6190# a_31172_6374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4288 a_28550_n6744# d0 a_29352_n6372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4289 a_22034_n7279# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4290 a_18476_n2814# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4291 a_21976_7462# d0 a_22451_7367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4292 a_7707_1299# a_7711_1122# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4293 gnd d1 a_33135_n4737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4294 a_8757_196# a_8539_196# a_4309_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4295 a_20790_5605# a_21043_5592# a_19993_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4296 vdd d4 a_15496_n6355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4297 vdd d0 a_12468_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4298 a_16289_n3319# a_16284_n3919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4299 a_19790_n5701# a_20047_n5717# a_19695_n5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4300 a_624_1840# d1 a_1409_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4301 gnd d0 a_21025_4162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4302 a_24987_n7978# a_25244_n7994# a_24194_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4303 gnd d0 a_34202_8684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4304 a_31082_1284# a_30864_1284# a_30607_1379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4305 a_33016_6023# d1 a_33115_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4306 a_18015_2870# a_17797_2870# a_17524_2683# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4307 a_14328_3124# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4308 a_33131_7628# d0 a_33929_7444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4309 a_32899_n5551# a_33152_n5755# a_32800_n5141# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4310 a_1487_2476# a_1285_1460# a_1409_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4311 a_19727_n7327# d1 a_19809_n6719# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4312 vdd d2 a_2830_7996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4313 a_32614_n6163# a_32867_n6367# a_32552_n10615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4314 a_19736_n2647# a_19993_n2663# a_19654_n3255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4315 a_11162_2946# d2 a_11245_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4316 a_10099_5557# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4317 a_9458_6955# a_9240_6955# a_8969_7061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4318 a_697_5912# d1 a_1482_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4319 a_9295_n9315# a_9077_n9315# a_8804_n9121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4320 a_29291_n3918# a_29295_n3730# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4321 a_6750_n3478# a_7003_n3682# a_6651_n3068# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4322 a_13766_3914# d1 a_14551_3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4323 a_26111_n5378# d0 a_26592_n5667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4324 a_7003_6396# d0 a_7796_6801# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4325 a_2455_n7725# a_2712_n7741# a_2360_n7127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4326 a_17670_n7266# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4327 a_4880_7961# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4328 a_4825_5319# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4329 a_30537_n8628# d0 a_31012_n8734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4330 a_18014_3282# a_17796_3282# a_17539_3377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4331 a_19813_n6531# d0 a_20610_n6759# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4332 a_30511_n7427# d0 a_30992_n7716# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4333 a_20735_2139# a_20730_2728# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4334 a_32841_n2685# d0 a_33643_n2313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4335 a_4346_n4336# a_4352_n4519# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4336 a_18611_4116# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4337 a_33079_4397# d0 a_33872_4802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4338 a_23042_n3666# a_22840_n2827# a_22964_n2827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4339 a_11208_1926# a_11461_1913# a_11158_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4340 a_4388_n6555# d0 a_4863_n6661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4341 gnd d0 a_12271_n8600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4342 a_10105_n5877# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4343 a_26756_2895# d1 a_27553_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4344 a_18756_n7902# a_18586_n8922# a_18710_n8922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4345 a_9874_n9543# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4346 a_22913_n6899# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4347 a_23456_271# d5 a_21581_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4348 a_133_1847# a_135_1946# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4349 gnd d0 a_7981_2127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4350 vdd d0 a_16598_n6577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4351 a_10220_n7915# d4 a_10323_n5877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4352 a_33822_1571# a_34075_1558# a_33025_1343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4353 a_28533_2958# d2 a_28612_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4354 a_19546_n10577# a_21579_n10680# a_21421_n10664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4355 a_2283_n3243# d1 a_2365_n2635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4356 a_11958_n5530# a_12215_n5546# a_11160_n5714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4357 a_24235_4139# a_24492_3949# a_24156_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4358 a_33950_8285# a_33945_8874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4359 a_20043_8608# a_20300_8418# a_19948_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4360 a_29333_n5354# a_29586_n5558# a_28531_n5726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4361 a_17586_6248# a_17592_6431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4362 gnd d0 a_8037_5181# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4363 a_17029_133# d8 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4364 a_14546_3124# a_14328_3124# a_13748_3308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4365 gnd d1 a_15907_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4366 a_24334_4549# d0 a_25132_4365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4367 gnd d2 a_24565_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4368 a_15547_n6557# d0 a_16344_n6785# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4369 a_26260_2384# d0 a_26735_2289# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4370 gnd d0 a_34113_3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4371 a_16358_n7579# a_16615_n7595# a_15560_n7763# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4372 a_3400_4575# a_3653_4562# a_2603_4347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4373 a_10301_6573# a_10099_5557# a_10223_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4374 vdd d0 a_3689_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4375 a_22272_n8297# a_22054_n8297# a_21783_n8202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4376 a_5043_5319# a_4825_5319# a_4568_5414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4377 a_13320_6274# d0 a_13801_6362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4378 a_22975_4129# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4379 a_6854_7183# d2 a_6900_6163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4380 a_n8_n5123# d0 a_481_n5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4381 a_15723_5580# a_15980_5390# a_15641_6188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4382 a_31173_5962# a_30955_5962# a_30684_6068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4383 a_26320_6055# d0 a_26809_5949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4384 a_6746_n3666# d0 a_7548_n3294# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4385 a_18104_8372# a_17886_8372# a_17623_8284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4386 a_26138_n7097# d0 a_26629_n7291# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4387 a_10916_n10590# d5 a_10817_n10590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4388 gnd d0 a_3492_n6951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4389 a_17849_6336# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4390 a_6802_n6720# d0 a_7604_n6348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4391 a_7783_5606# a_7797_6389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4392 a_19944_8198# d1 a_20030_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4393 a_14592_2514# a_14390_1498# a_14509_1088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4394 a_26628_7985# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4395 a_5744_n7726# a_5542_n6887# a_5666_n6887# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4396 a_11123_n3678# d0 a_11925_n3306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4397 a_26310_5255# d0 a_26791_5343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4398 a_15470_n2673# d0 a_16268_n2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4399 a_22161_2883# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4400 a_15392_n3093# a_15645_n3297# a_15342_n4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4401 a_20591_n5741# a_20844_n5945# a_19794_n5513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4402 a_13801_6362# d1 a_14587_5689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4403 a_13080_n4143# d0 a_13569_n4238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4404 a_4555_5013# d0 a_5044_4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4405 a_23212_5147# d2 a_23295_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4406 a_13320_6274# a_13326_6457# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4407 vdd d0 a_21025_4162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4408 a_10260_7712# a_10054_8201# a_9475_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4409 a_12030_n10014# a_12287_n10030# a_11237_n9598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4410 vdd d0 a_34202_8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4411 a_17346_n4117# a_17353_n4335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4412 a_23020_1485# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4413 a_27470_5569# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4414 a_33131_7628# d0 a_33933_7267# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4415 a_13188_n9958# a_16651_n10043# a_15601_n9611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4416 a_22160_3295# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4417 a_16344_n6785# a_16358_n7579# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4418 a_16326_n5355# a_16321_n5955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4419 a_26791_5343# d1 a_27589_5159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4420 vdd d3 a_28859_7017# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4421 gnd d1 a_33351_5402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4422 a_22468_8385# a_22250_8385# a_21987_8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4423 a_11363_5390# d0 a_12160_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4424 a_9184_n3619# d1 a_9970_n2827# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4425 a_9420_5331# a_9202_5331# a_8939_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4426 a_27352_4141# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4427 a_16325_n5767# a_16578_n5971# a_15528_n5539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4428 a_7003_6396# d0 a_7800_6624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4429 a_23227_2620# a_23057_3521# a_23176_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4430 a_8949_6043# a_8956_6261# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4431 a_3290_n9577# a_3547_n9593# a_2492_n9761# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4432 a_31136_4338# d1 a_31922_3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4433 gnd d2 a_7084_1901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4434 a_16469_2165# a_16464_2754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4435 a_22468_8385# d1 a_23254_7712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4436 a_33079_4397# d0 a_33876_4625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4437 a_189_4901# d0 a_680_4894# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4438 a_17513_2176# d0 a_17994_2264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4439 a_27419_n3678# d3 a_27518_n3855# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4440 vdd d0 a_33913_n3535# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4441 a_15474_n2485# d0 a_16271_n2713# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4442 a_2577_8009# a_2830_7996# a_2494_6993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4443 a_16341_n6561# a_16345_n6373# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4444 gnd d2 a_6977_n7344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4445 a_1224_n2625# a_1006_n2392# a_427_n2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4446 a_8950_n2189# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4447 a_4319_n3100# d0 a_4808_n3195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4448 a_32790_n8197# d2 a_32869_n9401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4449 a_7585_n5330# a_7838_n5534# a_6783_n5702# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4450 a_5950_2489# d4 a_6090_378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4451 gnd d2 a_11354_n7356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4452 a_32878_n4721# d0 a_33680_n4349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4453 a_13294_4939# d0 a_13785_4932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4454 a_11147_n4508# d0 a_11940_n4924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4455 a_25150_5795# a_25407_5605# a_24357_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4456 a_31209_8410# a_30991_8410# a_30734_8505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4457 a_2402_n4671# d0 a_3200_n4487# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4458 a_17539_3377# a_17541_3895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4459 vdd d0 a_8037_5181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4460 a_9365_1865# d1 a_10150_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4461 a_29295_n3730# a_29548_n3934# a_28498_n3502# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4462 a_24334_4549# d0 a_25136_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4463 vdd d2 a_24565_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4464 a_9060_n8297# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4465 a_16541_6649# a_16558_7432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4466 a_19191_258# a_18973_258# a_19092_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4467 a_3384_3145# a_3379_3734# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4468 a_17833_4906# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4469 a_4900_n8697# d1 a_5698_n8746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4470 vdd d0 a_34113_3182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4471 a_19861_7182# d2 a_19911_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4472 a_10400_6573# a_10182_6573# a_10301_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4473 a_30431_n3137# a_30438_n3355# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4474 a_23972_n4288# d2 a_24022_n3080# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4475 gnd d0 a_3437_n3485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4476 a_3396_4752# a_3653_4562# a_2603_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4477 a_27558_3652# a_27352_4141# a_26772_4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4478 a_4570_5932# d0 a_5061_5925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4479 a_4570_5932# a_4572_6031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4480 a_1297_n6697# a_1079_n6464# a_499_n6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4481 a_15528_n5539# d0 a_16325_n5767# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4482 a_21877_2189# d0 a_22358_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4483 a_11245_3962# d1 a_11340_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4484 a_20803_6800# a_20807_6623# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4485 a_3235_n6935# a_3239_n6747# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4486 a_26237_1183# a_26243_1366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4487 a_6757_n9364# a_7014_n9380# a_6678_n8160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4488 a_24374_6408# d0 a_25167_6813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4489 a_22251_7973# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4490 a_18595_n2637# a_18377_n2404# a_17798_n2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4491 a_6909_1483# d0 a_7711_1122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4492 gnd d7 a_25872_n10681# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4493 a_20771_4587# a_20787_5370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4494 a_19834_2090# a_20091_1900# a_19788_3110# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4495 gnd d0 a_16758_4600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4496 a_18051_4906# d1 a_18848_5134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4497 a_28509_n9200# a_28762_n9404# a_28426_n8184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4498 a_13067_n3343# a_13073_n3526# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4499 vdd d2 a_19948_n5307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4500 a_25131_4777# a_25135_4600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4501 a_26648_n8721# a_26430_n8721# a_26173_n8615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4502 a_2622_5365# a_2875_5352# a_2536_6150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4503 a_31815_n8960# d2 a_31861_n7940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4504 a_7580_n5930# a_7837_n5946# a_6787_n5514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4505 a_9022_n6673# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4506 a_19695_n5103# a_19948_n5307# a_19612_n4087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4507 a_10467_390# d5 a_10561_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4508 a_23300_6692# d3 a_23394_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4509 a_5846_5664# a_5640_6153# a_5060_6337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4510 a_26175_n9133# d0 a_26666_n9327# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4511 a_19826_n7737# d0 a_20628_n7365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4512 a_11097_n7340# d1 a_11179_n6732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4513 gnd d0 a_29748_3581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4514 gnd d2 a_33053_n5345# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4515 a_24898_n2476# a_25155_n2492# a_24100_n2660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4516 a_11106_n2660# a_11363_n2676# a_11024_n3268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4517 a_9956_n8935# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4518 a_14485_n7751# a_14283_n6912# a_14402_n6735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4519 a_26447_n9739# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4520 vdd d0 a_3436_n3897# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4521 a_1820_246# d6 a_4309_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4522 a_18668_n6709# a_18450_n6476# a_17870_n6660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4523 a_33732_n7815# a_33749_n8609# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4524 gnd d2 a_6904_n3272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4525 a_21688_n3013# a_21690_n3112# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4526 a_30449_n4056# a_30451_n4155# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4527 a_7621_n7366# a_7616_n7966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4528 a_26808_6361# a_26590_6361# a_26333_6456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4529 a_12210_8849# a_12467_8659# a_11417_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4530 a_27656_4547# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4531 a_63_n9096# a_65_n9195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4532 a_20771_4587# a_21024_4574# a_19974_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4533 a_27553_6585# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4534 a_13093_n4544# a_13095_n5062# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4535 a_5061_5925# a_4843_5925# a_4570_5932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4536 a_20555_n3293# a_20808_n3497# a_19753_n3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4537 gnd d0 a_20901_n8587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4538 a_8956_6261# a_8962_6444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4539 a_32036_6598# d3 a_32135_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4540 a_5810_3628# d2 a_5856_2608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4541 a_29984_n2069# d0 a_30903_n2214# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4542 a_28591_n8592# d0 a_29388_n8820# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4543 a_23032_n6722# a_22814_n6489# a_22235_n6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4544 a_30939_n4662# a_30721_n4662# a_30464_n4556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4545 a_12692_n10677# d5 a_14687_n5890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4546 a_9240_6955# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4547 a_24280_1495# d0 a_25078_1311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4548 a_27594_5688# a_27388_6177# a_26809_5949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4549 a_13346_7475# a_13348_7993# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4550 a_15678_8224# d1 a_15760_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4551 a_4789_3283# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4552 a_1296_7158# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4553 a_19612_n4087# d2 a_19695_n5103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4554 a_24177_n6544# d0 a_24974_n6772# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4555 gnd d0 a_7837_n5946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4556 a_18710_n8922# a_18504_n9530# a_17924_n9714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4557 a_24045_n8360# d2 a_24095_n7152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4558 a_4405_n7573# a_4410_n8091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4559 a_1178_n6874# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4560 a_30956_n5680# a_30738_n5680# a_30475_n5391# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4561 a_22831_n7507# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4562 gnd d0 a_20880_n7981# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4563 a_30738_n5680# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4564 a_28571_n7574# a_28824_n7778# a_28472_n7164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4565 a_14826_284# d4 a_15423_4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4566 a_500_n6236# a_282_n6236# a_11_n6141# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4567 a_33913_6249# a_33908_6838# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4568 gnd d0 a_3673_5168# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4569 a_4862_7355# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4570 a_697_5912# a_479_5912# a_208_6018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4571 gnd d0 a_16742_3170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4572 a_17412_n7572# d0 a_17887_n7678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4573 a_13177_n9451# d0 a_13658_n9740# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4574 gnd d1 a_33115_n3719# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4575 a_27838_402# a_27656_4547# a_27771_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4576 a_32836_n7177# d1 a_32935_n7587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4577 a_31662_1100# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4578 a_19865_7005# d2 a_19944_8198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4579 a_226_6743# a_228_7036# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4580 a_1385_n7890# a_1215_n8910# a_1334_n8733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4581 a_24897_n2888# a_24901_n2700# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4582 a_3453_7394# a_3457_7217# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4583 a_3235_n6935# a_3492_n6951# a_2442_n6519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4584 a_13168_n9134# a_13170_n9233# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4585 a_19753_n3665# d0 a_20555_n3293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4586 a_7783_5606# a_8036_5593# a_6986_5378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4587 a_11907_n2700# a_12160_n2904# a_11110_n2472# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4588 a_12121_3347# a_12378_3157# a_11323_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4589 a_17871_n6248# a_17653_n6248# a_17380_n6054# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4590 a_5025_3889# a_4807_3889# a_4534_3896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4591 a_2438_n6707# a_2695_n6723# a_2356_n7315# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4592 a_24374_6408# d0 a_25171_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4593 gnd d0 a_8018_4163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4594 a_4844_n5643# a_4626_n5643# a_4369_n5537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4595 a_25607_n2057# a_26050_n2106# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4596 a_9965_n2650# d2 a_10048_n3666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4597 a_14707_284# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4598 a_33859_3607# a_34112_3594# a_33062_3379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4599 a_33659_n3743# a_33912_n3947# a_32862_n3515# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4600 a_26374_n5667# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4601 a_14584_n7928# d4 a_14687_n5890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4602 a_1514_7158# a_1296_7158# a_716_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4603 a_24132_n9188# d1 a_24231_n9598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4604 a_2421_2921# d2 a_2504_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4605 a_2618_5542# a_2875_5352# a_2536_6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4606 a_19948_8021# a_20201_8008# a_19865_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4607 a_26117_n5561# d0 a_26592_n5667# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4608 a_26792_4931# a_26574_4931# a_26303_5037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4609 a_17670_n7266# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4610 gnd d1 a_33208_n8809# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4611 a_12194_7419# a_12451_7229# a_11396_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4612 a_32717_n4125# a_32970_n4329# a_32610_n6351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4613 a_12613_n2057# a_13043_n2107# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4614 a_6733_n2460# a_6986_n2664# a_6647_n3256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4615 a_26177_n9232# a_26184_n9450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4616 a_30517_n7610# d0 a_30992_n7716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4617 vdd d0 a_29748_3581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4618 gnd d1 a_28968_4371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4619 a_29528_5395# a_29532_5218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4620 a_11941_n4512# a_12198_n4528# a_11143_n4696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4621 a_23042_n3666# a_22840_n2827# a_22959_n2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4622 a_21703_n3513# d0 a_22178_n3619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4623 a_31082_1284# d1 a_31880_1100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4624 a_5805_3099# a_5587_3099# a_5008_2871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4625 a_18756_n7902# a_18586_n8922# a_18705_n8745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4626 a_24955_n5754# a_25208_n5958# a_24158_n5526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4627 a_10105_n5877# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4628 a_26338_n3219# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4629 a_1477_5122# d2 a_1560_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4630 a_24154_n5714# d0 a_24952_n5530# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4631 gnd d0 a_12251_n7582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4632 a_31155_5356# a_30937_5356# a_30674_5268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4633 gnd d0 a_12357_2551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4634 a_17886_8372# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4635 a_28518_n4520# a_28771_n4724# a_28432_n5316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4636 a_2540_5973# d1 a_2635_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4637 a_8857_854# d0 a_9348_847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4638 a_21897_3207# a_21903_3390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4639 a_20767_4764# a_21024_4574# a_19974_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4640 a_8956_6261# d0 a_9437_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4641 a_5625_n4674# d2 a_5676_n3831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4642 gnd d0 a_20807_n3909# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4643 a_13839_7986# a_13621_7986# a_13348_7993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4644 a_14687_n5890# a_15438_n10619# a_12692_n10677# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4645 gnd d2 a_19984_n7343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4646 a_29532_5218# a_29785_5205# a_28730_5579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4647 a_24280_1495# d0 a_25082_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4648 a_19777_n4495# d0 a_20570_n4911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4649 a_21770_n7402# d0 a_22251_n7691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4650 a_30811_n9752# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4651 gnd d3 a_19865_n4291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4652 a_22252_n7279# a_22034_n7279# a_21763_n7184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4653 a_1261_n7890# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4654 a_18684_8188# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4655 a_15678_8224# d1 a_15764_7439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4656 gnd d0 a_29839_8259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4657 a_26628_n7703# d1 a_27414_n6911# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4658 gnd d1 a_7113_n9790# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4659 a_1312_n3818# a_1142_n4838# a_1261_n4661# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4660 a_7797_6389# a_7801_6212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4661 a_9401_4313# a_9183_4313# a_8920_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4662 a_26829_6967# a_26611_6967# a_26338_6780# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4663 a_5649_1473# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4664 a_19993_5377# a_20246_5364# a_19907_6162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4665 a_26282_3920# a_26284_4019# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4666 gnd d3 a_24409_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4667 a_13838_8398# a_13620_8398# a_13363_8493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4668 a_17524_2683# a_17526_2976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4669 a_33855_3784# a_33859_3607# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4670 a_13348_7993# a_13350_8092# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4671 a_24353_5567# d0 a_25155_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4672 gnd d1 a_33405_8456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4673 a_17614_7967# d0 a_18105_7960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4674 a_24158_n5526# d0 a_24955_n5754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4675 a_9927_1075# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4676 vdd d0 a_16742_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4677 a_26370_8492# a_25208_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4678 a_14619_7196# a_14401_7196# a_13822_6968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4679 a_12692_n10677# a_12949_n10693# a_8244_n10653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4680 a_6937_8199# d1 a_7023_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4681 a_19937_2323# d0 a_20730_2728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4682 a_11976_n6960# a_11980_n6772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4683 a_13060_n3125# d0 a_13549_n3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4684 a_29385_n8596# a_29389_n8408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4685 gnd d0 a_33950_n5571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4686 a_24059_n5116# d1 a_24158_n5526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4687 a_5722_5545# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4688 a_13294_4939# a_13296_5038# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4689 a_5043_5319# d1 a_5841_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4690 a_19993_5377# d0 a_20786_5782# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4691 a_13275_3921# d0 a_13766_3914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4692 vdd d0 a_8018_4163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4693 gnd d0 a_7801_n3498# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4694 a_10000_5147# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4695 a_21725_n5049# a_21727_n5148# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4696 vdd d0 a_3510_n7557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4697 a_26719_859# a_26501_859# a_26228_866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4698 a_19861_7182# a_20118_6992# a_19689_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4699 a_30919_n3644# d1 a_31705_n2852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4700 a_23031_7183# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4701 a_3166_n2675# a_3180_n3469# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4702 a_14587_5689# d2 a_14665_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4703 a_13238_1885# d0 a_13729_1878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4704 a_17814_3888# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4705 gnd d2 a_11534_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4706 a_26265_2708# d0 a_26756_2895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4707 gnd d0 a_20971_1108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4708 a_18729_5544# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4709 a_29311_n4936# a_29315_n4748# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4710 a_17870_6942# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4711 vdd d1 a_28968_4371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4712 a_28604_n9798# d0 a_29406_n9426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4713 a_17359_n4518# a_17361_n5036# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4714 a_21717_n4348# d0 a_22198_n4637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4715 a_27424_n3855# d3 a_27518_n3855# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4716 a_11051_n8360# d2 a_11097_n7340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4717 a_13749_2896# a_13531_2896# a_13260_3002# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4718 a_33643_n2313# a_33896_n2517# a_32841_n2685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4719 a_3163_n2451# a_3167_n2263# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4720 a_11024_n3268# a_11281_n3284# a_10978_n4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4721 gnd d1 a_24537_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4722 a_12160_5618# a_12174_6401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4723 vdd d0 a_12357_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4724 a_18953_n5864# a_19704_n10593# a_19546_n10577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4725 a_2540_5973# d1 a_2639_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4726 a_2603_4347# a_2856_4334# a_2504_3937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4727 a_5424_n5459# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4728 a_17148_133# d8 a_17217_n720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4729 a_11127_n3490# d0 a_11920_n3906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4730 a_11413_8621# d0 a_12215_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4731 a_10182_3111# a_9964_3111# a_9384_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4732 a_2382_n3653# d0 a_3180_n3469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4733 a_1203_2068# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4734 a_33025_1343# d0 a_33818_1748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4735 a_9846_n2827# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4736 gnd d1 a_7183_2311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4737 a_10080_n8935# a_9874_n9543# a_9294_n9727# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4738 a_4880_n7679# d1 a_5666_n6887# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4739 a_1659_6548# a_1441_6548# a_1560_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4740 a_29984_n2069# a_29275_n2488# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4741 a_13785_4932# d1 a_14582_5160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4742 a_15568_2116# a_15825_1926# a_15522_3136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4743 a_1297_n6697# a_1079_n6464# a_500_n6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4744 a_18931_6560# a_18729_5544# a_18853_5663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4745 gnd d2 a_28725_n7368# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4746 a_13290_4421# a_13294_4939# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4747 a_20787_5370# a_20791_5193# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4748 vdd d0 a_29532_n2504# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4749 a_15595_7208# d2 a_15641_6188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4750 a_19989_5554# a_20246_5364# a_19907_6162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4751 a_11981_n6360# a_12234_n6564# a_11179_n6732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4752 a_n10_n5024# d0 a_481_n5218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4753 a_16977_n2070# a_16268_n2489# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4754 a_18780_1591# d2 a_18858_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4755 a_4918_n9303# a_4700_n9303# a_4429_n9208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4756 a_16321_n5955# a_16325_n5767# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4757 a_25205_8437# a_25462_8247# a_24407_8621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4758 a_22379_2883# d1 a_23176_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4759 vdd d1 a_33405_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4760 a_30444_n3538# a_30449_n4056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4761 a_4970_1247# a_4752_1247# a_4489_1159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4762 a_30991_8410# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4763 a_3346_1521# a_3599_1508# a_2549_1293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4764 a_22451_7367# a_22233_7367# a_21976_7462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4765 a_26648_n8721# a_26430_n8721# a_26167_n8432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4766 vdd d6 a_4208_n10668# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4767 a_32041_6717# a_31871_7618# a_31990_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4768 a_26628_n7703# a_26410_n7703# a_26153_n7597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4769 a_6827_2091# a_7084_1901# a_6781_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4770 a_26177_n9232# d0 a_26666_n9327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4771 a_13078_n4044# d0 a_13569_n4238# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4772 vdd d3 a_24482_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4773 a_4482_941# a_4489_1159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4774 a_17776_2264# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4775 a_2386_n3465# d0 a_3183_n3693# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4776 a_9956_n8935# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4777 a_2490_7170# a_2747_6980# a_2318_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4778 a_32794_5009# d3 a_32966_7220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4779 a_19911_5985# d1 a_20006_6572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4780 a_5908_4523# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4781 a_478_6324# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4782 a_30940_n4250# d1 a_31737_n4711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4783 a_16488_3595# a_16741_3582# a_15691_3367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4784 a_18668_n6709# a_18450_n6476# a_17871_n6248# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4785 a_118_928# a_125_1146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4786 vdd d1 a_11490_n9802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4787 a_2134_n6301# d3 a_2241_n4075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4788 a_26518_1877# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4789 a_7641_n8384# a_7894_n8588# a_6839_n8756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4790 a_7567_n4724# a_7581_n5518# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4791 a_10218_5147# a_10000_5147# a_9421_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4792 a_10817_n10590# a_11074_n10606# a_10916_n10590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4793 a_11976_n6960# a_12233_n6976# a_11183_n6544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4794 a_15461_n7353# d1 a_15547_n6557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4795 a_679_5306# a_461_5306# a_198_5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4796 a_13583_6362# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4797 a_6678_5149# a_6935_4959# a_6085_259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4798 a_30956_n5680# d1 a_31742_n4888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4799 a_30414_n2119# d0 a_30903_n2214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4800 a_7764_4588# a_8017_4575# a_6967_4360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4801 a_30939_n4662# a_30721_n4662# a_30458_n4373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4802 a_27409_n6734# d2 a_27492_n7750# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4803 a_26517_2289# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4804 a_26591_5949# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4805 a_30919_n3644# a_30701_n3644# a_30444_n3538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4806 a_20718_1121# a_20713_1710# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4807 a_31922_3665# a_31716_4154# a_31137_3926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4808 a_3415_5770# a_3419_5593# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4809 a_21914_4225# a_21920_4408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4810 a_24338_4372# d0 a_25135_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4811 a_2455_n7725# d0 a_3253_n7541# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4812 a_30485_n6092# a_30487_n6191# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4813 a_13784_5344# a_13566_5344# a_13303_5256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4814 a_16271_n2713# a_16524_n2917# a_15474_n2485# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4815 a_26573_5343# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4816 a_17577_5931# a_17579_6030# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4817 a_27298_1087# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4818 a_17994_2264# a_17776_2264# a_17519_2359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4819 a_26576_n4237# d1 a_27373_n4698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4820 a_2599_4524# a_2856_4334# a_2504_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4821 a_14381_6178# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4822 a_31880_1100# d2 a_31963_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4823 a_24_n6542# d0 a_499_n6648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4824 a_26228_866# a_29455_1323# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4825 a_26773_3913# a_26555_3913# a_26284_4019# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4826 a_6605_n4088# d2 a_6684_n5292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4827 vdd d0 a_25265_n8600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4828 a_500_n6236# a_282_n6236# a_9_n6042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4829 a_15474_n2485# a_15727_n2689# a_15388_n3281# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4830 a_23093_5557# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4831 a_19505_n6313# d3 a_19612_n4087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4832 a_32943_1951# d1 a_33038_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4833 vdd d1 a_7183_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4834 a_26736_1877# a_26518_1877# a_26247_1983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4835 a_17569_5230# a_17575_5413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4836 a_7658_n9402# a_7653_n10002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4837 a_30485_n6092# d0 a_30976_n6286# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4838 a_21970_7279# a_21976_7462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4839 a_17434_n9108# d0 a_17925_n9302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4840 a_27371_5159# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4841 vdd d2 a_20164_5972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4842 a_33012_6200# d1 a_33094_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4843 a_19030_6560# a_18812_6560# a_18931_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4844 a_26575_n4649# a_26357_n4649# a_26094_n4360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4845 a_17560_4913# d0 a_18051_4906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4846 gnd d0 a_12468_8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4847 a_11233_n9786# a_11490_n9802# a_11138_n9188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4848 a_26555_n3631# a_26337_n3631# a_26080_n3525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4849 a_9239_7367# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4850 a_28353_n4112# a_28606_n4316# a_28246_n6338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4851 a_31700_n2675# d2 a_31783_n3691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4852 a_14469_n5890# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4853 a_335_n9702# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4854 a_30063_n10689# d5 a_32058_n5902# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4855 a_4844_n5643# a_4626_n5643# a_4363_n5354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4856 a_1492_2595# a_1322_3496# a_1441_3086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4857 gnd d0 a_29585_n5970# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4858 a_9970_n2827# d2 a_10048_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4859 a_26374_n5667# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4860 a_33818_1748# a_33822_1571# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4861 a_15528_n5539# a_15781_n5743# a_15429_n5129# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4862 a_462_4894# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4863 a_29513_4200# a_29766_4187# a_28711_4561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4864 a_30607_1379# a_30609_1897# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4865 a_31810_n8783# d2 a_31861_n7940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4866 a_11061_n5304# d1 a_11143_n4696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4867 a_13423_n8722# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4868 gnd d1 a_33188_n7791# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4869 gnd d1 a_7059_n6736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4870 a_172_3982# a_179_4200# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4871 a_3256_n7765# a_3273_n8559# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4872 a_33908_6838# a_34165_6648# a_33115_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4873 a_8945_5426# a_8947_5944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4874 a_32794_5009# d3 a_32970_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4875 a_19974_4359# a_20227_4346# a_19875_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4876 a_19911_5985# d1 a_20010_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4877 a_21725_n5049# d0 a_22216_n5243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4878 a_25910_208# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4879 a_11921_n3494# a_12178_n3510# a_11123_n3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4880 vdd d0 a_3456_n4915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4881 a_7748_3158# a_8001_3145# a_6946_3519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4882 a_16484_3772# a_16741_3582# a_15691_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4883 vdd d1 a_15997_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4884 a_24934_n4924# a_24938_n4736# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4885 a_5506_n4851# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4886 a_28529_3135# d2 a_28579_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4887 a_12083_1723# a_12087_1546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4888 a_2406_n4483# a_2659_n4687# a_2320_n5279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4889 a_20804_6388# a_21061_6198# a_20006_6572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4890 a_7603_n6760# a_7856_n6964# a_6806_n6532# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4891 a_5630_n4851# d2 a_5676_n3831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4892 a_20047_8431# a_20300_8418# a_19948_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4893 a_20575_n4311# a_20828_n4515# a_19773_n4683# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4894 a_26190_n9633# a_26195_n9957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4895 a_18051_4906# a_17833_4906# a_17560_4913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4896 a_2672_8596# d0 a_3470_8412# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4897 vdd d0 a_25192_n4528# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4898 vdd d1 a_28987_5389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4899 a_19764_n9363# d1 a_19850_n8567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4900 a_3199_n4899# a_3203_n4711# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4901 a_7760_4765# a_8017_4575# a_6967_4360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4902 a_19974_4359# d0 a_20767_4764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4903 a_27208_n7519# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4904 a_30811_n9752# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4905 a_170_3883# d0 a_661_3876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4906 a_2639_6383# d0 a_3432_6788# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4907 a_6783_n5702# a_7040_n5718# a_6688_n5104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4908 a_9981_4129# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4909 a_5856_2608# a_5686_3509# a_5805_3099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4910 a_15708_4385# d0 a_16501_4790# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4911 a_13078_n4044# a_13080_n4143# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4912 a_13273_3403# d0 a_13748_3308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4913 a_13531_n2614# d1 a_14329_n2663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4914 a_17322_n2482# d0 a_17797_n2588# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4915 a_12087_1546# a_12340_1533# a_11290_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4916 a_245_8054# a_252_8272# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4917 a_31968_2645# d3 a_32062_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4918 a_6678_5149# d3 a_6781_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4919 a_10462_271# d4 a_11059_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4920 a_28591_n8592# a_28844_n8796# a_28505_n9388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4921 vdd d1 a_20030_n4699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4922 a_29491_3771# a_29495_3594# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4923 a_28698_3366# d0 a_29491_3771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4924 a_6986_5378# a_7239_5365# a_6900_6163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4925 a_13604_6968# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4926 a_18766_7580# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4927 a_24275_5998# d1 a_24374_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4928 a_17432_n8590# d0 a_17907_n8696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4929 a_24141_n4508# d0 a_24938_n4736# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4930 a_2320_n5279# d1 a_2406_n4483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4931 a_26087_n4142# a_26094_n4360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4932 a_23279_4535# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4933 gnd d0 a_25444_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4934 a_33062_3379# a_33315_3366# a_32976_4164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4935 a_1385_n7890# a_1215_n8910# a_1339_n8910# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4936 a_643_3270# a_425_3270# a_168_3365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4937 a_20570_n4911# a_20827_n4927# a_19777_n4495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4938 a_30684_n2626# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4939 a_19773_n4683# d0 a_20575_n4311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4940 a_19097_377# a_18915_4522# a_19030_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4941 a_31499_n3460# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4942 a_32058_n5902# a_32809_n10631# a_30063_n10689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4943 gnd d1 a_6986_n2664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4944 a_17871_n6248# a_17653_n6248# a_17382_n6153# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4945 a_25132_4365# a_25136_4188# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4946 a_24049_5161# a_24306_4971# a_23456_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4947 gnd d3 a_28859_7017# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4948 a_33679_n4761# a_33932_n4965# a_32882_n4533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4949 vdd d0 a_25352_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4950 a_29352_n6372# a_29347_n6972# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4951 a_23217_5676# a_23011_6165# a_22432_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4952 gnd d4 a_33047_4996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4953 a_6986_5378# d0 a_7779_5783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4954 a_14670_6705# a_14500_7606# a_14619_7196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4955 a_17309_n2081# a_17316_n2299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4956 a_33062_3379# d0 a_33855_3784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4957 a_4326_n3318# a_4332_n3501# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4958 a_27507_7605# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4959 a_26539_n2201# a_26321_n2201# a_26050_n2106# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4960 a_2545_1470# d0 a_3343_1286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4961 a_18068_5924# a_17850_5924# a_17579_6030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4962 gnd d1 a_11560_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4963 a_19970_4536# a_20227_4346# a_19875_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4964 a_21723_n4531# d0 a_22198_n4637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4965 a_25615_n10665# d6 a_28287_n10602# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4966 gnd d0 a_29569_n4540# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4967 a_19691_n5291# d1 a_19777_n4495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4968 a_21697_n3330# d0 a_22178_n3619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4969 a_7744_3335# a_8001_3145# a_6946_3519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4970 a_19953_3518# d0 a_20751_3334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4971 a_20648_n8383# a_20901_n8587# a_19846_n8755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4972 a_23461_390# a_23279_4535# a_23394_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4973 a_24091_n7340# d1 a_24177_n6544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4974 a_26338_n3219# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4975 vdd d0 a_16542_n3523# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4976 a_8947_5944# a_8949_6043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4977 gnd d4 a_6755_n6330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4978 a_26121_n6079# a_26123_n6178# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4979 a_9348_847# a_9130_847# a_8859_953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4980 a_17616_8066# d0 a_18105_7960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4981 a_28250_n6150# a_28503_n6354# a_28188_n10602# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4982 a_2672_8596# d0 a_3474_8235# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4983 a_3951_n10652# d5 a_5946_n5865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4984 a_9846_n2827# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4985 a_6864_4127# a_7121_3937# a_6785_2934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4986 a_19974_4359# d0 a_20771_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4987 a_30531_n8445# a_30537_n8628# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4988 a_27228_n8537# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4989 a_10080_n8935# a_9874_n9543# a_9295_n9315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4990 a_28422_n8372# d2 a_28468_n7352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4991 a_20627_n7777# a_20880_n7981# a_19830_n7549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4992 a_28477_n2672# d0 a_29279_n2300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4993 a_28395_n3280# a_28652_n3296# a_28349_n4300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4994 a_3400_4575# a_3416_5358# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4995 vdd d1 a_11380_n3694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X4996 a_8889_2372# d0 a_9364_2277# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4997 a_20587_n5929# a_20591_n5741# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X4998 a_33716_n6385# a_33969_n6589# a_32914_n6757# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4999 a_28678_2348# a_28931_2335# a_28579_1938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5000 a_26629_n7291# d1 a_27414_n6911# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5001 a_12083_1723# a_12340_1533# a_11290_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5002 a_3359_2716# a_3363_2539# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5003 a_27518_n3855# d4 a_27694_n5889# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5004 a_1312_n3818# a_1142_n4838# a_1266_n4838# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5005 vdd d0 a_25371_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5006 a_14509_1088# d2 a_14592_2514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5007 a_7723_2729# a_7980_2539# a_6930_2324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5008 a_4682_n8697# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5009 a_31737_n7940# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5010 a_10187_3640# a_9981_4129# a_9402_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5011 a_553_n9702# d1 a_1339_n8910# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5012 a_4918_n9303# a_4700_n9303# a_4427_n9109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5013 a_18087_7354# d1 a_18885_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5014 a_6720_n7328# a_6977_n7344# a_6674_n8348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5015 a_28698_3366# d0 a_29495_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5016 a_21753_n6384# a_21759_n6567# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5017 a_19863_n9773# a_20120_n9789# a_19768_n9175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5018 a_9146_2277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5019 a_6982_5555# a_7239_5365# a_6900_6163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5020 vdd d0 a_12270_n9012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5021 a_31840_n5902# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5022 a_10255_7183# a_10037_7183# a_9458_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5023 a_21980_8079# d0 a_22469_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5024 a_9919_n6899# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5025 a_29279_n2300# a_29274_n2900# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5026 a_9040_n7279# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5027 a_26628_n7703# a_26410_n7703# a_26147_n7414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5028 a_2318_4959# a_2571_4946# a_1721_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5029 vdd d0 a_25444_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5030 a_33058_3556# a_33315_3366# a_32976_4164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5031 a_15641_6188# d1 a_15723_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5032 a_30691_6286# a_30697_6469# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5033 a_13765_4326# a_13547_4326# a_13284_4238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5034 a_13058_n3026# d0 a_13549_n3220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5035 a_26554_4325# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5036 a_679_5306# d1 a_1477_5122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5037 a_14444_n8948# d2 a_14490_n7928# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5038 a_29328_n5954# a_29585_n5970# a_28535_n5538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5039 a_9347_1259# a_9129_1259# a_8866_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5040 a_7747_3570# a_7761_4353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5041 a_31519_n4478# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5042 a_4646_n6249# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5043 a_24158_n5526# a_24411_n5730# a_24059_n5116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5044 a_32713_n4313# d2 a_32759_n3293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5045 a_30655_4250# d0 a_31136_4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5046 gnd d0 a_16561_n4953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5047 vdd d0 a_3474_n5521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5048 gnd d0 a_7821_n4516# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5049 gnd d0 a_20970_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5050 a_21987_8297# d0 a_22468_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5051 vdd d0 a_3530_n8575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5052 a_11961_n5754# a_11977_n6548# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5053 a_7833_8837# a_7837_8660# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5054 a_30920_n3232# d1 a_31705_n2852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5055 a_6904_5986# d1 a_6999_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5056 a_26755_3307# a_26537_3307# a_26274_3219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5057 a_32931_n7775# a_33188_n7791# a_32836_n7177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5058 a_13586_n5256# d1 a_14371_n4876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5059 a_13712_860# a_13494_860# a_13221_867# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5060 a_7621_n7366# a_7874_n7570# a_6819_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5061 gnd d0 a_33896_n2517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5062 a_17978_834# a_17760_834# a_17487_841# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5063 a_12214_8672# a_12467_8659# a_11417_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5064 a_32914_n6757# d0 a_33716_n6385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5065 a_22451_7367# d1 a_23249_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5066 a_32980_3987# d1 a_33075_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5067 vdd d0 a_3600_1096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5068 a_26431_n8309# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5069 a_4843_5925# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5070 a_17382_n6153# d0 a_17871_n6248# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5071 vdd d1 a_11560_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5072 a_29984_n2069# a_30414_n2119# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5073 a_25082_1134# a_25077_1723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5074 a_72_n9413# a_78_n9596# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5075 a_15423_4997# d3 a_15599_7031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5076 gnd d0 a_16794_6636# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5077 a_27414_n6911# d2 a_27492_n7750# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5078 a_33765_n10039# a_30559_n9970# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5079 a_25098_2564# a_25351_2551# a_24301_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5080 a_5625_n4674# a_5407_n4441# a_4827_n4625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5081 a_24049_5161# d3 a_24152_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5082 a_30919_n3644# a_30701_n3644# a_30438_n3355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5083 a_10228_2501# d3 a_10327_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5084 a_13585_n5668# a_13367_n5668# a_13104_n5379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5085 gnd d3 a_2674_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5086 a_27155_n4465# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5087 a_12613_n2057# d0 a_13532_n2202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5088 a_19953_3518# d0 a_20755_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5089 vdd d1 a_11616_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5090 a_24210_n8768# d0 a_25012_n8396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5091 a_9348_847# d1 a_10145_1075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5092 a_26575_n4649# d1 a_27373_n4698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5093 vdd d2 a_2720_1888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5094 a_29527_5807# a_29784_5617# a_28734_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5095 vdd d1 a_11633_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5096 a_46_n8078# d0 a_537_n8272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5097 a_7585_n5330# a_7580_n5930# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5098 a_26556_n3219# d1 a_27341_n2839# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5099 a_22958_3111# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5100 a_5424_n5459# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5101 a_10400_6573# d4 a_10467_390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5102 a_17217_n720# a_17029_133# a_8757_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5103 a_2324_n5091# a_2577_n5295# a_2241_n4075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5104 vdd d0 a_29766_4187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5105 vdd d1 a_11453_n7766# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5106 vdd d0 a_25245_n7582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5107 a_31193_6980# d1 a_31990_7208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5108 gnd d1 a_15800_n6761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5109 vdd d0 a_7820_n4928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5110 a_31664_n3868# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5111 a_406_1840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5112 a_5623_5135# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5113 a_6647_n3256# a_6904_n3272# a_6601_n4276# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5114 a_17436_n9207# d0 a_17925_n9302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5115 a_65_n9195# d0 a_554_n9290# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5116 a_32970_7043# d2 a_33049_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5117 vdd d2 a_7194_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5118 a_10561_271# a_10343_271# a_10462_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5119 a_21243_n2044# a_20534_n2463# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5120 a_30722_n4250# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5121 a_21888_2696# d0 a_22379_2883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5122 a_28674_2525# a_28931_2335# a_28579_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5123 a_14463_5570# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5124 a_26555_n3631# a_26337_n3631# a_26074_n3342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5125 gnd d0 a_33968_n7001# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5126 a_30702_n3232# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5127 a_18973_258# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5128 a_13511_1878# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5129 a_29508_4789# a_29512_4612# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5130 a_33856_3372# a_33860_3195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5131 a_4971_835# a_4753_835# a_4482_941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5132 a_31705_n2852# d2 a_31783_n3691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5133 vdd d2 a_7157_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5134 a_335_n9702# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5135 a_12125_3170# a_12378_3157# a_11323_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5136 a_20828_7229# a_20823_7818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5137 a_33697_n5367# a_33950_n5571# a_32895_n5739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5138 a_13153_n8215# d0 a_13642_n8310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5139 gnd d2 a_15898_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5140 vdd d2 a_33233_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5141 a_33115_6433# a_33368_6420# a_33016_6023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5142 a_18858_2488# a_18656_1472# a_18775_1062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5143 a_32858_n3703# a_33115_n3719# a_32763_n3105# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5144 a_7548_n3294# a_7801_n3498# a_6746_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5145 gnd d0 a_7894_n8588# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5146 a_15691_3367# a_15944_3354# a_15605_4152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5147 a_13423_n8722# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5148 a_27932_283# a_27714_283# a_27833_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5149 a_12198_7242# a_12451_7229# a_11396_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5150 a_11028_n3080# d1 a_11123_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5151 a_13403_n7704# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5152 a_12031_n9602# a_12035_n9414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5153 a_2406_n4483# d0 a_3203_n4711# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5154 a_24095_n7152# a_24348_n7356# a_24045_n8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5155 a_20734_2551# a_20751_3334# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5156 a_5841_5135# a_5623_5135# a_5043_5319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5157 a_21727_n5148# d0 a_22216_n5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5158 a_6781_3111# d2 a_6831_1914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5159 a_4526_3195# a_4532_3378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5160 vdd d0 a_20970_1520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5161 a_15522_3136# d2 a_15568_2116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5162 a_5506_n4851# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5163 gnd d4 a_15676_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5164 a_6904_5986# d1 a_7003_6396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5165 a_30937_5356# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5166 a_18647_6152# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5167 a_20823_7818# a_20827_7641# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5168 a_13073_n3526# a_13078_n4044# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5169 a_12120_3759# a_12124_3582# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5170 a_11220_n8580# d0 a_12013_n8996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5171 a_4683_n8285# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5172 a_2386_n3465# a_2639_n3669# a_2287_n3055# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5173 a_15601_n9611# a_15854_n9815# a_15502_n9201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5174 gnd d0 a_7873_n7982# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5175 a_21462_184# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5176 a_13223_966# a_13230_1184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5177 a_27599_2513# a_27397_1497# a_27521_1616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5178 a_32980_3987# d1 a_33079_4397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5179 a_48_n8177# a_55_n8395# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5180 a_10126_n7915# a_9956_n8935# a_10080_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5181 a_22289_n9315# d1 a_23074_n8935# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5182 a_5666_n6887# d2 a_5744_n7726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5183 a_7797_6389# a_8054_6199# a_6999_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5184 a_1482_5651# a_1276_6140# a_697_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5185 vdd d0 a_21043_5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5186 a_26393_n6685# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5187 a_18848_5134# a_18630_5134# a_18051_4906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5188 vdd d0 a_16794_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5189 a_33696_n5779# a_33712_n6573# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5190 a_19731_n7139# d1 a_19830_n7549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5191 a_25094_2741# a_25351_2551# a_24301_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5192 a_32955_n8605# d0 a_33748_n9021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5193 a_17579_n2588# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5194 a_33873_4390# a_34130_4200# a_33075_4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5195 a_3276_n8783# a_3529_n8987# a_2479_n8555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5196 a_17363_n5135# d0 a_17852_n5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5197 a_6757_n9364# d1 a_6839_n8756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5198 a_24970_n6960# a_24974_n6772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5199 a_2475_n8743# d0 a_3273_n8559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5200 a_142_2164# a_148_2347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5201 a_2397_n9163# a_2650_n9367# a_2314_n8147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5202 a_15522_3136# a_15779_2946# a_15419_5174# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5203 a_6967_4360# d0 a_7760_4765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5204 a_17344_n4018# d0 a_17835_n4212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5205 a_2318_4959# d3 a_2490_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5206 a_18_n6359# d0 a_499_n6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5207 gnd d2 a_2757_3924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5208 a_262_n5630# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5209 gnd d0 a_34166_6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5210 vdd d1 a_20010_n3681# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5211 a_31963_2526# a_31761_1510# a_31885_1629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5212 a_22140_2277# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5213 a_116_829# a_3343_1286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5214 a_32970_7043# d2 a_33053_8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5215 a_20538_n2275# a_20791_n2479# a_19736_n2647# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5216 a_13114_n6080# a_13116_n6179# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5217 a_2287_n3055# d1 a_2386_n3465# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5218 a_30607_1379# d0 a_31082_1284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5219 a_26575_n4649# a_26357_n4649# a_26100_n4543# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5220 a_30684_n2626# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5221 a_2175_n10565# d5 a_2076_n10565# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5222 a_13350_n4650# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5223 a_25150_5795# a_25154_5618# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5224 a_20550_n3893# a_20807_n3909# a_19757_n3477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5225 vdd d0 a_20900_n8999# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5226 gnd d0 a_16579_n5559# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5227 a_13802_5950# a_13584_5950# a_13313_6056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5228 a_22214_5937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5229 a_10038_n6722# a_9820_n6489# a_9240_n6673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5230 a_33111_6610# a_33368_6420# a_33016_6023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5231 a_30667_5050# d0 a_31156_4944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5232 a_2479_n8555# d0 a_3276_n8783# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5233 a_245_8054# d0 a_734_7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5234 a_22196_5331# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5235 gnd d0 a_25191_n4940# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5236 a_26100_n4543# a_26102_n5061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5237 a_15687_3544# a_15944_3354# a_15605_4152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5238 a_26539_n2201# a_26321_n2201# a_25607_n2057# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5239 a_22396_3901# a_22178_3901# a_21907_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5240 gnd d2 a_24312_n5320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5241 a_18885_7170# d2 a_18936_6679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5242 a_235_7254# d0 a_716_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5243 a_11241_4139# a_11498_3949# a_11162_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5244 a_19092_258# d5 a_19191_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5245 a_14238_n9556# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5246 a_5008_2871# d1 a_5805_3099# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5247 a_4790_n2589# a_4572_n2589# a_4309_n2300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5248 a_16468_2577# a_16485_3360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5249 a_30757_n6698# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5250 vdd d2 a_20091_1900# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5251 a_17706_n9714# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5252 a_11340_4549# d0 a_12138_4365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5253 a_6770_n4496# d0 a_7563_n4912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5254 gnd d2 a_11571_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5255 gnd d0 a_20917_n10017# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5256 a_15487_n3691# d0 a_16289_n3319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5257 a_443_n3594# d1 a_1229_n2802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5258 a_13659_n9328# a_13441_n9328# a_13168_n9134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5259 gnd d0 a_29549_n3522# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5260 a_19658_n3067# d1 a_19757_n3477# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5261 a_15461_n7353# a_15718_n7369# a_15415_n8373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5262 a_6440_n10578# d4 a_6498_n6314# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5263 a_4497_1860# a_4499_1959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5264 a_33115_6433# d0 a_33912_6661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5265 a_14546_3124# d2 a_14597_2633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5266 a_6684_n5292# d1 a_6766_n4684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5267 a_16557_7844# a_16561_7667# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5268 a_17125_n10728# a_17382_n10744# a_17212_n839# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5269 a_15342_n4301# a_15599_n4317# a_15239_n6339# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5270 a_27409_n6734# a_27191_n6501# a_26611_n6685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5271 a_10817_n10590# d4 a_10875_n6326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5272 a_8913_4007# d0 a_9402_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5273 a_31012_n8734# a_30794_n8734# a_30537_n8628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5274 a_15609_3975# d1 a_15704_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5275 a_31815_n8960# a_31609_n9568# a_31030_n9340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5276 a_11413_8621# d0 a_12211_8437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5277 a_18693_3508# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5278 a_4585_6432# a_4590_6756# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5279 a_660_4288# d1 a_1446_3615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5280 gnd d0 a_12413_5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5281 a_28616_3974# a_28869_3961# a_28533_2958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5282 a_20006_6572# d0 a_20808_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5283 a_3416_5358# a_3420_5181# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5284 a_27228_n8537# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5285 gnd d0 a_21081_7216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5286 a_4616_8285# d0 a_5097_8373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5287 a_4863_n6661# a_4645_n6661# a_4388_n6555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5288 a_5946_n5865# a_5728_n5865# a_5843_n7903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5289 a_27208_n7519# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5290 vdd d5 a_6697_n10594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5291 a_25136_4188# a_25389_4175# a_24334_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5292 a_27476_n5889# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5293 a_23139_1075# a_22921_1075# a_22341_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5294 a_9384_3295# a_9166_3295# a_8903_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5295 a_28612_4151# d1 a_28694_3543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5296 a_6967_4360# d0 a_7764_4588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5297 a_26175_n9133# a_26177_n9232# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5298 a_13532_n2202# d1 a_14329_n2663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5299 a_33932_7679# a_33946_8462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5300 a_21997_n5655# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5301 a_7744_3335# a_7748_3158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5302 a_6950_3342# d0 a_7747_3570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5303 a_28689_8046# a_28942_8033# a_28606_7030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5304 gnd d1 a_24647_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5305 a_24938_n4736# a_25191_n4940# a_24141_n4508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5306 a_4662_n7679# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5307 a_11055_n8172# d2 a_11138_n9188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5308 vdd d0 a_34166_6236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5309 a_13822_6968# d1 a_14619_7196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5310 a_5097_8373# d1 a_5883_7700# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5311 a_19092_258# d4 a_19689_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5312 a_9458_6955# a_9240_6955# a_8967_6768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5313 a_25209_8260# a_25462_8247# a_24407_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5314 a_23212_5147# a_22994_5147# a_22414_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5315 a_31840_n5902# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5316 a_29365_n7578# a_29369_n7390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5317 a_24141_n4508# a_24394_n4712# a_24055_n5304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5318 a_24152_3123# d2 a_24202_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5319 vdd d0 a_12250_n7994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5320 a_4806_4301# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5321 a_4880_7961# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5322 vdd d1 a_11597_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5323 a_13441_n9328# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5324 vdd d1 a_28751_n3706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5325 a_17397_n7072# a_17399_n7171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5326 a_33693_n5555# a_33697_n5367# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5327 a_2419_n5689# d0 a_3221_n5317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5328 a_15346_n4113# d2 a_15425_n5317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5329 a_15760_7616# d0 a_16558_7432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5330 a_2566_2311# d0 a_3359_2716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5331 a_29508_4789# a_29765_4599# a_28715_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5332 a_21807_n9438# a_21813_n9621# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5333 a_31499_n3460# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5334 a_21753_n6384# d0 a_22234_n6673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5335 a_14165_n5484# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5336 a_246_n4200# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5337 a_33819_1336# a_33823_1159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5338 gnd d0 a_16541_n3935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5339 a_515_8360# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5340 a_22053_n8709# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5341 vdd d1 a_28861_n9814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5342 vdd d2 a_33016_n3309# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5343 a_5604_4117# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5344 a_20772_4175# a_20767_4764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5345 a_29348_n6560# a_29352_n6372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5346 a_28426_5173# d3 a_28533_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5347 a_1492_2595# d3 a_1586_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5348 a_33094_5592# d0 a_33896_5231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5349 a_5660_7171# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5350 a_12014_n8584# a_12271_n8600# a_11216_n8768# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5351 a_17339_n3500# a_17344_n4018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5352 a_26411_n7291# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5353 a_13314_n2202# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5354 a_8945_5426# d0 a_9420_5331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5355 a_4534_3896# d0 a_5025_3889# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5356 a_5625_n4674# a_5407_n4441# a_4828_n4213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5357 a_11340_4549# d0 a_12142_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5358 vdd d2 a_11571_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5359 a_5593_n2815# a_5387_n3423# a_4807_n3607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5360 a_27155_n4465# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5361 a_13043_n2107# d0 a_13532_n2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5362 gnd d2 a_20128_3936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5363 a_11981_n6360# a_11976_n6960# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5364 a_8709_n3513# d0 a_9184_n3619# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5365 gnd d2 a_2540_n3259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5366 a_5846_5664# d2 a_5924_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5367 a_319_n8272# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5368 gnd d2 a_15755_n9405# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5369 a_16309_n4337# a_16562_n4541# a_15507_n4709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5370 a_31099_2302# a_30881_2302# a_30624_2397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5371 a_31173_5962# a_30955_5962# a_30682_5969# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5372 vdd d0 a_33949_n5983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5373 a_4808_n3195# a_4590_n3195# a_4319_n3100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5374 gnd d2 a_15862_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5375 a_11101_n7152# d1 a_11200_n7562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5376 a_24190_n7750# d0 a_24992_n7378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5377 a_48_n8177# d0 a_537_n8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5378 a_8789_n8202# a_8796_n8420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5379 a_26555_n3631# d1 a_27341_n2839# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5380 a_31922_3665# d2 a_31968_2645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5381 a_26_n7060# d0 a_517_n7254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5382 a_15609_3975# d1 a_15708_4385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5383 a_23130_7593# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5384 a_3416_5358# a_3673_5168# a_2618_5542# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5385 a_1441_6548# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5386 a_11286_1495# a_11543_1305# a_11204_2103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5387 vdd d0 a_7800_n3910# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5388 a_5810_3628# a_5604_4117# a_5024_4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5389 a_2659_7401# a_2912_7388# a_2573_8186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5390 a_10982_n4100# d2 a_11065_n5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5391 a_13605_n6274# d1 a_14402_n6735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5392 vdd d0 a_21081_7216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5393 a_14418_8214# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5394 a_25132_4365# a_25389_4175# a_24334_4549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5395 a_29292_n3506# a_29296_n3318# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5396 a_26593_n5255# a_26375_n5255# a_26104_n5160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5397 a_28612_4151# d1 a_28698_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5398 a_13114_n6080# d0 a_13605_n6274# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5399 vdd d3 a_6858_n4292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5400 a_30702_n3232# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5401 a_17502_1341# a_17504_1859# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5402 a_30918_4338# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5403 a_6785_2934# d2 a_6868_3950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5404 a_8776_n7402# d0 a_9257_n7691# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5405 a_10306_6692# d3 a_10400_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5406 a_30758_n6286# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5407 a_29492_3359# a_29496_3182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5408 a_28685_8223# a_28942_8033# a_28606_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5409 a_10145_1075# d2 a_10228_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5410 a_5732_2489# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5411 a_26773_3913# d1 a_27558_3652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5412 a_4337_n4019# a_4339_n4118# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5413 vdd d1 a_24647_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5414 vdd d3 a_11235_n4304# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5415 a_30974_7392# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5416 a_131_1329# d0 a_606_1234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5417 a_31737_n7940# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5418 a_554_n9290# d1 a_1339_n8910# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5419 a_11208_1926# d1 a_11303_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5420 gnd d0 a_34023_n9643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5421 a_20574_n4723# a_20588_n5517# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5422 a_31788_n3868# a_31618_n4888# a_31737_n4711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5423 a_18817_3627# a_18611_4116# a_18032_3888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5424 a_1312_n3818# d3 a_1406_n3818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5425 a_32078_296# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5426 a_27604_2632# a_27434_3533# a_27558_3652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5427 a_31592_n8550# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5428 a_31572_n7532# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5429 a_15498_n9389# d1 a_15580_n8781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5430 a_20538_n2275# a_20533_n2875# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5431 a_24156_2946# d2 a_24235_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5432 a_18885_7170# a_18667_7170# a_18088_6942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5433 a_26846_7985# d1 a_27631_7724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5434 a_13403_n7704# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5435 gnd d0 a_34130_4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5436 a_15760_7616# d0 a_16562_7255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5437 a_14439_n8771# d2 a_14490_n7928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5438 a_2566_2311# d0 a_3363_2539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5439 a_33912_6661# a_34165_6648# a_33115_6433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5440 a_4646_n6249# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5441 a_2549_1293# d0 a_3346_1521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5442 a_20791_5193# a_21044_5180# a_19989_5554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5443 a_9944_2093# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5444 a_14624_7725# a_14418_8214# a_13838_8398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5445 a_5843_n7903# a_5625_n7903# a_5749_n7903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5446 a_4512_2360# d0 a_4987_2265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5447 a_13296_5038# d0 a_13785_4932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5448 a_15740_6598# a_15997_6408# a_15645_6011# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5449 a_27373_n7927# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5450 a_24301_2336# a_24554_2323# a_24202_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5451 gnd d0 a_34203_8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5452 a_11200_n7562# d0 a_11993_n7978# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5453 a_10126_n7915# a_9956_n8935# a_10075_n8758# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5454 a_32786_n8385# a_33043_n8401# a_32614_n6163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5455 a_22288_n9727# d1 a_23074_n8935# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5456 a_17833_4906# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5457 a_26431_n8309# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5458 a_17380_n6054# d0 a_17871_n6248# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5459 a_n47_n2988# d0 a_444_n3182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5460 a_27626_7195# a_27408_7195# a_26828_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5461 a_14546_6586# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5462 a_18683_n3830# d3 a_18777_n3830# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5463 a_28477_n2672# a_28734_n2688# a_28395_n3280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5464 a_24321_3354# d0 a_25118_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5465 a_28730_5579# a_28987_5389# a_28648_6187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5466 a_14390_1498# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5467 a_13253_2385# a_13258_2709# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5468 a_4572_6031# d0 a_5061_5925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5469 a_17617_n4212# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5470 a_1186_1050# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5471 a_32935_n7587# d0 a_33728_n8003# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5472 a_19790_n5701# d0 a_20588_n5517# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5473 a_13585_n5668# a_13367_n5668# a_13110_n5562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5474 vdd d0 a_8036_5593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5475 a_8723_n4348# d0 a_9204_n4637# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5476 a_3256_n7765# a_3509_n7969# a_2459_n7537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5477 a_6724_n7140# d1 a_6819_n7738# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5478 a_28287_n10602# a_30320_n10705# a_25615_n10665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5479 a_225_n3594# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5480 vdd d1 a_33225_n9827# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5481 a_17346_n4117# d0 a_17835_n4212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5482 a_22251_7973# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5483 a_22177_4313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5484 vdd d0 a_34112_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5485 a_33752_n8833# a_33766_n9627# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5486 a_17978_834# d1 a_18775_1062# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5487 a_2314_n8147# a_2567_n8351# a_2138_n6113# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5488 a_16520_5808# a_16524_5631# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5489 vdd d1 a_11473_n8784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5490 a_31664_n3868# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5491 a_13309_5439# a_13311_5957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5492 a_33716_n6385# a_33711_n6985# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5493 a_19788_3110# d2 a_19834_2090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5494 a_27672_6585# a_27470_5569# a_27589_5159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5495 a_5946_n5865# a_6697_n10594# a_3951_n10652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5496 a_22162_n2189# d1 a_22959_n2650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5497 a_33823_1159# a_34076_1146# a_33021_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5498 a_26_n7060# a_28_n7159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5499 a_4091_172# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5500 a_7636_n8984# a_7893_n9000# a_6843_n8568# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5501 a_13549_n3220# a_13331_n3220# a_13058_n3026# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5502 a_3360_2304# a_3364_2127# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5503 a_17908_n8284# d1 a_18705_n8745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5504 a_22250_8385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5505 gnd d1 a_2749_n9777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5506 a_9365_1865# a_9147_1865# a_8876_1971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5507 gnd d0 a_20864_n6551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5508 a_30722_n4250# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5509 a_19695_n5103# d1 a_19790_n5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5510 gnd d1 a_15764_n4725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5511 a_5370_n2405# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5512 vdd d2 a_2793_5960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5513 a_29496_3182# a_29491_3771# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5514 a_14366_n4699# d2 a_14417_n3856# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5515 a_17533_3194# a_17539_3377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5516 a_3401_4163# a_3654_4150# a_2599_4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5517 a_4573_n2177# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5518 a_13151_n8116# d0 a_13642_n8310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5519 a_14439_n8771# a_14221_n8538# a_13642_n8310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5520 a_11208_1926# d1 a_11307_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5521 gnd d0 a_12394_4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5522 gnd d0 a_25352_2139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5523 a_3951_n10652# a_4208_n10668# a_4050_n10652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5524 a_15601_n9611# d0 a_16394_n10027# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5525 a_5044_4907# a_4826_4907# a_4555_5013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5526 a_2577_8009# d1 a_2672_8596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5527 a_16377_n9009# a_16381_n8821# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5528 a_17443_n9425# a_17449_n9608# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5529 a_30682_5969# a_30684_6068# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5530 a_23976_n4100# d2 a_24055_n5304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5531 a_5770_n3831# a_5552_n3831# a_5676_n3831# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5532 a_2459_n7537# d0 a_3256_n7765# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5533 vdd d3 a_19938_n8363# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5534 a_30468_n5173# a_30475_n5391# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5535 a_21924_4926# a_21926_5025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5536 vdd d0 a_12161_n2492# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5537 a_3239_n6747# a_3253_n7541# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5538 a_7568_n4312# a_7821_n4516# a_6766_n4684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5539 a_19685_n8159# a_19938_n8363# a_19509_n6125# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5540 a_8750_n6067# d0 a_9241_n6261# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5541 a_14238_n9556# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5542 gnd d1 a_7276_7401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5543 a_2417_3098# d2 a_2467_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5544 a_17706_n9714# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5545 a_29278_n2712# a_29531_n2916# a_28481_n2484# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5546 a_32800_n5141# d1 a_32895_n5739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5547 a_30594_978# d0 a_31083_872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5548 a_623_2252# a_405_2252# a_142_2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5549 a_20787_5370# a_21044_5180# a_19989_5554# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5550 gnd d4 a_11312_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5551 a_8769_n7184# d0 a_9258_n7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5552 a_23181_3640# a_22975_4129# a_22395_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5553 a_24297_2513# a_24554_2323# a_24202_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5554 a_27409_n6734# a_27191_n6501# a_26612_n6273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5555 a_14764_6586# d4 a_14831_403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5556 vdd d0 a_34203_8272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5557 a_3236_n6523# a_3240_n6335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5558 a_31012_n8734# a_30794_n8734# a_30531_n8445# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5559 vdd d1 a_7023_n4700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5560 a_30992_n7716# a_30774_n7716# a_30517_n7610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5561 a_22161_2883# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5562 a_21673_n2094# d0 a_22162_n2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5563 a_24353_5567# a_24610_5377# a_24271_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5564 vdd d4 a_11132_n6342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5565 a_697_5912# a_479_5912# a_206_5919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5566 gnd d2 a_24385_n9392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5567 a_7564_n4500# a_7568_n4312# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5568 a_13058_n3026# a_13060_n3125# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5569 a_18574_2080# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5570 a_4863_n6661# a_4645_n6661# a_4382_n6372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5571 a_5946_n5865# a_5728_n5865# a_5770_n3831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5572 a_11359_5567# d0 a_12161_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5573 a_463_n4612# a_245_n4612# a_n12_n4506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5574 a_6999_6573# d0 a_7801_6212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5575 a_116_829# d0 a_607_822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5576 a_17361_n5036# d0 a_17852_n5230# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5577 a_7563_n4912# a_7820_n4928# a_6770_n4496# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5578 a_11158_3123# a_11415_2933# a_11055_5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5579 a_15547_n6557# a_15800_n6761# a_15461_n7353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5580 a_13363_8493# d0 a_13838_8398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5581 a_13802_5950# a_13584_5950# a_13311_5957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5582 a_19509_n6125# d3 a_19685_n8159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5583 a_21997_n5655# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5584 a_11059_4984# d3 a_11231_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5585 a_6498_n6314# a_6755_n6330# a_6440_n10578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5586 a_33075_4574# d0 a_33877_4213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5587 gnd d0 a_25371_3569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5588 a_22288_n9727# a_22070_n9727# a_21813_n9621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5589 a_7727_2552# a_7980_2539# a_6930_2324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5590 a_24918_n3718# a_25171_n3922# a_24121_n3490# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5591 gnd d0 a_29802_6223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5592 a_262_n5630# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5593 a_8926_4408# d0 a_9401_4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5594 a_26067_n3124# a_26074_n3342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5595 a_26353_7474# d0 a_26828_7379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5596 a_28652_6010# d1 a_28751_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5597 a_17519_2359# a_17524_2683# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5598 a_26792_4931# a_26574_4931# a_26301_4938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5599 a_25209_8260# a_25204_8849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5600 a_24121_n3490# a_24374_n3694# a_24022_n3080# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5601 a_33819_1336# a_34076_1146# a_33021_1520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5602 a_21920_4408# a_21924_4926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5603 a_n8_n5123# a_n1_n5341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5604 a_29509_4377# a_29513_4200# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5605 a_14514_1617# a_14308_2106# a_13729_1878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5606 vdd d5 a_28445_n10618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5607 a_4399_n7390# a_4405_n7573# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5608 a_27315_2105# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5609 a_25151_5383# a_25408_5193# a_24353_5567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5610 a_23222_2501# a_23020_1485# a_23144_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5611 a_13350_n4650# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5612 gnd a_n62_n2069# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5613 a_14582_5160# a_14364_5160# a_13785_4932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5614 a_5883_7700# d2 a_5929_6680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5615 a_21759_n6567# d0 a_22234_n6673# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5616 a_24229_7018# a_24482_7005# a_24053_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5617 a_3397_4340# a_3654_4150# a_2599_4524# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5618 a_25011_n8808# a_25264_n9012# a_24214_n8580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5619 a_226_n3182# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5620 a_19191_258# d6 a_21680_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5621 a_32939_2128# a_33196_1938# a_32893_3148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5622 a_191_5000# a_198_5218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5623 a_26357_8091# a_26364_8309# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5624 a_29565_7431# a_29569_7254# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5625 vdd d0 a_29621_n8006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5626 a_23069_n8758# d2 a_23120_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5627 gnd d2 a_33269_6010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5628 a_24370_6585# d0 a_25168_6401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5629 a_11994_n7566# a_12251_n7582# a_11196_n7750# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5630 a_4879_8373# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5631 vdd d3 a_28679_n8388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5632 a_13314_n2202# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5633 a_15419_n8185# d2 a_15498_n9389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5634 a_16541_6649# a_16794_6636# a_15744_6421# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5635 a_2479_n8555# a_2732_n8759# a_2393_n9351# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5636 a_31679_2118# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5637 a_15423_4997# d3 a_15595_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5638 a_29402_n9614# a_29406_n9426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5639 a_15425_n5317# a_15682_n5333# a_15346_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5640 a_5593_n2815# a_5387_n3423# a_4808_n3195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5641 a_8949_n2601# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5642 a_12121_3347# a_12125_3170# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5643 a_18936_6679# a_18766_7580# a_18890_7699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5644 a_8731_n5049# d0 a_9222_n5243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5645 a_26085_n4043# a_26087_n4142# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5646 a_444_n3182# d1 a_1229_n2802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5647 a_319_n8272# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5648 a_13659_n9328# a_13441_n9328# a_13170_n9233# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5649 gnd d1 a_11616_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5650 a_299_n7254# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5651 a_16289_n3319# a_16542_n3523# a_15487_n3691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5652 a_2438_n6707# d0 a_3240_n6335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5653 a_12951_197# a_14707_284# a_14831_403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5654 gnd d0 a_29821_7653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5655 a_4790_2871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5656 a_168_3365# d0 a_643_3270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5657 gnd d2 a_7121_3937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5658 a_29531_5630# a_29784_5617# a_28734_5402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5659 a_28_n7159# d0 a_517_n7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5660 vdd d5 a_24068_n10606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5661 a_14184_n6502# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5662 a_31752_6190# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5663 a_21870_1971# a_21877_2189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5664 a_17550_4212# d0 a_18031_4300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5665 a_443_3876# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5666 a_31815_n8960# a_31609_n9568# a_31029_n9752# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5667 a_27378_n4875# a_27172_n5483# a_26593_n5255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5668 a_6864_4127# d1 a_6950_3342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5669 a_13604_n6686# d1 a_14402_n6735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5670 a_13387_n6274# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5671 a_29328_n5954# a_29332_n5766# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5672 a_12211_8437# a_12468_8247# a_11413_8621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5673 a_13238_1885# a_13240_1984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5674 a_17606_7266# d0 a_18087_7354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5675 a_20772_4175# a_21025_4162# a_19970_4536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5676 gnd d1 a_2875_5352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5677 a_26593_n5255# a_26375_n5255# a_26102_n5061# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5678 a_5666_n6887# a_5460_n7495# a_4880_n7679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5679 a_13116_n6179# d0 a_13605_n6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5680 a_33949_8697# a_34202_8684# a_33152_8469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5681 vdd d1 a_20103_n8771# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5682 a_10875_n6326# d3 a_10982_n4100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5683 a_22415_4919# a_22197_4919# a_21926_5025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5684 a_13277_4020# d0 a_13766_3914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5685 a_16382_n8409# a_16635_n8613# a_15580_n8781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5686 a_28246_n6338# d3 a_28349_n4300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5687 a_17797_2870# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5688 a_25025_n9602# a_25029_n9414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5689 a_8802_n8603# a_8804_n9121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5690 a_442_4288# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5691 vdd d3 a_11488_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5692 a_1285_1460# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5693 vdd d1 a_33295_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5694 a_1188_n3818# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5695 vdd d0 a_29802_6223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5696 a_9458_6955# d1 a_10255_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5697 vdd d0 a_29568_n4952# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5698 vdd d0 a_8000_3557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5699 a_15645_6011# a_15898_5998# a_15595_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5700 a_20643_n8983# a_20900_n8999# a_19850_n8567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5701 vdd d4 a_19942_4958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5702 a_27451_n8947# a_27245_n9555# a_26665_n9739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5703 a_11235_7018# d2 a_11314_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5704 a_17796_3282# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5705 a_17870_6942# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5706 a_31572_n7532# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5707 vdd d1 a_28771_n4724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5708 a_25151_5383# a_25155_5206# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5709 a_5883_7700# a_5677_8189# a_5098_7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5710 a_23321_2501# a_23103_2501# a_23222_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5711 a_15465_n7165# d1 a_15560_n7763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5712 a_13441_n9328# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5713 a_13277_4020# a_13284_4238# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5714 vdd d1 a_33171_n6773# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5715 a_15487_n3691# a_15744_n3707# a_15392_n3093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5716 vdd d1 a_15837_n8797# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5717 a_21970_7279# d0 a_22451_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5718 a_6678_n8160# d2 a_6761_n9176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5719 a_13748_3308# d1 a_14546_3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5720 vdd d3 a_28606_n4316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5721 a_29352_n6372# a_29605_n6576# a_28550_n6744# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5722 a_3221_n5317# a_3474_n5521# a_2419_n5689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5723 vdd d0 a_20791_n2479# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5724 a_5843_n7903# a_5625_n7903# a_5744_n7726# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5725 a_10121_n7738# a_9919_n6899# a_10043_n6899# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5726 a_29459_1146# a_29454_1735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5727 a_20592_n5329# a_20587_n5929# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5728 a_22053_n8709# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5729 a_27373_n7927# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5730 a_26845_8397# a_26627_8397# a_26364_8309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5731 a_24235_4139# d1 a_24317_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5732 a_31861_n7940# a_31691_n8960# a_31810_n8783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5733 a_26364_8309# a_26370_8492# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5734 a_33711_n6985# a_33968_n7001# a_32918_n6569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5735 a_11344_4372# d0 a_12141_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5736 a_7784_5194# a_8037_5181# a_6982_5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5737 vdd d2 a_33269_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5738 a_31030_n9340# a_30812_n9340# a_30539_n9146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5739 a_2365_n2635# d0 a_3167_n2263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5740 a_14328_3124# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5741 a_18559_n3830# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5742 a_536_n8684# d1 a_1334_n8733# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5743 a_24370_6585# d0 a_25172_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5744 a_24312_8034# a_24565_8021# a_24229_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5745 a_n47_n2988# a_n45_n3087# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5746 a_24100_n2660# d0 a_24902_n2288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5747 a_33860_3195# a_34113_3182# a_33058_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5748 a_1406_n3818# d4 a_1582_n5852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5749 a_10099_5557# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5750 a_16537_6826# a_16794_6636# a_15744_6421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5751 a_31742_n4888# a_31536_n5496# a_30956_n5680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5752 a_5080_7355# a_4862_7355# a_4599_7267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5753 a_32873_n9213# d1 a_32972_n9623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5754 vdd d1 a_28807_n6760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5755 a_17617_n4212# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5756 a_26310_5255# a_26316_5438# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5757 a_4825_5319# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5758 a_16558_7432# a_16562_7255# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5759 a_8729_n4531# d0 a_9204_n4637# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5760 a_14401_7196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5761 a_11977_n6548# a_11981_n6360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5762 a_8703_n3330# d0 a_9184_n3619# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5763 a_5025_3889# a_4807_3889# a_4536_3995# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5764 a_11920_n3906# a_11924_n3718# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5765 vdd d0 a_29749_3169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5766 a_30901_3320# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5767 vdd d0 a_29821_7653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5768 a_11134_n9376# d1 a_11220_n8580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5769 a_17326_n3099# d0 a_17815_n3194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5770 a_24128_n9376# a_24385_n9392# a_24049_n8172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5771 vdd d1 a_7076_n7754# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5772 a_10017_6165# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5773 a_25131_4777# a_25388_4587# a_24338_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5774 a_8819_n9621# a_8824_n9945# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5775 a_4339_n4118# a_4346_n4336# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5776 a_29347_n6972# a_29604_n6988# a_28554_n6556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5777 a_30903_n2214# a_30685_n2214# a_30414_n2119# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5778 a_10879_n6138# d3 a_11055_n8172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5779 a_18487_n8512# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5780 a_21877_2189# a_21883_2372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5781 vdd d1 a_20210_3328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5782 a_28250_n6150# d3 a_28422_n8372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5783 a_31968_2645# a_31798_3546# a_31917_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5784 a_18812_3098# a_18594_3098# a_18014_3282# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5785 a_22161_n2601# d1 a_22959_n2650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5786 a_536_n8684# a_318_n8684# a_55_n8395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5787 a_15425_n5317# d1 a_15507_n4709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5788 vdd d1 a_2875_5352# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5789 a_10054_8201# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5790 a_17907_n8696# d1 a_18705_n8745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5791 a_17029_133# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5792 a_20768_4352# a_21025_4162# a_19970_4536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5793 a_8947_5944# d0 a_9438_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5794 a_7616_n7966# a_7873_n7982# a_6823_n7550# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5795 a_33945_8874# a_34202_8684# a_33152_8469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5796 a_20588_n5517# a_20845_n5533# a_19790_n5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5797 a_5370_n2405# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5798 a_8824_n9945# a_12287_n10030# a_11237_n9598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5799 vdd d1 a_33098_n2701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5800 vdd d1 a_20283_7400# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5801 a_28751_6420# d0 a_29544_6825# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5802 a_33770_n9439# a_33765_n10039# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5803 a_14371_n4876# d2 a_14417_n3856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5804 a_22199_n4225# a_21981_n4225# a_21710_n4130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5805 gnd d0 a_21061_6198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5806 gnd d2 a_24275_n3284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5807 a_5856_2608# d3 a_5950_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5808 a_30644_3415# d0 a_31119_3320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5809 a_9202_5331# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5810 a_14407_n6912# a_14201_n7520# a_13622_n7292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5811 a_5770_n3831# a_5552_n3831# a_5671_n3654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5812 a_17887_n7678# a_17669_n7678# a_17406_n7389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5813 a_23057_3521# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5814 a_19838_1913# d1 a_19933_2500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5815 a_11235_7018# d2 a_11318_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5816 a_1307_n3641# d3 a_1406_n3818# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5817 a_18104_8372# a_17886_8372# a_17629_8467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5818 a_31592_n8550# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5819 a_6733_n2460# d0 a_7526_n2876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5820 a_1446_3615# d2 a_1492_2595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5821 gnd d0 a_3636_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5822 a_13839_7986# a_13621_7986# a_13350_8092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5823 a_8752_n6166# d0 a_9241_n6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5824 a_28604_n9798# a_28861_n9814# a_28509_n9200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5825 a_22778_n4453# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5826 a_5671_n3654# a_5469_n2815# a_5593_n2815# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5827 gnd d1 a_24627_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5828 a_11110_n2472# d0 a_11903_n2888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5829 a_13802_5950# d1 a_14587_5689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5830 a_19846_n8755# d0 a_20644_n8571# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5831 a_10260_7712# a_10054_8201# a_9474_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5832 a_24190_n7750# a_24447_n7766# a_24095_n7152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5833 a_1519_7687# d2 a_1565_6667# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5834 vdd d1 a_33152_n5755# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5835 a_28518_n4520# d0 a_29311_n4936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5836 a_33115_6433# d0 a_33908_6838# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5837 a_24235_4139# d1 a_24321_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5838 a_19867_n9585# d0 a_17454_n9932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5839 a_17502_1341# d0 a_17977_1246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5840 a_26773_3913# a_26555_3913# a_26282_3920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5841 a_14665_6586# a_14463_5570# a_14587_5689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5842 a_30594_978# a_30601_1196# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5843 a_7780_5371# a_8037_5181# a_6982_5555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5844 a_4436_n9426# d0 a_4917_n9715# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5845 a_19989_5554# d0 a_20787_5370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5846 a_28188_n10602# d4 a_28246_n6338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5847 a_26792_4931# d1 a_27589_5159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5848 a_n45_n3087# a_n38_n3305# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5849 a_24308_8211# a_24565_8021# a_24229_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5850 a_24055_n5304# a_24312_n5320# a_23976_n4100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5851 a_30992_n7716# a_30774_n7716# a_30511_n7427# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5852 vdd d1 a_7003_n3682# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5853 a_4987_2265# a_4769_2265# a_4506_2177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5854 a_n27_n4006# d0 a_464_n4200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5855 a_17614_7967# a_17616_8066# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5856 a_33856_3372# a_34113_3182# a_33058_3556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5857 a_10182_6573# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5858 a_16322_n5543# a_16326_n5355# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5859 a_32972_n9623# d0 a_33765_n10039# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5860 a_14551_3653# a_14345_4142# a_13766_3914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5861 a_28602_7207# d2 a_28648_6187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5862 a_9420_5331# a_9202_5331# a_8945_5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5863 a_33711_n6985# a_33715_n6797# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5864 a_4901_n8285# a_4683_n8285# a_4412_n8190# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5865 a_27352_4141# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5866 a_18678_n3653# d3 a_18777_n3830# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5867 a_23227_2620# a_23057_3521# a_23181_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5868 a_17562_5012# d0 a_18051_4906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5869 a_29292_n3506# a_29549_n3522# a_28494_n3690# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5870 a_463_n4612# a_245_n4612# a_n18_n4323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5871 a_31137_3926# d1 a_31922_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5872 a_22469_7973# d1 a_23254_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5873 a_26611_n6685# a_26393_n6685# a_26136_n6579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5874 a_7543_n3894# a_7800_n3910# a_6750_n3478# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5875 vdd d0 a_7893_n9000# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5876 gnd d0 a_12450_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5877 a_3436_6611# a_3689_6598# a_2639_6383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5878 a_27553_3123# a_27335_3123# a_26756_2895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5879 a_22288_n9727# a_22070_n9727# a_21807_n9438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5880 a_6950_3342# d0 a_7743_3747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5881 a_16505_4613# a_16758_4600# a_15708_4385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5882 a_6502_n6126# d3 a_6674_n8348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5883 a_31654_n6924# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5884 a_1726_365# a_1544_4510# a_1659_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5885 a_12035_n9414# a_12288_n9618# a_11233_n9786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5886 vdd d0 a_12358_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5887 a_13549_n3220# a_13331_n3220# a_13060_n3125# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5888 a_29495_3594# a_29748_3581# a_28698_3366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5889 gnd d1 a_11597_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5890 gnd d0 a_34092_2576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5891 a_16578_8685# a_16831_8672# a_15781_8457# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5892 a_28591_n8592# d0 a_29384_n9008# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5893 a_19191_258# a_18973_258# a_19097_377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5894 a_6085_259# d4 a_6678_5149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5895 a_33021_1520# d0 a_33819_1336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5896 a_10400_6573# a_10182_6573# a_10306_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5897 a_8894_2696# a_8896_2989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5898 a_23249_7183# a_23031_7183# a_22451_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5899 a_28751_6420# d0 a_29548_6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5900 gnd d4 a_15496_n6355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5901 a_5950_2489# a_5732_2489# a_5856_2608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5902 a_24991_n7790# a_25244_n7994# a_24194_n7562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5903 a_22071_n9315# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5904 a_26080_n3525# a_26085_n4043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5905 a_14439_n8771# a_14221_n8538# a_13641_n8722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5906 a_22124_847# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5907 a_8982_7462# a_8984_7980# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5908 a_29568_7666# a_29821_7653# a_28771_7438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5909 a_33729_n7591# a_33986_n7607# a_32931_n7775# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5910 a_23074_n8935# d2 a_23120_n7915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5911 a_19838_1913# d1 a_19937_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5912 vdd d0 a_3636_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5913 vdd d2 a_15645_n3297# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5914 a_25114_3759# a_25118_3582# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5915 gnd d1 a_2856_4334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5916 a_33094_5592# d0 a_33892_5408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5917 a_4363_n5354# d0 a_4844_n5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5918 a_21903_3390# a_21905_3908# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5919 a_28436_n5128# a_28689_n5332# a_28353_n4112# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5920 a_19740_n2459# a_19993_n2663# a_19654_n3255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5921 a_17629_8467# a_16578_8685# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5922 a_27388_6177# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5923 a_10462_271# d5 a_10561_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5924 a_23295_6573# d3 a_23394_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5925 a_22452_6955# a_22234_6955# a_21963_7061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5926 a_2459_n7537# a_2712_n7741# a_2360_n7127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5927 a_8949_n2601# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5928 a_8733_n5148# d0 a_9222_n5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5929 a_3474_8235# a_3469_8824# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5930 a_19813_n6531# d0 a_20606_n6947# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5931 a_8789_n8202# d0 a_9278_n8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5932 a_8896_2989# d0 a_9385_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5933 vdd d2 a_15825_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5934 a_299_n7254# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5935 a_20533_n2875# a_20790_n2891# a_19740_n2459# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5936 a_13097_n5161# a_13104_n5379# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5937 a_22033_n7691# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5938 a_19989_5554# d0 a_20791_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5939 a_14184_n6502# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5940 gnd d2 a_24455_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5941 a_4210_172# d6 a_4309_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5942 vdd d0 a_16578_n5971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5943 a_26327_6273# a_26333_6456# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5944 a_3420_5181# a_3673_5168# a_2618_5542# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5945 vdd d0 a_7838_n5534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5946 a_479_5912# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5947 a_16489_3183# a_16742_3170# a_15687_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5948 gnd d0 a_16598_n6577# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5949 a_6601_n4276# d2 a_6651_n3068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5950 a_14831_403# a_14649_4548# a_14691_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5951 a_12013_n8996# a_12017_n8808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5952 a_13387_n6274# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5953 a_24938_n4736# a_24952_n5530# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5954 a_8903_3207# d0 a_9384_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5955 a_27656_4547# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5956 a_14764_6586# a_14546_6586# a_14670_6705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5957 a_5_n5524# a_9_n6042# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5958 a_32062_2526# d4 a_32202_415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5959 a_14584_n7928# a_14366_n7928# a_14485_n7751# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5960 a_10121_n7738# d3 a_10220_n7915# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5961 a_5805_3099# d2 a_5856_2608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5962 a_15547_n6557# d0 a_16340_n6973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5963 vdd d1 a_20083_n7753# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5964 a_4807_3889# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5965 a_16521_5396# a_16525_5219# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5966 vdd d0 a_12450_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5967 a_16362_n7391# a_16615_n7595# a_15560_n7763# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5968 a_7765_4176# a_8018_4163# a_6963_4537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5969 a_31735_5172# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5970 gnd d0 a_21007_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5971 a_27594_5688# a_27388_6177# a_26808_6361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5972 a_13642_n8310# a_13424_n8310# a_13151_n8116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5973 a_32951_n8793# d0 a_33749_n8609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5974 a_6090_378# a_5908_4523# a_5950_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5975 a_1296_7158# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5976 a_26138_n7097# a_26140_n7196# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5977 a_26574_4931# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5978 a_27451_n8947# a_27245_n9555# a_26666_n9327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5979 a_14366_n4699# a_14148_n4466# a_13568_n4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5980 a_6746_n3666# d0 a_7544_n3482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5981 a_18068_5924# a_17850_5924# a_17577_5931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5982 gnd d0 a_16652_n9631# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5983 a_6802_n6720# d0 a_7600_n6536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5984 a_29491_3771# a_29748_3581# a_28698_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5985 a_7801_6212# a_7796_6801# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5986 a_4392_n7172# a_4399_n7390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5987 a_17412_n7572# a_17417_n8090# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5988 a_30548_n9463# a_30554_n9646# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5989 vdd d0 a_34092_2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5990 a_18817_3627# d2 a_18863_2607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5991 a_16574_8862# a_16831_8672# a_15781_8457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5992 a_17419_n8189# a_17426_n8407# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5993 a_7527_n2464# a_7784_n2480# a_6729_n2648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5994 a_11123_n3678# d0 a_11921_n3494# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5995 vdd d4 a_6935_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5996 a_33021_1520# d0 a_33823_1159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5997 a_4862_7355# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X5998 a_4536_3995# a_4543_4213# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X5999 vdd d1 a_15817_n7779# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6000 a_5587_3099# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6001 a_2314_5136# d3 a_2421_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6002 a_27419_n3678# a_27217_n2839# a_27336_n2662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6003 a_17524_2683# d0 a_18015_2870# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6004 a_22358_2277# a_22140_2277# a_21877_2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6005 a_12104_2564# a_12357_2551# a_11307_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6006 a_11055_5161# d3 a_11158_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6007 a_29564_7843# a_29821_7653# a_28771_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6008 a_1116_n8500# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6009 vdd d0 a_29641_n9024# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6010 a_28788_8456# a_29041_8443# a_28689_8046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6011 a_5929_6680# a_5759_7581# a_5878_7171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6012 a_9167_n2601# a_8949_n2601# a_8692_n2495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6013 vdd d2 a_28762_n9404# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6014 vdd d1 a_2856_4334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6015 a_1364_n5852# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6016 a_16357_n7991# a_16614_n8007# a_15564_n7575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6017 a_7833_8837# a_8090_8647# a_7040_8432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6018 a_32893_3148# d2 a_32943_1951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6019 a_516_n7666# d1 a_1302_n6874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6020 a_13620_8398# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6021 a_1479_n7890# d4 a_1582_n5852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6022 a_17869_7354# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6023 a_32955_n8605# d0 a_33752_n8833# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6024 a_2467_1901# a_2720_1888# a_2417_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6025 a_8984_7980# d0 a_9475_7973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6026 a_12177_6636# a_12430_6623# a_11380_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6027 vdd d2 a_24348_n7356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6028 a_24321_3354# d0 a_25114_3759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6029 a_15415_n8373# a_15672_n8389# a_15243_n6151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6030 a_30611_1996# a_30618_2214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6031 a_481_n5218# a_263_n5218# a_n10_n5024# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6032 a_17597_n3194# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6033 a_3294_n9389# a_3547_n9593# a_2492_n9761# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6034 a_8769_n7184# a_8776_n7402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6035 a_9183_4313# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6036 a_28788_8456# d0 a_29581_8861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6037 a_26610_7379# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6038 a_24156_2946# a_24409_2933# a_24049_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6039 a_10048_n3666# d3 a_10147_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6040 a_4410_n8091# a_4412_n8190# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6041 a_18431_n5458# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6042 a_33152_8469# a_33405_8456# a_33053_8059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6043 a_31155_5356# a_30937_5356# a_30680_5451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6044 a_30903_n2214# a_30685_n2214# a_29984_n2069# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6045 a_16485_3360# a_16742_3170# a_15687_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6046 a_18487_n8512# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6047 a_733_8360# a_515_8360# a_258_8455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6048 a_32878_n4721# d0 a_33676_n4537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6049 a_32897_2971# a_33150_2958# a_32790_5186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6050 a_8752_n6166# a_8759_n6384# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6051 a_17887_n7678# d1 a_18673_n6886# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6052 a_4317_n3001# a_4319_n3100# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6053 a_19757_n3477# d0 a_20554_n3705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6054 a_28505_n9388# d1 a_28591_n8592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6055 gnd d0 a_16778_5206# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6056 a_23972_n4288# d2 a_24018_n3268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6057 vdd d0 a_20918_n9605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6058 a_11204_2103# d1 a_11286_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6059 vdd d0 a_21007_3556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6060 a_7761_4353# a_8018_4163# a_6963_4537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6061 a_19970_4536# d0 a_20768_4352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6062 a_32966_7220# d2 a_33012_6200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6063 a_2536_6150# a_2793_5960# a_2490_7170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6064 a_31773_n6747# a_31555_n6514# a_30975_n6698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6065 a_4352_n4519# a_4354_n5037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6066 a_9003_n5655# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6067 a_22199_n4225# a_21981_n4225# a_21708_n4031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6068 a_2635_6560# d0 a_3433_6376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6069 a_13604_n6686# a_13386_n6686# a_13123_n6397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6070 a_1188_n3818# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6071 a_22179_n3207# a_21961_n3207# a_21690_n3112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6072 a_15528_n5539# d0 a_16321_n5955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6073 a_11281_5998# a_11534_5985# a_11231_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6074 a_29512_4612# a_29528_5395# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6075 gnd d1 a_7040_n5718# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6076 a_30976_n6286# a_30758_n6286# a_30487_n6191# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6077 a_427_n2164# d1 a_1224_n2625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6078 a_17925_n9302# a_17707_n9302# a_17436_n9207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6079 a_11957_n5942# a_11961_n5754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6080 a_9401_4313# a_9183_4313# a_8926_4408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6081 a_22034_n7279# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6082 a_6761_n9176# a_7014_n9380# a_6678_n8160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6083 a_16304_n4937# a_16561_n4953# a_15511_n4521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6084 a_12088_1134# a_12341_1121# a_11286_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6085 a_29471_2753# a_29475_2576# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6086 a_26353_7474# a_26355_7992# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6087 gnd d0 a_25209_n5546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6088 gnd d1 a_11417_n5730# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6089 a_15239_n6339# a_15496_n6355# a_15181_n10603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6090 a_13494_860# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6091 a_20791_5193# a_20786_5782# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6092 a_22778_n4453# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6093 a_15507_n4709# a_15764_n4725# a_15425_n5317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6094 a_21987_8297# a_21993_8480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6095 a_5671_n3654# a_5469_n2815# a_5588_n2638# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6096 gnd d2 a_19948_n5307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6097 a_22758_n3435# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6098 a_9927_1075# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6099 a_23069_n8758# a_22851_n8525# a_22271_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6100 a_30522_n8128# a_30524_n8227# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6101 a_6783_n5702# d0 a_7581_n5518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6102 a_24284_1318# a_24537_1305# a_24198_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6103 a_19826_n7737# d0 a_20624_n7553# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6104 a_32552_n10615# d4 a_32614_n6163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6105 a_12100_2741# a_12357_2551# a_11307_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6106 a_5044_4907# d1 a_5841_5135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6107 a_20588_n5517# a_20592_n5329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6108 a_27521_1616# d2 a_27599_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6109 a_24902_n2288# a_25155_n2492# a_24100_n2660# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6110 a_28784_8633# a_29041_8443# a_28689_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6111 a_20607_n6535# a_20864_n6551# a_19809_n6719# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6112 a_28498_n3502# d0 a_29291_n3918# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6113 a_4442_n9609# d0 a_4917_n9715# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6114 a_33859_3607# a_33873_4390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6115 a_31861_n7940# a_31691_n8960# a_31815_n8960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6116 a_33638_n2913# a_33642_n2725# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6117 a_25098_2564# a_25115_3347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6118 a_1380_n7713# d3 a_1479_n7890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6119 a_31030_n9340# a_30812_n9340# a_30541_n9245# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6120 gnd d0 a_3436_n3897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6121 a_10000_5147# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6122 a_26719_859# a_26501_859# a_26230_965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6123 a_4489_1159# a_4495_1342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6124 a_18559_n3830# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6125 a_426_n2576# a_208_n2576# a_n49_n2470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6126 a_28399_n3092# d1 a_28494_n3690# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6127 a_206_5919# a_208_6018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6128 gnd d2 a_2613_n7331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6129 a_24357_5390# a_24610_5377# a_24271_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6130 a_6982_5555# d0 a_7780_5371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6131 a_12173_6813# a_12430_6623# a_11380_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6132 a_33945_8874# a_33949_8697# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6133 vdd d0 a_25461_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6134 a_21866_1354# a_21868_1872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6135 a_4881_n7267# a_4663_n7267# a_4392_n7172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6136 vdd d0 a_34022_n10055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6137 a_23972_n4288# a_24229_n4304# a_23869_n6326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6138 a_18729_5544# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6139 a_32197_296# d5 a_30322_209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6140 a_17148_133# a_25910_208# a_26029_208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6141 a_33058_3556# d0 a_33856_3372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6142 a_32972_n9623# a_33225_n9827# a_32873_n9213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6143 vdd d0 a_25208_n5958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6144 a_28788_8456# d0 a_29585_8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6145 a_28531_n5726# d0 a_29333_n5354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6146 a_16341_n6561# a_16598_n6577# a_15543_n6745# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6147 a_33891_5820# a_33895_5643# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6148 a_1560_6548# a_1358_5532# a_1477_5122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6149 vdd d1 a_24411_n5730# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6150 a_33148_8646# a_33405_8456# a_33053_8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6151 a_4752_1247# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6152 a_31654_n6924# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6153 a_19612_n4087# d2 a_19691_n5291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6154 a_9437_6349# a_9219_6349# a_8956_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6155 a_6688_n5104# d1 a_6787_n5514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6156 a_3294_n9389# a_3289_n9989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6157 a_11_n6141# a_18_n6359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6158 gnd d0 a_21060_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6159 a_23032_n6722# d2 a_23115_n7738# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6160 a_19970_4536# d0 a_20772_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6161 a_32966_7220# d2 a_33016_6023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6162 a_1659_6548# a_1441_6548# a_1565_6667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6163 a_22996_n7915# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6164 a_13273_3403# a_13275_3921# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6165 a_16357_n7991# a_16361_n7803# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6166 a_32836_n7177# d1 a_32931_n7775# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6167 a_33766_n9627# a_33770_n9439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6168 gnd d0 a_25282_n9618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6169 a_2635_6560# d0 a_3437_6199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6170 a_3239_n6747# a_3492_n6951# a_2442_n6519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6171 a_135_1946# d0 a_624_1840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6172 a_1404_1050# a_1186_1050# a_606_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6173 a_22071_n9315# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6174 a_15342_n4301# d2 a_15392_n3093# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6175 vdd d0 a_29659_n9630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6176 a_19794_n5513# d0 a_20591_n5741# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6177 a_19753_n3665# d0 a_20551_n3481# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6178 a_17907_n8696# a_17689_n8696# a_17426_n8407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6179 a_5542_n6887# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6180 a_14407_n6912# a_14201_n7520# a_13621_n7704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6181 a_12084_1311# a_12341_1121# a_11286_1495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6182 a_18775_1062# d2 a_18858_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6183 a_3457_7217# a_3710_7204# a_2655_7578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6184 a_14687_n5890# a_14469_n5890# a_14584_n7928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6185 a_9929_n3843# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6186 a_7724_2317# a_7981_2127# a_6926_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6187 a_4369_n5537# d0 a_4844_n5643# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6188 a_n32_n3488# a_n27_n4006# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6189 a_19865_7005# d2 a_19948_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6190 a_4346_n4336# d0 a_4827_n4625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6191 a_4970_1247# a_4752_1247# a_4495_1342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6192 a_28694_3543# d0 a_29496_3182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6193 a_31716_4154# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6194 a_24132_n9188# d1 a_24227_n9786# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6195 a_32041_6717# a_31871_7618# a_31995_7737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6196 a_16505_4613# a_16521_5396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6197 a_33692_n5967# a_33696_n5779# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6198 a_13566_5344# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6199 a_24210_n8768# a_24467_n8784# a_24128_n9376# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6200 vdd d0 a_25445_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6201 a_16464_2754# a_16468_2577# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6202 a_17776_2264# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6203 a_19871_4126# d1 a_19957_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6204 a_26555_3913# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6205 vdd d0 a_20863_n6963# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6206 a_19944_8198# a_20201_8008# a_19865_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6207 a_24045_n8360# a_24302_n8376# a_23873_n6138# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6208 a_7530_n2688# a_7544_n3482# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6209 a_30638_3232# a_30644_3415# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6210 a_30646_3933# d0 a_31137_3926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6211 a_5908_4523# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6212 a_9220_5937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6213 a_7544_n3482# a_7548_n3294# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6214 a_13729_1878# a_13511_1878# a_13238_1885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6215 a_179_4200# a_185_4383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6216 a_26518_1877# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6217 a_26301_4938# a_26303_5037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6218 vdd d1 a_20066_n6735# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6219 a_17977_1246# a_17759_1246# a_17496_1158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6220 a_27604_2632# d3 a_27698_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6221 a_6982_5555# d0 a_7784_5194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6222 gnd d0 a_34148_5630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6223 a_16382_n8409# a_16377_n9009# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6224 a_19907_6162# a_20164_5972# a_19861_7182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6225 a_6864_4127# d1 a_6946_3519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6226 a_18812_6560# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6227 a_12215_8260# a_12468_8247# a_11413_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6228 a_10218_5147# a_10000_5147# a_9420_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6229 a_679_5306# a_461_5306# a_204_5401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6230 a_33058_3556# d0 a_33860_3195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6231 a_30541_n9245# d0 a_31030_n9340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6232 a_10126_n7915# d3 a_10220_n7915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6233 a_25205_8437# a_25209_8260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6234 a_13728_2290# a_13510_2290# a_13253_2385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6235 gnd d0 a_29785_5205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6236 gnd d1 a_24357_n2676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6237 a_1322_3496# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6238 gnd d0 a_16795_6224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6239 a_7527_n2464# a_7531_n2276# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6240 a_31922_3665# a_31716_4154# a_31136_4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6241 a_12951_197# d6 a_8658_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6242 a_4572_6031# a_4579_6249# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6243 a_13622_n7292# a_13404_n7292# a_13131_n7098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6244 gnd d1 a_33295_2348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6245 a_13784_5344# a_13566_5344# a_13309_5439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6246 a_21680_184# a_21462_184# a_21581_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6247 a_14509_1088# a_14291_1088# a_13712_860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6248 a_15597_n9799# d0 a_16395_n9615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6249 gnd d0 a_8000_3557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6250 a_14381_6178# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6251 a_14366_n4699# a_14148_n4466# a_13569_n4238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6252 a_22396_3901# a_22178_3901# a_21905_3908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6253 a_33895_5643# a_33909_6426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6254 a_21981_n4225# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6255 vdd d0 a_21060_6610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6256 a_8982_7462# d0 a_9457_7367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6257 vdd d0 a_33986_n7607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6258 a_24158_n5526# d0 a_24951_n5942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6259 vdd d0 a_7857_n6552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6260 a_8236_n2045# d0 a_9168_n2189# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6261 a_10916_n10590# a_12949_n10693# a_8244_n10653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6262 a_22921_1075# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6263 a_27371_5159# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6264 vdd d0 a_12234_n6564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6265 a_18780_1591# a_18574_2080# a_17994_2264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6266 a_28426_5173# a_28683_4983# a_27833_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6267 a_28426_n8184# d2 a_28509_n9200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6268 a_23869_n6326# a_24126_n6342# a_23811_n10590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6269 a_1006_n2392# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6270 a_9239_7367# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6271 a_24971_n6548# a_24975_n6360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6272 a_9167_n2601# a_8949_n2601# a_8686_n2312# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6273 a_28_n7159# a_35_n7377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6274 a_6858_7006# a_7111_6993# a_6682_4972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6275 a_20808_6211# a_20803_6800# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6276 a_1096_n7482# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6277 a_1364_n5852# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6278 gnd d0 a_3510_n7557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6279 a_23176_3111# a_22958_3111# a_22379_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6280 a_444_n3182# a_226_n3182# a_n45_n3087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6281 a_21322_n10664# d5 a_23317_n5877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6282 a_22251_n7691# a_22033_n7691# a_21776_n7585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6283 a_26297_4420# a_26301_4938# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6284 gnd d0 a_16759_4188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6285 a_11400_7426# d0 a_12193_7831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6286 a_10136_7593# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6287 a_26065_n3025# a_26067_n3124# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6288 a_21851_854# a_25078_1311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6289 a_31917_6598# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6290 a_n38_n3305# a_n32_n3488# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6291 a_5686_3509# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6292 a_20717_1533# a_20731_2316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6293 gnd d5 a_11074_n10606# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6294 a_30468_n5173# d0 a_30957_n5268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6295 a_10053_n3843# d3 a_10147_n3843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6296 a_11303_2513# d0 a_12105_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6297 gnd d0 a_29749_3169# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6298 a_29385_n8596# a_29642_n8612# a_28587_n8780# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6299 a_2549_1293# a_2802_1280# a_2463_2078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6300 a_11028_n3080# a_11281_n3284# a_10978_n4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6301 gnd d4 a_19762_n6329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6302 vdd d0 a_20971_1108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6303 a_33822_1571# a_33836_2354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6304 a_30697_6469# d0 a_31172_6374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6305 a_1266_n4838# a_1060_n5446# a_480_n5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6306 a_12178_6224# a_12173_6813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6307 vdd d0 a_34148_5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6308 a_18467_n7494# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6309 a_30609_1897# a_30611_1996# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6310 gnd d1 a_20210_3328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6311 a_32858_n3703# d0 a_33656_n3519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6312 a_26809_5949# a_26591_5949# a_26320_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6313 a_25191_7654# a_25444_7641# a_24394_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6314 gnd d2 a_33126_n9417# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6315 a_13260_3002# d0 a_13749_2896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6316 vdd d0 a_33933_n4553# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6317 a_425_3270# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6318 a_33908_6838# a_33912_6661# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6319 a_8782_n7585# a_8787_n8103# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6320 gnd d1 a_15944_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6321 a_14584_n7928# a_14366_n7928# a_14490_n7928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6322 a_30697_6469# a_30702_6793# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6323 a_28472_n7164# d1 a_28571_n7574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6324 vdd d0 a_16795_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6325 a_31773_n6747# a_31555_n6514# a_30976_n6286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6326 vdd d0 a_7784_n2480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6327 a_25095_2329# a_25352_2139# a_24297_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6328 a_17543_3994# a_17550_4212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6329 a_9981_4129# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6330 a_13160_n8433# d0 a_13641_n8722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6331 a_30738_n5680# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6332 a_9003_n5655# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6333 a_32794_5009# a_33047_4996# a_32197_296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6334 a_9278_n8297# d1 a_10075_n8758# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6335 a_12087_1546# a_12101_2329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6336 a_5856_2608# a_5686_3509# a_5810_3628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6337 a_4410_n8091# d0 a_4901_n8285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6338 a_13642_n8310# a_13424_n8310# a_13153_n8215# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6339 a_22179_n3207# a_21961_n3207# a_21688_n3013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6340 a_30881_2302# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6341 a_13267_3220# d0 a_13748_3308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6342 a_9294_n9727# a_9076_n9727# a_8819_n9621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6343 vdd d1 a_15727_n2689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6344 a_11065_n5116# d1 a_11160_n5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6345 a_17925_n9302# a_17707_n9302# a_17434_n9108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6346 a_4519_2977# d0 a_5008_2871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6347 gnd d0 a_29532_n2504# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6348 a_31963_2526# d3 a_32062_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6349 a_19727_n7327# a_19984_n7343# a_19681_n8347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6350 a_28188_n10602# a_28445_n10618# a_28287_n10602# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6351 a_8765_n6567# a_8767_n7085# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6352 a_12173_6813# a_12177_6636# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6353 a_17489_940# a_17496_1158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6354 a_30541_n9245# a_30548_n9463# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6355 a_22758_n3435# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6356 a_23069_n8758# a_22851_n8525# a_22272_n8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6357 gnd d6 a_4208_n10668# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6358 a_15595_7208# d2 a_15645_6011# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6359 a_7036_8609# a_7293_8419# a_6941_8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6360 a_4526_3195# d0 a_5007_3283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6361 a_23279_4535# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6362 a_32862_n3515# d0 a_33659_n3743# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6363 a_11055_n8172# a_11308_n8376# a_10879_n6138# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6364 a_27419_n3678# a_27217_n2839# a_27341_n2839# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6365 a_11327_3354# d0 a_12124_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6366 a_14210_n2840# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6367 a_2386_n3465# d0 a_3179_n3881# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6368 a_32763_n3105# d1 a_32862_n3515# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6369 a_19685_5148# d3 a_19788_3110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6370 a_3342_1698# a_3599_1508# a_2549_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6371 a_2310_n8335# d2 a_2356_n7315# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6372 a_3162_n2863# a_3419_n2879# a_2369_n2447# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6373 a_18015_2870# a_17797_2870# a_17526_2976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6374 a_26828_7379# d1 a_27626_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6375 a_6647_n3256# d1 a_6733_n2460# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6376 a_16377_n9009# a_16634_n9025# a_15584_n8593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6377 a_2283_n3243# a_2540_n3259# a_2237_n4263# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6378 a_17212_n839# d8 a_8343_n10653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6379 a_9474_8385# a_9256_8385# a_8993_8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6380 gnd d1 a_11490_n9802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6381 a_2134_n6301# d3 a_2237_n4263# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6382 a_426_n2576# a_208_n2576# a_n55_n2287# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6383 a_23217_5676# a_23011_6165# a_22431_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6384 a_28689_8046# d1 a_28784_8633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6385 a_n62_n2069# a_n55_n2287# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6386 a_11400_7426# d0 a_12197_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6387 a_20555_n3293# a_20550_n3893# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6388 a_29581_8861# a_29585_8684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6389 a_10026_1485# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6390 a_7040_8432# d0 a_7837_8660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6391 a_14670_6705# a_14500_7606# a_14624_7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6392 a_4881_n7267# a_4663_n7267# a_4390_n7073# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6393 a_15461_n7353# d1 a_15543_n6745# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6394 a_6856_n9774# d0 a_7654_n9590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6395 a_481_n5218# a_263_n5218# a_n8_n5123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6396 a_3347_1109# a_3342_1698# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6397 a_23811_n10590# a_24068_n10606# a_21322_n10664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6398 a_26318_5956# a_26320_6055# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6399 vdd d1 a_2659_n4687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6400 a_28571_n7574# d0 a_29364_n7990# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6401 a_13160_n8433# a_13166_n8616# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6402 a_21798_n9121# a_21800_n9220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6403 a_2545_1470# a_2802_1280# a_2463_2078# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6404 a_21421_n10664# d6 a_19546_n10577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6405 a_26190_n9633# d0 a_26665_n9739# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6406 a_22235_n6261# a_22017_n6261# a_21746_n6166# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6407 a_18431_n5458# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6408 a_4210_172# a_5966_259# a_6085_259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6409 a_25187_7831# a_25444_7641# a_24394_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6410 gnd d0 a_12358_2139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6411 a_17852_n5230# a_17634_n5230# a_17361_n5036# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6412 a_4599_7267# a_4605_7450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6413 gnd d0 a_25265_n8600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6414 a_29384_n9008# a_29388_n8820# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6415 a_2419_n5689# a_2676_n5705# a_2324_n5091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6416 a_19654_n3255# a_19911_n3271# a_19608_n4275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6417 a_17887_7960# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6418 a_10007_n4863# a_9801_n5471# a_9221_n5655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6419 a_19505_n6313# d3 a_19608_n4275# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6420 a_9129_1259# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6421 vdd d1 a_15944_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6422 a_1261_n7890# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6423 a_22252_n7279# a_22034_n7279# a_21761_n7085# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6424 a_32790_5186# d3 a_32893_3148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6425 gnd d0 a_12414_5193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6426 a_1142_n4838# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6427 a_22996_n7915# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6428 a_660_4288# a_442_4288# a_179_4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6429 a_21734_n5366# a_21740_n5549# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6430 a_4607_7968# d0 a_5098_7961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6431 a_8883_2189# d0 a_9364_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6432 a_11237_n9598# a_11490_n9802# a_11138_n9188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6433 a_19834_2090# d1 a_19916_1482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6434 a_13296_5038# a_13303_5256# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6435 a_6860_n9586# d0 a_4447_n9933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6436 gnd d0 a_34129_4612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6437 a_22233_7367# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6438 a_4609_n4625# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6439 a_9929_n3843# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6440 a_10187_3640# a_9981_4129# a_9401_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6441 vdd d1 a_24430_n6748# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6442 a_2676_8419# a_2929_8406# a_2577_8009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6443 a_30674_5268# a_30680_5451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6444 a_4352_n4519# d0 a_4827_n4625# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6445 gnd d2 a_28869_3961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6446 a_4326_n3318# d0 a_4807_n3607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6447 a_2421_2921# a_2674_2908# a_2314_5136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6448 a_11359_5567# a_11616_5377# a_11277_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6449 a_25007_n8996# a_25011_n8808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6450 a_21746_n6166# a_21753_n6384# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6451 a_21723_n4531# a_21725_n5049# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6452 a_13116_n6179# a_13123_n6397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6453 a_18105_7960# d1 a_18890_7699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6454 a_6720_n7328# d1 a_6806_n6532# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6455 a_26756_2895# a_26538_2895# a_26265_2708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6456 a_3162_n2863# a_3166_n2675# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6457 a_13765_4326# a_13547_4326# a_13290_4421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6458 a_680_4894# d1 a_1477_5122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6459 a_11908_n2288# a_11903_n2888# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6460 a_9347_1259# a_9129_1259# a_8872_1354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6461 a_16501_4790# a_16505_4613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6462 a_11376_6585# a_11633_6395# a_11281_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6463 a_18513_n4850# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6464 a_11925_n3306# a_12178_n3510# a_11123_n3678# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6465 a_2562_2488# d0 a_3360_2304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6466 a_29509_4377# a_29766_4187# a_28711_4561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6467 a_2490_7170# d2 a_2536_6150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6468 gnd d2 a_28942_8033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6469 gnd d0 a_3456_n4915# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6470 a_8716_n4130# a_8723_n4348# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6471 a_30322_209# a_32078_296# a_32197_296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6472 a_17690_n8284# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6473 a_28689_8046# d1 a_28788_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6474 a_26755_3307# a_26537_3307# a_26280_3402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6475 a_10228_2501# a_10026_1485# a_10145_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6476 a_25024_n10014# a_25281_n10030# a_24231_n9598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6477 a_17978_834# a_17760_834# a_17489_940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6478 a_15723_5580# d0 a_16521_5396# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6479 a_18673_n6886# d2 a_18751_n7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6480 a_4970_1247# d1 a_5768_1063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6481 a_13253_2385# d0 a_13728_2290# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6482 a_9437_6349# d1 a_10223_5676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6483 a_19689_4971# d3 a_19865_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6484 a_24018_n3268# d1 a_24100_n2660# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6485 a_221_6419# d0 a_696_6324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6486 a_19764_n9363# d1 a_19846_n8755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6487 a_427_n2164# a_209_n2164# gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6488 a_6900_6163# a_7157_5973# a_6854_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6489 a_16267_n2901# a_16271_n2713# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6490 a_33752_n8833# a_34005_n9037# a_32955_n8605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6491 a_7548_n3294# a_7543_n3894# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6492 a_17797_n2588# a_17579_n2588# a_17322_n2482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6493 a_26243_1366# d0 a_26718_1271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6494 a_32976_4164# a_33233_3974# a_32897_2971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6495 a_5044_4907# a_4826_4907# a_4553_4914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6496 a_18656_1472# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6497 vdd d4 a_28503_n6354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6498 gnd d0 a_20827_n4927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6499 a_11235_7018# a_11488_7005# a_11059_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6500 a_19850_n8567# d0 a_20647_n8795# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6501 vdd d0 a_16777_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6502 gnd d2 a_33306_8046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6503 a_23144_1604# d2 a_23222_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6504 gnd d0 a_25334_1533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6505 a_22958_3111# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6506 a_23047_n3843# a_22877_n4863# a_23001_n4863# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6507 a_21981_n4225# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6508 a_10327_2501# d4 a_10467_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6509 gnd d1 a_20030_n4699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6510 a_2639_6383# d0 a_3436_6611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6511 a_21961_n3207# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6512 a_5623_5135# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6513 gnd d0 a_25227_n6976# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6514 a_11179_n6732# d0 a_11981_n6360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6515 a_11097_n7340# a_11354_n7356# a_11051_n8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6516 a_28550_n6744# d0 a_29348_n6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6517 a_24898_n2476# a_24902_n2288# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6518 a_2076_n10565# d4 a_2134_n6301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6519 a_24141_n4508# d0 a_24934_n4924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6520 a_2320_n5279# d1 a_2402_n4671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6521 a_10561_271# a_10343_271# a_10467_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6522 a_15423_4997# a_15676_4984# a_14826_284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6523 a_29472_2341# a_29476_2164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6524 a_30511_n7427# a_30517_n7610# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6525 a_18973_258# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6526 a_9205_n4225# a_8987_n4225# a_8716_n4130# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6527 a_19773_n4683# d0 a_20571_n4499# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6528 vdd d0 a_34129_4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6529 a_22851_n8525# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6530 a_27397_1497# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6531 a_24411_8444# d0 a_25208_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6532 a_21978_7980# a_21980_8079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6533 a_16395_n9615# a_16652_n9631# a_15597_n9799# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6534 gnd d1 a_2695_n6723# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6535 a_1276_6140# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6536 a_20786_5782# a_21043_5592# a_19993_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6537 a_7837_8660# a_8090_8647# a_7040_8432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6538 a_18858_2488# a_18656_1472# a_18780_1591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6539 a_168_3365# a_170_3883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6540 a_30592_879# a_30594_978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6541 gnd d1 a_2912_7388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6542 a_9784_n4453# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6543 vdd d0 a_29605_n6576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6544 a_30494_n6409# a_30500_n6592# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6545 a_30500_n6592# a_30502_n7110# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6546 a_6839_n8756# d0 a_7641_n8384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6547 a_1602_246# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6548 a_30939_n4662# d1 a_31737_n4711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6549 a_31136_4338# a_30918_4338# a_30655_4250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6550 a_19447_n10577# d4 a_19505_n6313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6551 a_21853_953# d0 a_22342_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6552 gnd d0 a_29658_n10042# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6553 a_17506_1958# d0 a_17995_1852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6554 gnd d0 a_12198_n4528# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6555 a_25615_n10665# d6 a_30063_n10689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6556 a_19691_n5291# d1 a_19773_n4683# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6557 a_2562_2488# d0 a_3364_2127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6558 a_2504_3937# a_2757_3924# a_2421_2921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6559 vdd d2 a_28942_8033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6560 a_28554_n6556# d0 a_29351_n6784# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6561 a_33913_6249# a_34166_6236# a_33111_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6562 a_33946_8462# a_33950_8285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6563 a_31192_7392# a_30974_7392# a_30711_7304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6564 a_29365_n7578# a_29622_n7594# a_28567_n7762# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6565 a_24091_n7340# d1 a_24173_n6732# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6566 a_12084_1311# a_12088_1134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6567 a_30937_5356# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6568 a_1266_n4838# a_1060_n5446# a_481_n5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6569 a_2500_4114# d1 a_2582_3506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6570 a_16378_n8597# a_16382_n8409# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6571 a_24951_n5942# a_24955_n5754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6572 a_11962_n5342# a_12215_n5546# a_11160_n5714# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6573 a_3951_n10652# d5 a_6440_n10578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6574 a_33892_5408# a_33896_5231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6575 a_18848_5134# a_18630_5134# a_18050_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6576 a_30539_n9146# d0 a_31030_n9340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6577 gnd d0 a_12177_n3922# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6578 a_10327_2501# a_10109_2501# a_10228_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6579 a_13584_5950# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6580 a_3273_n8559# a_3277_n8371# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6581 a_15388_n3281# d1 a_15474_n2485# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6582 a_24317_3531# d0 a_25119_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6583 a_6941_8022# a_7194_8009# a_6858_7006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6584 a_5770_n3831# d4 a_5946_n5865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6585 a_13166_n8616# d0 a_13641_n8722# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6586 a_28477_n2672# d0 a_29275_n2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6587 a_9277_n8709# d1 a_10075_n8758# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6588 gnd d1 a_11380_n3694# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6589 a_13140_n7415# d0 a_13621_n7704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6590 a_3420_5181# a_3415_5770# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6591 a_9258_n7279# d1 a_10043_n6899# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6592 a_9294_n9727# a_9076_n9727# a_8813_n9438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6593 a_4616_8285# a_4622_8468# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6594 a_4390_n7073# d0 a_4881_n7267# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6595 a_21870_1971# d0 a_22359_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6596 vdd d2 a_2577_n5295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6597 vdd d2 a_33306_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6598 a_20030_7413# a_20283_7400# a_19944_8198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6599 a_5773_1592# a_5567_2081# a_4988_1853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6600 a_13095_n5062# a_13097_n5161# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6601 a_16304_n4937# a_16308_n4749# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6602 vdd d0 a_25334_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6603 a_4627_n5231# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6604 a_32845_n2497# d0 a_33642_n2725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6605 a_22178_3901# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6606 a_12210_8849# a_12214_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6607 a_33656_n3519# a_33913_n3535# a_32858_n3703# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6608 a_6724_n7140# a_6977_n7344# a_6674_n8348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6609 vdd d0 a_34006_n8625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6610 a_19867_n9585# a_20120_n9789# a_19768_n9175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6611 gnd d0 a_12270_n9012# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6612 a_13313_6056# a_13320_6274# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6613 a_26337_n3631# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6614 gnd d0 a_25281_n10030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6615 a_22140_2277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6616 a_23227_2620# d3 a_23321_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6617 vdd d0 a_16597_n6989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6618 a_9130_847# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6619 a_11957_n5942# a_12214_n5958# a_11164_n5526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6620 a_26136_n6579# d0 a_26611_n6685# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6621 a_29332_n5766# a_29585_n5970# a_28535_n5538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6622 a_15429_n5129# d1 a_15528_n5539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6623 a_11314_8211# d1 a_11396_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6624 a_27480_2513# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6625 a_6766_n4684# d0 a_7568_n4312# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6626 a_7765_4176# a_7760_4765# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6627 a_22341_1259# a_22123_1259# a_21860_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6628 a_11160_n5714# a_11417_n5730# a_11065_n5116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6629 a_4918_n9303# d1 a_5703_n8923# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6630 gnd d0 a_3530_n8575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6631 a_12160_5618# a_12413_5605# a_11363_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6632 a_30554_n9646# a_30559_n9970# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6633 a_28715_4384# d0 a_29508_4789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6634 a_28481_n2484# d0 a_29278_n2712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6635 a_32935_n7587# a_33188_n7791# a_32836_n7177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6636 vdd d0 a_25171_n3922# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6637 a_6682_4972# d3 a_6854_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6638 gnd d0 a_12395_4175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6639 a_32914_n6757# d0 a_33712_n6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6640 vdd d8 a_17382_n10744# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6641 a_9166_3295# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6642 gnd d0 a_25461_8659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6643 a_5_n5524# d0 a_480_n5630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6644 a_22415_4919# a_22197_4919# a_21924_4926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6645 a_18632_n4673# a_18414_n4440# a_17835_n4212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6646 a_10037_7183# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6647 a_25154_5618# a_25168_6401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6648 a_6750_n3478# d0 a_7547_n3706# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6649 a_4390_n7073# a_4392_n7172# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6650 a_18600_n2814# a_18394_n3422# a_17814_n3606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6651 vdd d1 a_33351_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6652 a_6806_n6532# d0 a_7603_n6760# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6653 a_4605_7450# d0 a_5080_7355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6654 a_1339_n8910# a_1133_n9518# a_554_n9290# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6655 a_24394_7426# a_24647_7413# a_24308_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6656 a_30466_n5074# d0 a_30957_n5268# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6657 a_31083_872# d1 a_31880_1100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6658 a_33909_6426# a_34166_6236# a_33111_6610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6659 a_17815_n3194# a_17597_n3194# a_17326_n3099# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6660 vdd d1 a_2639_n3669# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6661 a_32614_n6163# d3 a_32790_n8197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6662 a_27631_7724# d2 a_27677_6704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6663 a_18014_3282# d1 a_18812_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6664 a_22235_n6261# a_22017_n6261# a_21744_n6067# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6665 a_27833_283# d4 a_28426_5173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6666 a_2356_n7315# a_2613_n7331# a_2310_n8335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6667 a_13093_n4544# d0 a_13568_n4650# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6668 a_24210_n8768# d0 a_25008_n8584# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6669 vdd d0 a_29784_5617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6670 a_13067_n3343# d0 a_13548_n3632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6671 a_24935_n4512# a_25192_n4528# a_24137_n4696# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6672 a_2500_4114# d1 a_2586_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6673 a_10007_n4863# a_9801_n5471# a_9222_n5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6674 a_2573_8186# a_2830_7996# a_2494_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6675 gnd d0 a_25245_n7582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6676 a_661_3876# d1 a_1446_3615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6677 vdd d0 a_3529_n8987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6678 a_4332_n3501# a_4337_n4019# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6679 a_554_n9290# a_336_n9290# a_65_n9195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6680 a_33896_5231# a_33891_5820# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6681 a_6651_n3068# a_6904_n3272# a_6601_n4276# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6682 a_30631_3014# a_30638_3232# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6683 a_15605_4152# a_15862_3962# a_15526_2959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6684 a_1441_3086# a_1223_3086# a_644_2858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6685 a_22959_n2650# a_22741_n2417# a_22161_n2601# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6686 a_15704_4562# d0 a_16502_4378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6687 a_3289_n9989# a_3546_n10005# a_2496_n9573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6688 a_4609_n4625# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6689 a_32197_296# d4 a_32790_5186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6690 a_21673_n2094# a_21680_n2312# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6691 a_26147_n7414# a_26153_n7597# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6692 a_4589_n3607# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6693 a_7599_n6948# a_7603_n6760# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6694 a_7728_2140# a_7981_2127# a_6926_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6695 a_26291_4237# a_26297_4420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6696 a_5008_2871# a_4790_2871# a_4517_2684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6697 a_4332_n3501# d0 a_4807_n3607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6698 a_8903_3207# a_8909_3390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6699 a_1409_1579# d2 a_1487_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6700 a_28694_3543# d0 a_29492_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6701 a_19875_3949# a_20128_3936# a_19792_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6702 a_7584_n5742# a_7837_n5946# a_6787_n5514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6703 a_29329_n5542# a_29333_n5354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6704 a_32882_n4533# d0 a_33679_n4761# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6705 a_8750_n6067# a_8752_n6166# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6706 a_2406_n4483# d0 a_3199_n4899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6707 a_11314_8211# d1 a_11400_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6708 vdd d2 a_15898_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6709 gnd d0 a_25445_7229# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6710 a_14210_n2840# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6711 a_16485_3360# a_16489_3183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6712 vdd d0 a_16758_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6713 a_11110_n2472# a_11363_n2676# a_11024_n3268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6714 a_19871_4126# d1 a_19953_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6715 a_20755_3157# a_20750_3746# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6716 a_5007_3283# a_4789_3283# a_4532_3378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6717 a_26136_n6579# a_26138_n7097# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6718 gnd d3 a_20045_2920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6719 a_5604_4117# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6720 a_7834_8425# a_7838_8248# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6721 a_5744_n7726# d3 a_5843_n7903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6722 a_14582_5160# d2 a_14665_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6723 vdd d7 a_8501_n10669# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6724 a_26297_4420# d0 a_26772_4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6725 a_153_2671# a_155_2964# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6726 vdd d0 a_12395_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6727 a_9837_n7507# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6728 a_17887_7960# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6729 a_1487_2476# d3 a_1586_2476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6730 a_21759_n6567# a_21761_n7085# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6731 a_11962_n5342# a_11957_n5942# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6732 a_10306_6692# a_10136_7593# a_10260_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6733 a_8949_6043# d0 a_9438_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6734 a_5660_7171# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6735 a_15645_6011# d1 a_15740_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6736 a_716_7342# a_498_7342# a_235_7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6737 a_17606_7266# a_17612_7449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6738 gnd d3 a_28786_2945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6739 a_8939_5243# d0 a_9420_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6740 vdd d0 a_8090_8647# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6741 a_22741_n2417# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6742 a_23144_1604# a_22938_2093# a_22359_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6743 a_24390_7603# a_24647_7413# a_24308_8211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6744 a_19731_n7139# d1 a_19826_n7737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6745 a_16542_6237# a_16795_6224# a_15740_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6746 a_13153_n8215# a_13160_n8433# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6747 a_21944_n2189# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6748 a_28648_6187# d1 a_28730_5579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6749 a_5841_5135# d2 a_5924_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6750 a_13821_7380# a_13603_7380# a_13340_7292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6751 vdd d4 a_2391_n6317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6752 a_26184_n9450# d0 a_26665_n9739# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6753 a_19830_n7549# d0 a_20627_n7777# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6754 a_33909_6426# a_33913_6249# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6755 a_24177_n6544# d0 a_24970_n6960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6756 a_31917_3136# d2 a_31968_2645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6757 a_18667_7170# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6758 a_23047_n3843# a_22877_n4863# a_22996_n4686# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6759 a_24045_n8360# d2 a_24091_n7340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6760 a_24897_n2888# a_25154_n2904# a_24104_n2472# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6761 a_33643_n2313# a_33638_n2913# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6762 a_23249_7183# d2 a_23300_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6763 a_17852_n5230# a_17634_n5230# a_17363_n5135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6764 a_21796_n8603# d0 a_22271_n8709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6765 a_21961_n3207# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6766 a_22272_n8297# a_22054_n8297# a_21781_n8103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6767 gnd d1 a_20010_n3681# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6768 a_5097_8373# a_4879_8373# a_4616_8285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6769 a_32202_415# a_32020_4560# a_32062_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6770 a_24312_8034# d1 a_24407_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6771 a_27591_n7927# d4 a_27694_n5889# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6772 a_1142_n4838# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6773 a_24121_n3490# d0 a_24914_n3906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6774 a_14418_8214# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6775 a_17597_6755# d0 a_18088_6942# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6776 a_2287_n3055# d1 a_2382_n3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6777 a_26140_n7196# d0 a_26629_n7291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6778 a_30992_7998# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6779 a_8889_2372# a_8894_2696# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6780 a_30918_4338# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6781 a_10301_6573# d3 a_10400_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6782 a_9205_n4225# a_8987_n4225# a_8714_n4031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6783 a_13340_7292# a_13346_7475# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6784 a_29406_n9426# a_29659_n9630# a_28604_n9798# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6785 gnd d1 a_20173_1292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6786 a_33950_8285# a_34203_8272# a_33148_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6787 a_22851_n8525# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6788 a_20554_n3705# a_20807_n3909# a_19757_n3477# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6789 a_17580_n2176# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6790 a_2365_n2635# a_2622_n2651# a_2283_n3243# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6791 gnd d0 a_20900_n8999# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6792 a_9185_n3207# a_8967_n3207# a_8696_n3112# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6793 a_5744_n7726# a_5542_n6887# a_5661_n6710# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6794 gnd d2 a_24492_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6795 a_9919_n6899# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6796 a_30421_n2337# d0 a_30902_n2626# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6797 a_125_1146# d0 a_606_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6798 a_9040_n7279# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6799 a_27408_7195# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6800 a_18817_3627# a_18611_4116# a_18031_4300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6801 a_2479_n8555# d0 a_3272_n8971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6802 gnd d2 a_11461_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6803 a_17489_940# d0 a_17978_834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6804 a_33876_4625# a_33892_5408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6805 a_30991_8410# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6806 a_31519_n4478# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6807 a_9784_n4453# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6808 vdd d2 a_6941_n5308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6809 a_7779_5783# a_8036_5593# a_6986_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6810 a_9764_n3435# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6811 a_17504_1859# a_17506_1958# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6812 a_2134_n6301# a_2391_n6317# a_2076_n10565# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6813 a_8969_7061# a_8976_7279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6814 a_25077_1723# a_25081_1546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6815 a_6819_n7738# d0 a_7621_n7366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6816 vdd d2 a_11318_n5320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6817 a_11204_2103# a_11461_1913# a_11158_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6818 a_20534_n2463# a_20538_n2275# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6819 a_10147_n3843# a_9929_n3843# a_10053_n3843# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6820 a_33855_3784# a_34112_3594# a_33062_3379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6821 a_18739_2488# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6822 a_24357_5390# d0 a_25150_5795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6823 vdd d1 a_20300_8418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6824 a_9278_n8297# a_9060_n8297# a_8789_n8202# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6825 a_18890_7699# a_18684_8188# a_18104_8372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6826 a_16489_3183# a_16484_3772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6827 a_18513_n4850# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6828 a_11303_2513# d0 a_12101_2329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6829 a_17592_6431# a_17597_6755# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6830 a_19658_n3067# d1 a_19753_n3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6831 a_8658_196# a_12832_197# a_10561_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6832 a_29582_8449# a_29586_8272# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6833 a_15465_n7165# a_15718_n7369# a_15415_n8373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6834 a_7728_2140# a_7723_2729# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6835 a_14670_6705# d3 a_14764_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6836 a_28533_2958# d2 a_28616_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6837 a_16268_n2489# a_16525_n2505# a_15470_n2673# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6838 a_20824_7406# a_20828_7229# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6839 a_19813_n6531# a_20066_n6735# a_19727_n7327# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6840 a_4506_2177# d0 a_4987_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6841 a_8343_n10653# a_17382_n10744# a_17212_n839# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6842 a_21581_184# a_23337_271# a_23456_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6843 a_4436_n9426# a_4442_n9609# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6844 a_30702_6793# d0 a_31193_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6845 a_3200_n4487# a_3204_n4299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6846 a_17870_n6660# a_17652_n6660# a_17389_n6371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6847 a_9241_n6261# d1 a_10038_n6722# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6848 vdd d1 a_24484_n9802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6849 a_28579_1938# a_28832_1925# a_28529_3135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6850 a_31012_n8734# d1 a_31810_n8783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6851 a_30734_8505# d0 a_31209_8410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6852 vdd d0 a_16562_n4541# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6853 a_30993_n7304# d1 a_31778_n6924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6854 gnd d5 a_6697_n10594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6855 a_5929_6680# d3 a_6023_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6856 a_16345_n6373# a_16340_n6973# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6857 a_5843_n7903# d4 a_5946_n5865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6858 a_13712_860# d1 a_14509_1088# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6859 a_16538_6414# a_16795_6224# a_15740_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6860 a_2241_n4075# d2 a_2324_n5091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6861 gnd d0 a_3726_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6862 a_33715_n6797# a_33729_n7591# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6863 a_19505_n6313# a_19762_n6329# a_19447_n10577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6864 a_25099_2152# a_25352_2139# a_24297_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6865 a_13146_n7598# d0 a_13621_n7704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6866 a_4826_4907# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6867 a_9257_n7691# d1 a_10043_n6899# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6868 a_22379_2883# a_22161_2883# a_21888_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6869 a_6854_7183# d2 a_6904_5986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6870 a_4392_n7172# d0 a_4881_n7267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6871 a_11237_n9598# d0 a_12030_n10014# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6872 a_1544_4510# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6873 a_4770_1853# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6874 a_4590_6756# a_4592_7049# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6875 a_4425_n8591# a_4427_n9109# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6876 a_26067_n3124# d0 a_26556_n3219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6877 a_32869_n9401# a_33126_n9417# a_32790_n8197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6878 a_4627_n5231# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6879 a_30902_2908# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6880 a_11055_n8172# d2 a_11134_n9376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6881 a_29528_5395# a_29785_5205# a_28730_5579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6882 a_12194_7419# a_12198_7242# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6883 a_7023_7414# a_7276_7401# a_6937_8199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6884 a_17798_n2176# a_17580_n2176# a_16977_n2070# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6885 a_27492_n7750# d3 a_27591_n7927# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6886 a_1229_n2802# a_1023_n3410# a_444_n3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6887 a_26337_n3631# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6888 a_27672_6585# a_27470_5569# a_27594_5688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6889 a_15415_n8373# d2 a_15465_n7165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6890 a_24312_8034# d1 a_24411_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6891 gnd d0 a_12250_n7994# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6892 a_22378_3295# a_22160_3295# a_21903_3390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6893 a_22452_6955# a_22234_6955# a_21961_6768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6894 a_17592_6431# d0 a_18067_6336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6895 a_405_2252# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6896 a_32895_n5739# d0 a_33697_n5367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6897 a_33712_n6573# a_33716_n6385# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6898 vdd d1 a_33388_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6899 a_15239_n6339# d3 a_15346_n4113# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6900 a_27838_402# d5 a_27932_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6901 a_11059_4984# a_11312_4971# a_10462_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6902 a_7040_8432# a_7293_8419# a_6941_8022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6903 a_19030_6560# a_18812_6560# a_18936_6679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6904 a_10002_n7915# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6905 a_11327_3354# d0 a_12120_3759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6906 a_30504_n7209# a_30511_n7427# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6907 a_5497_n9531# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6908 a_33946_8462# a_34203_8272# a_33148_8646# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6909 a_5550_1063# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6910 a_3200_n4487# a_3457_n4503# a_2402_n4671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6911 a_13510_2290# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6912 a_4917_n9715# d1 a_5703_n8923# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6913 a_28747_6597# d0 a_29545_6413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6914 a_479_5912# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6915 a_32897_2971# d2 a_32976_4164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6916 gnd d1 a_28861_n9814# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6917 gnd d2 a_33016_n3309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6918 a_1302_n6874# a_1096_n7482# a_516_n7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6919 a_116_829# a_118_928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6920 a_12018_n8396# a_12271_n8600# a_11216_n8768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6921 a_15601_n9611# d0 a_13188_n9958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6922 a_19993_5377# d0 a_20790_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6923 a_17436_n9207# a_17443_n9425# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6924 a_7040_8432# d0 a_7833_8837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6925 a_26500_1271# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6926 a_18858_2488# d3 a_18957_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6927 gnd d0 a_3637_3132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6928 a_13584_5950# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6929 a_18600_n2814# a_18394_n3422# a_17815_n3194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6930 a_8976_7279# a_8982_7462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6931 a_15502_n9201# d1 a_15601_n9611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6932 a_30203_209# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6933 a_21939_5426# d0 a_22414_5331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6934 a_22342_847# a_22124_847# a_21851_854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6935 a_30592_879# d0 a_31083_872# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6936 a_623_2252# a_405_2252# a_148_2347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6937 vdd d2 a_20021_n9379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6938 a_29585_8684# a_29838_8671# a_28788_8456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6939 a_26574_4931# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6940 a_29586_8272# a_29581_8861# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6941 a_4791_n2177# d1 a_5588_n2638# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6942 a_6802_n6720# a_7059_n6736# a_6720_n7328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6943 gnd d0 a_33949_n5983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6944 a_13073_n3526# d0 a_13548_n3632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6945 a_17995_1852# a_17777_1852# a_17504_1859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6946 a_17623_8284# a_17629_8467# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6947 a_24190_n7750# d0 a_24988_n7566# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6948 a_14308_2106# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6949 a_14691_2514# d4 a_14831_403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6950 a_33111_6610# d0 a_33909_6426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6951 a_24915_n3494# a_25172_n3510# a_24117_n3678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6952 a_2314_n8147# d2 a_2397_n9163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6953 a_3872_n2032# d0 a_4791_n2177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6954 a_24971_n6548# a_25228_n6564# a_24173_n6732# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6955 a_11179_n6732# a_11436_n6748# a_11097_n7340# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6956 a_14364_5160# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6957 gnd d0 a_7800_n3910# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6958 a_18673_n6886# a_18467_n7494# a_17887_n7678# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6959 vdd d0 a_3509_n7969# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6960 vdd d1 a_24537_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6961 a_33933_7267# a_33928_7856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6962 a_30864_1284# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6963 a_22469_7973# a_22251_7973# a_21980_8079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6964 a_31788_n3868# d3 a_31882_n3868# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6965 vdd d0 a_3726_8634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6966 gnd d3 a_6858_n4292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6967 vdd d3 a_2567_n8351# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6968 a_22959_n2650# a_22741_n2417# a_22162_n2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6969 a_33016_6023# a_33269_6010# a_32966_7220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6970 a_26085_n4043# d0 a_26576_n4237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6971 a_6858_7006# d2 a_6937_8199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6972 a_2655_7578# a_2912_7388# a_2573_8186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6973 a_18775_1062# a_18557_1062# a_17978_834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6974 a_19736_n2647# d0 a_20538_n2275# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6975 gnd d3 a_11235_n4304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6976 a_4589_n3607# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6977 a_6946_3519# d0 a_7744_3335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6978 a_7796_6801# a_7800_6624# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6979 a_4844_n5643# d1 a_5630_n4851# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6980 a_8920_4225# d0 a_9401_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6981 a_27771_6585# a_27553_6585# a_27672_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6982 a_8986_8079# d0 a_9475_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6983 a_26347_7291# d0 a_26828_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6984 a_33642_n2725# a_33895_n2929# a_32845_n2497# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6985 a_12198_7242# a_12193_7831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6986 a_1726_365# d5 a_1820_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6987 a_20627_n7777# a_20644_n8571# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6988 a_18766_7580# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6989 a_7764_4588# a_7780_5371# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6990 a_14514_1617# a_14308_2106# a_13728_2290# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6991 a_11363_5390# a_11616_5377# a_11277_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6992 a_19685_n8159# d2 a_19768_n9175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6993 a_10038_n6722# a_9820_n6489# a_9241_n6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6994 gnd d0 a_34093_2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6995 a_16579_8273# a_16832_8260# a_15777_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X6996 a_8993_8297# d0 a_9474_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6997 a_23873_n6138# d3 a_24049_n8172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6998 a_21686_n2495# a_21688_n3013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X6999 a_32878_n4721# a_33135_n4737# a_32796_n5329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7000 a_28747_6597# d0 a_29549_6236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7001 a_27516_1087# a_27298_1087# a_26718_1271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7002 a_389_822# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7003 a_5749_n7903# d3 a_5843_n7903# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7004 a_9837_n7507# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7005 a_29569_7254# a_29822_7241# a_28767_7615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7006 a_30757_n6698# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7007 gnd d3 a_7038_2921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7008 gnd d0 a_21097_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7009 vdd d0 a_3637_3132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7010 a_16506_4201# a_16501_4790# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7011 a_22197_4919# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7012 a_11980_n6772# a_12233_n6976# a_11183_n6544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7013 a_32790_n8197# a_33043_n8401# a_32614_n6163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7014 a_10323_n5877# a_11074_n10606# a_10916_n10590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7015 a_26184_n9450# a_26190_n9633# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7016 a_n1_n5341# d0 a_480_n5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7017 a_4879_8373# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7018 a_7636_n8984# a_7640_n8796# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7019 a_18632_n4673# a_18414_n4440# a_17834_n4624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7020 a_22741_n2417# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7021 a_30539_n9146# a_30541_n9245# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7022 a_28481_n2484# a_28734_n2688# a_28395_n3280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7023 a_4917_n9715# a_4699_n9715# a_4442_n9609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7024 a_226_6743# d0 a_717_6930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7025 a_1339_n8910# a_1133_n9518# a_553_n9702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7026 a_12613_n2057# a_11904_n2476# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7027 a_29581_8861# a_29838_8671# a_28788_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7028 a_16452_1147# a_16447_1736# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7029 a_29364_n7990# a_29368_n7802# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7030 a_13087_n4361# d0 a_13568_n4650# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7031 a_32759_n3293# d1 a_32845_n2497# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7032 a_21853_953# a_21860_1171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7033 a_9964_3111# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7034 a_2622_5365# d0 a_3415_5770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7035 gnd d0 a_16777_5618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7036 a_33111_6610# d0 a_33913_6249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7037 a_13331_6781# d0 a_13822_6968# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7038 vdd d3 a_2494_n4279# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7039 a_23103_2501# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7040 a_5677_8189# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7041 a_26057_n2324# a_26063_n2507# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7042 a_1307_n3641# a_1105_n2802# a_1229_n2802# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7043 a_4645_n6661# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7044 gnd d1 a_11473_n8784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7045 a_443_3876# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7046 a_27476_n5889# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7047 a_21776_n7585# d0 a_22251_n7691# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7048 vout a_17093_n839# a_17217_n720# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7049 a_5966_259# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7050 a_13530_3308# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7051 a_22814_n6489# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7052 a_7640_n8796# a_7893_n9000# a_6843_n8568# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7053 a_20718_1121# a_20971_1108# a_19916_1482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7054 a_8894_2696# d0 a_9385_2883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7055 a_13166_n8616# a_13168_n9134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7056 a_4662_n7679# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7057 a_2467_1901# d1 a_2562_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7058 a_26627_8397# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7059 a_644_2858# a_426_2858# a_153_2671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7060 a_24055_n5304# d1 a_24141_n4508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7061 a_5698_n8746# d2 a_5749_n7903# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7062 a_33012_6200# a_33269_6010# a_32966_7220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7063 a_12211_8437# a_12215_8260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7064 gnd d2 a_20201_8008# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7065 a_26430_n8721# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7066 a_9185_n3207# a_8967_n3207# a_8694_n3013# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7067 a_27434_3533# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7068 a_20807_6623# a_20824_7406# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7069 vdd d0 a_12451_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7070 a_30427_n2520# d0 a_30902_n2626# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7071 a_24411_8444# d0 a_25204_8849# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7072 a_8539_196# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7073 gnd d0 a_21008_3144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7074 a_6946_3519# d0 a_7748_3158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7075 vdd d1 a_24374_n3694# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7076 a_20767_4764# a_20771_4587# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7077 gnd d1 a_7166_1293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7078 gnd d0 a_34185_7666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7079 a_18088_6942# d1 a_18885_7170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7080 a_2175_n10565# a_4208_n10668# a_4050_n10652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7081 a_33012_6200# d1 a_33098_5415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7082 a_23456_271# d4 a_24049_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7083 gnd d3 a_19938_n8363# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7084 a_2459_n7537# d0 a_3252_n7953# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7085 a_18678_n3653# a_18476_n2814# a_18600_n2814# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7086 gnd d0 a_12161_n2492# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7087 a_9764_n3435# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7088 a_23321_2501# a_23103_2501# a_23227_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7089 a_29389_n8408# a_29384_n9008# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7090 a_18450_n6476# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7091 a_4807_3889# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7092 a_29492_3359# a_29749_3169# a_28694_3543# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7093 a_32058_n5902# a_31840_n5902# a_31955_n7940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7094 vdd d0 a_34093_2164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7095 vdd d0 a_12394_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7096 a_16575_8450# a_16832_8260# a_15777_8634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7097 vdd d0 a_25264_n9012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7098 a_10147_n3843# a_9929_n3843# a_10048_n3666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7099 a_13749_2896# d1 a_14546_3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7100 a_4863_6943# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7101 a_32036_6598# a_31834_5582# a_31958_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7102 a_9258_n7279# a_9040_n7279# a_8769_n7184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7103 a_30494_n6409# d0 a_30975_n6698# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7104 a_17443_n9425# d0 a_17924_n9714# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7105 a_15526_2959# d2 a_15605_4152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7106 a_72_n9413# d0 a_553_n9702# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7107 a_31798_3546# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7108 a_18594_3098# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7109 a_30721_n4662# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7110 a_13712_860# a_13494_860# a_13223_966# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7111 a_29565_7431# a_29822_7241# a_28767_7615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7112 a_22162_n2189# a_21944_n2189# a_21673_n2094# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7113 a_26538_n2613# d1 a_27336_n2662# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7114 vdd d0 a_21097_8646# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7115 a_11281_5998# d1 a_11376_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7116 a_11958_n5530# a_11962_n5342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7117 gnd d1 a_7023_n4700# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7118 vdd d1 a_2732_n8759# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7119 a_15507_n4709# d0 a_16309_n4337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7120 a_33642_n2725# a_33656_n3519# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7121 gnd d4 a_11132_n6342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7122 a_17389_n6371# a_17395_n6554# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7123 a_5080_7355# a_4862_7355# a_4605_7450# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7124 a_31871_7618# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7125 a_30992_n7716# d1 a_31778_n6924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7126 a_12178_6224# a_12431_6211# a_11376_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7127 a_21744_n6067# a_21746_n6166# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7128 a_24317_3531# d0 a_25115_3347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7129 gnd d1 a_15980_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7130 a_8939_5243# a_8945_5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7131 gnd d0 a_29728_2563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7132 a_25187_7831# a_25191_7654# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7133 a_3167_n2263# a_3162_n2863# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7134 a_26357_8091# d0 a_26846_7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7135 a_19509_n6125# d3 a_19681_n8347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7136 vdd d3 a_24409_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7137 a_3383_3557# a_3636_3544# a_2586_3329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7138 a_2622_5365# d0 a_3419_5593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7139 a_9241_n6261# a_9023_n6261# a_8752_n6166# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7140 a_8857_854# a_12084_1311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7141 a_10017_6165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7142 a_29549_6236# a_29544_6825# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7143 gnd d0 a_12287_n10030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7144 a_21734_n5366# d0 a_22215_n5655# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7145 a_33639_n2501# a_33643_n2313# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X7146 a_24374_6408# a_24627_6395# a_24275_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7147 a_27497_n7927# d3 a_27591_n7927# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7148 a_21790_n8420# d0 a_22271_n8709# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7149 a_11920_n3906# a_12177_n3922# a_11127_n3490# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7150 a_9147_1865# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7151 a_5773_1592# d2 a_5851_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7152 a_15708_4385# d0 a_16505_4613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7153 a_31156_4944# a_30938_4944# a_30667_5050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7154 a_31968_2645# a_31798_3546# a_31922_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7155 a_18087_7354# a_17869_7354# a_17606_7266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7156 a_734_7948# a_516_7948# a_245_8054# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7157 a_26364_8309# d0 a_26845_8397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7158 vdd d0 a_3420_n2467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7159 a_21920_4408# d0 a_22395_4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X7160 vdd d0 a_16635_n8613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7161 a_10054_8201# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
C0 d4 gnd 2.53fF
C1 a_23456_271# a_23461_390# 5.60fF
C2 a_18953_n5864# a_19447_n10577# 5.60fF
C3 d2 gnd 10.12fF
C4 a_10462_271# a_10467_390# 5.60fF
C5 a_14826_284# a_14831_403# 5.60fF
C6 a_23317_n5877# a_23811_n10590# 5.60fF
C7 d0 vdd 14.44fF
C8 a_6085_259# a_6090_378# 5.60fF
C9 d0 gnd 38.17fF
C10 a_27833_283# a_27838_402# 5.60fF
C11 a_1721_246# a_1726_365# 5.60fF
C12 d3 vdd 3.07fF
C13 a_32197_296# a_32202_415# 5.60fF
C14 a_32058_n5902# a_32552_n10615# 5.60fF
C15 a_27694_n5889# a_28188_n10602# 5.60fF
C16 d3 gnd 5.06fF
C17 a_5946_n5865# a_6440_n10578# 5.60fF
C18 vdd gnd 19.42fF
C19 a_10323_n5877# a_10817_n10590# 5.60fF
C20 a_19092_258# a_19097_377# 5.60fF
C21 d1 vdd 8.55fF
C22 d1 gnd 20.24fF
C23 a_2076_n10565# a_1582_n5852# 5.60fF
C24 a_14687_n5890# a_15181_n10603# 5.60fF
C25 d2 vdd 7.47fF
C26 gnd SUB 218.71fF
C27 vdd SUB 982.54fF
C28 a_30063_n10689# SUB 3.77fF
C29 d6 SUB 4.89fF
C30 d5 SUB 11.92fF
C31 a_28287_n10602# SUB 3.15fF
C32 a_25615_n10665# SUB 5.69fF
C33 d7 SUB 3.23fF
C34 a_21322_n10664# SUB 3.77fF
C35 a_21421_n10664# SUB 5.73fF
C36 a_17125_n10728# SUB 9.23fF
C37 a_19546_n10577# SUB 3.15fF
C38 a_12692_n10677# SUB 3.77fF
C39 a_10916_n10590# SUB 3.15fF
C40 a_8244_n10653# SUB 5.69fF
C41 a_8343_n10653# SUB 9.57fF
C42 a_3951_n10652# SUB 3.77fF
C43 a_4050_n10652# SUB 5.68fF
C44 a_2175_n10565# SUB 3.15fF
C45 a_30559_n9970# SUB 5.34fF
C46 d0 SUB 338.31fF
C47 a_26195_n9957# SUB 5.34fF
C48 a_21818_n9945# SUB 5.34fF
C49 a_32972_n9623# SUB 2.21fF
C50 d1 SUB 182.57fF
C51 a_32968_n9811# SUB 2.30fF
C52 a_17454_n9932# SUB 5.34fF
C53 a_13188_n9958# SUB 5.34fF
C54 a_28608_n9610# SUB 2.21fF
C55 a_31029_n9752# SUB 2.30fF
C56 a_28604_n9798# SUB 2.30fF
C57 a_24231_n9598# SUB 2.21fF
C58 a_8824_n9945# SUB 5.34fF
C59 a_26665_n9739# SUB 2.30fF
C60 a_24227_n9786# SUB 2.30fF
C61 a_19867_n9585# SUB 2.21fF
C62 d2 SUB 91.78fF
C63 a_31030_n9340# SUB 2.21fF
C64 a_22288_n9727# SUB 2.30fF
C65 a_19863_n9773# SUB 2.30fF
C66 a_4447_n9933# SUB 5.34fF
C67 a_15601_n9611# SUB 2.21fF
C68 a_15597_n9799# SUB 2.30fF
C69 a_83_n9920# SUB 5.34fF
C70 a_11237_n9598# SUB 2.21fF
C71 a_17924_n9714# SUB 2.30fF
C72 a_22289_n9315# SUB 2.21fF
C73 a_13658_n9740# SUB 2.30fF
C74 a_11233_n9786# SUB 2.30fF
C75 a_6860_n9586# SUB 2.21fF
C76 a_9294_n9727# SUB 2.30fF
C77 a_2496_n9573# SUB 2.21fF
C78 a_17925_n9302# SUB 2.21fF
C79 a_13659_n9328# SUB 2.21fF
C80 a_4917_n9715# SUB 2.30fF
C81 a_2492_n9761# SUB 2.30fF
C82 a_9295_n9315# SUB 2.21fF
C83 a_553_n9702# SUB 2.30fF
C84 a_554_n9290# SUB 2.21fF
C85 a_32955_n8605# SUB 2.21fF
C86 a_32951_n8793# SUB 2.30fF
C87 a_28591_n8592# SUB 2.21fF
C88 a_31012_n8734# SUB 2.30fF
C89 a_28587_n8780# SUB 2.30fF
C90 a_24214_n8580# SUB 2.21fF
C91 a_24210_n8768# SUB 2.30fF
C92 a_19850_n8567# SUB 2.21fF
C93 a_32790_n8197# SUB 2.37fF
C94 d3 SUB 45.68fF
C95 a_31013_n8322# SUB 2.21fF
C96 a_22271_n8709# SUB 2.30fF
C97 a_19846_n8755# SUB 2.30fF
C98 a_15584_n8593# SUB 2.21fF
C99 a_15580_n8781# SUB 2.30fF
C100 a_11220_n8580# SUB 2.21fF
C101 a_28426_n8184# SUB 2.37fF
C102 a_26649_n8309# SUB 2.21fF
C103 a_17907_n8696# SUB 2.30fF
C104 a_24049_n8172# SUB 2.37fF
C105 a_22272_n8297# SUB 2.21fF
C106 a_13641_n8722# SUB 2.30fF
C107 a_11216_n8768# SUB 2.30fF
C108 a_6843_n8568# SUB 2.21fF
C109 a_19685_n8159# SUB 2.37fF
C110 a_9277_n8709# SUB 2.30fF
C111 a_6839_n8756# SUB 2.30fF
C112 a_2479_n8555# SUB 2.21fF
C113 a_15419_n8185# SUB 2.37fF
C114 a_17908_n8284# SUB 2.21fF
C115 a_13642_n8310# SUB 2.21fF
C116 a_2475_n8743# SUB 2.30fF
C117 a_11055_n8172# SUB 2.37fF
C118 a_9278_n8297# SUB 2.21fF
C119 a_536_n8684# SUB 2.30fF
C120 a_6678_n8160# SUB 2.37fF
C121 a_2314_n8147# SUB 2.37fF
C122 a_537_n8272# SUB 2.21fF
C123 a_32935_n7587# SUB 2.21fF
C124 a_32931_n7775# SUB 2.30fF
C125 a_28571_n7574# SUB 2.21fF
C126 a_30992_n7716# SUB 2.30fF
C127 a_28567_n7762# SUB 2.30fF
C128 a_24194_n7562# SUB 2.21fF
C129 a_24190_n7750# SUB 2.30fF
C130 a_19830_n7549# SUB 2.21fF
C131 a_30993_n7304# SUB 2.21fF
C132 a_22251_n7691# SUB 2.30fF
C133 a_19826_n7737# SUB 2.30fF
C134 a_15564_n7575# SUB 2.21fF
C135 a_15560_n7763# SUB 2.30fF
C136 a_11200_n7562# SUB 2.21fF
C137 a_17887_n7678# SUB 2.30fF
C138 a_22252_n7279# SUB 2.21fF
C139 a_13621_n7704# SUB 2.30fF
C140 a_11196_n7750# SUB 2.30fF
C141 a_6823_n7550# SUB 2.21fF
C142 a_9257_n7691# SUB 2.30fF
C143 a_6819_n7738# SUB 2.30fF
C144 a_2459_n7537# SUB 2.21fF
C145 a_17888_n7266# SUB 2.21fF
C146 a_13622_n7292# SUB 2.21fF
C147 a_2455_n7725# SUB 2.30fF
C148 a_9258_n7279# SUB 2.21fF
C149 a_516_n7666# SUB 2.30fF
C150 a_517_n7254# SUB 2.21fF
C151 a_31856_n7763# SUB 2.63fF
C152 a_32918_n6569# SUB 2.21fF
C153 a_27492_n7750# SUB 2.63fF
C154 a_32914_n6757# SUB 2.30fF
C155 a_28554_n6556# SUB 2.21fF
C156 a_23115_n7738# SUB 2.63fF
C157 a_30975_n6698# SUB 2.30fF
C158 a_28550_n6744# SUB 2.30fF
C159 a_24177_n6544# SUB 2.21fF
C160 a_18751_n7725# SUB 2.63fF
C161 a_32552_n10615# SUB 5.00fF
C162 a_24173_n6732# SUB 2.30fF
C163 a_14485_n7751# SUB 2.63fF
C164 a_19813_n6531# SUB 2.21fF
C165 a_32614_n6163# SUB 4.04fF
C166 d4 SUB 22.85fF
C167 a_28188_n10602# SUB 5.00fF
C168 a_22234_n6673# SUB 2.30fF
C169 a_19809_n6719# SUB 2.30fF
C170 a_15547_n6557# SUB 2.21fF
C171 a_10121_n7738# SUB 2.63fF
C172 a_15543_n6745# SUB 2.30fF
C173 a_11183_n6544# SUB 2.21fF
C174 a_28250_n6150# SUB 4.04fF
C175 a_30976_n6286# SUB 2.21fF
C176 a_23811_n10590# SUB 5.00fF
C177 a_17870_n6660# SUB 2.30fF
C178 a_5744_n7726# SUB 2.63fF
C179 a_23873_n6138# SUB 4.04fF
C180 a_19447_n10577# SUB 5.00fF
C181 a_13604_n6686# SUB 2.30fF
C182 a_11179_n6732# SUB 2.30fF
C183 a_6806_n6532# SUB 2.21fF
C184 a_1380_n7713# SUB 2.63fF
C185 a_19509_n6125# SUB 4.04fF
C186 a_22235_n6261# SUB 2.21fF
C187 a_15181_n10603# SUB 5.00fF
C188 a_9240_n6673# SUB 2.30fF
C189 a_6802_n6720# SUB 2.30fF
C190 a_2442_n6519# SUB 2.21fF
C191 a_15243_n6151# SUB 4.04fF
C192 a_10817_n10590# SUB 5.00fF
C193 a_4863_n6661# SUB 2.30fF
C194 a_2438_n6707# SUB 2.30fF
C195 a_10879_n6138# SUB 4.04fF
C196 a_17871_n6248# SUB 2.21fF
C197 a_13605_n6274# SUB 2.21fF
C198 a_6440_n10578# SUB 5.00fF
C199 a_499_n6648# SUB 2.30fF
C200 a_6502_n6126# SUB 4.04fF
C201 a_9241_n6261# SUB 2.21fF
C202 a_2076_n10565# SUB 5.00fF
C203 a_2138_n6113# SUB 4.04fF
C204 a_4864_n6249# SUB 2.21fF
C205 a_500_n6236# SUB 2.21fF
C206 a_31955_n7940# SUB 2.94fF
C207 a_32058_n5902# SUB 5.75fF
C208 a_32899_n5551# SUB 2.21fF
C209 a_27591_n7927# SUB 2.94fF
C210 a_27694_n5889# SUB 5.75fF
C211 a_32895_n5739# SUB 2.30fF
C212 a_28535_n5538# SUB 2.21fF
C213 a_23214_n7915# SUB 2.94fF
C214 a_23317_n5877# SUB 5.75fF
C215 a_30956_n5680# SUB 2.30fF
C216 a_28531_n5726# SUB 2.30fF
C217 a_24158_n5526# SUB 2.21fF
C218 a_18850_n7902# SUB 2.94fF
C219 a_18953_n5864# SUB 5.75fF
C220 a_24154_n5714# SUB 2.30fF
C221 a_14584_n7928# SUB 2.94fF
C222 a_14687_n5890# SUB 5.75fF
C223 a_19794_n5513# SUB 2.21fF
C224 a_30957_n5268# SUB 2.21fF
C225 a_22215_n5655# SUB 2.30fF
C226 a_19790_n5701# SUB 2.30fF
C227 a_15528_n5539# SUB 2.21fF
C228 a_10220_n7915# SUB 2.94fF
C229 a_10323_n5877# SUB 5.75fF
C230 a_15524_n5727# SUB 2.30fF
C231 a_11164_n5526# SUB 2.21fF
C232 a_17851_n5642# SUB 2.30fF
C233 a_5843_n7903# SUB 2.94fF
C234 a_5946_n5865# SUB 5.75fF
C235 a_22216_n5243# SUB 2.21fF
C236 a_13585_n5668# SUB 2.30fF
C237 a_11160_n5714# SUB 2.30fF
C238 a_6787_n5514# SUB 2.21fF
C239 a_1479_n7890# SUB 2.94fF
C240 a_1582_n5852# SUB 5.75fF
C241 a_9221_n5655# SUB 2.30fF
C242 a_6783_n5702# SUB 2.30fF
C243 a_2423_n5501# SUB 2.21fF
C244 a_17852_n5230# SUB 2.21fF
C245 a_13586_n5256# SUB 2.21fF
C246 a_4844_n5643# SUB 2.30fF
C247 a_2419_n5689# SUB 2.30fF
C248 a_9222_n5243# SUB 2.21fF
C249 a_480_n5630# SUB 2.30fF
C250 a_4845_n5231# SUB 2.21fF
C251 a_481_n5218# SUB 2.21fF
C252 a_32882_n4533# SUB 2.21fF
C253 a_32878_n4721# SUB 2.30fF
C254 a_28518_n4520# SUB 2.21fF
C255 a_30939_n4662# SUB 2.30fF
C256 a_28514_n4708# SUB 2.30fF
C257 a_24141_n4508# SUB 2.21fF
C258 a_32610_n6351# SUB 2.94fF
C259 a_24137_n4696# SUB 2.30fF
C260 a_19777_n4495# SUB 2.21fF
C261 a_32717_n4125# SUB 2.63fF
C262 a_30940_n4250# SUB 2.21fF
C263 a_28246_n6338# SUB 2.94fF
C264 a_22198_n4637# SUB 2.30fF
C265 a_19773_n4683# SUB 2.30fF
C266 a_15511_n4521# SUB 2.21fF
C267 a_15507_n4709# SUB 2.30fF
C268 a_11147_n4508# SUB 2.21fF
C269 a_28353_n4112# SUB 2.63fF
C270 a_23869_n6326# SUB 2.94fF
C271 a_17834_n4624# SUB 2.30fF
C272 a_23976_n4100# SUB 2.63fF
C273 a_22199_n4225# SUB 2.21fF
C274 a_19505_n6313# SUB 2.94fF
C275 a_13568_n4650# SUB 2.30fF
C276 a_11143_n4696# SUB 2.30fF
C277 a_6770_n4496# SUB 2.21fF
C278 a_19612_n4087# SUB 2.63fF
C279 a_15239_n6339# SUB 2.94fF
C280 a_9204_n4637# SUB 2.30fF
C281 a_6766_n4684# SUB 2.30fF
C282 a_2406_n4483# SUB 2.21fF
C283 a_15346_n4113# SUB 2.63fF
C284 a_17835_n4212# SUB 2.21fF
C285 a_13569_n4238# SUB 2.21fF
C286 a_10875_n6326# SUB 2.94fF
C287 a_4827_n4625# SUB 2.30fF
C288 a_2402_n4671# SUB 2.30fF
C289 a_10982_n4100# SUB 2.63fF
C290 a_9205_n4225# SUB 2.21fF
C291 a_6498_n6314# SUB 2.94fF
C292 a_463_n4612# SUB 2.30fF
C293 a_6605_n4088# SUB 2.63fF
C294 a_4828_n4213# SUB 2.21fF
C295 a_2134_n6301# SUB 2.94fF
C296 a_2241_n4075# SUB 2.63fF
C297 a_464_n4200# SUB 2.21fF
C298 a_31882_n3868# SUB 4.03fF
C299 a_32862_n3515# SUB 2.21fF
C300 a_27518_n3855# SUB 4.03fF
C301 a_32858_n3703# SUB 2.30fF
C302 a_28498_n3502# SUB 2.21fF
C303 a_23141_n3843# SUB 4.03fF
C304 a_30919_n3644# SUB 2.30fF
C305 a_28494_n3690# SUB 2.30fF
C306 a_24121_n3490# SUB 2.21fF
C307 a_18777_n3830# SUB 4.03fF
C308 a_26555_n3631# SUB 2.30fF
C309 a_24117_n3678# SUB 2.30fF
C310 a_14511_n3856# SUB 4.03fF
C311 a_19757_n3477# SUB 2.21fF
C312 a_30920_n3232# SUB 2.21fF
C313 a_22178_n3619# SUB 2.30fF
C314 a_19753_n3665# SUB 2.30fF
C315 a_15491_n3503# SUB 2.21fF
C316 a_10147_n3843# SUB 4.03fF
C317 a_15487_n3691# SUB 2.30fF
C318 a_11127_n3490# SUB 2.21fF
C319 a_26556_n3219# SUB 2.21fF
C320 a_17814_n3606# SUB 2.30fF
C321 a_5770_n3831# SUB 4.03fF
C322 a_22179_n3207# SUB 2.21fF
C323 a_13548_n3632# SUB 2.30fF
C324 a_11123_n3678# SUB 2.30fF
C325 a_6750_n3478# SUB 2.21fF
C326 a_1406_n3818# SUB 4.03fF
C327 a_9184_n3619# SUB 2.30fF
C328 a_6746_n3666# SUB 2.30fF
C329 a_2386_n3465# SUB 2.21fF
C330 a_17815_n3194# SUB 2.21fF
C331 a_13549_n3220# SUB 2.21fF
C332 a_4807_n3607# SUB 2.30fF
C333 a_2382_n3653# SUB 2.30fF
C334 a_443_n3594# SUB 2.30fF
C335 a_4808_n3195# SUB 2.21fF
C336 a_444_n3182# SUB 2.21fF
C337 a_31783_n3691# SUB 2.37fF
C338 a_32845_n2497# SUB 2.21fF
C339 a_27419_n3678# SUB 2.37fF
C340 a_32841_n2685# SUB 2.30fF
C341 a_28481_n2484# SUB 2.21fF
C342 a_23042_n3666# SUB 2.37fF
C343 a_30902_n2626# SUB 2.30fF
C344 a_28477_n2672# SUB 2.30fF
C345 a_24104_n2472# SUB 2.21fF
C346 a_18678_n3653# SUB 2.37fF
C347 a_26538_n2613# SUB 2.30fF
C348 a_24100_n2660# SUB 2.30fF
C349 a_14412_n3679# SUB 2.37fF
C350 a_19740_n2459# SUB 2.21fF
C351 a_22161_n2601# SUB 2.30fF
C352 a_19736_n2647# SUB 2.30fF
C353 a_15474_n2485# SUB 2.21fF
C354 a_10048_n3666# SUB 2.37fF
C355 a_15470_n2673# SUB 2.30fF
C356 a_11110_n2472# SUB 2.21fF
C357 a_30903_n2214# SUB 2.21fF
C358 a_17797_n2588# SUB 2.30fF
C359 a_5671_n3654# SUB 2.37fF
C360 a_13531_n2614# SUB 2.30fF
C361 a_11106_n2660# SUB 2.30fF
C362 a_6733_n2460# SUB 2.21fF
C363 a_1307_n3641# SUB 2.37fF
C364 a_29984_n2069# SUB 2.31fF
C365 a_26539_n2201# SUB 2.21fF
C366 a_6729_n2648# SUB 2.30fF
C367 a_2369_n2447# SUB 2.21fF
C368 a_25607_n2057# SUB 2.54fF
C369 a_22162_n2189# SUB 2.21fF
C370 a_4790_n2589# SUB 2.30fF
C371 a_2365_n2635# SUB 2.30fF
C372 a_21243_n2044# SUB 2.31fF
C373 a_17798_n2176# SUB 2.21fF
C374 a_13532_n2202# SUB 2.21fF
C375 a_426_n2576# SUB 2.30fF
C376 a_12613_n2057# SUB 2.31fF
C377 a_16977_n2070# SUB 2.37fF
C378 a_8236_n2045# SUB 2.54fF
C379 a_4791_n2177# SUB 2.21fF
C380 a_3872_n2032# SUB 2.31fF
C381 a_427_n2164# SUB 2.21fF
C382 a_17212_n839# SUB 10.33fF
C383 a_30322_209# SUB 3.15fF
C384 a_27932_283# SUB 3.77fF
C385 a_21581_184# SUB 3.15fF
C386 a_21680_184# SUB 5.69fF
C387 a_17148_133# SUB 9.57fF
C388 a_17217_n720# SUB 2.02fF
C389 a_19191_258# SUB 3.77fF
C390 a_12951_197# SUB 3.15fF
C391 a_10561_271# SUB 3.77fF
C392 a_8658_196# SUB 5.73fF
C393 a_8757_196# SUB 9.23fF
C394 a_1820_246# SUB 3.77fF
C395 a_30592_879# SUB 5.34fF
C396 a_26228_866# SUB 5.34fF
C397 a_21851_854# SUB 5.34fF
C398 a_17487_841# SUB 5.34fF
C399 a_13221_867# SUB 5.34fF
C400 a_31083_872# SUB 2.21fF
C401 a_26719_859# SUB 2.21fF
C402 a_31082_1284# SUB 2.30fF
C403 a_22342_847# SUB 2.21fF
C404 a_8857_854# SUB 5.34fF
C405 a_4480_842# SUB 5.34fF
C406 a_116_829# SUB 5.34fF
C407 a_33021_1520# SUB 2.30fF
C408 a_26718_1271# SUB 2.30fF
C409 a_17978_834# SUB 2.21fF
C410 a_28657_1507# SUB 2.30fF
C411 a_22341_1259# SUB 2.30fF
C412 a_13712_860# SUB 2.21fF
C413 a_24280_1495# SUB 2.30fF
C414 a_17977_1246# SUB 2.30fF
C415 a_9348_847# SUB 2.21fF
C416 a_33025_1343# SUB 2.21fF
C417 a_19916_1482# SUB 2.30fF
C418 a_13711_1272# SUB 2.30fF
C419 a_4971_835# SUB 2.21fF
C420 a_28661_1330# SUB 2.21fF
C421 a_15650_1508# SUB 2.30fF
C422 a_9347_1259# SUB 2.30fF
C423 a_607_822# SUB 2.21fF
C424 a_24284_1318# SUB 2.21fF
C425 a_11286_1495# SUB 2.30fF
C426 a_19920_1305# SUB 2.21fF
C427 a_6909_1483# SUB 2.30fF
C428 a_606_1234# SUB 2.30fF
C429 a_15654_1331# SUB 2.21fF
C430 a_2545_1470# SUB 2.30fF
C431 a_11290_1318# SUB 2.21fF
C432 a_6913_1306# SUB 2.21fF
C433 a_2549_1293# SUB 2.21fF
C434 a_31100_1890# SUB 2.21fF
C435 a_26736_1877# SUB 2.21fF
C436 a_31099_2302# SUB 2.30fF
C437 a_22359_1865# SUB 2.21fF
C438 a_26735_2289# SUB 2.30fF
C439 a_17995_1852# SUB 2.21fF
C440 a_33038_2538# SUB 2.30fF
C441 a_22358_2277# SUB 2.30fF
C442 a_13729_1878# SUB 2.21fF
C443 a_28674_2525# SUB 2.30fF
C444 a_31963_2526# SUB 2.37fF
C445 a_17994_2264# SUB 2.30fF
C446 a_9365_1865# SUB 2.21fF
C447 a_24297_2513# SUB 2.30fF
C448 a_33042_2361# SUB 2.21fF
C449 a_27599_2513# SUB 2.37fF
C450 a_13728_2290# SUB 2.30fF
C451 a_19933_2500# SUB 2.30fF
C452 a_28678_2348# SUB 2.21fF
C453 a_23222_2501# SUB 2.37fF
C454 a_9364_2277# SUB 2.30fF
C455 a_624_1840# SUB 2.21fF
C456 a_15667_2526# SUB 2.30fF
C457 a_24301_2336# SUB 2.21fF
C458 a_18858_2488# SUB 2.37fF
C459 a_4987_2265# SUB 2.30fF
C460 a_11303_2513# SUB 2.30fF
C461 a_19937_2323# SUB 2.21fF
C462 a_14592_2514# SUB 2.37fF
C463 a_623_2252# SUB 2.30fF
C464 a_6926_2501# SUB 2.30fF
C465 a_15671_2349# SUB 2.21fF
C466 a_10228_2501# SUB 2.37fF
C467 a_2562_2488# SUB 2.30fF
C468 a_11307_2336# SUB 2.21fF
C469 a_5851_2489# SUB 2.37fF
C470 a_6930_2324# SUB 2.21fF
C471 a_1487_2476# SUB 2.37fF
C472 a_2566_2311# SUB 2.21fF
C473 a_31120_2908# SUB 2.21fF
C474 a_26756_2895# SUB 2.21fF
C475 a_31119_3320# SUB 2.30fF
C476 a_22379_2883# SUB 2.21fF
C477 a_33058_3556# SUB 2.30fF
C478 a_26755_3307# SUB 2.30fF
C479 a_18015_2870# SUB 2.21fF
C480 a_28694_3543# SUB 2.30fF
C481 a_13749_2896# SUB 2.21fF
C482 a_24317_3531# SUB 2.30fF
C483 a_18014_3282# SUB 2.30fF
C484 a_9385_2883# SUB 2.21fF
C485 a_33062_3379# SUB 2.21fF
C486 a_19953_3518# SUB 2.30fF
C487 a_13748_3308# SUB 2.30fF
C488 a_5008_2871# SUB 2.21fF
C489 a_28698_3366# SUB 2.21fF
C490 a_15687_3544# SUB 2.30fF
C491 a_9384_3295# SUB 2.30fF
C492 a_644_2858# SUB 2.21fF
C493 a_24321_3354# SUB 2.21fF
C494 a_11323_3531# SUB 2.30fF
C495 a_5007_3283# SUB 2.30fF
C496 a_19957_3341# SUB 2.21fF
C497 a_6946_3519# SUB 2.30fF
C498 a_643_3270# SUB 2.30fF
C499 a_15691_3367# SUB 2.21fF
C500 a_2582_3506# SUB 2.30fF
C501 a_11327_3354# SUB 2.21fF
C502 a_6950_3342# SUB 2.21fF
C503 a_2586_3329# SUB 2.21fF
C504 a_32897_2971# SUB 2.63fF
C505 a_28533_2958# SUB 2.63fF
C506 a_31137_3926# SUB 2.21fF
C507 a_24156_2946# SUB 2.63fF
C508 a_26773_3913# SUB 2.21fF
C509 a_19792_2933# SUB 2.63fF
C510 a_31136_4338# SUB 2.30fF
C511 a_15526_2959# SUB 2.63fF
C512 a_26772_4325# SUB 2.30fF
C513 a_18032_3888# SUB 2.21fF
C514 a_11162_2946# SUB 2.63fF
C515 a_33075_4574# SUB 2.30fF
C516 a_22395_4313# SUB 2.30fF
C517 a_13766_3914# SUB 2.21fF
C518 a_6785_2934# SUB 2.63fF
C519 a_28711_4561# SUB 2.30fF
C520 a_32062_2526# SUB 4.04fF
C521 a_32202_415# SUB 5.00fF
C522 a_18031_4300# SUB 2.30fF
C523 a_9402_3901# SUB 2.21fF
C524 a_2421_2921# SUB 2.63fF
C525 a_24334_4549# SUB 2.30fF
C526 a_33079_4397# SUB 2.21fF
C527 a_27698_2513# SUB 4.04fF
C528 a_27838_402# SUB 5.00fF
C529 a_19970_4536# SUB 2.30fF
C530 a_28715_4384# SUB 2.21fF
C531 a_23321_2501# SUB 4.04fF
C532 a_23461_390# SUB 5.00fF
C533 a_13765_4326# SUB 2.30fF
C534 a_5025_3889# SUB 2.21fF
C535 a_9401_4313# SUB 2.30fF
C536 a_661_3876# SUB 2.21fF
C537 a_15704_4562# SUB 2.30fF
C538 a_24338_4372# SUB 2.21fF
C539 a_18957_2488# SUB 4.04fF
C540 a_19097_377# SUB 5.00fF
C541 a_5024_4301# SUB 2.30fF
C542 a_11340_4549# SUB 2.30fF
C543 a_19974_4359# SUB 2.21fF
C544 a_14691_2514# SUB 4.04fF
C545 a_14831_403# SUB 5.00fF
C546 a_660_4288# SUB 2.30fF
C547 a_6963_4537# SUB 2.30fF
C548 a_15708_4385# SUB 2.21fF
C549 a_10327_2501# SUB 4.04fF
C550 a_10467_390# SUB 5.00fF
C551 a_2599_4524# SUB 2.30fF
C552 a_11344_4372# SUB 2.21fF
C553 a_5950_2489# SUB 4.04fF
C554 a_6090_378# SUB 5.00fF
C555 a_6967_4360# SUB 2.21fF
C556 a_1586_2476# SUB 4.04fF
C557 a_1726_365# SUB 5.00fF
C558 a_2603_4347# SUB 2.21fF
C559 a_32197_296# SUB 5.75fF
C560 a_32790_5186# SUB 2.94fF
C561 a_27833_283# SUB 5.75fF
C562 a_28426_5173# SUB 2.94fF
C563 a_31156_4944# SUB 2.21fF
C564 a_23456_271# SUB 5.75fF
C565 a_24049_5161# SUB 2.94fF
C566 a_26792_4931# SUB 2.21fF
C567 a_19092_258# SUB 5.75fF
C568 a_19685_5148# SUB 2.94fF
C569 a_31155_5356# SUB 2.30fF
C570 a_22415_4919# SUB 2.21fF
C571 a_14826_284# SUB 5.75fF
C572 a_15419_5174# SUB 2.94fF
C573 a_33094_5592# SUB 2.30fF
C574 a_26791_5343# SUB 2.30fF
C575 a_18051_4906# SUB 2.21fF
C576 a_10462_271# SUB 5.75fF
C577 a_11055_5161# SUB 2.94fF
C578 a_28730_5579# SUB 2.30fF
C579 a_13785_4932# SUB 2.21fF
C580 a_6085_259# SUB 5.75fF
C581 a_6678_5149# SUB 2.94fF
C582 a_24353_5567# SUB 2.30fF
C583 a_18050_5318# SUB 2.30fF
C584 a_9421_4919# SUB 2.21fF
C585 a_1721_246# SUB 5.75fF
C586 a_2314_5136# SUB 2.94fF
C587 a_33098_5415# SUB 2.21fF
C588 a_19989_5554# SUB 2.30fF
C589 a_13784_5344# SUB 2.30fF
C590 a_5044_4907# SUB 2.21fF
C591 a_28734_5402# SUB 2.21fF
C592 a_15723_5580# SUB 2.30fF
C593 a_9420_5331# SUB 2.30fF
C594 a_680_4894# SUB 2.21fF
C595 a_24357_5390# SUB 2.21fF
C596 a_11359_5567# SUB 2.30fF
C597 a_5043_5319# SUB 2.30fF
C598 a_19993_5377# SUB 2.21fF
C599 a_6982_5555# SUB 2.30fF
C600 a_15727_5403# SUB 2.21fF
C601 a_2618_5542# SUB 2.30fF
C602 a_11363_5390# SUB 2.21fF
C603 a_6986_5378# SUB 2.21fF
C604 a_2622_5365# SUB 2.21fF
C605 a_31173_5962# SUB 2.21fF
C606 a_26809_5949# SUB 2.21fF
C607 a_31172_6374# SUB 2.30fF
C608 a_26808_6361# SUB 2.30fF
C609 a_18068_5924# SUB 2.21fF
C610 a_33111_6610# SUB 2.30fF
C611 a_22431_6349# SUB 2.30fF
C612 a_13802_5950# SUB 2.21fF
C613 a_28747_6597# SUB 2.30fF
C614 a_32036_6598# SUB 2.63fF
C615 a_32135_6598# SUB 2.94fF
C616 a_18067_6336# SUB 2.30fF
C617 a_9438_5937# SUB 2.21fF
C618 a_24370_6585# SUB 2.30fF
C619 a_33115_6433# SUB 2.21fF
C620 a_27672_6585# SUB 2.63fF
C621 a_27771_6585# SUB 2.94fF
C622 a_13801_6362# SUB 2.30fF
C623 a_5061_5925# SUB 2.21fF
C624 a_20006_6572# SUB 2.30fF
C625 a_28751_6420# SUB 2.21fF
C626 a_23295_6573# SUB 2.63fF
C627 a_23394_6573# SUB 2.94fF
C628 a_9437_6349# SUB 2.30fF
C629 a_15740_6598# SUB 2.30fF
C630 a_24374_6408# SUB 2.21fF
C631 a_18931_6560# SUB 2.63fF
C632 a_19030_6560# SUB 2.94fF
C633 a_5060_6337# SUB 2.30fF
C634 a_11376_6585# SUB 2.30fF
C635 a_20010_6395# SUB 2.21fF
C636 a_14665_6586# SUB 2.63fF
C637 a_14764_6586# SUB 2.94fF
C638 a_6999_6573# SUB 2.30fF
C639 a_15744_6421# SUB 2.21fF
C640 a_10301_6573# SUB 2.63fF
C641 a_10400_6573# SUB 2.94fF
C642 a_2635_6560# SUB 2.30fF
C643 a_11380_6408# SUB 2.21fF
C644 a_5924_6561# SUB 2.63fF
C645 a_6023_6561# SUB 2.94fF
C646 a_7003_6396# SUB 2.21fF
C647 a_1560_6548# SUB 2.63fF
C648 a_1659_6548# SUB 2.94fF
C649 a_2639_6383# SUB 2.21fF
C650 a_32794_5009# SUB 4.03fF
C651 a_28430_4996# SUB 4.03fF
C652 a_31193_6980# SUB 2.21fF
C653 a_24053_4984# SUB 4.03fF
C654 a_26829_6967# SUB 2.21fF
C655 a_19689_4971# SUB 4.03fF
C656 a_31192_7392# SUB 2.30fF
C657 a_22452_6955# SUB 2.21fF
C658 a_15423_4997# SUB 4.03fF
C659 a_33131_7628# SUB 2.30fF
C660 a_26828_7379# SUB 2.30fF
C661 a_18088_6942# SUB 2.21fF
C662 a_11059_4984# SUB 4.03fF
C663 a_28767_7615# SUB 2.30fF
C664 a_13822_6968# SUB 2.21fF
C665 a_6682_4972# SUB 4.03fF
C666 a_24390_7603# SUB 2.30fF
C667 a_18087_7354# SUB 2.30fF
C668 a_9458_6955# SUB 2.21fF
C669 a_2318_4959# SUB 4.03fF
C670 a_33135_7451# SUB 2.21fF
C671 a_20026_7590# SUB 2.30fF
C672 a_13821_7380# SUB 2.30fF
C673 a_5081_6943# SUB 2.21fF
C674 a_28771_7438# SUB 2.21fF
C675 a_15760_7616# SUB 2.30fF
C676 a_9457_7367# SUB 2.30fF
C677 a_24394_7426# SUB 2.21fF
C678 a_11396_7603# SUB 2.30fF
C679 a_5080_7355# SUB 2.30fF
C680 a_20030_7413# SUB 2.21fF
C681 a_7019_7591# SUB 2.30fF
C682 a_15764_7439# SUB 2.21fF
C683 a_2655_7578# SUB 2.30fF
C684 a_11400_7426# SUB 2.21fF
C685 a_7023_7414# SUB 2.21fF
C686 a_2659_7401# SUB 2.21fF
C687 a_32970_7043# SUB 2.37fF
C688 a_28606_7030# SUB 2.37fF
C689 a_31210_7998# SUB 2.21fF
C690 a_24229_7018# SUB 2.37fF
C691 a_26846_7985# SUB 2.21fF
C692 a_19865_7005# SUB 2.37fF
C693 a_31209_8410# SUB 2.30fF
C694 a_15599_7031# SUB 2.37fF
C695 a_26845_8397# SUB 2.30fF
C696 a_18105_7960# SUB 2.21fF
C697 a_11235_7018# SUB 2.37fF
C698 a_22468_8385# SUB 2.30fF
C699 a_13839_7986# SUB 2.21fF
C700 a_6858_7006# SUB 2.37fF
C701 a_18104_8372# SUB 2.30fF
C702 a_9475_7973# SUB 2.21fF
C703 a_2494_6993# SUB 2.37fF
C704 a_33148_8646# SUB 2.30fF
C705 a_28784_8633# SUB 2.30fF
C706 a_24407_8621# SUB 2.30fF
C707 a_33949_8697# SUB 13.95fF
C708 a_33152_8469# SUB 2.21fF
C709 a_20043_8608# SUB 2.30fF
C710 a_13838_8398# SUB 2.30fF
C711 a_5098_7961# SUB 2.21fF
C712 a_9474_8385# SUB 2.30fF
C713 a_5097_8373# SUB 2.30fF
C714 a_733_8360# SUB 2.30fF
C715 a_29585_8684# SUB 2.31fF
C716 a_28788_8456# SUB 2.21fF
C717 a_15777_8634# SUB 2.30fF
C718 a_24411_8444# SUB 2.21fF
C719 a_11413_8621# SUB 2.30fF
C720 a_20844_8659# SUB 2.31fF
C721 a_20047_8431# SUB 2.21fF
C722 a_7036_8609# SUB 2.30fF
C723 a_16578_8685# SUB 2.37fF
C724 a_15781_8457# SUB 2.21fF
C725 a_2672_8596# SUB 2.30fF
C726 a_12214_8672# SUB 2.31fF
C727 a_11417_8444# SUB 2.21fF
C728 a_7837_8660# SUB 2.54fF
C729 a_7040_8432# SUB 2.21fF
C730 a_3473_8647# SUB 2.31fF
C731 a_2676_8419# SUB 2.21fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40ns 80ns)
Vd4 d4 0 pulse(0 1.8 0ns 0.1ns 0.1ns 80ns 160ns)
Vd5 d5 0 pulse(0 1.8 0ns 0.1ns 0.1ns 160ns 320ns)
Vd6 d6 0 pulse(0 1.8 0ns 0.1ns 0.1ns 320ns 640ns)
Vd7 d7 0 pulse(0 1.8 0ns 0.1ns 0.1ns 640ns 1280ns)
Vd8 d8 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1280ns 2560ns)
Vd9 d9 0 pulse(0 1.8 0ns 0.1ns 0.1ns 2560ns 5120ns)


.tran 10ns 5120ns
.control
run
plot V(vout) 
.endc
.end

magic
tech sky130A
timestamp 1616086429
<< nwell >>
rect 274 594 882 744
rect 1136 410 1744 560
rect 275 182 883 332
rect 1218 -198 1826 -48
rect 257 -424 865 -274
rect 1119 -608 1727 -458
rect 258 -836 866 -686
<< nmos >>
rect 338 493 388 535
rect 556 493 606 535
rect 764 493 814 535
rect 1200 309 1250 351
rect 1418 309 1468 351
rect 1626 309 1676 351
rect 339 81 389 123
rect 557 81 607 123
rect 765 81 815 123
rect 1282 -299 1332 -257
rect 1500 -299 1550 -257
rect 1708 -299 1758 -257
rect 321 -525 371 -483
rect 539 -525 589 -483
rect 747 -525 797 -483
rect 1183 -709 1233 -667
rect 1401 -709 1451 -667
rect 1609 -709 1659 -667
rect 322 -937 372 -895
rect 540 -937 590 -895
rect 748 -937 798 -895
<< pmos >>
rect 338 612 388 712
rect 556 612 606 712
rect 764 612 814 712
rect 1200 428 1250 528
rect 1418 428 1468 528
rect 1626 428 1676 528
rect 339 200 389 300
rect 557 200 607 300
rect 765 200 815 300
rect 1282 -180 1332 -80
rect 1500 -180 1550 -80
rect 1708 -180 1758 -80
rect 321 -406 371 -306
rect 539 -406 589 -306
rect 747 -406 797 -306
rect 1183 -590 1233 -490
rect 1401 -590 1451 -490
rect 1609 -590 1659 -490
rect 322 -818 372 -718
rect 540 -818 590 -718
rect 748 -818 798 -718
<< ndiff >>
rect 289 525 338 535
rect 289 505 300 525
rect 320 505 338 525
rect 289 493 338 505
rect 388 529 432 535
rect 388 509 403 529
rect 423 509 432 529
rect 388 493 432 509
rect 507 525 556 535
rect 507 505 518 525
rect 538 505 556 525
rect 507 493 556 505
rect 606 529 650 535
rect 606 509 621 529
rect 641 509 650 529
rect 606 493 650 509
rect 720 529 764 535
rect 720 509 729 529
rect 749 509 764 529
rect 720 493 764 509
rect 814 525 863 535
rect 814 505 832 525
rect 852 505 863 525
rect 814 493 863 505
rect 1151 341 1200 351
rect 1151 321 1162 341
rect 1182 321 1200 341
rect 1151 309 1200 321
rect 1250 345 1294 351
rect 1250 325 1265 345
rect 1285 325 1294 345
rect 1250 309 1294 325
rect 1369 341 1418 351
rect 1369 321 1380 341
rect 1400 321 1418 341
rect 1369 309 1418 321
rect 1468 345 1512 351
rect 1468 325 1483 345
rect 1503 325 1512 345
rect 1468 309 1512 325
rect 1582 345 1626 351
rect 1582 325 1591 345
rect 1611 325 1626 345
rect 1582 309 1626 325
rect 1676 341 1725 351
rect 1676 321 1694 341
rect 1714 321 1725 341
rect 1676 309 1725 321
rect 290 113 339 123
rect 290 93 301 113
rect 321 93 339 113
rect 290 81 339 93
rect 389 117 433 123
rect 389 97 404 117
rect 424 97 433 117
rect 389 81 433 97
rect 508 113 557 123
rect 508 93 519 113
rect 539 93 557 113
rect 508 81 557 93
rect 607 117 651 123
rect 607 97 622 117
rect 642 97 651 117
rect 607 81 651 97
rect 721 117 765 123
rect 721 97 730 117
rect 750 97 765 117
rect 721 81 765 97
rect 815 113 864 123
rect 815 93 833 113
rect 853 93 864 113
rect 815 81 864 93
rect 1233 -267 1282 -257
rect 1233 -287 1244 -267
rect 1264 -287 1282 -267
rect 1233 -299 1282 -287
rect 1332 -263 1376 -257
rect 1332 -283 1347 -263
rect 1367 -283 1376 -263
rect 1332 -299 1376 -283
rect 1451 -267 1500 -257
rect 1451 -287 1462 -267
rect 1482 -287 1500 -267
rect 1451 -299 1500 -287
rect 1550 -263 1594 -257
rect 1550 -283 1565 -263
rect 1585 -283 1594 -263
rect 1550 -299 1594 -283
rect 1664 -263 1708 -257
rect 1664 -283 1673 -263
rect 1693 -283 1708 -263
rect 1664 -299 1708 -283
rect 1758 -267 1807 -257
rect 1758 -287 1776 -267
rect 1796 -287 1807 -267
rect 1758 -299 1807 -287
rect 272 -493 321 -483
rect 272 -513 283 -493
rect 303 -513 321 -493
rect 272 -525 321 -513
rect 371 -489 415 -483
rect 371 -509 386 -489
rect 406 -509 415 -489
rect 371 -525 415 -509
rect 490 -493 539 -483
rect 490 -513 501 -493
rect 521 -513 539 -493
rect 490 -525 539 -513
rect 589 -489 633 -483
rect 589 -509 604 -489
rect 624 -509 633 -489
rect 589 -525 633 -509
rect 703 -489 747 -483
rect 703 -509 712 -489
rect 732 -509 747 -489
rect 703 -525 747 -509
rect 797 -493 846 -483
rect 797 -513 815 -493
rect 835 -513 846 -493
rect 797 -525 846 -513
rect 1134 -677 1183 -667
rect 1134 -697 1145 -677
rect 1165 -697 1183 -677
rect 1134 -709 1183 -697
rect 1233 -673 1277 -667
rect 1233 -693 1248 -673
rect 1268 -693 1277 -673
rect 1233 -709 1277 -693
rect 1352 -677 1401 -667
rect 1352 -697 1363 -677
rect 1383 -697 1401 -677
rect 1352 -709 1401 -697
rect 1451 -673 1495 -667
rect 1451 -693 1466 -673
rect 1486 -693 1495 -673
rect 1451 -709 1495 -693
rect 1565 -673 1609 -667
rect 1565 -693 1574 -673
rect 1594 -693 1609 -673
rect 1565 -709 1609 -693
rect 1659 -677 1708 -667
rect 1659 -697 1677 -677
rect 1697 -697 1708 -677
rect 1659 -709 1708 -697
rect 273 -905 322 -895
rect 273 -925 284 -905
rect 304 -925 322 -905
rect 273 -937 322 -925
rect 372 -901 416 -895
rect 372 -921 387 -901
rect 407 -921 416 -901
rect 372 -937 416 -921
rect 491 -905 540 -895
rect 491 -925 502 -905
rect 522 -925 540 -905
rect 491 -937 540 -925
rect 590 -901 634 -895
rect 590 -921 605 -901
rect 625 -921 634 -901
rect 590 -937 634 -921
rect 704 -901 748 -895
rect 704 -921 713 -901
rect 733 -921 748 -901
rect 704 -937 748 -921
rect 798 -905 847 -895
rect 798 -925 816 -905
rect 836 -925 847 -905
rect 798 -937 847 -925
<< pdiff >>
rect 294 674 338 712
rect 294 654 306 674
rect 326 654 338 674
rect 294 612 338 654
rect 388 674 430 712
rect 388 654 402 674
rect 422 654 430 674
rect 388 612 430 654
rect 512 674 556 712
rect 512 654 524 674
rect 544 654 556 674
rect 512 612 556 654
rect 606 674 648 712
rect 606 654 620 674
rect 640 654 648 674
rect 606 612 648 654
rect 722 674 764 712
rect 722 654 730 674
rect 750 654 764 674
rect 722 612 764 654
rect 814 681 859 712
rect 814 674 858 681
rect 814 654 826 674
rect 846 654 858 674
rect 814 612 858 654
rect 1156 490 1200 528
rect 1156 470 1168 490
rect 1188 470 1200 490
rect 1156 428 1200 470
rect 1250 490 1292 528
rect 1250 470 1264 490
rect 1284 470 1292 490
rect 1250 428 1292 470
rect 1374 490 1418 528
rect 1374 470 1386 490
rect 1406 470 1418 490
rect 1374 428 1418 470
rect 1468 490 1510 528
rect 1468 470 1482 490
rect 1502 470 1510 490
rect 1468 428 1510 470
rect 1584 490 1626 528
rect 1584 470 1592 490
rect 1612 470 1626 490
rect 1584 428 1626 470
rect 1676 497 1721 528
rect 1676 490 1720 497
rect 1676 470 1688 490
rect 1708 470 1720 490
rect 1676 428 1720 470
rect 295 262 339 300
rect 295 242 307 262
rect 327 242 339 262
rect 295 200 339 242
rect 389 262 431 300
rect 389 242 403 262
rect 423 242 431 262
rect 389 200 431 242
rect 513 262 557 300
rect 513 242 525 262
rect 545 242 557 262
rect 513 200 557 242
rect 607 262 649 300
rect 607 242 621 262
rect 641 242 649 262
rect 607 200 649 242
rect 723 262 765 300
rect 723 242 731 262
rect 751 242 765 262
rect 723 200 765 242
rect 815 269 860 300
rect 815 262 859 269
rect 815 242 827 262
rect 847 242 859 262
rect 815 200 859 242
rect 1238 -118 1282 -80
rect 1238 -138 1250 -118
rect 1270 -138 1282 -118
rect 1238 -180 1282 -138
rect 1332 -118 1374 -80
rect 1332 -138 1346 -118
rect 1366 -138 1374 -118
rect 1332 -180 1374 -138
rect 1456 -118 1500 -80
rect 1456 -138 1468 -118
rect 1488 -138 1500 -118
rect 1456 -180 1500 -138
rect 1550 -118 1592 -80
rect 1550 -138 1564 -118
rect 1584 -138 1592 -118
rect 1550 -180 1592 -138
rect 1666 -118 1708 -80
rect 1666 -138 1674 -118
rect 1694 -138 1708 -118
rect 1666 -180 1708 -138
rect 1758 -111 1803 -80
rect 1758 -118 1802 -111
rect 1758 -138 1770 -118
rect 1790 -138 1802 -118
rect 1758 -180 1802 -138
rect 277 -344 321 -306
rect 277 -364 289 -344
rect 309 -364 321 -344
rect 277 -406 321 -364
rect 371 -344 413 -306
rect 371 -364 385 -344
rect 405 -364 413 -344
rect 371 -406 413 -364
rect 495 -344 539 -306
rect 495 -364 507 -344
rect 527 -364 539 -344
rect 495 -406 539 -364
rect 589 -344 631 -306
rect 589 -364 603 -344
rect 623 -364 631 -344
rect 589 -406 631 -364
rect 705 -344 747 -306
rect 705 -364 713 -344
rect 733 -364 747 -344
rect 705 -406 747 -364
rect 797 -337 842 -306
rect 797 -344 841 -337
rect 797 -364 809 -344
rect 829 -364 841 -344
rect 797 -406 841 -364
rect 1139 -528 1183 -490
rect 1139 -548 1151 -528
rect 1171 -548 1183 -528
rect 1139 -590 1183 -548
rect 1233 -528 1275 -490
rect 1233 -548 1247 -528
rect 1267 -548 1275 -528
rect 1233 -590 1275 -548
rect 1357 -528 1401 -490
rect 1357 -548 1369 -528
rect 1389 -548 1401 -528
rect 1357 -590 1401 -548
rect 1451 -528 1493 -490
rect 1451 -548 1465 -528
rect 1485 -548 1493 -528
rect 1451 -590 1493 -548
rect 1567 -528 1609 -490
rect 1567 -548 1575 -528
rect 1595 -548 1609 -528
rect 1567 -590 1609 -548
rect 1659 -521 1704 -490
rect 1659 -528 1703 -521
rect 1659 -548 1671 -528
rect 1691 -548 1703 -528
rect 1659 -590 1703 -548
rect 278 -756 322 -718
rect 278 -776 290 -756
rect 310 -776 322 -756
rect 278 -818 322 -776
rect 372 -756 414 -718
rect 372 -776 386 -756
rect 406 -776 414 -756
rect 372 -818 414 -776
rect 496 -756 540 -718
rect 496 -776 508 -756
rect 528 -776 540 -756
rect 496 -818 540 -776
rect 590 -756 632 -718
rect 590 -776 604 -756
rect 624 -776 632 -756
rect 590 -818 632 -776
rect 706 -756 748 -718
rect 706 -776 714 -756
rect 734 -776 748 -756
rect 706 -818 748 -776
rect 798 -749 843 -718
rect 798 -756 842 -749
rect 798 -776 810 -756
rect 830 -776 842 -756
rect 798 -818 842 -776
<< ndiffc >>
rect 136 912 154 930
rect 134 813 152 831
rect 131 588 149 606
rect 129 489 147 507
rect 300 505 320 525
rect 403 509 423 529
rect 518 505 538 525
rect 621 509 641 529
rect 729 509 749 529
rect 832 505 852 525
rect 125 405 143 423
rect 123 306 141 324
rect 1162 321 1182 341
rect 1265 325 1285 345
rect 1380 321 1400 341
rect 1483 325 1503 345
rect 1591 325 1611 345
rect 1694 321 1714 341
rect 118 187 136 205
rect 116 88 134 106
rect 301 93 321 113
rect 404 97 424 117
rect 519 93 539 113
rect 622 97 642 117
rect 730 97 750 117
rect 833 93 853 113
rect 119 -106 137 -88
rect 117 -205 135 -187
rect 1244 -287 1264 -267
rect 1347 -283 1367 -263
rect 1462 -287 1482 -267
rect 1565 -283 1585 -263
rect 1673 -283 1693 -263
rect 1776 -287 1796 -267
rect 114 -430 132 -412
rect 112 -529 130 -511
rect 283 -513 303 -493
rect 386 -509 406 -489
rect 501 -513 521 -493
rect 604 -509 624 -489
rect 712 -509 732 -489
rect 815 -513 835 -493
rect 108 -613 126 -595
rect 106 -712 124 -694
rect 1145 -697 1165 -677
rect 1248 -693 1268 -673
rect 1363 -697 1383 -677
rect 1466 -693 1486 -673
rect 1574 -693 1594 -673
rect 1677 -697 1697 -677
rect 101 -831 119 -813
rect 99 -930 117 -912
rect 284 -925 304 -905
rect 387 -921 407 -901
rect 502 -925 522 -905
rect 605 -921 625 -901
rect 713 -921 733 -901
rect 816 -925 836 -905
<< pdiffc >>
rect 306 654 326 674
rect 402 654 422 674
rect 524 654 544 674
rect 620 654 640 674
rect 730 654 750 674
rect 826 654 846 674
rect 1168 470 1188 490
rect 1264 470 1284 490
rect 1386 470 1406 490
rect 1482 470 1502 490
rect 1592 470 1612 490
rect 1688 470 1708 490
rect 307 242 327 262
rect 403 242 423 262
rect 525 242 545 262
rect 621 242 641 262
rect 731 242 751 262
rect 827 242 847 262
rect 1250 -138 1270 -118
rect 1346 -138 1366 -118
rect 1468 -138 1488 -118
rect 1564 -138 1584 -118
rect 1674 -138 1694 -118
rect 1770 -138 1790 -118
rect 289 -364 309 -344
rect 385 -364 405 -344
rect 507 -364 527 -344
rect 603 -364 623 -344
rect 713 -364 733 -344
rect 809 -364 829 -344
rect 1151 -548 1171 -528
rect 1247 -548 1267 -528
rect 1369 -548 1389 -528
rect 1465 -548 1485 -528
rect 1575 -548 1595 -528
rect 1671 -548 1691 -528
rect 290 -776 310 -756
rect 386 -776 406 -756
rect 508 -776 528 -756
rect 604 -776 624 -756
rect 714 -776 734 -756
rect 810 -776 830 -756
<< poly >>
rect 338 712 388 725
rect 556 712 606 725
rect 764 712 814 725
rect 338 584 388 612
rect 338 564 351 584
rect 371 564 388 584
rect 338 535 388 564
rect 556 587 606 612
rect 556 567 569 587
rect 589 567 606 587
rect 556 535 606 567
rect 764 585 814 612
rect 764 565 787 585
rect 807 565 814 585
rect 764 535 814 565
rect 1200 528 1250 541
rect 1418 528 1468 541
rect 1626 528 1676 541
rect 338 477 388 493
rect 556 477 606 493
rect 764 477 814 493
rect 1200 400 1250 428
rect 1200 380 1213 400
rect 1233 380 1250 400
rect 1200 351 1250 380
rect 1418 403 1468 428
rect 1418 383 1431 403
rect 1451 383 1468 403
rect 1418 351 1468 383
rect 1626 401 1676 428
rect 1626 381 1649 401
rect 1669 381 1676 401
rect 1626 351 1676 381
rect 339 300 389 313
rect 557 300 607 313
rect 765 300 815 313
rect 1200 293 1250 309
rect 1418 293 1468 309
rect 1626 293 1676 309
rect 339 172 389 200
rect 339 152 352 172
rect 372 152 389 172
rect 339 123 389 152
rect 557 175 607 200
rect 557 155 570 175
rect 590 155 607 175
rect 557 123 607 155
rect 765 173 815 200
rect 765 153 788 173
rect 808 153 815 173
rect 765 123 815 153
rect 339 65 389 81
rect 557 65 607 81
rect 765 65 815 81
rect 1282 -80 1332 -67
rect 1500 -80 1550 -67
rect 1708 -80 1758 -67
rect 1282 -208 1332 -180
rect 1282 -228 1295 -208
rect 1315 -228 1332 -208
rect 1282 -257 1332 -228
rect 1500 -205 1550 -180
rect 1500 -225 1513 -205
rect 1533 -225 1550 -205
rect 1500 -257 1550 -225
rect 1708 -207 1758 -180
rect 1708 -227 1731 -207
rect 1751 -227 1758 -207
rect 1708 -257 1758 -227
rect 321 -306 371 -293
rect 539 -306 589 -293
rect 747 -306 797 -293
rect 1282 -315 1332 -299
rect 1500 -315 1550 -299
rect 1708 -315 1758 -299
rect 321 -434 371 -406
rect 321 -454 334 -434
rect 354 -454 371 -434
rect 321 -483 371 -454
rect 539 -431 589 -406
rect 539 -451 552 -431
rect 572 -451 589 -431
rect 539 -483 589 -451
rect 747 -433 797 -406
rect 747 -453 770 -433
rect 790 -453 797 -433
rect 747 -483 797 -453
rect 1183 -490 1233 -477
rect 1401 -490 1451 -477
rect 1609 -490 1659 -477
rect 321 -541 371 -525
rect 539 -541 589 -525
rect 747 -541 797 -525
rect 1183 -618 1233 -590
rect 1183 -638 1196 -618
rect 1216 -638 1233 -618
rect 1183 -667 1233 -638
rect 1401 -615 1451 -590
rect 1401 -635 1414 -615
rect 1434 -635 1451 -615
rect 1401 -667 1451 -635
rect 1609 -617 1659 -590
rect 1609 -637 1632 -617
rect 1652 -637 1659 -617
rect 1609 -667 1659 -637
rect 322 -718 372 -705
rect 540 -718 590 -705
rect 748 -718 798 -705
rect 1183 -725 1233 -709
rect 1401 -725 1451 -709
rect 1609 -725 1659 -709
rect 322 -846 372 -818
rect 322 -866 335 -846
rect 355 -866 372 -846
rect 322 -895 372 -866
rect 540 -843 590 -818
rect 540 -863 553 -843
rect 573 -863 590 -843
rect 540 -895 590 -863
rect 748 -845 798 -818
rect 748 -865 771 -845
rect 791 -865 798 -845
rect 748 -895 798 -865
rect 322 -953 372 -937
rect 540 -953 590 -937
rect 748 -953 798 -937
<< polycont >>
rect 351 564 371 584
rect 569 567 589 587
rect 787 565 807 585
rect 1213 380 1233 400
rect 1431 383 1451 403
rect 1649 381 1669 401
rect 352 152 372 172
rect 570 155 590 175
rect 788 153 808 173
rect 1295 -228 1315 -208
rect 1513 -225 1533 -205
rect 1731 -227 1751 -207
rect 334 -454 354 -434
rect 552 -451 572 -431
rect 770 -453 790 -433
rect 1196 -638 1216 -618
rect 1414 -635 1434 -615
rect 1632 -637 1652 -617
rect 335 -866 355 -846
rect 553 -863 573 -843
rect 771 -865 791 -845
<< ndiffres >>
rect 113 934 174 950
rect 18 930 174 934
rect 18 912 136 930
rect 154 912 174 930
rect 18 891 174 912
rect 18 890 118 891
rect 19 854 61 890
rect 19 831 170 854
rect 19 816 134 831
rect 113 813 134 816
rect 152 813 170 831
rect 113 794 170 813
rect 108 610 169 626
rect 13 606 169 610
rect 13 588 131 606
rect 149 588 169 606
rect 13 567 169 588
rect 13 566 113 567
rect 14 530 56 566
rect 14 507 165 530
rect 14 492 129 507
rect 108 489 129 492
rect 147 489 165 507
rect 108 470 165 489
rect 102 427 163 443
rect 7 423 163 427
rect 7 405 125 423
rect 143 405 163 423
rect 7 384 163 405
rect 7 383 107 384
rect 8 347 50 383
rect 8 324 159 347
rect 8 309 123 324
rect 102 306 123 309
rect 141 306 159 324
rect 102 287 159 306
rect 95 209 156 225
rect 0 205 156 209
rect 0 187 118 205
rect 136 187 156 205
rect 0 166 156 187
rect 0 165 100 166
rect 1 129 43 165
rect 1 106 152 129
rect 1 91 116 106
rect 95 88 116 91
rect 134 88 152 106
rect 95 69 152 88
rect 96 -84 157 -68
rect 1 -88 157 -84
rect 1 -106 119 -88
rect 137 -106 157 -88
rect 1 -127 157 -106
rect 1 -128 101 -127
rect 2 -164 44 -128
rect 2 -187 153 -164
rect 2 -202 117 -187
rect 96 -205 117 -202
rect 135 -205 153 -187
rect 96 -224 153 -205
rect 91 -408 152 -392
rect -4 -412 152 -408
rect -4 -430 114 -412
rect 132 -430 152 -412
rect -4 -451 152 -430
rect -4 -452 96 -451
rect -3 -488 39 -452
rect -3 -511 148 -488
rect -3 -526 112 -511
rect 91 -529 112 -526
rect 130 -529 148 -511
rect 91 -548 148 -529
rect 85 -591 146 -575
rect -10 -595 146 -591
rect -10 -613 108 -595
rect 126 -613 146 -595
rect -10 -634 146 -613
rect -10 -635 90 -634
rect -9 -671 33 -635
rect -9 -694 142 -671
rect -9 -709 106 -694
rect 85 -712 106 -709
rect 124 -712 142 -694
rect 85 -731 142 -712
rect 78 -809 139 -793
rect -17 -813 139 -809
rect -17 -831 101 -813
rect 119 -831 139 -813
rect -17 -852 139 -831
rect -17 -853 83 -852
rect -16 -889 26 -853
rect -16 -912 135 -889
rect -16 -927 99 -912
rect 78 -930 99 -927
rect 117 -930 135 -912
rect 78 -949 135 -930
<< locali >>
rect 126 930 173 1046
rect 126 912 136 930
rect 154 912 173 930
rect 126 908 173 912
rect 127 903 164 908
rect 115 841 167 843
rect 113 837 546 841
rect 113 831 552 837
rect 113 813 134 831
rect 152 813 552 831
rect 113 795 552 813
rect 115 606 167 795
rect 513 770 552 795
rect 297 745 484 769
rect 513 750 908 770
rect 928 750 931 770
rect 513 745 931 750
rect 297 674 334 745
rect 513 744 856 745
rect 513 741 552 744
rect 818 743 855 744
rect 449 684 480 685
rect 297 654 306 674
rect 326 654 334 674
rect 297 644 334 654
rect 393 674 480 684
rect 393 654 402 674
rect 422 654 480 674
rect 393 645 480 654
rect 393 644 430 645
rect 115 588 131 606
rect 149 588 167 606
rect 449 594 480 645
rect 515 674 552 741
rect 667 684 703 685
rect 515 654 524 674
rect 544 654 552 674
rect 515 644 552 654
rect 611 674 759 684
rect 859 681 955 683
rect 611 654 620 674
rect 640 654 730 674
rect 750 654 759 674
rect 611 645 759 654
rect 817 674 955 681
rect 817 654 826 674
rect 846 654 955 674
rect 817 645 955 654
rect 611 644 648 645
rect 341 591 382 592
rect 115 570 167 588
rect 233 584 382 591
rect 233 564 292 584
rect 312 564 351 584
rect 371 564 382 584
rect 233 556 382 564
rect 449 587 606 594
rect 449 567 569 587
rect 589 567 606 587
rect 449 557 606 567
rect 449 556 484 557
rect 449 535 480 556
rect 667 535 703 645
rect 722 644 759 645
rect 818 644 855 645
rect 778 585 868 591
rect 778 565 787 585
rect 807 583 868 585
rect 807 565 832 583
rect 778 563 832 565
rect 852 563 868 583
rect 778 557 868 563
rect 292 534 329 535
rect 291 525 329 534
rect 119 507 159 517
rect 119 489 129 507
rect 147 489 159 507
rect 291 505 300 525
rect 320 505 329 525
rect 291 497 329 505
rect 395 529 480 535
rect 510 534 547 535
rect 395 509 403 529
rect 423 509 480 529
rect 395 501 480 509
rect 509 525 547 534
rect 509 505 518 525
rect 538 505 547 525
rect 395 500 431 501
rect 509 497 547 505
rect 613 529 757 535
rect 613 509 621 529
rect 641 509 674 529
rect 694 509 729 529
rect 749 509 757 529
rect 613 501 757 509
rect 613 500 649 501
rect 721 500 757 501
rect 823 534 860 535
rect 823 533 861 534
rect 823 525 887 533
rect 823 505 832 525
rect 852 511 887 525
rect 907 511 910 531
rect 852 506 910 511
rect 852 505 887 506
rect 119 433 159 489
rect 292 468 329 497
rect 293 466 329 468
rect 293 444 484 466
rect 510 465 547 497
rect 823 493 887 505
rect 927 467 954 645
rect 786 465 954 467
rect 510 455 954 465
rect 1159 561 1346 585
rect 1377 566 1770 586
rect 1790 566 1793 586
rect 1377 561 1793 566
rect 1159 490 1196 561
rect 1377 560 1718 561
rect 1311 500 1342 501
rect 1159 470 1168 490
rect 1188 470 1196 490
rect 1159 460 1196 470
rect 1255 490 1342 500
rect 1255 470 1264 490
rect 1284 470 1342 490
rect 1255 461 1342 470
rect 1255 460 1292 461
rect 116 428 159 433
rect 507 439 954 455
rect 507 433 535 439
rect 786 438 954 439
rect 116 425 266 428
rect 507 425 534 433
rect 116 423 534 425
rect 116 405 125 423
rect 143 405 534 423
rect 1311 410 1342 461
rect 1377 490 1414 560
rect 1680 559 1717 560
rect 1529 500 1565 501
rect 1377 470 1386 490
rect 1406 470 1414 490
rect 1377 460 1414 470
rect 1473 490 1621 500
rect 1721 497 1817 499
rect 1473 470 1482 490
rect 1502 470 1592 490
rect 1612 470 1621 490
rect 1473 461 1621 470
rect 1679 490 1817 497
rect 1679 470 1688 490
rect 1708 470 1817 490
rect 1679 461 1817 470
rect 1473 460 1510 461
rect 1203 407 1244 408
rect 116 402 534 405
rect 116 396 159 402
rect 119 393 159 396
rect 1095 400 1244 407
rect 516 384 556 385
rect 227 367 556 384
rect 1095 380 1154 400
rect 1174 380 1213 400
rect 1233 380 1244 400
rect 1095 372 1244 380
rect 1311 403 1468 410
rect 1311 383 1431 403
rect 1451 383 1468 403
rect 1311 373 1468 383
rect 1311 372 1346 373
rect 111 324 154 335
rect 111 306 123 324
rect 141 306 154 324
rect 111 280 154 306
rect 227 280 254 367
rect 516 358 556 367
rect 111 259 254 280
rect 298 332 332 348
rect 516 338 909 358
rect 929 338 932 358
rect 1311 351 1342 372
rect 1529 351 1565 461
rect 1584 460 1621 461
rect 1680 460 1717 461
rect 1640 401 1730 407
rect 1640 381 1649 401
rect 1669 399 1730 401
rect 1669 381 1694 399
rect 1640 379 1694 381
rect 1714 379 1730 399
rect 1640 373 1730 379
rect 1154 350 1191 351
rect 516 333 932 338
rect 1153 341 1191 350
rect 516 332 857 333
rect 298 262 335 332
rect 450 272 481 273
rect 111 257 248 259
rect 111 215 154 257
rect 298 242 307 262
rect 327 242 335 262
rect 298 232 335 242
rect 394 262 481 272
rect 394 242 403 262
rect 423 242 481 262
rect 394 233 481 242
rect 394 232 431 233
rect 109 205 154 215
rect 109 187 118 205
rect 136 187 154 205
rect 109 181 154 187
rect 450 182 481 233
rect 516 262 553 332
rect 819 331 856 332
rect 1153 321 1162 341
rect 1182 321 1191 341
rect 1153 313 1191 321
rect 1257 345 1342 351
rect 1372 350 1409 351
rect 1257 325 1265 345
rect 1285 325 1342 345
rect 1257 317 1342 325
rect 1371 341 1409 350
rect 1371 321 1380 341
rect 1400 321 1409 341
rect 1257 316 1293 317
rect 1371 313 1409 321
rect 1475 345 1619 351
rect 1475 325 1483 345
rect 1503 326 1535 345
rect 1556 326 1591 345
rect 1503 325 1591 326
rect 1611 325 1619 345
rect 1475 317 1619 325
rect 1475 316 1511 317
rect 1583 316 1619 317
rect 1685 350 1722 351
rect 1685 349 1723 350
rect 1685 341 1749 349
rect 1685 321 1694 341
rect 1714 327 1749 341
rect 1769 327 1772 347
rect 1714 322 1772 327
rect 1714 321 1749 322
rect 1154 284 1191 313
rect 1155 282 1191 284
rect 668 272 704 273
rect 516 242 525 262
rect 545 242 553 262
rect 516 232 553 242
rect 612 262 760 272
rect 860 269 956 271
rect 612 242 621 262
rect 641 242 731 262
rect 751 242 760 262
rect 612 233 760 242
rect 818 262 956 269
rect 818 242 827 262
rect 847 242 956 262
rect 1155 260 1346 282
rect 1372 281 1409 313
rect 1685 309 1749 321
rect 1789 283 1816 461
rect 1648 281 1816 283
rect 1372 255 1816 281
rect 818 233 956 242
rect 612 232 649 233
rect 109 178 146 181
rect 342 179 383 180
rect 234 172 383 179
rect 234 152 293 172
rect 313 152 352 172
rect 372 152 383 172
rect 234 144 383 152
rect 450 175 607 182
rect 450 155 570 175
rect 590 155 607 175
rect 450 145 607 155
rect 450 144 485 145
rect 450 123 481 144
rect 668 123 704 233
rect 723 232 760 233
rect 819 232 856 233
rect 779 173 869 179
rect 779 153 788 173
rect 808 171 869 173
rect 808 153 833 171
rect 779 151 833 153
rect 853 151 869 171
rect 779 145 869 151
rect 293 122 330 123
rect 106 114 143 116
rect 106 106 148 114
rect 106 88 116 106
rect 134 88 148 106
rect 106 79 148 88
rect 292 113 330 122
rect 292 93 301 113
rect 321 93 330 113
rect 292 85 330 93
rect 396 117 481 123
rect 511 122 548 123
rect 396 97 404 117
rect 424 97 481 117
rect 396 89 481 97
rect 510 113 548 122
rect 510 93 519 113
rect 539 93 548 113
rect 396 88 432 89
rect 510 85 548 93
rect 614 121 758 123
rect 614 117 666 121
rect 614 97 622 117
rect 642 101 666 117
rect 686 117 758 121
rect 686 101 730 117
rect 642 97 730 101
rect 750 97 758 117
rect 614 89 758 97
rect 614 88 650 89
rect 722 88 758 89
rect 824 122 861 123
rect 824 121 862 122
rect 824 113 888 121
rect 824 93 833 113
rect 853 99 888 113
rect 908 99 911 119
rect 853 94 911 99
rect 853 93 888 94
rect 107 54 148 79
rect 293 54 330 85
rect 511 54 548 85
rect 824 81 888 93
rect 928 55 955 233
rect 107 27 156 54
rect 292 28 341 54
rect 510 53 591 54
rect 787 53 955 55
rect 510 28 955 53
rect 511 27 955 28
rect 109 -6 156 27
rect 512 -6 552 27
rect 787 26 955 27
rect 1482 31 1522 255
rect 1648 254 1816 255
rect 1482 9 1490 31
rect 1514 9 1522 31
rect 1482 1 1522 9
rect 109 -45 552 -6
rect 109 -88 156 -45
rect 512 -50 552 -45
rect 1241 -47 1428 -23
rect 1459 -42 1852 -22
rect 1872 -42 1875 -22
rect 1459 -47 1875 -42
rect 109 -106 119 -88
rect 137 -106 156 -88
rect 109 -110 156 -106
rect 110 -115 147 -110
rect 1241 -118 1278 -47
rect 1459 -48 1800 -47
rect 1393 -108 1424 -107
rect 1241 -138 1250 -118
rect 1270 -138 1278 -118
rect 1241 -148 1278 -138
rect 1337 -118 1424 -108
rect 1337 -138 1346 -118
rect 1366 -138 1424 -118
rect 1337 -147 1424 -138
rect 1337 -148 1374 -147
rect 98 -177 150 -175
rect 96 -181 529 -177
rect 96 -187 535 -181
rect 96 -205 117 -187
rect 135 -205 535 -187
rect 1393 -198 1424 -147
rect 1459 -118 1496 -48
rect 1762 -49 1799 -48
rect 1611 -108 1647 -107
rect 1459 -138 1468 -118
rect 1488 -138 1496 -118
rect 1459 -148 1496 -138
rect 1555 -118 1703 -108
rect 1803 -111 1899 -109
rect 1555 -138 1564 -118
rect 1584 -138 1674 -118
rect 1694 -138 1703 -118
rect 1555 -147 1703 -138
rect 1761 -118 1899 -111
rect 1761 -138 1770 -118
rect 1790 -138 1899 -118
rect 1761 -147 1899 -138
rect 1555 -148 1592 -147
rect 1285 -201 1326 -200
rect 96 -223 535 -205
rect 98 -412 150 -223
rect 496 -248 535 -223
rect 1177 -208 1326 -201
rect 1177 -228 1236 -208
rect 1256 -228 1295 -208
rect 1315 -228 1326 -208
rect 1177 -236 1326 -228
rect 1393 -205 1550 -198
rect 1393 -225 1513 -205
rect 1533 -225 1550 -205
rect 1393 -235 1550 -225
rect 1393 -236 1428 -235
rect 280 -273 467 -249
rect 496 -268 891 -248
rect 911 -268 914 -248
rect 1393 -257 1424 -236
rect 1611 -257 1647 -147
rect 1666 -148 1703 -147
rect 1762 -148 1799 -147
rect 1722 -207 1812 -201
rect 1722 -227 1731 -207
rect 1751 -209 1812 -207
rect 1751 -227 1776 -209
rect 1722 -229 1776 -227
rect 1796 -229 1812 -209
rect 1722 -235 1812 -229
rect 1236 -258 1273 -257
rect 496 -273 914 -268
rect 1235 -267 1273 -258
rect 280 -344 317 -273
rect 496 -274 839 -273
rect 496 -277 535 -274
rect 801 -275 838 -274
rect 432 -334 463 -333
rect 280 -364 289 -344
rect 309 -364 317 -344
rect 280 -374 317 -364
rect 376 -344 463 -334
rect 376 -364 385 -344
rect 405 -364 463 -344
rect 376 -373 463 -364
rect 376 -374 413 -373
rect 98 -430 114 -412
rect 132 -430 150 -412
rect 432 -424 463 -373
rect 498 -344 535 -277
rect 1235 -287 1244 -267
rect 1264 -287 1273 -267
rect 1235 -295 1273 -287
rect 1339 -263 1424 -257
rect 1454 -258 1491 -257
rect 1339 -283 1347 -263
rect 1367 -283 1424 -263
rect 1339 -291 1424 -283
rect 1453 -267 1491 -258
rect 1453 -287 1462 -267
rect 1482 -287 1491 -267
rect 1339 -292 1375 -291
rect 1453 -295 1491 -287
rect 1557 -263 1701 -257
rect 1557 -283 1565 -263
rect 1585 -283 1673 -263
rect 1693 -283 1701 -263
rect 1557 -291 1701 -283
rect 1557 -292 1593 -291
rect 1665 -292 1701 -291
rect 1767 -258 1804 -257
rect 1767 -259 1805 -258
rect 1767 -267 1831 -259
rect 1767 -287 1776 -267
rect 1796 -281 1831 -267
rect 1851 -281 1854 -261
rect 1796 -286 1854 -281
rect 1796 -287 1831 -286
rect 1236 -324 1273 -295
rect 1237 -326 1273 -324
rect 650 -334 686 -333
rect 498 -364 507 -344
rect 527 -364 535 -344
rect 498 -374 535 -364
rect 594 -344 742 -334
rect 842 -337 938 -335
rect 594 -364 603 -344
rect 623 -364 713 -344
rect 733 -364 742 -344
rect 594 -373 742 -364
rect 800 -344 938 -337
rect 800 -364 809 -344
rect 829 -364 938 -344
rect 1237 -348 1428 -326
rect 1454 -327 1491 -295
rect 1767 -299 1831 -287
rect 1871 -325 1898 -147
rect 1730 -327 1898 -325
rect 1454 -341 1898 -327
rect 1454 -353 1901 -341
rect 1497 -355 1530 -353
rect 800 -373 938 -364
rect 594 -374 631 -373
rect 324 -427 365 -426
rect 98 -448 150 -430
rect 216 -434 365 -427
rect 216 -454 275 -434
rect 295 -454 334 -434
rect 354 -454 365 -434
rect 216 -462 365 -454
rect 432 -431 589 -424
rect 432 -451 552 -431
rect 572 -451 589 -431
rect 432 -461 589 -451
rect 432 -462 467 -461
rect 432 -483 463 -462
rect 650 -483 686 -373
rect 705 -374 742 -373
rect 801 -374 838 -373
rect 761 -433 851 -427
rect 761 -453 770 -433
rect 790 -435 851 -433
rect 790 -453 815 -435
rect 761 -455 815 -453
rect 835 -455 851 -435
rect 761 -461 851 -455
rect 275 -484 312 -483
rect 274 -493 312 -484
rect 102 -511 142 -501
rect 102 -529 112 -511
rect 130 -529 142 -511
rect 274 -513 283 -493
rect 303 -513 312 -493
rect 274 -521 312 -513
rect 378 -489 463 -483
rect 493 -484 530 -483
rect 378 -509 386 -489
rect 406 -509 463 -489
rect 378 -517 463 -509
rect 492 -493 530 -484
rect 492 -513 501 -493
rect 521 -513 530 -493
rect 378 -518 414 -517
rect 492 -521 530 -513
rect 596 -489 740 -483
rect 596 -509 604 -489
rect 624 -509 657 -489
rect 677 -509 712 -489
rect 732 -509 740 -489
rect 596 -517 740 -509
rect 596 -518 632 -517
rect 704 -518 740 -517
rect 806 -484 843 -483
rect 806 -485 844 -484
rect 806 -493 870 -485
rect 806 -513 815 -493
rect 835 -507 870 -493
rect 890 -507 893 -487
rect 835 -512 893 -507
rect 835 -513 870 -512
rect 102 -585 142 -529
rect 275 -550 312 -521
rect 276 -552 312 -550
rect 276 -574 467 -552
rect 493 -553 530 -521
rect 806 -525 870 -513
rect 910 -551 937 -373
rect 1859 -398 1901 -353
rect 769 -553 937 -551
rect 493 -563 937 -553
rect 1142 -457 1329 -433
rect 1360 -452 1753 -432
rect 1773 -452 1776 -432
rect 1360 -457 1776 -452
rect 1142 -528 1179 -457
rect 1360 -458 1701 -457
rect 1294 -518 1325 -517
rect 1142 -548 1151 -528
rect 1171 -548 1179 -528
rect 1142 -558 1179 -548
rect 1238 -528 1325 -518
rect 1238 -548 1247 -528
rect 1267 -548 1325 -528
rect 1238 -557 1325 -548
rect 1238 -558 1275 -557
rect 99 -590 142 -585
rect 490 -579 937 -563
rect 490 -585 518 -579
rect 769 -580 937 -579
rect 99 -593 249 -590
rect 490 -593 517 -585
rect 99 -595 517 -593
rect 99 -613 108 -595
rect 126 -613 517 -595
rect 1294 -608 1325 -557
rect 1360 -528 1397 -458
rect 1663 -459 1700 -458
rect 1512 -518 1548 -517
rect 1360 -548 1369 -528
rect 1389 -548 1397 -528
rect 1360 -558 1397 -548
rect 1456 -528 1604 -518
rect 1704 -521 1800 -519
rect 1456 -548 1465 -528
rect 1485 -548 1575 -528
rect 1595 -548 1604 -528
rect 1456 -557 1604 -548
rect 1662 -528 1800 -521
rect 1662 -548 1671 -528
rect 1691 -548 1800 -528
rect 1662 -557 1800 -548
rect 1456 -558 1493 -557
rect 1186 -611 1227 -610
rect 99 -616 517 -613
rect 99 -622 142 -616
rect 102 -625 142 -622
rect 1078 -618 1227 -611
rect 499 -634 539 -633
rect 210 -651 539 -634
rect 1078 -638 1137 -618
rect 1157 -638 1196 -618
rect 1216 -638 1227 -618
rect 1078 -646 1227 -638
rect 1294 -615 1451 -608
rect 1294 -635 1414 -615
rect 1434 -635 1451 -615
rect 1294 -645 1451 -635
rect 1294 -646 1329 -645
rect 94 -694 137 -683
rect 94 -712 106 -694
rect 124 -712 137 -694
rect 94 -738 137 -712
rect 210 -738 237 -651
rect 499 -660 539 -651
rect 94 -759 237 -738
rect 281 -686 315 -670
rect 499 -680 892 -660
rect 912 -680 915 -660
rect 1294 -667 1325 -646
rect 1512 -667 1548 -557
rect 1567 -558 1604 -557
rect 1663 -558 1700 -557
rect 1623 -617 1713 -611
rect 1623 -637 1632 -617
rect 1652 -619 1713 -617
rect 1652 -637 1677 -619
rect 1623 -639 1677 -637
rect 1697 -639 1713 -619
rect 1623 -645 1713 -639
rect 1137 -668 1174 -667
rect 499 -685 915 -680
rect 1136 -677 1174 -668
rect 499 -686 840 -685
rect 281 -756 318 -686
rect 433 -746 464 -745
rect 94 -761 231 -759
rect 94 -803 137 -761
rect 281 -776 290 -756
rect 310 -776 318 -756
rect 281 -786 318 -776
rect 377 -756 464 -746
rect 377 -776 386 -756
rect 406 -776 464 -756
rect 377 -785 464 -776
rect 377 -786 414 -785
rect 92 -813 137 -803
rect 92 -831 101 -813
rect 119 -831 137 -813
rect 92 -837 137 -831
rect 433 -836 464 -785
rect 499 -756 536 -686
rect 802 -687 839 -686
rect 1136 -697 1145 -677
rect 1165 -697 1174 -677
rect 1136 -705 1174 -697
rect 1240 -673 1325 -667
rect 1355 -668 1392 -667
rect 1240 -693 1248 -673
rect 1268 -693 1325 -673
rect 1240 -701 1325 -693
rect 1354 -677 1392 -668
rect 1354 -697 1363 -677
rect 1383 -697 1392 -677
rect 1240 -702 1276 -701
rect 1354 -705 1392 -697
rect 1458 -673 1602 -667
rect 1458 -693 1466 -673
rect 1486 -676 1574 -673
rect 1486 -693 1521 -676
rect 1458 -694 1521 -693
rect 1540 -693 1574 -676
rect 1594 -693 1602 -673
rect 1540 -694 1602 -693
rect 1458 -701 1602 -694
rect 1458 -702 1494 -701
rect 1566 -702 1602 -701
rect 1668 -668 1705 -667
rect 1668 -669 1706 -668
rect 1728 -669 1755 -665
rect 1668 -671 1755 -669
rect 1668 -677 1732 -671
rect 1668 -697 1677 -677
rect 1697 -691 1732 -677
rect 1752 -691 1755 -671
rect 1697 -696 1755 -691
rect 1697 -697 1732 -696
rect 1137 -734 1174 -705
rect 1138 -736 1174 -734
rect 651 -746 687 -745
rect 499 -776 508 -756
rect 528 -776 536 -756
rect 499 -786 536 -776
rect 595 -756 743 -746
rect 843 -749 939 -747
rect 595 -776 604 -756
rect 624 -776 714 -756
rect 734 -776 743 -756
rect 595 -785 743 -776
rect 801 -756 939 -749
rect 801 -776 810 -756
rect 830 -776 939 -756
rect 1138 -758 1329 -736
rect 1355 -737 1392 -705
rect 1668 -709 1732 -697
rect 1772 -735 1799 -557
rect 1631 -737 1799 -735
rect 1355 -763 1799 -737
rect 801 -785 939 -776
rect 595 -786 632 -785
rect 92 -840 129 -837
rect 325 -839 366 -838
rect 217 -846 366 -839
rect 217 -866 276 -846
rect 296 -866 335 -846
rect 355 -866 366 -846
rect 217 -874 366 -866
rect 433 -843 590 -836
rect 433 -863 553 -843
rect 573 -863 590 -843
rect 433 -873 590 -863
rect 433 -874 468 -873
rect 433 -895 464 -874
rect 651 -895 687 -785
rect 706 -786 743 -785
rect 802 -786 839 -785
rect 762 -845 852 -839
rect 762 -865 771 -845
rect 791 -847 852 -845
rect 791 -865 816 -847
rect 762 -867 816 -865
rect 836 -867 852 -847
rect 762 -873 852 -867
rect 276 -896 313 -895
rect 89 -904 126 -902
rect 89 -912 131 -904
rect 89 -930 99 -912
rect 117 -930 131 -912
rect 89 -939 131 -930
rect 275 -905 313 -896
rect 275 -925 284 -905
rect 304 -925 313 -905
rect 275 -933 313 -925
rect 379 -901 464 -895
rect 494 -896 531 -895
rect 379 -921 387 -901
rect 407 -921 464 -901
rect 379 -929 464 -921
rect 493 -905 531 -896
rect 493 -925 502 -905
rect 522 -925 531 -905
rect 379 -930 415 -929
rect 493 -933 531 -925
rect 597 -897 741 -895
rect 597 -901 649 -897
rect 597 -921 605 -901
rect 625 -917 649 -901
rect 669 -901 741 -897
rect 669 -917 713 -901
rect 625 -921 713 -917
rect 733 -921 741 -901
rect 597 -929 741 -921
rect 597 -930 633 -929
rect 705 -930 741 -929
rect 807 -896 844 -895
rect 807 -897 845 -896
rect 807 -905 871 -897
rect 807 -925 816 -905
rect 836 -919 871 -905
rect 891 -919 894 -899
rect 836 -924 894 -919
rect 836 -925 871 -924
rect 90 -964 131 -939
rect 276 -964 313 -933
rect 494 -964 531 -933
rect 807 -937 871 -925
rect 911 -963 938 -785
rect 90 -965 574 -964
rect 770 -965 938 -963
rect 90 -990 938 -965
rect 90 -991 131 -990
rect 494 -991 938 -990
rect 770 -992 938 -991
rect 1465 -987 1505 -763
rect 1631 -764 1799 -763
rect 1863 -731 1896 -398
rect 1863 -739 1900 -731
rect 1863 -758 1871 -739
rect 1892 -758 1900 -739
rect 1863 -764 1900 -758
rect 1465 -1009 1473 -987
rect 1497 -1009 1505 -987
rect 1465 -1017 1505 -1009
<< viali >>
rect 908 750 928 770
rect 292 564 312 584
rect 832 563 852 583
rect 674 509 694 529
rect 887 511 907 531
rect 1770 566 1790 586
rect 1154 380 1174 400
rect 909 338 929 358
rect 1694 379 1714 399
rect 1535 326 1556 345
rect 1749 327 1769 347
rect 293 152 313 172
rect 833 151 853 171
rect 666 101 686 121
rect 888 99 908 119
rect 1490 9 1514 31
rect 1852 -42 1872 -22
rect 1236 -228 1256 -208
rect 891 -268 911 -248
rect 1776 -229 1796 -209
rect 1831 -281 1851 -261
rect 275 -454 295 -434
rect 815 -455 835 -435
rect 657 -509 677 -489
rect 870 -507 890 -487
rect 1753 -452 1773 -432
rect 1137 -638 1157 -618
rect 892 -680 912 -660
rect 1677 -639 1697 -619
rect 1521 -694 1540 -676
rect 1732 -691 1752 -671
rect 276 -866 296 -846
rect 816 -867 836 -847
rect 649 -917 669 -897
rect 871 -919 891 -899
rect 1871 -758 1892 -739
rect 1473 -1009 1497 -987
<< metal1 >>
rect 904 775 936 776
rect 901 770 936 775
rect 901 750 908 770
rect 928 750 936 770
rect 901 742 936 750
rect 283 584 868 592
rect 283 564 292 584
rect 312 583 868 584
rect 312 564 832 583
rect 283 563 832 564
rect 852 563 868 583
rect 283 557 868 563
rect 902 536 936 742
rect 666 529 701 536
rect 666 509 674 529
rect 694 509 701 529
rect 666 436 701 509
rect 880 531 936 536
rect 880 511 887 531
rect 907 511 936 531
rect 880 504 936 511
rect 971 638 1001 640
rect 1764 638 1797 639
rect 971 612 1798 638
rect 880 503 915 504
rect 971 437 1001 612
rect 1764 591 1798 612
rect 1763 586 1798 591
rect 1763 566 1770 586
rect 1790 566 1798 586
rect 1763 558 1798 566
rect 966 436 1001 437
rect 665 409 1001 436
rect 971 408 1001 409
rect 1145 400 1730 408
rect 1145 380 1154 400
rect 1174 399 1730 400
rect 1174 380 1694 399
rect 1145 379 1694 380
rect 1714 379 1730 399
rect 1145 373 1730 379
rect 905 363 937 364
rect 902 358 937 363
rect 902 338 909 358
rect 929 338 937 358
rect 1764 352 1798 558
rect 902 330 937 338
rect 284 172 869 180
rect 284 152 293 172
rect 313 171 869 172
rect 313 152 833 171
rect 284 151 833 152
rect 853 151 869 171
rect 284 145 869 151
rect 658 121 697 125
rect 903 124 937 330
rect 1530 345 1565 351
rect 1530 326 1535 345
rect 1556 326 1565 345
rect 1530 317 1565 326
rect 1742 347 1798 352
rect 1742 327 1749 347
rect 1769 327 1798 347
rect 1742 320 1798 327
rect 1742 319 1777 320
rect 1534 249 1563 317
rect 1534 215 1880 249
rect 658 101 666 121
rect 686 101 697 121
rect 658 26 697 101
rect 881 119 937 124
rect 881 99 888 119
rect 908 99 937 119
rect 881 92 937 99
rect 881 91 916 92
rect 1485 31 1524 44
rect 1485 26 1490 31
rect 658 9 1490 26
rect 1514 26 1524 31
rect 1514 9 1525 26
rect 658 1 1525 9
rect 660 0 946 1
rect 1841 -22 1880 215
rect 1841 -34 1852 -22
rect 1845 -42 1852 -34
rect 1872 -42 1880 -22
rect 1845 -50 1880 -42
rect 1227 -208 1812 -200
rect 1227 -228 1236 -208
rect 1256 -209 1812 -208
rect 1256 -228 1776 -209
rect 1227 -229 1776 -228
rect 1796 -229 1812 -209
rect 1227 -235 1812 -229
rect 887 -243 919 -242
rect 884 -248 919 -243
rect 884 -268 891 -248
rect 911 -268 919 -248
rect 1846 -256 1880 -50
rect 884 -276 919 -268
rect 266 -434 851 -426
rect 266 -454 275 -434
rect 295 -435 851 -434
rect 295 -454 815 -435
rect 266 -455 815 -454
rect 835 -455 851 -435
rect 266 -461 851 -455
rect 885 -482 919 -276
rect 1824 -261 1880 -256
rect 1824 -281 1831 -261
rect 1851 -281 1880 -261
rect 1824 -288 1880 -281
rect 1824 -289 1859 -288
rect 649 -489 684 -482
rect 649 -509 657 -489
rect 677 -509 684 -489
rect 649 -582 684 -509
rect 863 -487 919 -482
rect 863 -507 870 -487
rect 890 -507 919 -487
rect 863 -514 919 -507
rect 954 -380 984 -378
rect 1747 -380 1780 -379
rect 954 -406 1781 -380
rect 863 -515 898 -514
rect 954 -581 984 -406
rect 1747 -427 1781 -406
rect 1746 -432 1781 -427
rect 1746 -452 1753 -432
rect 1773 -452 1781 -432
rect 1746 -460 1781 -452
rect 949 -582 984 -581
rect 648 -609 984 -582
rect 954 -610 984 -609
rect 1128 -618 1713 -610
rect 1128 -638 1137 -618
rect 1157 -619 1713 -618
rect 1157 -638 1677 -619
rect 1128 -639 1677 -638
rect 1697 -639 1713 -619
rect 1128 -645 1713 -639
rect 888 -655 920 -654
rect 885 -660 920 -655
rect 885 -680 892 -660
rect 912 -680 920 -660
rect 1747 -666 1781 -460
rect 885 -688 920 -680
rect 267 -846 852 -838
rect 267 -866 276 -846
rect 296 -847 852 -846
rect 296 -866 816 -847
rect 267 -867 816 -866
rect 836 -867 852 -847
rect 267 -873 852 -867
rect 641 -897 680 -893
rect 886 -894 920 -688
rect 1514 -676 1548 -668
rect 1514 -694 1521 -676
rect 1540 -694 1548 -676
rect 1514 -701 1548 -694
rect 1725 -671 1781 -666
rect 1725 -691 1732 -671
rect 1752 -691 1781 -671
rect 1725 -698 1781 -691
rect 1725 -699 1760 -698
rect 1518 -731 1547 -701
rect 1518 -739 1900 -731
rect 1518 -758 1871 -739
rect 1892 -758 1900 -739
rect 1518 -763 1900 -758
rect 641 -917 649 -897
rect 669 -917 680 -897
rect 641 -992 680 -917
rect 864 -899 920 -894
rect 864 -919 871 -899
rect 891 -919 920 -899
rect 864 -926 920 -919
rect 864 -927 899 -926
rect 1468 -987 1507 -974
rect 1468 -992 1473 -987
rect 641 -1009 1473 -992
rect 1497 -992 1507 -987
rect 1497 -1009 1508 -992
rect 641 -1017 1508 -1009
rect 643 -1018 929 -1017
<< labels >>
rlabel locali 246 566 268 581 1 d0
rlabel locali 300 754 329 760 1 vdd
rlabel locali 297 455 326 461 1 gnd
rlabel space 403 473 432 482 1 gnd
rlabel nwell 435 731 458 734 1 vdd
rlabel locali 247 154 269 169 1 d0
rlabel locali 301 342 330 348 1 vdd
rlabel locali 298 43 327 49 1 gnd
rlabel space 404 61 433 70 1 gnd
rlabel nwell 436 319 459 322 1 vdd
rlabel locali 1162 570 1191 576 1 vdd
rlabel locali 1159 271 1188 277 1 gnd
rlabel space 1265 289 1294 298 1 gnd
rlabel nwell 1297 547 1320 550 1 vdd
rlabel locali 1102 378 1124 395 1 d1
rlabel locali 137 999 161 1029 1 vref
rlabel locali 229 -452 251 -437 1 d0
rlabel locali 283 -264 312 -258 1 vdd
rlabel locali 280 -563 309 -557 1 gnd
rlabel space 386 -545 415 -536 1 gnd
rlabel nwell 418 -287 441 -284 1 vdd
rlabel locali 230 -864 252 -849 1 d0
rlabel locali 284 -676 313 -670 1 vdd
rlabel locali 281 -975 310 -969 1 gnd
rlabel space 387 -957 416 -948 1 gnd
rlabel nwell 419 -699 442 -696 1 vdd
rlabel locali 1145 -448 1174 -442 1 vdd
rlabel locali 1142 -747 1171 -741 1 gnd
rlabel space 1248 -729 1277 -720 1 gnd
rlabel nwell 1280 -471 1303 -468 1 vdd
rlabel locali 1085 -640 1107 -623 1 d1
rlabel locali 96 -976 124 -958 1 gnd
rlabel locali 1244 -38 1273 -32 1 vdd
rlabel locali 1241 -337 1270 -331 1 gnd
rlabel space 1347 -319 1376 -310 1 gnd
rlabel nwell 1379 -61 1402 -58 1 vdd
rlabel locali 1617 -191 1639 -176 1 vout
rlabel locali 1186 -230 1206 -206 1 d2
<< end >>

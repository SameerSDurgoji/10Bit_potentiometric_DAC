magic
tech sky130A
timestamp 1616092942
<< nwell >>
rect 3450 7874 4058 8024
rect 401 7720 1009 7870
rect 1199 7536 1807 7686
rect 2653 7646 3261 7796
rect 3451 7462 4059 7612
rect 402 7308 1010 7458
rect 2554 7236 3162 7386
rect 1281 6928 1889 7078
rect 3433 6856 4041 7006
rect 384 6702 992 6852
rect 1182 6518 1790 6668
rect 2636 6628 3244 6778
rect 3434 6444 4042 6594
rect 385 6290 993 6440
rect 2471 6220 3079 6370
rect 1327 5908 1935 6058
rect 3413 5838 4021 5988
rect 364 5684 972 5834
rect 1162 5500 1770 5650
rect 2616 5610 3224 5760
rect 3414 5426 4022 5576
rect 365 5272 973 5422
rect 2517 5200 3125 5350
rect 1244 4892 1852 5042
rect 3396 4820 4004 4970
rect 347 4666 955 4816
rect 1145 4482 1753 4632
rect 2599 4592 3207 4742
rect 3397 4408 4005 4558
rect 348 4254 956 4404
rect 2295 4186 2903 4336
rect 1430 3870 2038 4020
rect 3377 3802 3985 3952
rect 328 3648 936 3798
rect 1126 3464 1734 3614
rect 2580 3574 3188 3724
rect 3378 3390 3986 3540
rect 329 3236 937 3386
rect 2481 3164 3089 3314
rect 1208 2856 1816 3006
rect 3360 2784 3968 2934
rect 311 2630 919 2780
rect 1109 2446 1717 2596
rect 2563 2556 3171 2706
rect 3361 2372 3969 2522
rect 312 2218 920 2368
rect 2398 2148 3006 2298
rect 1254 1836 1862 1986
rect 3340 1766 3948 1916
rect 291 1612 899 1762
rect 1089 1428 1697 1578
rect 2543 1538 3151 1688
rect 3341 1354 3949 1504
rect 292 1200 900 1350
rect 2444 1128 3052 1278
rect 1171 820 1779 970
rect 3323 748 3931 898
rect 274 594 882 744
rect 1072 410 1680 560
rect 2526 520 3134 670
rect 3324 336 3932 486
rect 275 182 883 332
rect 1488 -394 2096 -244
<< nmos >>
rect 3518 8083 3568 8125
rect 3726 8083 3776 8125
rect 3944 8083 3994 8125
rect 2721 7855 2771 7897
rect 2929 7855 2979 7897
rect 3147 7855 3197 7897
rect 465 7619 515 7661
rect 683 7619 733 7661
rect 891 7619 941 7661
rect 3519 7671 3569 7713
rect 3727 7671 3777 7713
rect 3945 7671 3995 7713
rect 1263 7435 1313 7477
rect 1481 7435 1531 7477
rect 1689 7435 1739 7477
rect 2622 7445 2672 7487
rect 2830 7445 2880 7487
rect 3048 7445 3098 7487
rect 466 7207 516 7249
rect 684 7207 734 7249
rect 892 7207 942 7249
rect 3501 7065 3551 7107
rect 3709 7065 3759 7107
rect 3927 7065 3977 7107
rect 1345 6827 1395 6869
rect 1563 6827 1613 6869
rect 1771 6827 1821 6869
rect 2704 6837 2754 6879
rect 2912 6837 2962 6879
rect 3130 6837 3180 6879
rect 448 6601 498 6643
rect 666 6601 716 6643
rect 874 6601 924 6643
rect 3502 6653 3552 6695
rect 3710 6653 3760 6695
rect 3928 6653 3978 6695
rect 1246 6417 1296 6459
rect 1464 6417 1514 6459
rect 1672 6417 1722 6459
rect 2539 6429 2589 6471
rect 2747 6429 2797 6471
rect 2965 6429 3015 6471
rect 449 6189 499 6231
rect 667 6189 717 6231
rect 875 6189 925 6231
rect 3481 6047 3531 6089
rect 3689 6047 3739 6089
rect 3907 6047 3957 6089
rect 1391 5807 1441 5849
rect 1609 5807 1659 5849
rect 1817 5807 1867 5849
rect 2684 5819 2734 5861
rect 2892 5819 2942 5861
rect 3110 5819 3160 5861
rect 428 5583 478 5625
rect 646 5583 696 5625
rect 854 5583 904 5625
rect 3482 5635 3532 5677
rect 3690 5635 3740 5677
rect 3908 5635 3958 5677
rect 1226 5399 1276 5441
rect 1444 5399 1494 5441
rect 1652 5399 1702 5441
rect 2585 5409 2635 5451
rect 2793 5409 2843 5451
rect 3011 5409 3061 5451
rect 429 5171 479 5213
rect 647 5171 697 5213
rect 855 5171 905 5213
rect 3464 5029 3514 5071
rect 3672 5029 3722 5071
rect 3890 5029 3940 5071
rect 1308 4791 1358 4833
rect 1526 4791 1576 4833
rect 1734 4791 1784 4833
rect 2667 4801 2717 4843
rect 2875 4801 2925 4843
rect 3093 4801 3143 4843
rect 411 4565 461 4607
rect 629 4565 679 4607
rect 837 4565 887 4607
rect 3465 4617 3515 4659
rect 3673 4617 3723 4659
rect 3891 4617 3941 4659
rect 1209 4381 1259 4423
rect 1427 4381 1477 4423
rect 1635 4381 1685 4423
rect 2363 4395 2413 4437
rect 2571 4395 2621 4437
rect 2789 4395 2839 4437
rect 412 4153 462 4195
rect 630 4153 680 4195
rect 838 4153 888 4195
rect 3445 4011 3495 4053
rect 3653 4011 3703 4053
rect 3871 4011 3921 4053
rect 1494 3769 1544 3811
rect 1712 3769 1762 3811
rect 1920 3769 1970 3811
rect 2648 3783 2698 3825
rect 2856 3783 2906 3825
rect 3074 3783 3124 3825
rect 392 3547 442 3589
rect 610 3547 660 3589
rect 818 3547 868 3589
rect 3446 3599 3496 3641
rect 3654 3599 3704 3641
rect 3872 3599 3922 3641
rect 1190 3363 1240 3405
rect 1408 3363 1458 3405
rect 1616 3363 1666 3405
rect 2549 3373 2599 3415
rect 2757 3373 2807 3415
rect 2975 3373 3025 3415
rect 393 3135 443 3177
rect 611 3135 661 3177
rect 819 3135 869 3177
rect 3428 2993 3478 3035
rect 3636 2993 3686 3035
rect 3854 2993 3904 3035
rect 1272 2755 1322 2797
rect 1490 2755 1540 2797
rect 1698 2755 1748 2797
rect 2631 2765 2681 2807
rect 2839 2765 2889 2807
rect 3057 2765 3107 2807
rect 375 2529 425 2571
rect 593 2529 643 2571
rect 801 2529 851 2571
rect 3429 2581 3479 2623
rect 3637 2581 3687 2623
rect 3855 2581 3905 2623
rect 1173 2345 1223 2387
rect 1391 2345 1441 2387
rect 1599 2345 1649 2387
rect 2466 2357 2516 2399
rect 2674 2357 2724 2399
rect 2892 2357 2942 2399
rect 376 2117 426 2159
rect 594 2117 644 2159
rect 802 2117 852 2159
rect 3408 1975 3458 2017
rect 3616 1975 3666 2017
rect 3834 1975 3884 2017
rect 1318 1735 1368 1777
rect 1536 1735 1586 1777
rect 1744 1735 1794 1777
rect 2611 1747 2661 1789
rect 2819 1747 2869 1789
rect 3037 1747 3087 1789
rect 355 1511 405 1553
rect 573 1511 623 1553
rect 781 1511 831 1553
rect 3409 1563 3459 1605
rect 3617 1563 3667 1605
rect 3835 1563 3885 1605
rect 1153 1327 1203 1369
rect 1371 1327 1421 1369
rect 1579 1327 1629 1369
rect 2512 1337 2562 1379
rect 2720 1337 2770 1379
rect 2938 1337 2988 1379
rect 356 1099 406 1141
rect 574 1099 624 1141
rect 782 1099 832 1141
rect 3391 957 3441 999
rect 3599 957 3649 999
rect 3817 957 3867 999
rect 1235 719 1285 761
rect 1453 719 1503 761
rect 1661 719 1711 761
rect 2594 729 2644 771
rect 2802 729 2852 771
rect 3020 729 3070 771
rect 338 493 388 535
rect 556 493 606 535
rect 764 493 814 535
rect 3392 545 3442 587
rect 3600 545 3650 587
rect 3818 545 3868 587
rect 1136 309 1186 351
rect 1354 309 1404 351
rect 1562 309 1612 351
rect 339 81 389 123
rect 557 81 607 123
rect 765 81 815 123
rect 1552 -495 1602 -453
rect 1770 -495 1820 -453
rect 1978 -495 2028 -453
<< pmos >>
rect 3518 7906 3568 8006
rect 3726 7906 3776 8006
rect 3944 7906 3994 8006
rect 465 7738 515 7838
rect 683 7738 733 7838
rect 891 7738 941 7838
rect 2721 7678 2771 7778
rect 2929 7678 2979 7778
rect 3147 7678 3197 7778
rect 1263 7554 1313 7654
rect 1481 7554 1531 7654
rect 1689 7554 1739 7654
rect 3519 7494 3569 7594
rect 3727 7494 3777 7594
rect 3945 7494 3995 7594
rect 466 7326 516 7426
rect 684 7326 734 7426
rect 892 7326 942 7426
rect 2622 7268 2672 7368
rect 2830 7268 2880 7368
rect 3048 7268 3098 7368
rect 1345 6946 1395 7046
rect 1563 6946 1613 7046
rect 1771 6946 1821 7046
rect 3501 6888 3551 6988
rect 3709 6888 3759 6988
rect 3927 6888 3977 6988
rect 448 6720 498 6820
rect 666 6720 716 6820
rect 874 6720 924 6820
rect 2704 6660 2754 6760
rect 2912 6660 2962 6760
rect 3130 6660 3180 6760
rect 1246 6536 1296 6636
rect 1464 6536 1514 6636
rect 1672 6536 1722 6636
rect 3502 6476 3552 6576
rect 3710 6476 3760 6576
rect 3928 6476 3978 6576
rect 449 6308 499 6408
rect 667 6308 717 6408
rect 875 6308 925 6408
rect 2539 6252 2589 6352
rect 2747 6252 2797 6352
rect 2965 6252 3015 6352
rect 1391 5926 1441 6026
rect 1609 5926 1659 6026
rect 1817 5926 1867 6026
rect 3481 5870 3531 5970
rect 3689 5870 3739 5970
rect 3907 5870 3957 5970
rect 428 5702 478 5802
rect 646 5702 696 5802
rect 854 5702 904 5802
rect 2684 5642 2734 5742
rect 2892 5642 2942 5742
rect 3110 5642 3160 5742
rect 1226 5518 1276 5618
rect 1444 5518 1494 5618
rect 1652 5518 1702 5618
rect 3482 5458 3532 5558
rect 3690 5458 3740 5558
rect 3908 5458 3958 5558
rect 429 5290 479 5390
rect 647 5290 697 5390
rect 855 5290 905 5390
rect 2585 5232 2635 5332
rect 2793 5232 2843 5332
rect 3011 5232 3061 5332
rect 1308 4910 1358 5010
rect 1526 4910 1576 5010
rect 1734 4910 1784 5010
rect 3464 4852 3514 4952
rect 3672 4852 3722 4952
rect 3890 4852 3940 4952
rect 411 4684 461 4784
rect 629 4684 679 4784
rect 837 4684 887 4784
rect 2667 4624 2717 4724
rect 2875 4624 2925 4724
rect 3093 4624 3143 4724
rect 1209 4500 1259 4600
rect 1427 4500 1477 4600
rect 1635 4500 1685 4600
rect 3465 4440 3515 4540
rect 3673 4440 3723 4540
rect 3891 4440 3941 4540
rect 412 4272 462 4372
rect 630 4272 680 4372
rect 838 4272 888 4372
rect 2363 4218 2413 4318
rect 2571 4218 2621 4318
rect 2789 4218 2839 4318
rect 1494 3888 1544 3988
rect 1712 3888 1762 3988
rect 1920 3888 1970 3988
rect 3445 3834 3495 3934
rect 3653 3834 3703 3934
rect 3871 3834 3921 3934
rect 392 3666 442 3766
rect 610 3666 660 3766
rect 818 3666 868 3766
rect 2648 3606 2698 3706
rect 2856 3606 2906 3706
rect 3074 3606 3124 3706
rect 1190 3482 1240 3582
rect 1408 3482 1458 3582
rect 1616 3482 1666 3582
rect 3446 3422 3496 3522
rect 3654 3422 3704 3522
rect 3872 3422 3922 3522
rect 393 3254 443 3354
rect 611 3254 661 3354
rect 819 3254 869 3354
rect 2549 3196 2599 3296
rect 2757 3196 2807 3296
rect 2975 3196 3025 3296
rect 1272 2874 1322 2974
rect 1490 2874 1540 2974
rect 1698 2874 1748 2974
rect 3428 2816 3478 2916
rect 3636 2816 3686 2916
rect 3854 2816 3904 2916
rect 375 2648 425 2748
rect 593 2648 643 2748
rect 801 2648 851 2748
rect 2631 2588 2681 2688
rect 2839 2588 2889 2688
rect 3057 2588 3107 2688
rect 1173 2464 1223 2564
rect 1391 2464 1441 2564
rect 1599 2464 1649 2564
rect 3429 2404 3479 2504
rect 3637 2404 3687 2504
rect 3855 2404 3905 2504
rect 376 2236 426 2336
rect 594 2236 644 2336
rect 802 2236 852 2336
rect 2466 2180 2516 2280
rect 2674 2180 2724 2280
rect 2892 2180 2942 2280
rect 1318 1854 1368 1954
rect 1536 1854 1586 1954
rect 1744 1854 1794 1954
rect 3408 1798 3458 1898
rect 3616 1798 3666 1898
rect 3834 1798 3884 1898
rect 355 1630 405 1730
rect 573 1630 623 1730
rect 781 1630 831 1730
rect 2611 1570 2661 1670
rect 2819 1570 2869 1670
rect 3037 1570 3087 1670
rect 1153 1446 1203 1546
rect 1371 1446 1421 1546
rect 1579 1446 1629 1546
rect 3409 1386 3459 1486
rect 3617 1386 3667 1486
rect 3835 1386 3885 1486
rect 356 1218 406 1318
rect 574 1218 624 1318
rect 782 1218 832 1318
rect 2512 1160 2562 1260
rect 2720 1160 2770 1260
rect 2938 1160 2988 1260
rect 1235 838 1285 938
rect 1453 838 1503 938
rect 1661 838 1711 938
rect 3391 780 3441 880
rect 3599 780 3649 880
rect 3817 780 3867 880
rect 338 612 388 712
rect 556 612 606 712
rect 764 612 814 712
rect 2594 552 2644 652
rect 2802 552 2852 652
rect 3020 552 3070 652
rect 1136 428 1186 528
rect 1354 428 1404 528
rect 1562 428 1612 528
rect 3392 368 3442 468
rect 3600 368 3650 468
rect 3818 368 3868 468
rect 339 200 389 300
rect 557 200 607 300
rect 765 200 815 300
rect 1552 -376 1602 -276
rect 1770 -376 1820 -276
rect 1978 -376 2028 -276
<< ndiff >>
rect 3469 8113 3518 8125
rect 3469 8093 3480 8113
rect 3500 8093 3518 8113
rect 3469 8083 3518 8093
rect 3568 8109 3612 8125
rect 3568 8089 3583 8109
rect 3603 8089 3612 8109
rect 3568 8083 3612 8089
rect 3682 8109 3726 8125
rect 3682 8089 3691 8109
rect 3711 8089 3726 8109
rect 3682 8083 3726 8089
rect 3776 8113 3825 8125
rect 3776 8093 3794 8113
rect 3814 8093 3825 8113
rect 3776 8083 3825 8093
rect 3900 8109 3944 8125
rect 3900 8089 3909 8109
rect 3929 8089 3944 8109
rect 3900 8083 3944 8089
rect 3994 8113 4043 8125
rect 3994 8093 4012 8113
rect 4032 8093 4043 8113
rect 3994 8083 4043 8093
rect 2672 7885 2721 7897
rect 2672 7865 2683 7885
rect 2703 7865 2721 7885
rect 2672 7855 2721 7865
rect 2771 7881 2815 7897
rect 2771 7861 2786 7881
rect 2806 7861 2815 7881
rect 2771 7855 2815 7861
rect 2885 7881 2929 7897
rect 2885 7861 2894 7881
rect 2914 7861 2929 7881
rect 2885 7855 2929 7861
rect 2979 7885 3028 7897
rect 2979 7865 2997 7885
rect 3017 7865 3028 7885
rect 2979 7855 3028 7865
rect 3103 7881 3147 7897
rect 3103 7861 3112 7881
rect 3132 7861 3147 7881
rect 3103 7855 3147 7861
rect 3197 7885 3246 7897
rect 3197 7865 3215 7885
rect 3235 7865 3246 7885
rect 3197 7855 3246 7865
rect 3470 7701 3519 7713
rect 3470 7681 3481 7701
rect 3501 7681 3519 7701
rect 416 7651 465 7661
rect 416 7631 427 7651
rect 447 7631 465 7651
rect 416 7619 465 7631
rect 515 7655 559 7661
rect 515 7635 530 7655
rect 550 7635 559 7655
rect 515 7619 559 7635
rect 634 7651 683 7661
rect 634 7631 645 7651
rect 665 7631 683 7651
rect 634 7619 683 7631
rect 733 7655 777 7661
rect 733 7635 748 7655
rect 768 7635 777 7655
rect 733 7619 777 7635
rect 847 7655 891 7661
rect 847 7635 856 7655
rect 876 7635 891 7655
rect 847 7619 891 7635
rect 941 7651 990 7661
rect 3470 7671 3519 7681
rect 3569 7697 3613 7713
rect 3569 7677 3584 7697
rect 3604 7677 3613 7697
rect 3569 7671 3613 7677
rect 3683 7697 3727 7713
rect 3683 7677 3692 7697
rect 3712 7677 3727 7697
rect 3683 7671 3727 7677
rect 3777 7701 3826 7713
rect 3777 7681 3795 7701
rect 3815 7681 3826 7701
rect 3777 7671 3826 7681
rect 3901 7697 3945 7713
rect 3901 7677 3910 7697
rect 3930 7677 3945 7697
rect 3901 7671 3945 7677
rect 3995 7701 4044 7713
rect 3995 7681 4013 7701
rect 4033 7681 4044 7701
rect 3995 7671 4044 7681
rect 941 7631 959 7651
rect 979 7631 990 7651
rect 941 7619 990 7631
rect 1214 7467 1263 7477
rect 1214 7447 1225 7467
rect 1245 7447 1263 7467
rect 1214 7435 1263 7447
rect 1313 7471 1357 7477
rect 1313 7451 1328 7471
rect 1348 7451 1357 7471
rect 1313 7435 1357 7451
rect 1432 7467 1481 7477
rect 1432 7447 1443 7467
rect 1463 7447 1481 7467
rect 1432 7435 1481 7447
rect 1531 7471 1575 7477
rect 1531 7451 1546 7471
rect 1566 7451 1575 7471
rect 1531 7435 1575 7451
rect 1645 7471 1689 7477
rect 1645 7451 1654 7471
rect 1674 7451 1689 7471
rect 1645 7435 1689 7451
rect 1739 7467 1788 7477
rect 1739 7447 1757 7467
rect 1777 7447 1788 7467
rect 1739 7435 1788 7447
rect 2573 7475 2622 7487
rect 2573 7455 2584 7475
rect 2604 7455 2622 7475
rect 2573 7445 2622 7455
rect 2672 7471 2716 7487
rect 2672 7451 2687 7471
rect 2707 7451 2716 7471
rect 2672 7445 2716 7451
rect 2786 7471 2830 7487
rect 2786 7451 2795 7471
rect 2815 7451 2830 7471
rect 2786 7445 2830 7451
rect 2880 7475 2929 7487
rect 2880 7455 2898 7475
rect 2918 7455 2929 7475
rect 2880 7445 2929 7455
rect 3004 7471 3048 7487
rect 3004 7451 3013 7471
rect 3033 7451 3048 7471
rect 3004 7445 3048 7451
rect 3098 7475 3147 7487
rect 3098 7455 3116 7475
rect 3136 7455 3147 7475
rect 3098 7445 3147 7455
rect 417 7239 466 7249
rect 417 7219 428 7239
rect 448 7219 466 7239
rect 417 7207 466 7219
rect 516 7243 560 7249
rect 516 7223 531 7243
rect 551 7223 560 7243
rect 516 7207 560 7223
rect 635 7239 684 7249
rect 635 7219 646 7239
rect 666 7219 684 7239
rect 635 7207 684 7219
rect 734 7243 778 7249
rect 734 7223 749 7243
rect 769 7223 778 7243
rect 734 7207 778 7223
rect 848 7243 892 7249
rect 848 7223 857 7243
rect 877 7223 892 7243
rect 848 7207 892 7223
rect 942 7239 991 7249
rect 942 7219 960 7239
rect 980 7219 991 7239
rect 942 7207 991 7219
rect 3452 7095 3501 7107
rect 3452 7075 3463 7095
rect 3483 7075 3501 7095
rect 3452 7065 3501 7075
rect 3551 7091 3595 7107
rect 3551 7071 3566 7091
rect 3586 7071 3595 7091
rect 3551 7065 3595 7071
rect 3665 7091 3709 7107
rect 3665 7071 3674 7091
rect 3694 7071 3709 7091
rect 3665 7065 3709 7071
rect 3759 7095 3808 7107
rect 3759 7075 3777 7095
rect 3797 7075 3808 7095
rect 3759 7065 3808 7075
rect 3883 7091 3927 7107
rect 3883 7071 3892 7091
rect 3912 7071 3927 7091
rect 3883 7065 3927 7071
rect 3977 7095 4026 7107
rect 3977 7075 3995 7095
rect 4015 7075 4026 7095
rect 3977 7065 4026 7075
rect 1296 6859 1345 6869
rect 1296 6839 1307 6859
rect 1327 6839 1345 6859
rect 1296 6827 1345 6839
rect 1395 6863 1439 6869
rect 1395 6843 1410 6863
rect 1430 6843 1439 6863
rect 1395 6827 1439 6843
rect 1514 6859 1563 6869
rect 1514 6839 1525 6859
rect 1545 6839 1563 6859
rect 1514 6827 1563 6839
rect 1613 6863 1657 6869
rect 1613 6843 1628 6863
rect 1648 6843 1657 6863
rect 1613 6827 1657 6843
rect 1727 6863 1771 6869
rect 1727 6843 1736 6863
rect 1756 6843 1771 6863
rect 1727 6827 1771 6843
rect 1821 6859 1870 6869
rect 1821 6839 1839 6859
rect 1859 6839 1870 6859
rect 1821 6827 1870 6839
rect 2655 6867 2704 6879
rect 2655 6847 2666 6867
rect 2686 6847 2704 6867
rect 2655 6837 2704 6847
rect 2754 6863 2798 6879
rect 2754 6843 2769 6863
rect 2789 6843 2798 6863
rect 2754 6837 2798 6843
rect 2868 6863 2912 6879
rect 2868 6843 2877 6863
rect 2897 6843 2912 6863
rect 2868 6837 2912 6843
rect 2962 6867 3011 6879
rect 2962 6847 2980 6867
rect 3000 6847 3011 6867
rect 2962 6837 3011 6847
rect 3086 6863 3130 6879
rect 3086 6843 3095 6863
rect 3115 6843 3130 6863
rect 3086 6837 3130 6843
rect 3180 6867 3229 6879
rect 3180 6847 3198 6867
rect 3218 6847 3229 6867
rect 3180 6837 3229 6847
rect 3453 6683 3502 6695
rect 3453 6663 3464 6683
rect 3484 6663 3502 6683
rect 399 6633 448 6643
rect 399 6613 410 6633
rect 430 6613 448 6633
rect 399 6601 448 6613
rect 498 6637 542 6643
rect 498 6617 513 6637
rect 533 6617 542 6637
rect 498 6601 542 6617
rect 617 6633 666 6643
rect 617 6613 628 6633
rect 648 6613 666 6633
rect 617 6601 666 6613
rect 716 6637 760 6643
rect 716 6617 731 6637
rect 751 6617 760 6637
rect 716 6601 760 6617
rect 830 6637 874 6643
rect 830 6617 839 6637
rect 859 6617 874 6637
rect 830 6601 874 6617
rect 924 6633 973 6643
rect 3453 6653 3502 6663
rect 3552 6679 3596 6695
rect 3552 6659 3567 6679
rect 3587 6659 3596 6679
rect 3552 6653 3596 6659
rect 3666 6679 3710 6695
rect 3666 6659 3675 6679
rect 3695 6659 3710 6679
rect 3666 6653 3710 6659
rect 3760 6683 3809 6695
rect 3760 6663 3778 6683
rect 3798 6663 3809 6683
rect 3760 6653 3809 6663
rect 3884 6679 3928 6695
rect 3884 6659 3893 6679
rect 3913 6659 3928 6679
rect 3884 6653 3928 6659
rect 3978 6683 4027 6695
rect 3978 6663 3996 6683
rect 4016 6663 4027 6683
rect 3978 6653 4027 6663
rect 924 6613 942 6633
rect 962 6613 973 6633
rect 924 6601 973 6613
rect 2490 6459 2539 6471
rect 1197 6449 1246 6459
rect 1197 6429 1208 6449
rect 1228 6429 1246 6449
rect 1197 6417 1246 6429
rect 1296 6453 1340 6459
rect 1296 6433 1311 6453
rect 1331 6433 1340 6453
rect 1296 6417 1340 6433
rect 1415 6449 1464 6459
rect 1415 6429 1426 6449
rect 1446 6429 1464 6449
rect 1415 6417 1464 6429
rect 1514 6453 1558 6459
rect 1514 6433 1529 6453
rect 1549 6433 1558 6453
rect 1514 6417 1558 6433
rect 1628 6453 1672 6459
rect 1628 6433 1637 6453
rect 1657 6433 1672 6453
rect 1628 6417 1672 6433
rect 1722 6449 1771 6459
rect 1722 6429 1740 6449
rect 1760 6429 1771 6449
rect 2490 6439 2501 6459
rect 2521 6439 2539 6459
rect 2490 6429 2539 6439
rect 2589 6455 2633 6471
rect 2589 6435 2604 6455
rect 2624 6435 2633 6455
rect 2589 6429 2633 6435
rect 2703 6455 2747 6471
rect 2703 6435 2712 6455
rect 2732 6435 2747 6455
rect 2703 6429 2747 6435
rect 2797 6459 2846 6471
rect 2797 6439 2815 6459
rect 2835 6439 2846 6459
rect 2797 6429 2846 6439
rect 2921 6455 2965 6471
rect 2921 6435 2930 6455
rect 2950 6435 2965 6455
rect 2921 6429 2965 6435
rect 3015 6459 3064 6471
rect 3015 6439 3033 6459
rect 3053 6439 3064 6459
rect 3015 6429 3064 6439
rect 1722 6417 1771 6429
rect 400 6221 449 6231
rect 400 6201 411 6221
rect 431 6201 449 6221
rect 400 6189 449 6201
rect 499 6225 543 6231
rect 499 6205 514 6225
rect 534 6205 543 6225
rect 499 6189 543 6205
rect 618 6221 667 6231
rect 618 6201 629 6221
rect 649 6201 667 6221
rect 618 6189 667 6201
rect 717 6225 761 6231
rect 717 6205 732 6225
rect 752 6205 761 6225
rect 717 6189 761 6205
rect 831 6225 875 6231
rect 831 6205 840 6225
rect 860 6205 875 6225
rect 831 6189 875 6205
rect 925 6221 974 6231
rect 925 6201 943 6221
rect 963 6201 974 6221
rect 925 6189 974 6201
rect 3432 6077 3481 6089
rect 3432 6057 3443 6077
rect 3463 6057 3481 6077
rect 3432 6047 3481 6057
rect 3531 6073 3575 6089
rect 3531 6053 3546 6073
rect 3566 6053 3575 6073
rect 3531 6047 3575 6053
rect 3645 6073 3689 6089
rect 3645 6053 3654 6073
rect 3674 6053 3689 6073
rect 3645 6047 3689 6053
rect 3739 6077 3788 6089
rect 3739 6057 3757 6077
rect 3777 6057 3788 6077
rect 3739 6047 3788 6057
rect 3863 6073 3907 6089
rect 3863 6053 3872 6073
rect 3892 6053 3907 6073
rect 3863 6047 3907 6053
rect 3957 6077 4006 6089
rect 3957 6057 3975 6077
rect 3995 6057 4006 6077
rect 3957 6047 4006 6057
rect 2635 5849 2684 5861
rect 1342 5839 1391 5849
rect 1342 5819 1353 5839
rect 1373 5819 1391 5839
rect 1342 5807 1391 5819
rect 1441 5843 1485 5849
rect 1441 5823 1456 5843
rect 1476 5823 1485 5843
rect 1441 5807 1485 5823
rect 1560 5839 1609 5849
rect 1560 5819 1571 5839
rect 1591 5819 1609 5839
rect 1560 5807 1609 5819
rect 1659 5843 1703 5849
rect 1659 5823 1674 5843
rect 1694 5823 1703 5843
rect 1659 5807 1703 5823
rect 1773 5843 1817 5849
rect 1773 5823 1782 5843
rect 1802 5823 1817 5843
rect 1773 5807 1817 5823
rect 1867 5839 1916 5849
rect 1867 5819 1885 5839
rect 1905 5819 1916 5839
rect 2635 5829 2646 5849
rect 2666 5829 2684 5849
rect 2635 5819 2684 5829
rect 2734 5845 2778 5861
rect 2734 5825 2749 5845
rect 2769 5825 2778 5845
rect 2734 5819 2778 5825
rect 2848 5845 2892 5861
rect 2848 5825 2857 5845
rect 2877 5825 2892 5845
rect 2848 5819 2892 5825
rect 2942 5849 2991 5861
rect 2942 5829 2960 5849
rect 2980 5829 2991 5849
rect 2942 5819 2991 5829
rect 3066 5845 3110 5861
rect 3066 5825 3075 5845
rect 3095 5825 3110 5845
rect 3066 5819 3110 5825
rect 3160 5849 3209 5861
rect 3160 5829 3178 5849
rect 3198 5829 3209 5849
rect 3160 5819 3209 5829
rect 1867 5807 1916 5819
rect 3433 5665 3482 5677
rect 3433 5645 3444 5665
rect 3464 5645 3482 5665
rect 379 5615 428 5625
rect 379 5595 390 5615
rect 410 5595 428 5615
rect 379 5583 428 5595
rect 478 5619 522 5625
rect 478 5599 493 5619
rect 513 5599 522 5619
rect 478 5583 522 5599
rect 597 5615 646 5625
rect 597 5595 608 5615
rect 628 5595 646 5615
rect 597 5583 646 5595
rect 696 5619 740 5625
rect 696 5599 711 5619
rect 731 5599 740 5619
rect 696 5583 740 5599
rect 810 5619 854 5625
rect 810 5599 819 5619
rect 839 5599 854 5619
rect 810 5583 854 5599
rect 904 5615 953 5625
rect 3433 5635 3482 5645
rect 3532 5661 3576 5677
rect 3532 5641 3547 5661
rect 3567 5641 3576 5661
rect 3532 5635 3576 5641
rect 3646 5661 3690 5677
rect 3646 5641 3655 5661
rect 3675 5641 3690 5661
rect 3646 5635 3690 5641
rect 3740 5665 3789 5677
rect 3740 5645 3758 5665
rect 3778 5645 3789 5665
rect 3740 5635 3789 5645
rect 3864 5661 3908 5677
rect 3864 5641 3873 5661
rect 3893 5641 3908 5661
rect 3864 5635 3908 5641
rect 3958 5665 4007 5677
rect 3958 5645 3976 5665
rect 3996 5645 4007 5665
rect 3958 5635 4007 5645
rect 904 5595 922 5615
rect 942 5595 953 5615
rect 904 5583 953 5595
rect 1177 5431 1226 5441
rect 1177 5411 1188 5431
rect 1208 5411 1226 5431
rect 1177 5399 1226 5411
rect 1276 5435 1320 5441
rect 1276 5415 1291 5435
rect 1311 5415 1320 5435
rect 1276 5399 1320 5415
rect 1395 5431 1444 5441
rect 1395 5411 1406 5431
rect 1426 5411 1444 5431
rect 1395 5399 1444 5411
rect 1494 5435 1538 5441
rect 1494 5415 1509 5435
rect 1529 5415 1538 5435
rect 1494 5399 1538 5415
rect 1608 5435 1652 5441
rect 1608 5415 1617 5435
rect 1637 5415 1652 5435
rect 1608 5399 1652 5415
rect 1702 5431 1751 5441
rect 1702 5411 1720 5431
rect 1740 5411 1751 5431
rect 1702 5399 1751 5411
rect 2536 5439 2585 5451
rect 2536 5419 2547 5439
rect 2567 5419 2585 5439
rect 2536 5409 2585 5419
rect 2635 5435 2679 5451
rect 2635 5415 2650 5435
rect 2670 5415 2679 5435
rect 2635 5409 2679 5415
rect 2749 5435 2793 5451
rect 2749 5415 2758 5435
rect 2778 5415 2793 5435
rect 2749 5409 2793 5415
rect 2843 5439 2892 5451
rect 2843 5419 2861 5439
rect 2881 5419 2892 5439
rect 2843 5409 2892 5419
rect 2967 5435 3011 5451
rect 2967 5415 2976 5435
rect 2996 5415 3011 5435
rect 2967 5409 3011 5415
rect 3061 5439 3110 5451
rect 3061 5419 3079 5439
rect 3099 5419 3110 5439
rect 3061 5409 3110 5419
rect 380 5203 429 5213
rect 380 5183 391 5203
rect 411 5183 429 5203
rect 380 5171 429 5183
rect 479 5207 523 5213
rect 479 5187 494 5207
rect 514 5187 523 5207
rect 479 5171 523 5187
rect 598 5203 647 5213
rect 598 5183 609 5203
rect 629 5183 647 5203
rect 598 5171 647 5183
rect 697 5207 741 5213
rect 697 5187 712 5207
rect 732 5187 741 5207
rect 697 5171 741 5187
rect 811 5207 855 5213
rect 811 5187 820 5207
rect 840 5187 855 5207
rect 811 5171 855 5187
rect 905 5203 954 5213
rect 905 5183 923 5203
rect 943 5183 954 5203
rect 905 5171 954 5183
rect 3415 5059 3464 5071
rect 3415 5039 3426 5059
rect 3446 5039 3464 5059
rect 3415 5029 3464 5039
rect 3514 5055 3558 5071
rect 3514 5035 3529 5055
rect 3549 5035 3558 5055
rect 3514 5029 3558 5035
rect 3628 5055 3672 5071
rect 3628 5035 3637 5055
rect 3657 5035 3672 5055
rect 3628 5029 3672 5035
rect 3722 5059 3771 5071
rect 3722 5039 3740 5059
rect 3760 5039 3771 5059
rect 3722 5029 3771 5039
rect 3846 5055 3890 5071
rect 3846 5035 3855 5055
rect 3875 5035 3890 5055
rect 3846 5029 3890 5035
rect 3940 5059 3989 5071
rect 3940 5039 3958 5059
rect 3978 5039 3989 5059
rect 3940 5029 3989 5039
rect 1259 4823 1308 4833
rect 1259 4803 1270 4823
rect 1290 4803 1308 4823
rect 1259 4791 1308 4803
rect 1358 4827 1402 4833
rect 1358 4807 1373 4827
rect 1393 4807 1402 4827
rect 1358 4791 1402 4807
rect 1477 4823 1526 4833
rect 1477 4803 1488 4823
rect 1508 4803 1526 4823
rect 1477 4791 1526 4803
rect 1576 4827 1620 4833
rect 1576 4807 1591 4827
rect 1611 4807 1620 4827
rect 1576 4791 1620 4807
rect 1690 4827 1734 4833
rect 1690 4807 1699 4827
rect 1719 4807 1734 4827
rect 1690 4791 1734 4807
rect 1784 4823 1833 4833
rect 1784 4803 1802 4823
rect 1822 4803 1833 4823
rect 1784 4791 1833 4803
rect 2618 4831 2667 4843
rect 2618 4811 2629 4831
rect 2649 4811 2667 4831
rect 2618 4801 2667 4811
rect 2717 4827 2761 4843
rect 2717 4807 2732 4827
rect 2752 4807 2761 4827
rect 2717 4801 2761 4807
rect 2831 4827 2875 4843
rect 2831 4807 2840 4827
rect 2860 4807 2875 4827
rect 2831 4801 2875 4807
rect 2925 4831 2974 4843
rect 2925 4811 2943 4831
rect 2963 4811 2974 4831
rect 2925 4801 2974 4811
rect 3049 4827 3093 4843
rect 3049 4807 3058 4827
rect 3078 4807 3093 4827
rect 3049 4801 3093 4807
rect 3143 4831 3192 4843
rect 3143 4811 3161 4831
rect 3181 4811 3192 4831
rect 3143 4801 3192 4811
rect 3416 4647 3465 4659
rect 3416 4627 3427 4647
rect 3447 4627 3465 4647
rect 362 4597 411 4607
rect 362 4577 373 4597
rect 393 4577 411 4597
rect 362 4565 411 4577
rect 461 4601 505 4607
rect 461 4581 476 4601
rect 496 4581 505 4601
rect 461 4565 505 4581
rect 580 4597 629 4607
rect 580 4577 591 4597
rect 611 4577 629 4597
rect 580 4565 629 4577
rect 679 4601 723 4607
rect 679 4581 694 4601
rect 714 4581 723 4601
rect 679 4565 723 4581
rect 793 4601 837 4607
rect 793 4581 802 4601
rect 822 4581 837 4601
rect 793 4565 837 4581
rect 887 4597 936 4607
rect 3416 4617 3465 4627
rect 3515 4643 3559 4659
rect 3515 4623 3530 4643
rect 3550 4623 3559 4643
rect 3515 4617 3559 4623
rect 3629 4643 3673 4659
rect 3629 4623 3638 4643
rect 3658 4623 3673 4643
rect 3629 4617 3673 4623
rect 3723 4647 3772 4659
rect 3723 4627 3741 4647
rect 3761 4627 3772 4647
rect 3723 4617 3772 4627
rect 3847 4643 3891 4659
rect 3847 4623 3856 4643
rect 3876 4623 3891 4643
rect 3847 4617 3891 4623
rect 3941 4647 3990 4659
rect 3941 4627 3959 4647
rect 3979 4627 3990 4647
rect 3941 4617 3990 4627
rect 887 4577 905 4597
rect 925 4577 936 4597
rect 887 4565 936 4577
rect 2314 4425 2363 4437
rect 1160 4413 1209 4423
rect 1160 4393 1171 4413
rect 1191 4393 1209 4413
rect 1160 4381 1209 4393
rect 1259 4417 1303 4423
rect 1259 4397 1274 4417
rect 1294 4397 1303 4417
rect 1259 4381 1303 4397
rect 1378 4413 1427 4423
rect 1378 4393 1389 4413
rect 1409 4393 1427 4413
rect 1378 4381 1427 4393
rect 1477 4417 1521 4423
rect 1477 4397 1492 4417
rect 1512 4397 1521 4417
rect 1477 4381 1521 4397
rect 1591 4417 1635 4423
rect 1591 4397 1600 4417
rect 1620 4397 1635 4417
rect 1591 4381 1635 4397
rect 1685 4413 1734 4423
rect 1685 4393 1703 4413
rect 1723 4393 1734 4413
rect 2314 4405 2325 4425
rect 2345 4405 2363 4425
rect 2314 4395 2363 4405
rect 2413 4421 2457 4437
rect 2413 4401 2428 4421
rect 2448 4401 2457 4421
rect 2413 4395 2457 4401
rect 2527 4421 2571 4437
rect 2527 4401 2536 4421
rect 2556 4401 2571 4421
rect 2527 4395 2571 4401
rect 2621 4425 2670 4437
rect 2621 4405 2639 4425
rect 2659 4405 2670 4425
rect 2621 4395 2670 4405
rect 2745 4421 2789 4437
rect 2745 4401 2754 4421
rect 2774 4401 2789 4421
rect 2745 4395 2789 4401
rect 2839 4425 2888 4437
rect 2839 4405 2857 4425
rect 2877 4405 2888 4425
rect 2839 4395 2888 4405
rect 1685 4381 1734 4393
rect 363 4185 412 4195
rect 363 4165 374 4185
rect 394 4165 412 4185
rect 363 4153 412 4165
rect 462 4189 506 4195
rect 462 4169 477 4189
rect 497 4169 506 4189
rect 462 4153 506 4169
rect 581 4185 630 4195
rect 581 4165 592 4185
rect 612 4165 630 4185
rect 581 4153 630 4165
rect 680 4189 724 4195
rect 680 4169 695 4189
rect 715 4169 724 4189
rect 680 4153 724 4169
rect 794 4189 838 4195
rect 794 4169 803 4189
rect 823 4169 838 4189
rect 794 4153 838 4169
rect 888 4185 937 4195
rect 888 4165 906 4185
rect 926 4165 937 4185
rect 888 4153 937 4165
rect 3396 4041 3445 4053
rect 3396 4021 3407 4041
rect 3427 4021 3445 4041
rect 3396 4011 3445 4021
rect 3495 4037 3539 4053
rect 3495 4017 3510 4037
rect 3530 4017 3539 4037
rect 3495 4011 3539 4017
rect 3609 4037 3653 4053
rect 3609 4017 3618 4037
rect 3638 4017 3653 4037
rect 3609 4011 3653 4017
rect 3703 4041 3752 4053
rect 3703 4021 3721 4041
rect 3741 4021 3752 4041
rect 3703 4011 3752 4021
rect 3827 4037 3871 4053
rect 3827 4017 3836 4037
rect 3856 4017 3871 4037
rect 3827 4011 3871 4017
rect 3921 4041 3970 4053
rect 3921 4021 3939 4041
rect 3959 4021 3970 4041
rect 3921 4011 3970 4021
rect 2599 3813 2648 3825
rect 1445 3801 1494 3811
rect 1445 3781 1456 3801
rect 1476 3781 1494 3801
rect 1445 3769 1494 3781
rect 1544 3805 1588 3811
rect 1544 3785 1559 3805
rect 1579 3785 1588 3805
rect 1544 3769 1588 3785
rect 1663 3801 1712 3811
rect 1663 3781 1674 3801
rect 1694 3781 1712 3801
rect 1663 3769 1712 3781
rect 1762 3805 1806 3811
rect 1762 3785 1777 3805
rect 1797 3785 1806 3805
rect 1762 3769 1806 3785
rect 1876 3805 1920 3811
rect 1876 3785 1885 3805
rect 1905 3785 1920 3805
rect 1876 3769 1920 3785
rect 1970 3801 2019 3811
rect 1970 3781 1988 3801
rect 2008 3781 2019 3801
rect 2599 3793 2610 3813
rect 2630 3793 2648 3813
rect 2599 3783 2648 3793
rect 2698 3809 2742 3825
rect 2698 3789 2713 3809
rect 2733 3789 2742 3809
rect 2698 3783 2742 3789
rect 2812 3809 2856 3825
rect 2812 3789 2821 3809
rect 2841 3789 2856 3809
rect 2812 3783 2856 3789
rect 2906 3813 2955 3825
rect 2906 3793 2924 3813
rect 2944 3793 2955 3813
rect 2906 3783 2955 3793
rect 3030 3809 3074 3825
rect 3030 3789 3039 3809
rect 3059 3789 3074 3809
rect 3030 3783 3074 3789
rect 3124 3813 3173 3825
rect 3124 3793 3142 3813
rect 3162 3793 3173 3813
rect 3124 3783 3173 3793
rect 1970 3769 2019 3781
rect 3397 3629 3446 3641
rect 3397 3609 3408 3629
rect 3428 3609 3446 3629
rect 343 3579 392 3589
rect 343 3559 354 3579
rect 374 3559 392 3579
rect 343 3547 392 3559
rect 442 3583 486 3589
rect 442 3563 457 3583
rect 477 3563 486 3583
rect 442 3547 486 3563
rect 561 3579 610 3589
rect 561 3559 572 3579
rect 592 3559 610 3579
rect 561 3547 610 3559
rect 660 3583 704 3589
rect 660 3563 675 3583
rect 695 3563 704 3583
rect 660 3547 704 3563
rect 774 3583 818 3589
rect 774 3563 783 3583
rect 803 3563 818 3583
rect 774 3547 818 3563
rect 868 3579 917 3589
rect 3397 3599 3446 3609
rect 3496 3625 3540 3641
rect 3496 3605 3511 3625
rect 3531 3605 3540 3625
rect 3496 3599 3540 3605
rect 3610 3625 3654 3641
rect 3610 3605 3619 3625
rect 3639 3605 3654 3625
rect 3610 3599 3654 3605
rect 3704 3629 3753 3641
rect 3704 3609 3722 3629
rect 3742 3609 3753 3629
rect 3704 3599 3753 3609
rect 3828 3625 3872 3641
rect 3828 3605 3837 3625
rect 3857 3605 3872 3625
rect 3828 3599 3872 3605
rect 3922 3629 3971 3641
rect 3922 3609 3940 3629
rect 3960 3609 3971 3629
rect 3922 3599 3971 3609
rect 868 3559 886 3579
rect 906 3559 917 3579
rect 868 3547 917 3559
rect 1141 3395 1190 3405
rect 1141 3375 1152 3395
rect 1172 3375 1190 3395
rect 1141 3363 1190 3375
rect 1240 3399 1284 3405
rect 1240 3379 1255 3399
rect 1275 3379 1284 3399
rect 1240 3363 1284 3379
rect 1359 3395 1408 3405
rect 1359 3375 1370 3395
rect 1390 3375 1408 3395
rect 1359 3363 1408 3375
rect 1458 3399 1502 3405
rect 1458 3379 1473 3399
rect 1493 3379 1502 3399
rect 1458 3363 1502 3379
rect 1572 3399 1616 3405
rect 1572 3379 1581 3399
rect 1601 3379 1616 3399
rect 1572 3363 1616 3379
rect 1666 3395 1715 3405
rect 1666 3375 1684 3395
rect 1704 3375 1715 3395
rect 1666 3363 1715 3375
rect 2500 3403 2549 3415
rect 2500 3383 2511 3403
rect 2531 3383 2549 3403
rect 2500 3373 2549 3383
rect 2599 3399 2643 3415
rect 2599 3379 2614 3399
rect 2634 3379 2643 3399
rect 2599 3373 2643 3379
rect 2713 3399 2757 3415
rect 2713 3379 2722 3399
rect 2742 3379 2757 3399
rect 2713 3373 2757 3379
rect 2807 3403 2856 3415
rect 2807 3383 2825 3403
rect 2845 3383 2856 3403
rect 2807 3373 2856 3383
rect 2931 3399 2975 3415
rect 2931 3379 2940 3399
rect 2960 3379 2975 3399
rect 2931 3373 2975 3379
rect 3025 3403 3074 3415
rect 3025 3383 3043 3403
rect 3063 3383 3074 3403
rect 3025 3373 3074 3383
rect 344 3167 393 3177
rect 344 3147 355 3167
rect 375 3147 393 3167
rect 344 3135 393 3147
rect 443 3171 487 3177
rect 443 3151 458 3171
rect 478 3151 487 3171
rect 443 3135 487 3151
rect 562 3167 611 3177
rect 562 3147 573 3167
rect 593 3147 611 3167
rect 562 3135 611 3147
rect 661 3171 705 3177
rect 661 3151 676 3171
rect 696 3151 705 3171
rect 661 3135 705 3151
rect 775 3171 819 3177
rect 775 3151 784 3171
rect 804 3151 819 3171
rect 775 3135 819 3151
rect 869 3167 918 3177
rect 869 3147 887 3167
rect 907 3147 918 3167
rect 869 3135 918 3147
rect 3379 3023 3428 3035
rect 3379 3003 3390 3023
rect 3410 3003 3428 3023
rect 3379 2993 3428 3003
rect 3478 3019 3522 3035
rect 3478 2999 3493 3019
rect 3513 2999 3522 3019
rect 3478 2993 3522 2999
rect 3592 3019 3636 3035
rect 3592 2999 3601 3019
rect 3621 2999 3636 3019
rect 3592 2993 3636 2999
rect 3686 3023 3735 3035
rect 3686 3003 3704 3023
rect 3724 3003 3735 3023
rect 3686 2993 3735 3003
rect 3810 3019 3854 3035
rect 3810 2999 3819 3019
rect 3839 2999 3854 3019
rect 3810 2993 3854 2999
rect 3904 3023 3953 3035
rect 3904 3003 3922 3023
rect 3942 3003 3953 3023
rect 3904 2993 3953 3003
rect 1223 2787 1272 2797
rect 1223 2767 1234 2787
rect 1254 2767 1272 2787
rect 1223 2755 1272 2767
rect 1322 2791 1366 2797
rect 1322 2771 1337 2791
rect 1357 2771 1366 2791
rect 1322 2755 1366 2771
rect 1441 2787 1490 2797
rect 1441 2767 1452 2787
rect 1472 2767 1490 2787
rect 1441 2755 1490 2767
rect 1540 2791 1584 2797
rect 1540 2771 1555 2791
rect 1575 2771 1584 2791
rect 1540 2755 1584 2771
rect 1654 2791 1698 2797
rect 1654 2771 1663 2791
rect 1683 2771 1698 2791
rect 1654 2755 1698 2771
rect 1748 2787 1797 2797
rect 1748 2767 1766 2787
rect 1786 2767 1797 2787
rect 1748 2755 1797 2767
rect 2582 2795 2631 2807
rect 2582 2775 2593 2795
rect 2613 2775 2631 2795
rect 2582 2765 2631 2775
rect 2681 2791 2725 2807
rect 2681 2771 2696 2791
rect 2716 2771 2725 2791
rect 2681 2765 2725 2771
rect 2795 2791 2839 2807
rect 2795 2771 2804 2791
rect 2824 2771 2839 2791
rect 2795 2765 2839 2771
rect 2889 2795 2938 2807
rect 2889 2775 2907 2795
rect 2927 2775 2938 2795
rect 2889 2765 2938 2775
rect 3013 2791 3057 2807
rect 3013 2771 3022 2791
rect 3042 2771 3057 2791
rect 3013 2765 3057 2771
rect 3107 2795 3156 2807
rect 3107 2775 3125 2795
rect 3145 2775 3156 2795
rect 3107 2765 3156 2775
rect 3380 2611 3429 2623
rect 3380 2591 3391 2611
rect 3411 2591 3429 2611
rect 326 2561 375 2571
rect 326 2541 337 2561
rect 357 2541 375 2561
rect 326 2529 375 2541
rect 425 2565 469 2571
rect 425 2545 440 2565
rect 460 2545 469 2565
rect 425 2529 469 2545
rect 544 2561 593 2571
rect 544 2541 555 2561
rect 575 2541 593 2561
rect 544 2529 593 2541
rect 643 2565 687 2571
rect 643 2545 658 2565
rect 678 2545 687 2565
rect 643 2529 687 2545
rect 757 2565 801 2571
rect 757 2545 766 2565
rect 786 2545 801 2565
rect 757 2529 801 2545
rect 851 2561 900 2571
rect 3380 2581 3429 2591
rect 3479 2607 3523 2623
rect 3479 2587 3494 2607
rect 3514 2587 3523 2607
rect 3479 2581 3523 2587
rect 3593 2607 3637 2623
rect 3593 2587 3602 2607
rect 3622 2587 3637 2607
rect 3593 2581 3637 2587
rect 3687 2611 3736 2623
rect 3687 2591 3705 2611
rect 3725 2591 3736 2611
rect 3687 2581 3736 2591
rect 3811 2607 3855 2623
rect 3811 2587 3820 2607
rect 3840 2587 3855 2607
rect 3811 2581 3855 2587
rect 3905 2611 3954 2623
rect 3905 2591 3923 2611
rect 3943 2591 3954 2611
rect 3905 2581 3954 2591
rect 851 2541 869 2561
rect 889 2541 900 2561
rect 851 2529 900 2541
rect 2417 2387 2466 2399
rect 1124 2377 1173 2387
rect 1124 2357 1135 2377
rect 1155 2357 1173 2377
rect 1124 2345 1173 2357
rect 1223 2381 1267 2387
rect 1223 2361 1238 2381
rect 1258 2361 1267 2381
rect 1223 2345 1267 2361
rect 1342 2377 1391 2387
rect 1342 2357 1353 2377
rect 1373 2357 1391 2377
rect 1342 2345 1391 2357
rect 1441 2381 1485 2387
rect 1441 2361 1456 2381
rect 1476 2361 1485 2381
rect 1441 2345 1485 2361
rect 1555 2381 1599 2387
rect 1555 2361 1564 2381
rect 1584 2361 1599 2381
rect 1555 2345 1599 2361
rect 1649 2377 1698 2387
rect 1649 2357 1667 2377
rect 1687 2357 1698 2377
rect 2417 2367 2428 2387
rect 2448 2367 2466 2387
rect 2417 2357 2466 2367
rect 2516 2383 2560 2399
rect 2516 2363 2531 2383
rect 2551 2363 2560 2383
rect 2516 2357 2560 2363
rect 2630 2383 2674 2399
rect 2630 2363 2639 2383
rect 2659 2363 2674 2383
rect 2630 2357 2674 2363
rect 2724 2387 2773 2399
rect 2724 2367 2742 2387
rect 2762 2367 2773 2387
rect 2724 2357 2773 2367
rect 2848 2383 2892 2399
rect 2848 2363 2857 2383
rect 2877 2363 2892 2383
rect 2848 2357 2892 2363
rect 2942 2387 2991 2399
rect 2942 2367 2960 2387
rect 2980 2367 2991 2387
rect 2942 2357 2991 2367
rect 1649 2345 1698 2357
rect 327 2149 376 2159
rect 327 2129 338 2149
rect 358 2129 376 2149
rect 327 2117 376 2129
rect 426 2153 470 2159
rect 426 2133 441 2153
rect 461 2133 470 2153
rect 426 2117 470 2133
rect 545 2149 594 2159
rect 545 2129 556 2149
rect 576 2129 594 2149
rect 545 2117 594 2129
rect 644 2153 688 2159
rect 644 2133 659 2153
rect 679 2133 688 2153
rect 644 2117 688 2133
rect 758 2153 802 2159
rect 758 2133 767 2153
rect 787 2133 802 2153
rect 758 2117 802 2133
rect 852 2149 901 2159
rect 852 2129 870 2149
rect 890 2129 901 2149
rect 852 2117 901 2129
rect 3359 2005 3408 2017
rect 3359 1985 3370 2005
rect 3390 1985 3408 2005
rect 3359 1975 3408 1985
rect 3458 2001 3502 2017
rect 3458 1981 3473 2001
rect 3493 1981 3502 2001
rect 3458 1975 3502 1981
rect 3572 2001 3616 2017
rect 3572 1981 3581 2001
rect 3601 1981 3616 2001
rect 3572 1975 3616 1981
rect 3666 2005 3715 2017
rect 3666 1985 3684 2005
rect 3704 1985 3715 2005
rect 3666 1975 3715 1985
rect 3790 2001 3834 2017
rect 3790 1981 3799 2001
rect 3819 1981 3834 2001
rect 3790 1975 3834 1981
rect 3884 2005 3933 2017
rect 3884 1985 3902 2005
rect 3922 1985 3933 2005
rect 3884 1975 3933 1985
rect 2562 1777 2611 1789
rect 1269 1767 1318 1777
rect 1269 1747 1280 1767
rect 1300 1747 1318 1767
rect 1269 1735 1318 1747
rect 1368 1771 1412 1777
rect 1368 1751 1383 1771
rect 1403 1751 1412 1771
rect 1368 1735 1412 1751
rect 1487 1767 1536 1777
rect 1487 1747 1498 1767
rect 1518 1747 1536 1767
rect 1487 1735 1536 1747
rect 1586 1771 1630 1777
rect 1586 1751 1601 1771
rect 1621 1751 1630 1771
rect 1586 1735 1630 1751
rect 1700 1771 1744 1777
rect 1700 1751 1709 1771
rect 1729 1751 1744 1771
rect 1700 1735 1744 1751
rect 1794 1767 1843 1777
rect 1794 1747 1812 1767
rect 1832 1747 1843 1767
rect 2562 1757 2573 1777
rect 2593 1757 2611 1777
rect 2562 1747 2611 1757
rect 2661 1773 2705 1789
rect 2661 1753 2676 1773
rect 2696 1753 2705 1773
rect 2661 1747 2705 1753
rect 2775 1773 2819 1789
rect 2775 1753 2784 1773
rect 2804 1753 2819 1773
rect 2775 1747 2819 1753
rect 2869 1777 2918 1789
rect 2869 1757 2887 1777
rect 2907 1757 2918 1777
rect 2869 1747 2918 1757
rect 2993 1773 3037 1789
rect 2993 1753 3002 1773
rect 3022 1753 3037 1773
rect 2993 1747 3037 1753
rect 3087 1777 3136 1789
rect 3087 1757 3105 1777
rect 3125 1757 3136 1777
rect 3087 1747 3136 1757
rect 1794 1735 1843 1747
rect 3360 1593 3409 1605
rect 3360 1573 3371 1593
rect 3391 1573 3409 1593
rect 306 1543 355 1553
rect 306 1523 317 1543
rect 337 1523 355 1543
rect 306 1511 355 1523
rect 405 1547 449 1553
rect 405 1527 420 1547
rect 440 1527 449 1547
rect 405 1511 449 1527
rect 524 1543 573 1553
rect 524 1523 535 1543
rect 555 1523 573 1543
rect 524 1511 573 1523
rect 623 1547 667 1553
rect 623 1527 638 1547
rect 658 1527 667 1547
rect 623 1511 667 1527
rect 737 1547 781 1553
rect 737 1527 746 1547
rect 766 1527 781 1547
rect 737 1511 781 1527
rect 831 1543 880 1553
rect 3360 1563 3409 1573
rect 3459 1589 3503 1605
rect 3459 1569 3474 1589
rect 3494 1569 3503 1589
rect 3459 1563 3503 1569
rect 3573 1589 3617 1605
rect 3573 1569 3582 1589
rect 3602 1569 3617 1589
rect 3573 1563 3617 1569
rect 3667 1593 3716 1605
rect 3667 1573 3685 1593
rect 3705 1573 3716 1593
rect 3667 1563 3716 1573
rect 3791 1589 3835 1605
rect 3791 1569 3800 1589
rect 3820 1569 3835 1589
rect 3791 1563 3835 1569
rect 3885 1593 3934 1605
rect 3885 1573 3903 1593
rect 3923 1573 3934 1593
rect 3885 1563 3934 1573
rect 831 1523 849 1543
rect 869 1523 880 1543
rect 831 1511 880 1523
rect 1104 1359 1153 1369
rect 1104 1339 1115 1359
rect 1135 1339 1153 1359
rect 1104 1327 1153 1339
rect 1203 1363 1247 1369
rect 1203 1343 1218 1363
rect 1238 1343 1247 1363
rect 1203 1327 1247 1343
rect 1322 1359 1371 1369
rect 1322 1339 1333 1359
rect 1353 1339 1371 1359
rect 1322 1327 1371 1339
rect 1421 1363 1465 1369
rect 1421 1343 1436 1363
rect 1456 1343 1465 1363
rect 1421 1327 1465 1343
rect 1535 1363 1579 1369
rect 1535 1343 1544 1363
rect 1564 1343 1579 1363
rect 1535 1327 1579 1343
rect 1629 1359 1678 1369
rect 1629 1339 1647 1359
rect 1667 1339 1678 1359
rect 1629 1327 1678 1339
rect 2463 1367 2512 1379
rect 2463 1347 2474 1367
rect 2494 1347 2512 1367
rect 2463 1337 2512 1347
rect 2562 1363 2606 1379
rect 2562 1343 2577 1363
rect 2597 1343 2606 1363
rect 2562 1337 2606 1343
rect 2676 1363 2720 1379
rect 2676 1343 2685 1363
rect 2705 1343 2720 1363
rect 2676 1337 2720 1343
rect 2770 1367 2819 1379
rect 2770 1347 2788 1367
rect 2808 1347 2819 1367
rect 2770 1337 2819 1347
rect 2894 1363 2938 1379
rect 2894 1343 2903 1363
rect 2923 1343 2938 1363
rect 2894 1337 2938 1343
rect 2988 1367 3037 1379
rect 2988 1347 3006 1367
rect 3026 1347 3037 1367
rect 2988 1337 3037 1347
rect 307 1131 356 1141
rect 307 1111 318 1131
rect 338 1111 356 1131
rect 307 1099 356 1111
rect 406 1135 450 1141
rect 406 1115 421 1135
rect 441 1115 450 1135
rect 406 1099 450 1115
rect 525 1131 574 1141
rect 525 1111 536 1131
rect 556 1111 574 1131
rect 525 1099 574 1111
rect 624 1135 668 1141
rect 624 1115 639 1135
rect 659 1115 668 1135
rect 624 1099 668 1115
rect 738 1135 782 1141
rect 738 1115 747 1135
rect 767 1115 782 1135
rect 738 1099 782 1115
rect 832 1131 881 1141
rect 832 1111 850 1131
rect 870 1111 881 1131
rect 832 1099 881 1111
rect 3342 987 3391 999
rect 3342 967 3353 987
rect 3373 967 3391 987
rect 3342 957 3391 967
rect 3441 983 3485 999
rect 3441 963 3456 983
rect 3476 963 3485 983
rect 3441 957 3485 963
rect 3555 983 3599 999
rect 3555 963 3564 983
rect 3584 963 3599 983
rect 3555 957 3599 963
rect 3649 987 3698 999
rect 3649 967 3667 987
rect 3687 967 3698 987
rect 3649 957 3698 967
rect 3773 983 3817 999
rect 3773 963 3782 983
rect 3802 963 3817 983
rect 3773 957 3817 963
rect 3867 987 3916 999
rect 3867 967 3885 987
rect 3905 967 3916 987
rect 3867 957 3916 967
rect 1186 751 1235 761
rect 1186 731 1197 751
rect 1217 731 1235 751
rect 1186 719 1235 731
rect 1285 755 1329 761
rect 1285 735 1300 755
rect 1320 735 1329 755
rect 1285 719 1329 735
rect 1404 751 1453 761
rect 1404 731 1415 751
rect 1435 731 1453 751
rect 1404 719 1453 731
rect 1503 755 1547 761
rect 1503 735 1518 755
rect 1538 735 1547 755
rect 1503 719 1547 735
rect 1617 755 1661 761
rect 1617 735 1626 755
rect 1646 735 1661 755
rect 1617 719 1661 735
rect 1711 751 1760 761
rect 1711 731 1729 751
rect 1749 731 1760 751
rect 1711 719 1760 731
rect 2545 759 2594 771
rect 2545 739 2556 759
rect 2576 739 2594 759
rect 2545 729 2594 739
rect 2644 755 2688 771
rect 2644 735 2659 755
rect 2679 735 2688 755
rect 2644 729 2688 735
rect 2758 755 2802 771
rect 2758 735 2767 755
rect 2787 735 2802 755
rect 2758 729 2802 735
rect 2852 759 2901 771
rect 2852 739 2870 759
rect 2890 739 2901 759
rect 2852 729 2901 739
rect 2976 755 3020 771
rect 2976 735 2985 755
rect 3005 735 3020 755
rect 2976 729 3020 735
rect 3070 759 3119 771
rect 3070 739 3088 759
rect 3108 739 3119 759
rect 3070 729 3119 739
rect 3343 575 3392 587
rect 3343 555 3354 575
rect 3374 555 3392 575
rect 289 525 338 535
rect 289 505 300 525
rect 320 505 338 525
rect 289 493 338 505
rect 388 529 432 535
rect 388 509 403 529
rect 423 509 432 529
rect 388 493 432 509
rect 507 525 556 535
rect 507 505 518 525
rect 538 505 556 525
rect 507 493 556 505
rect 606 529 650 535
rect 606 509 621 529
rect 641 509 650 529
rect 606 493 650 509
rect 720 529 764 535
rect 720 509 729 529
rect 749 509 764 529
rect 720 493 764 509
rect 814 525 863 535
rect 3343 545 3392 555
rect 3442 571 3486 587
rect 3442 551 3457 571
rect 3477 551 3486 571
rect 3442 545 3486 551
rect 3556 571 3600 587
rect 3556 551 3565 571
rect 3585 551 3600 571
rect 3556 545 3600 551
rect 3650 575 3699 587
rect 3650 555 3668 575
rect 3688 555 3699 575
rect 3650 545 3699 555
rect 3774 571 3818 587
rect 3774 551 3783 571
rect 3803 551 3818 571
rect 3774 545 3818 551
rect 3868 575 3917 587
rect 3868 555 3886 575
rect 3906 555 3917 575
rect 3868 545 3917 555
rect 814 505 832 525
rect 852 505 863 525
rect 814 493 863 505
rect 1087 341 1136 351
rect 1087 321 1098 341
rect 1118 321 1136 341
rect 1087 309 1136 321
rect 1186 345 1230 351
rect 1186 325 1201 345
rect 1221 325 1230 345
rect 1186 309 1230 325
rect 1305 341 1354 351
rect 1305 321 1316 341
rect 1336 321 1354 341
rect 1305 309 1354 321
rect 1404 345 1448 351
rect 1404 325 1419 345
rect 1439 325 1448 345
rect 1404 309 1448 325
rect 1518 345 1562 351
rect 1518 325 1527 345
rect 1547 325 1562 345
rect 1518 309 1562 325
rect 1612 341 1661 351
rect 1612 321 1630 341
rect 1650 321 1661 341
rect 1612 309 1661 321
rect 290 113 339 123
rect 290 93 301 113
rect 321 93 339 113
rect 290 81 339 93
rect 389 117 433 123
rect 389 97 404 117
rect 424 97 433 117
rect 389 81 433 97
rect 508 113 557 123
rect 508 93 519 113
rect 539 93 557 113
rect 508 81 557 93
rect 607 117 651 123
rect 607 97 622 117
rect 642 97 651 117
rect 607 81 651 97
rect 721 117 765 123
rect 721 97 730 117
rect 750 97 765 117
rect 721 81 765 97
rect 815 113 864 123
rect 815 93 833 113
rect 853 93 864 113
rect 815 81 864 93
rect 1503 -463 1552 -453
rect 1503 -483 1514 -463
rect 1534 -483 1552 -463
rect 1503 -495 1552 -483
rect 1602 -459 1646 -453
rect 1602 -479 1617 -459
rect 1637 -479 1646 -459
rect 1602 -495 1646 -479
rect 1721 -463 1770 -453
rect 1721 -483 1732 -463
rect 1752 -483 1770 -463
rect 1721 -495 1770 -483
rect 1820 -459 1864 -453
rect 1820 -479 1835 -459
rect 1855 -479 1864 -459
rect 1820 -495 1864 -479
rect 1934 -459 1978 -453
rect 1934 -479 1943 -459
rect 1963 -479 1978 -459
rect 1934 -495 1978 -479
rect 2028 -463 2077 -453
rect 2028 -483 2046 -463
rect 2066 -483 2077 -463
rect 2028 -495 2077 -483
<< pdiff >>
rect 3474 7964 3518 8006
rect 3474 7944 3486 7964
rect 3506 7944 3518 7964
rect 3474 7937 3518 7944
rect 3473 7906 3518 7937
rect 3568 7964 3610 8006
rect 3568 7944 3582 7964
rect 3602 7944 3610 7964
rect 3568 7906 3610 7944
rect 3684 7964 3726 8006
rect 3684 7944 3692 7964
rect 3712 7944 3726 7964
rect 3684 7906 3726 7944
rect 3776 7964 3820 8006
rect 3776 7944 3788 7964
rect 3808 7944 3820 7964
rect 3776 7906 3820 7944
rect 3902 7964 3944 8006
rect 3902 7944 3910 7964
rect 3930 7944 3944 7964
rect 3902 7906 3944 7944
rect 3994 7964 4038 8006
rect 3994 7944 4006 7964
rect 4026 7944 4038 7964
rect 3994 7906 4038 7944
rect 421 7800 465 7838
rect 421 7780 433 7800
rect 453 7780 465 7800
rect 421 7738 465 7780
rect 515 7800 557 7838
rect 515 7780 529 7800
rect 549 7780 557 7800
rect 515 7738 557 7780
rect 639 7800 683 7838
rect 639 7780 651 7800
rect 671 7780 683 7800
rect 639 7738 683 7780
rect 733 7800 775 7838
rect 733 7780 747 7800
rect 767 7780 775 7800
rect 733 7738 775 7780
rect 849 7800 891 7838
rect 849 7780 857 7800
rect 877 7780 891 7800
rect 849 7738 891 7780
rect 941 7807 986 7838
rect 941 7800 985 7807
rect 941 7780 953 7800
rect 973 7780 985 7800
rect 941 7738 985 7780
rect 2677 7736 2721 7778
rect 2677 7716 2689 7736
rect 2709 7716 2721 7736
rect 2677 7709 2721 7716
rect 2676 7678 2721 7709
rect 2771 7736 2813 7778
rect 2771 7716 2785 7736
rect 2805 7716 2813 7736
rect 2771 7678 2813 7716
rect 2887 7736 2929 7778
rect 2887 7716 2895 7736
rect 2915 7716 2929 7736
rect 2887 7678 2929 7716
rect 2979 7736 3023 7778
rect 2979 7716 2991 7736
rect 3011 7716 3023 7736
rect 2979 7678 3023 7716
rect 3105 7736 3147 7778
rect 3105 7716 3113 7736
rect 3133 7716 3147 7736
rect 3105 7678 3147 7716
rect 3197 7736 3241 7778
rect 3197 7716 3209 7736
rect 3229 7716 3241 7736
rect 3197 7678 3241 7716
rect 1219 7616 1263 7654
rect 1219 7596 1231 7616
rect 1251 7596 1263 7616
rect 1219 7554 1263 7596
rect 1313 7616 1355 7654
rect 1313 7596 1327 7616
rect 1347 7596 1355 7616
rect 1313 7554 1355 7596
rect 1437 7616 1481 7654
rect 1437 7596 1449 7616
rect 1469 7596 1481 7616
rect 1437 7554 1481 7596
rect 1531 7616 1573 7654
rect 1531 7596 1545 7616
rect 1565 7596 1573 7616
rect 1531 7554 1573 7596
rect 1647 7616 1689 7654
rect 1647 7596 1655 7616
rect 1675 7596 1689 7616
rect 1647 7554 1689 7596
rect 1739 7623 1784 7654
rect 1739 7616 1783 7623
rect 1739 7596 1751 7616
rect 1771 7596 1783 7616
rect 1739 7554 1783 7596
rect 3475 7552 3519 7594
rect 3475 7532 3487 7552
rect 3507 7532 3519 7552
rect 3475 7525 3519 7532
rect 3474 7494 3519 7525
rect 3569 7552 3611 7594
rect 3569 7532 3583 7552
rect 3603 7532 3611 7552
rect 3569 7494 3611 7532
rect 3685 7552 3727 7594
rect 3685 7532 3693 7552
rect 3713 7532 3727 7552
rect 3685 7494 3727 7532
rect 3777 7552 3821 7594
rect 3777 7532 3789 7552
rect 3809 7532 3821 7552
rect 3777 7494 3821 7532
rect 3903 7552 3945 7594
rect 3903 7532 3911 7552
rect 3931 7532 3945 7552
rect 3903 7494 3945 7532
rect 3995 7552 4039 7594
rect 3995 7532 4007 7552
rect 4027 7532 4039 7552
rect 3995 7494 4039 7532
rect 422 7388 466 7426
rect 422 7368 434 7388
rect 454 7368 466 7388
rect 422 7326 466 7368
rect 516 7388 558 7426
rect 516 7368 530 7388
rect 550 7368 558 7388
rect 516 7326 558 7368
rect 640 7388 684 7426
rect 640 7368 652 7388
rect 672 7368 684 7388
rect 640 7326 684 7368
rect 734 7388 776 7426
rect 734 7368 748 7388
rect 768 7368 776 7388
rect 734 7326 776 7368
rect 850 7388 892 7426
rect 850 7368 858 7388
rect 878 7368 892 7388
rect 850 7326 892 7368
rect 942 7395 987 7426
rect 942 7388 986 7395
rect 942 7368 954 7388
rect 974 7368 986 7388
rect 942 7326 986 7368
rect 2578 7326 2622 7368
rect 2578 7306 2590 7326
rect 2610 7306 2622 7326
rect 2578 7299 2622 7306
rect 2577 7268 2622 7299
rect 2672 7326 2714 7368
rect 2672 7306 2686 7326
rect 2706 7306 2714 7326
rect 2672 7268 2714 7306
rect 2788 7326 2830 7368
rect 2788 7306 2796 7326
rect 2816 7306 2830 7326
rect 2788 7268 2830 7306
rect 2880 7326 2924 7368
rect 2880 7306 2892 7326
rect 2912 7306 2924 7326
rect 2880 7268 2924 7306
rect 3006 7326 3048 7368
rect 3006 7306 3014 7326
rect 3034 7306 3048 7326
rect 3006 7268 3048 7306
rect 3098 7326 3142 7368
rect 3098 7306 3110 7326
rect 3130 7306 3142 7326
rect 3098 7268 3142 7306
rect 1301 7008 1345 7046
rect 1301 6988 1313 7008
rect 1333 6988 1345 7008
rect 1301 6946 1345 6988
rect 1395 7008 1437 7046
rect 1395 6988 1409 7008
rect 1429 6988 1437 7008
rect 1395 6946 1437 6988
rect 1519 7008 1563 7046
rect 1519 6988 1531 7008
rect 1551 6988 1563 7008
rect 1519 6946 1563 6988
rect 1613 7008 1655 7046
rect 1613 6988 1627 7008
rect 1647 6988 1655 7008
rect 1613 6946 1655 6988
rect 1729 7008 1771 7046
rect 1729 6988 1737 7008
rect 1757 6988 1771 7008
rect 1729 6946 1771 6988
rect 1821 7015 1866 7046
rect 1821 7008 1865 7015
rect 1821 6988 1833 7008
rect 1853 6988 1865 7008
rect 1821 6946 1865 6988
rect 3457 6946 3501 6988
rect 3457 6926 3469 6946
rect 3489 6926 3501 6946
rect 3457 6919 3501 6926
rect 3456 6888 3501 6919
rect 3551 6946 3593 6988
rect 3551 6926 3565 6946
rect 3585 6926 3593 6946
rect 3551 6888 3593 6926
rect 3667 6946 3709 6988
rect 3667 6926 3675 6946
rect 3695 6926 3709 6946
rect 3667 6888 3709 6926
rect 3759 6946 3803 6988
rect 3759 6926 3771 6946
rect 3791 6926 3803 6946
rect 3759 6888 3803 6926
rect 3885 6946 3927 6988
rect 3885 6926 3893 6946
rect 3913 6926 3927 6946
rect 3885 6888 3927 6926
rect 3977 6946 4021 6988
rect 3977 6926 3989 6946
rect 4009 6926 4021 6946
rect 3977 6888 4021 6926
rect 404 6782 448 6820
rect 404 6762 416 6782
rect 436 6762 448 6782
rect 404 6720 448 6762
rect 498 6782 540 6820
rect 498 6762 512 6782
rect 532 6762 540 6782
rect 498 6720 540 6762
rect 622 6782 666 6820
rect 622 6762 634 6782
rect 654 6762 666 6782
rect 622 6720 666 6762
rect 716 6782 758 6820
rect 716 6762 730 6782
rect 750 6762 758 6782
rect 716 6720 758 6762
rect 832 6782 874 6820
rect 832 6762 840 6782
rect 860 6762 874 6782
rect 832 6720 874 6762
rect 924 6789 969 6820
rect 924 6782 968 6789
rect 924 6762 936 6782
rect 956 6762 968 6782
rect 924 6720 968 6762
rect 2660 6718 2704 6760
rect 2660 6698 2672 6718
rect 2692 6698 2704 6718
rect 2660 6691 2704 6698
rect 2659 6660 2704 6691
rect 2754 6718 2796 6760
rect 2754 6698 2768 6718
rect 2788 6698 2796 6718
rect 2754 6660 2796 6698
rect 2870 6718 2912 6760
rect 2870 6698 2878 6718
rect 2898 6698 2912 6718
rect 2870 6660 2912 6698
rect 2962 6718 3006 6760
rect 2962 6698 2974 6718
rect 2994 6698 3006 6718
rect 2962 6660 3006 6698
rect 3088 6718 3130 6760
rect 3088 6698 3096 6718
rect 3116 6698 3130 6718
rect 3088 6660 3130 6698
rect 3180 6718 3224 6760
rect 3180 6698 3192 6718
rect 3212 6698 3224 6718
rect 3180 6660 3224 6698
rect 1202 6598 1246 6636
rect 1202 6578 1214 6598
rect 1234 6578 1246 6598
rect 1202 6536 1246 6578
rect 1296 6598 1338 6636
rect 1296 6578 1310 6598
rect 1330 6578 1338 6598
rect 1296 6536 1338 6578
rect 1420 6598 1464 6636
rect 1420 6578 1432 6598
rect 1452 6578 1464 6598
rect 1420 6536 1464 6578
rect 1514 6598 1556 6636
rect 1514 6578 1528 6598
rect 1548 6578 1556 6598
rect 1514 6536 1556 6578
rect 1630 6598 1672 6636
rect 1630 6578 1638 6598
rect 1658 6578 1672 6598
rect 1630 6536 1672 6578
rect 1722 6605 1767 6636
rect 1722 6598 1766 6605
rect 1722 6578 1734 6598
rect 1754 6578 1766 6598
rect 1722 6536 1766 6578
rect 3458 6534 3502 6576
rect 3458 6514 3470 6534
rect 3490 6514 3502 6534
rect 3458 6507 3502 6514
rect 3457 6476 3502 6507
rect 3552 6534 3594 6576
rect 3552 6514 3566 6534
rect 3586 6514 3594 6534
rect 3552 6476 3594 6514
rect 3668 6534 3710 6576
rect 3668 6514 3676 6534
rect 3696 6514 3710 6534
rect 3668 6476 3710 6514
rect 3760 6534 3804 6576
rect 3760 6514 3772 6534
rect 3792 6514 3804 6534
rect 3760 6476 3804 6514
rect 3886 6534 3928 6576
rect 3886 6514 3894 6534
rect 3914 6514 3928 6534
rect 3886 6476 3928 6514
rect 3978 6534 4022 6576
rect 3978 6514 3990 6534
rect 4010 6514 4022 6534
rect 3978 6476 4022 6514
rect 405 6370 449 6408
rect 405 6350 417 6370
rect 437 6350 449 6370
rect 405 6308 449 6350
rect 499 6370 541 6408
rect 499 6350 513 6370
rect 533 6350 541 6370
rect 499 6308 541 6350
rect 623 6370 667 6408
rect 623 6350 635 6370
rect 655 6350 667 6370
rect 623 6308 667 6350
rect 717 6370 759 6408
rect 717 6350 731 6370
rect 751 6350 759 6370
rect 717 6308 759 6350
rect 833 6370 875 6408
rect 833 6350 841 6370
rect 861 6350 875 6370
rect 833 6308 875 6350
rect 925 6377 970 6408
rect 925 6370 969 6377
rect 925 6350 937 6370
rect 957 6350 969 6370
rect 925 6308 969 6350
rect 2495 6310 2539 6352
rect 2495 6290 2507 6310
rect 2527 6290 2539 6310
rect 2495 6283 2539 6290
rect 2494 6252 2539 6283
rect 2589 6310 2631 6352
rect 2589 6290 2603 6310
rect 2623 6290 2631 6310
rect 2589 6252 2631 6290
rect 2705 6310 2747 6352
rect 2705 6290 2713 6310
rect 2733 6290 2747 6310
rect 2705 6252 2747 6290
rect 2797 6310 2841 6352
rect 2797 6290 2809 6310
rect 2829 6290 2841 6310
rect 2797 6252 2841 6290
rect 2923 6310 2965 6352
rect 2923 6290 2931 6310
rect 2951 6290 2965 6310
rect 2923 6252 2965 6290
rect 3015 6310 3059 6352
rect 3015 6290 3027 6310
rect 3047 6290 3059 6310
rect 3015 6252 3059 6290
rect 1347 5988 1391 6026
rect 1347 5968 1359 5988
rect 1379 5968 1391 5988
rect 1347 5926 1391 5968
rect 1441 5988 1483 6026
rect 1441 5968 1455 5988
rect 1475 5968 1483 5988
rect 1441 5926 1483 5968
rect 1565 5988 1609 6026
rect 1565 5968 1577 5988
rect 1597 5968 1609 5988
rect 1565 5926 1609 5968
rect 1659 5988 1701 6026
rect 1659 5968 1673 5988
rect 1693 5968 1701 5988
rect 1659 5926 1701 5968
rect 1775 5988 1817 6026
rect 1775 5968 1783 5988
rect 1803 5968 1817 5988
rect 1775 5926 1817 5968
rect 1867 5995 1912 6026
rect 1867 5988 1911 5995
rect 1867 5968 1879 5988
rect 1899 5968 1911 5988
rect 1867 5926 1911 5968
rect 3437 5928 3481 5970
rect 3437 5908 3449 5928
rect 3469 5908 3481 5928
rect 3437 5901 3481 5908
rect 3436 5870 3481 5901
rect 3531 5928 3573 5970
rect 3531 5908 3545 5928
rect 3565 5908 3573 5928
rect 3531 5870 3573 5908
rect 3647 5928 3689 5970
rect 3647 5908 3655 5928
rect 3675 5908 3689 5928
rect 3647 5870 3689 5908
rect 3739 5928 3783 5970
rect 3739 5908 3751 5928
rect 3771 5908 3783 5928
rect 3739 5870 3783 5908
rect 3865 5928 3907 5970
rect 3865 5908 3873 5928
rect 3893 5908 3907 5928
rect 3865 5870 3907 5908
rect 3957 5928 4001 5970
rect 3957 5908 3969 5928
rect 3989 5908 4001 5928
rect 3957 5870 4001 5908
rect 384 5764 428 5802
rect 384 5744 396 5764
rect 416 5744 428 5764
rect 384 5702 428 5744
rect 478 5764 520 5802
rect 478 5744 492 5764
rect 512 5744 520 5764
rect 478 5702 520 5744
rect 602 5764 646 5802
rect 602 5744 614 5764
rect 634 5744 646 5764
rect 602 5702 646 5744
rect 696 5764 738 5802
rect 696 5744 710 5764
rect 730 5744 738 5764
rect 696 5702 738 5744
rect 812 5764 854 5802
rect 812 5744 820 5764
rect 840 5744 854 5764
rect 812 5702 854 5744
rect 904 5771 949 5802
rect 904 5764 948 5771
rect 904 5744 916 5764
rect 936 5744 948 5764
rect 904 5702 948 5744
rect 2640 5700 2684 5742
rect 2640 5680 2652 5700
rect 2672 5680 2684 5700
rect 2640 5673 2684 5680
rect 2639 5642 2684 5673
rect 2734 5700 2776 5742
rect 2734 5680 2748 5700
rect 2768 5680 2776 5700
rect 2734 5642 2776 5680
rect 2850 5700 2892 5742
rect 2850 5680 2858 5700
rect 2878 5680 2892 5700
rect 2850 5642 2892 5680
rect 2942 5700 2986 5742
rect 2942 5680 2954 5700
rect 2974 5680 2986 5700
rect 2942 5642 2986 5680
rect 3068 5700 3110 5742
rect 3068 5680 3076 5700
rect 3096 5680 3110 5700
rect 3068 5642 3110 5680
rect 3160 5700 3204 5742
rect 3160 5680 3172 5700
rect 3192 5680 3204 5700
rect 3160 5642 3204 5680
rect 1182 5580 1226 5618
rect 1182 5560 1194 5580
rect 1214 5560 1226 5580
rect 1182 5518 1226 5560
rect 1276 5580 1318 5618
rect 1276 5560 1290 5580
rect 1310 5560 1318 5580
rect 1276 5518 1318 5560
rect 1400 5580 1444 5618
rect 1400 5560 1412 5580
rect 1432 5560 1444 5580
rect 1400 5518 1444 5560
rect 1494 5580 1536 5618
rect 1494 5560 1508 5580
rect 1528 5560 1536 5580
rect 1494 5518 1536 5560
rect 1610 5580 1652 5618
rect 1610 5560 1618 5580
rect 1638 5560 1652 5580
rect 1610 5518 1652 5560
rect 1702 5587 1747 5618
rect 1702 5580 1746 5587
rect 1702 5560 1714 5580
rect 1734 5560 1746 5580
rect 1702 5518 1746 5560
rect 3438 5516 3482 5558
rect 3438 5496 3450 5516
rect 3470 5496 3482 5516
rect 3438 5489 3482 5496
rect 3437 5458 3482 5489
rect 3532 5516 3574 5558
rect 3532 5496 3546 5516
rect 3566 5496 3574 5516
rect 3532 5458 3574 5496
rect 3648 5516 3690 5558
rect 3648 5496 3656 5516
rect 3676 5496 3690 5516
rect 3648 5458 3690 5496
rect 3740 5516 3784 5558
rect 3740 5496 3752 5516
rect 3772 5496 3784 5516
rect 3740 5458 3784 5496
rect 3866 5516 3908 5558
rect 3866 5496 3874 5516
rect 3894 5496 3908 5516
rect 3866 5458 3908 5496
rect 3958 5516 4002 5558
rect 3958 5496 3970 5516
rect 3990 5496 4002 5516
rect 3958 5458 4002 5496
rect 385 5352 429 5390
rect 385 5332 397 5352
rect 417 5332 429 5352
rect 385 5290 429 5332
rect 479 5352 521 5390
rect 479 5332 493 5352
rect 513 5332 521 5352
rect 479 5290 521 5332
rect 603 5352 647 5390
rect 603 5332 615 5352
rect 635 5332 647 5352
rect 603 5290 647 5332
rect 697 5352 739 5390
rect 697 5332 711 5352
rect 731 5332 739 5352
rect 697 5290 739 5332
rect 813 5352 855 5390
rect 813 5332 821 5352
rect 841 5332 855 5352
rect 813 5290 855 5332
rect 905 5359 950 5390
rect 905 5352 949 5359
rect 905 5332 917 5352
rect 937 5332 949 5352
rect 905 5290 949 5332
rect 2541 5290 2585 5332
rect 2541 5270 2553 5290
rect 2573 5270 2585 5290
rect 2541 5263 2585 5270
rect 2540 5232 2585 5263
rect 2635 5290 2677 5332
rect 2635 5270 2649 5290
rect 2669 5270 2677 5290
rect 2635 5232 2677 5270
rect 2751 5290 2793 5332
rect 2751 5270 2759 5290
rect 2779 5270 2793 5290
rect 2751 5232 2793 5270
rect 2843 5290 2887 5332
rect 2843 5270 2855 5290
rect 2875 5270 2887 5290
rect 2843 5232 2887 5270
rect 2969 5290 3011 5332
rect 2969 5270 2977 5290
rect 2997 5270 3011 5290
rect 2969 5232 3011 5270
rect 3061 5290 3105 5332
rect 3061 5270 3073 5290
rect 3093 5270 3105 5290
rect 3061 5232 3105 5270
rect 1264 4972 1308 5010
rect 1264 4952 1276 4972
rect 1296 4952 1308 4972
rect 1264 4910 1308 4952
rect 1358 4972 1400 5010
rect 1358 4952 1372 4972
rect 1392 4952 1400 4972
rect 1358 4910 1400 4952
rect 1482 4972 1526 5010
rect 1482 4952 1494 4972
rect 1514 4952 1526 4972
rect 1482 4910 1526 4952
rect 1576 4972 1618 5010
rect 1576 4952 1590 4972
rect 1610 4952 1618 4972
rect 1576 4910 1618 4952
rect 1692 4972 1734 5010
rect 1692 4952 1700 4972
rect 1720 4952 1734 4972
rect 1692 4910 1734 4952
rect 1784 4979 1829 5010
rect 1784 4972 1828 4979
rect 1784 4952 1796 4972
rect 1816 4952 1828 4972
rect 1784 4910 1828 4952
rect 3420 4910 3464 4952
rect 3420 4890 3432 4910
rect 3452 4890 3464 4910
rect 3420 4883 3464 4890
rect 3419 4852 3464 4883
rect 3514 4910 3556 4952
rect 3514 4890 3528 4910
rect 3548 4890 3556 4910
rect 3514 4852 3556 4890
rect 3630 4910 3672 4952
rect 3630 4890 3638 4910
rect 3658 4890 3672 4910
rect 3630 4852 3672 4890
rect 3722 4910 3766 4952
rect 3722 4890 3734 4910
rect 3754 4890 3766 4910
rect 3722 4852 3766 4890
rect 3848 4910 3890 4952
rect 3848 4890 3856 4910
rect 3876 4890 3890 4910
rect 3848 4852 3890 4890
rect 3940 4910 3984 4952
rect 3940 4890 3952 4910
rect 3972 4890 3984 4910
rect 3940 4852 3984 4890
rect 367 4746 411 4784
rect 367 4726 379 4746
rect 399 4726 411 4746
rect 367 4684 411 4726
rect 461 4746 503 4784
rect 461 4726 475 4746
rect 495 4726 503 4746
rect 461 4684 503 4726
rect 585 4746 629 4784
rect 585 4726 597 4746
rect 617 4726 629 4746
rect 585 4684 629 4726
rect 679 4746 721 4784
rect 679 4726 693 4746
rect 713 4726 721 4746
rect 679 4684 721 4726
rect 795 4746 837 4784
rect 795 4726 803 4746
rect 823 4726 837 4746
rect 795 4684 837 4726
rect 887 4753 932 4784
rect 887 4746 931 4753
rect 887 4726 899 4746
rect 919 4726 931 4746
rect 887 4684 931 4726
rect 2623 4682 2667 4724
rect 2623 4662 2635 4682
rect 2655 4662 2667 4682
rect 2623 4655 2667 4662
rect 2622 4624 2667 4655
rect 2717 4682 2759 4724
rect 2717 4662 2731 4682
rect 2751 4662 2759 4682
rect 2717 4624 2759 4662
rect 2833 4682 2875 4724
rect 2833 4662 2841 4682
rect 2861 4662 2875 4682
rect 2833 4624 2875 4662
rect 2925 4682 2969 4724
rect 2925 4662 2937 4682
rect 2957 4662 2969 4682
rect 2925 4624 2969 4662
rect 3051 4682 3093 4724
rect 3051 4662 3059 4682
rect 3079 4662 3093 4682
rect 3051 4624 3093 4662
rect 3143 4682 3187 4724
rect 3143 4662 3155 4682
rect 3175 4662 3187 4682
rect 3143 4624 3187 4662
rect 1165 4562 1209 4600
rect 1165 4542 1177 4562
rect 1197 4542 1209 4562
rect 1165 4500 1209 4542
rect 1259 4562 1301 4600
rect 1259 4542 1273 4562
rect 1293 4542 1301 4562
rect 1259 4500 1301 4542
rect 1383 4562 1427 4600
rect 1383 4542 1395 4562
rect 1415 4542 1427 4562
rect 1383 4500 1427 4542
rect 1477 4562 1519 4600
rect 1477 4542 1491 4562
rect 1511 4542 1519 4562
rect 1477 4500 1519 4542
rect 1593 4562 1635 4600
rect 1593 4542 1601 4562
rect 1621 4542 1635 4562
rect 1593 4500 1635 4542
rect 1685 4569 1730 4600
rect 1685 4562 1729 4569
rect 1685 4542 1697 4562
rect 1717 4542 1729 4562
rect 1685 4500 1729 4542
rect 3421 4498 3465 4540
rect 3421 4478 3433 4498
rect 3453 4478 3465 4498
rect 3421 4471 3465 4478
rect 3420 4440 3465 4471
rect 3515 4498 3557 4540
rect 3515 4478 3529 4498
rect 3549 4478 3557 4498
rect 3515 4440 3557 4478
rect 3631 4498 3673 4540
rect 3631 4478 3639 4498
rect 3659 4478 3673 4498
rect 3631 4440 3673 4478
rect 3723 4498 3767 4540
rect 3723 4478 3735 4498
rect 3755 4478 3767 4498
rect 3723 4440 3767 4478
rect 3849 4498 3891 4540
rect 3849 4478 3857 4498
rect 3877 4478 3891 4498
rect 3849 4440 3891 4478
rect 3941 4498 3985 4540
rect 3941 4478 3953 4498
rect 3973 4478 3985 4498
rect 3941 4440 3985 4478
rect 368 4334 412 4372
rect 368 4314 380 4334
rect 400 4314 412 4334
rect 368 4272 412 4314
rect 462 4334 504 4372
rect 462 4314 476 4334
rect 496 4314 504 4334
rect 462 4272 504 4314
rect 586 4334 630 4372
rect 586 4314 598 4334
rect 618 4314 630 4334
rect 586 4272 630 4314
rect 680 4334 722 4372
rect 680 4314 694 4334
rect 714 4314 722 4334
rect 680 4272 722 4314
rect 796 4334 838 4372
rect 796 4314 804 4334
rect 824 4314 838 4334
rect 796 4272 838 4314
rect 888 4341 933 4372
rect 888 4334 932 4341
rect 888 4314 900 4334
rect 920 4314 932 4334
rect 888 4272 932 4314
rect 2319 4276 2363 4318
rect 2319 4256 2331 4276
rect 2351 4256 2363 4276
rect 2319 4249 2363 4256
rect 2318 4218 2363 4249
rect 2413 4276 2455 4318
rect 2413 4256 2427 4276
rect 2447 4256 2455 4276
rect 2413 4218 2455 4256
rect 2529 4276 2571 4318
rect 2529 4256 2537 4276
rect 2557 4256 2571 4276
rect 2529 4218 2571 4256
rect 2621 4276 2665 4318
rect 2621 4256 2633 4276
rect 2653 4256 2665 4276
rect 2621 4218 2665 4256
rect 2747 4276 2789 4318
rect 2747 4256 2755 4276
rect 2775 4256 2789 4276
rect 2747 4218 2789 4256
rect 2839 4276 2883 4318
rect 2839 4256 2851 4276
rect 2871 4256 2883 4276
rect 2839 4218 2883 4256
rect 1450 3950 1494 3988
rect 1450 3930 1462 3950
rect 1482 3930 1494 3950
rect 1450 3888 1494 3930
rect 1544 3950 1586 3988
rect 1544 3930 1558 3950
rect 1578 3930 1586 3950
rect 1544 3888 1586 3930
rect 1668 3950 1712 3988
rect 1668 3930 1680 3950
rect 1700 3930 1712 3950
rect 1668 3888 1712 3930
rect 1762 3950 1804 3988
rect 1762 3930 1776 3950
rect 1796 3930 1804 3950
rect 1762 3888 1804 3930
rect 1878 3950 1920 3988
rect 1878 3930 1886 3950
rect 1906 3930 1920 3950
rect 1878 3888 1920 3930
rect 1970 3957 2015 3988
rect 1970 3950 2014 3957
rect 1970 3930 1982 3950
rect 2002 3930 2014 3950
rect 1970 3888 2014 3930
rect 3401 3892 3445 3934
rect 3401 3872 3413 3892
rect 3433 3872 3445 3892
rect 3401 3865 3445 3872
rect 3400 3834 3445 3865
rect 3495 3892 3537 3934
rect 3495 3872 3509 3892
rect 3529 3872 3537 3892
rect 3495 3834 3537 3872
rect 3611 3892 3653 3934
rect 3611 3872 3619 3892
rect 3639 3872 3653 3892
rect 3611 3834 3653 3872
rect 3703 3892 3747 3934
rect 3703 3872 3715 3892
rect 3735 3872 3747 3892
rect 3703 3834 3747 3872
rect 3829 3892 3871 3934
rect 3829 3872 3837 3892
rect 3857 3872 3871 3892
rect 3829 3834 3871 3872
rect 3921 3892 3965 3934
rect 3921 3872 3933 3892
rect 3953 3872 3965 3892
rect 3921 3834 3965 3872
rect 348 3728 392 3766
rect 348 3708 360 3728
rect 380 3708 392 3728
rect 348 3666 392 3708
rect 442 3728 484 3766
rect 442 3708 456 3728
rect 476 3708 484 3728
rect 442 3666 484 3708
rect 566 3728 610 3766
rect 566 3708 578 3728
rect 598 3708 610 3728
rect 566 3666 610 3708
rect 660 3728 702 3766
rect 660 3708 674 3728
rect 694 3708 702 3728
rect 660 3666 702 3708
rect 776 3728 818 3766
rect 776 3708 784 3728
rect 804 3708 818 3728
rect 776 3666 818 3708
rect 868 3735 913 3766
rect 868 3728 912 3735
rect 868 3708 880 3728
rect 900 3708 912 3728
rect 868 3666 912 3708
rect 2604 3664 2648 3706
rect 2604 3644 2616 3664
rect 2636 3644 2648 3664
rect 2604 3637 2648 3644
rect 2603 3606 2648 3637
rect 2698 3664 2740 3706
rect 2698 3644 2712 3664
rect 2732 3644 2740 3664
rect 2698 3606 2740 3644
rect 2814 3664 2856 3706
rect 2814 3644 2822 3664
rect 2842 3644 2856 3664
rect 2814 3606 2856 3644
rect 2906 3664 2950 3706
rect 2906 3644 2918 3664
rect 2938 3644 2950 3664
rect 2906 3606 2950 3644
rect 3032 3664 3074 3706
rect 3032 3644 3040 3664
rect 3060 3644 3074 3664
rect 3032 3606 3074 3644
rect 3124 3664 3168 3706
rect 3124 3644 3136 3664
rect 3156 3644 3168 3664
rect 3124 3606 3168 3644
rect 1146 3544 1190 3582
rect 1146 3524 1158 3544
rect 1178 3524 1190 3544
rect 1146 3482 1190 3524
rect 1240 3544 1282 3582
rect 1240 3524 1254 3544
rect 1274 3524 1282 3544
rect 1240 3482 1282 3524
rect 1364 3544 1408 3582
rect 1364 3524 1376 3544
rect 1396 3524 1408 3544
rect 1364 3482 1408 3524
rect 1458 3544 1500 3582
rect 1458 3524 1472 3544
rect 1492 3524 1500 3544
rect 1458 3482 1500 3524
rect 1574 3544 1616 3582
rect 1574 3524 1582 3544
rect 1602 3524 1616 3544
rect 1574 3482 1616 3524
rect 1666 3551 1711 3582
rect 1666 3544 1710 3551
rect 1666 3524 1678 3544
rect 1698 3524 1710 3544
rect 1666 3482 1710 3524
rect 3402 3480 3446 3522
rect 3402 3460 3414 3480
rect 3434 3460 3446 3480
rect 3402 3453 3446 3460
rect 3401 3422 3446 3453
rect 3496 3480 3538 3522
rect 3496 3460 3510 3480
rect 3530 3460 3538 3480
rect 3496 3422 3538 3460
rect 3612 3480 3654 3522
rect 3612 3460 3620 3480
rect 3640 3460 3654 3480
rect 3612 3422 3654 3460
rect 3704 3480 3748 3522
rect 3704 3460 3716 3480
rect 3736 3460 3748 3480
rect 3704 3422 3748 3460
rect 3830 3480 3872 3522
rect 3830 3460 3838 3480
rect 3858 3460 3872 3480
rect 3830 3422 3872 3460
rect 3922 3480 3966 3522
rect 3922 3460 3934 3480
rect 3954 3460 3966 3480
rect 3922 3422 3966 3460
rect 349 3316 393 3354
rect 349 3296 361 3316
rect 381 3296 393 3316
rect 349 3254 393 3296
rect 443 3316 485 3354
rect 443 3296 457 3316
rect 477 3296 485 3316
rect 443 3254 485 3296
rect 567 3316 611 3354
rect 567 3296 579 3316
rect 599 3296 611 3316
rect 567 3254 611 3296
rect 661 3316 703 3354
rect 661 3296 675 3316
rect 695 3296 703 3316
rect 661 3254 703 3296
rect 777 3316 819 3354
rect 777 3296 785 3316
rect 805 3296 819 3316
rect 777 3254 819 3296
rect 869 3323 914 3354
rect 869 3316 913 3323
rect 869 3296 881 3316
rect 901 3296 913 3316
rect 869 3254 913 3296
rect 2505 3254 2549 3296
rect 2505 3234 2517 3254
rect 2537 3234 2549 3254
rect 2505 3227 2549 3234
rect 2504 3196 2549 3227
rect 2599 3254 2641 3296
rect 2599 3234 2613 3254
rect 2633 3234 2641 3254
rect 2599 3196 2641 3234
rect 2715 3254 2757 3296
rect 2715 3234 2723 3254
rect 2743 3234 2757 3254
rect 2715 3196 2757 3234
rect 2807 3254 2851 3296
rect 2807 3234 2819 3254
rect 2839 3234 2851 3254
rect 2807 3196 2851 3234
rect 2933 3254 2975 3296
rect 2933 3234 2941 3254
rect 2961 3234 2975 3254
rect 2933 3196 2975 3234
rect 3025 3254 3069 3296
rect 3025 3234 3037 3254
rect 3057 3234 3069 3254
rect 3025 3196 3069 3234
rect 1228 2936 1272 2974
rect 1228 2916 1240 2936
rect 1260 2916 1272 2936
rect 1228 2874 1272 2916
rect 1322 2936 1364 2974
rect 1322 2916 1336 2936
rect 1356 2916 1364 2936
rect 1322 2874 1364 2916
rect 1446 2936 1490 2974
rect 1446 2916 1458 2936
rect 1478 2916 1490 2936
rect 1446 2874 1490 2916
rect 1540 2936 1582 2974
rect 1540 2916 1554 2936
rect 1574 2916 1582 2936
rect 1540 2874 1582 2916
rect 1656 2936 1698 2974
rect 1656 2916 1664 2936
rect 1684 2916 1698 2936
rect 1656 2874 1698 2916
rect 1748 2943 1793 2974
rect 1748 2936 1792 2943
rect 1748 2916 1760 2936
rect 1780 2916 1792 2936
rect 1748 2874 1792 2916
rect 3384 2874 3428 2916
rect 3384 2854 3396 2874
rect 3416 2854 3428 2874
rect 3384 2847 3428 2854
rect 3383 2816 3428 2847
rect 3478 2874 3520 2916
rect 3478 2854 3492 2874
rect 3512 2854 3520 2874
rect 3478 2816 3520 2854
rect 3594 2874 3636 2916
rect 3594 2854 3602 2874
rect 3622 2854 3636 2874
rect 3594 2816 3636 2854
rect 3686 2874 3730 2916
rect 3686 2854 3698 2874
rect 3718 2854 3730 2874
rect 3686 2816 3730 2854
rect 3812 2874 3854 2916
rect 3812 2854 3820 2874
rect 3840 2854 3854 2874
rect 3812 2816 3854 2854
rect 3904 2874 3948 2916
rect 3904 2854 3916 2874
rect 3936 2854 3948 2874
rect 3904 2816 3948 2854
rect 331 2710 375 2748
rect 331 2690 343 2710
rect 363 2690 375 2710
rect 331 2648 375 2690
rect 425 2710 467 2748
rect 425 2690 439 2710
rect 459 2690 467 2710
rect 425 2648 467 2690
rect 549 2710 593 2748
rect 549 2690 561 2710
rect 581 2690 593 2710
rect 549 2648 593 2690
rect 643 2710 685 2748
rect 643 2690 657 2710
rect 677 2690 685 2710
rect 643 2648 685 2690
rect 759 2710 801 2748
rect 759 2690 767 2710
rect 787 2690 801 2710
rect 759 2648 801 2690
rect 851 2717 896 2748
rect 851 2710 895 2717
rect 851 2690 863 2710
rect 883 2690 895 2710
rect 851 2648 895 2690
rect 2587 2646 2631 2688
rect 2587 2626 2599 2646
rect 2619 2626 2631 2646
rect 2587 2619 2631 2626
rect 2586 2588 2631 2619
rect 2681 2646 2723 2688
rect 2681 2626 2695 2646
rect 2715 2626 2723 2646
rect 2681 2588 2723 2626
rect 2797 2646 2839 2688
rect 2797 2626 2805 2646
rect 2825 2626 2839 2646
rect 2797 2588 2839 2626
rect 2889 2646 2933 2688
rect 2889 2626 2901 2646
rect 2921 2626 2933 2646
rect 2889 2588 2933 2626
rect 3015 2646 3057 2688
rect 3015 2626 3023 2646
rect 3043 2626 3057 2646
rect 3015 2588 3057 2626
rect 3107 2646 3151 2688
rect 3107 2626 3119 2646
rect 3139 2626 3151 2646
rect 3107 2588 3151 2626
rect 1129 2526 1173 2564
rect 1129 2506 1141 2526
rect 1161 2506 1173 2526
rect 1129 2464 1173 2506
rect 1223 2526 1265 2564
rect 1223 2506 1237 2526
rect 1257 2506 1265 2526
rect 1223 2464 1265 2506
rect 1347 2526 1391 2564
rect 1347 2506 1359 2526
rect 1379 2506 1391 2526
rect 1347 2464 1391 2506
rect 1441 2526 1483 2564
rect 1441 2506 1455 2526
rect 1475 2506 1483 2526
rect 1441 2464 1483 2506
rect 1557 2526 1599 2564
rect 1557 2506 1565 2526
rect 1585 2506 1599 2526
rect 1557 2464 1599 2506
rect 1649 2533 1694 2564
rect 1649 2526 1693 2533
rect 1649 2506 1661 2526
rect 1681 2506 1693 2526
rect 1649 2464 1693 2506
rect 3385 2462 3429 2504
rect 3385 2442 3397 2462
rect 3417 2442 3429 2462
rect 3385 2435 3429 2442
rect 3384 2404 3429 2435
rect 3479 2462 3521 2504
rect 3479 2442 3493 2462
rect 3513 2442 3521 2462
rect 3479 2404 3521 2442
rect 3595 2462 3637 2504
rect 3595 2442 3603 2462
rect 3623 2442 3637 2462
rect 3595 2404 3637 2442
rect 3687 2462 3731 2504
rect 3687 2442 3699 2462
rect 3719 2442 3731 2462
rect 3687 2404 3731 2442
rect 3813 2462 3855 2504
rect 3813 2442 3821 2462
rect 3841 2442 3855 2462
rect 3813 2404 3855 2442
rect 3905 2462 3949 2504
rect 3905 2442 3917 2462
rect 3937 2442 3949 2462
rect 3905 2404 3949 2442
rect 332 2298 376 2336
rect 332 2278 344 2298
rect 364 2278 376 2298
rect 332 2236 376 2278
rect 426 2298 468 2336
rect 426 2278 440 2298
rect 460 2278 468 2298
rect 426 2236 468 2278
rect 550 2298 594 2336
rect 550 2278 562 2298
rect 582 2278 594 2298
rect 550 2236 594 2278
rect 644 2298 686 2336
rect 644 2278 658 2298
rect 678 2278 686 2298
rect 644 2236 686 2278
rect 760 2298 802 2336
rect 760 2278 768 2298
rect 788 2278 802 2298
rect 760 2236 802 2278
rect 852 2305 897 2336
rect 852 2298 896 2305
rect 852 2278 864 2298
rect 884 2278 896 2298
rect 852 2236 896 2278
rect 2422 2238 2466 2280
rect 2422 2218 2434 2238
rect 2454 2218 2466 2238
rect 2422 2211 2466 2218
rect 2421 2180 2466 2211
rect 2516 2238 2558 2280
rect 2516 2218 2530 2238
rect 2550 2218 2558 2238
rect 2516 2180 2558 2218
rect 2632 2238 2674 2280
rect 2632 2218 2640 2238
rect 2660 2218 2674 2238
rect 2632 2180 2674 2218
rect 2724 2238 2768 2280
rect 2724 2218 2736 2238
rect 2756 2218 2768 2238
rect 2724 2180 2768 2218
rect 2850 2238 2892 2280
rect 2850 2218 2858 2238
rect 2878 2218 2892 2238
rect 2850 2180 2892 2218
rect 2942 2238 2986 2280
rect 2942 2218 2954 2238
rect 2974 2218 2986 2238
rect 2942 2180 2986 2218
rect 1274 1916 1318 1954
rect 1274 1896 1286 1916
rect 1306 1896 1318 1916
rect 1274 1854 1318 1896
rect 1368 1916 1410 1954
rect 1368 1896 1382 1916
rect 1402 1896 1410 1916
rect 1368 1854 1410 1896
rect 1492 1916 1536 1954
rect 1492 1896 1504 1916
rect 1524 1896 1536 1916
rect 1492 1854 1536 1896
rect 1586 1916 1628 1954
rect 1586 1896 1600 1916
rect 1620 1896 1628 1916
rect 1586 1854 1628 1896
rect 1702 1916 1744 1954
rect 1702 1896 1710 1916
rect 1730 1896 1744 1916
rect 1702 1854 1744 1896
rect 1794 1923 1839 1954
rect 1794 1916 1838 1923
rect 1794 1896 1806 1916
rect 1826 1896 1838 1916
rect 1794 1854 1838 1896
rect 3364 1856 3408 1898
rect 3364 1836 3376 1856
rect 3396 1836 3408 1856
rect 3364 1829 3408 1836
rect 3363 1798 3408 1829
rect 3458 1856 3500 1898
rect 3458 1836 3472 1856
rect 3492 1836 3500 1856
rect 3458 1798 3500 1836
rect 3574 1856 3616 1898
rect 3574 1836 3582 1856
rect 3602 1836 3616 1856
rect 3574 1798 3616 1836
rect 3666 1856 3710 1898
rect 3666 1836 3678 1856
rect 3698 1836 3710 1856
rect 3666 1798 3710 1836
rect 3792 1856 3834 1898
rect 3792 1836 3800 1856
rect 3820 1836 3834 1856
rect 3792 1798 3834 1836
rect 3884 1856 3928 1898
rect 3884 1836 3896 1856
rect 3916 1836 3928 1856
rect 3884 1798 3928 1836
rect 311 1692 355 1730
rect 311 1672 323 1692
rect 343 1672 355 1692
rect 311 1630 355 1672
rect 405 1692 447 1730
rect 405 1672 419 1692
rect 439 1672 447 1692
rect 405 1630 447 1672
rect 529 1692 573 1730
rect 529 1672 541 1692
rect 561 1672 573 1692
rect 529 1630 573 1672
rect 623 1692 665 1730
rect 623 1672 637 1692
rect 657 1672 665 1692
rect 623 1630 665 1672
rect 739 1692 781 1730
rect 739 1672 747 1692
rect 767 1672 781 1692
rect 739 1630 781 1672
rect 831 1699 876 1730
rect 831 1692 875 1699
rect 831 1672 843 1692
rect 863 1672 875 1692
rect 831 1630 875 1672
rect 2567 1628 2611 1670
rect 2567 1608 2579 1628
rect 2599 1608 2611 1628
rect 2567 1601 2611 1608
rect 2566 1570 2611 1601
rect 2661 1628 2703 1670
rect 2661 1608 2675 1628
rect 2695 1608 2703 1628
rect 2661 1570 2703 1608
rect 2777 1628 2819 1670
rect 2777 1608 2785 1628
rect 2805 1608 2819 1628
rect 2777 1570 2819 1608
rect 2869 1628 2913 1670
rect 2869 1608 2881 1628
rect 2901 1608 2913 1628
rect 2869 1570 2913 1608
rect 2995 1628 3037 1670
rect 2995 1608 3003 1628
rect 3023 1608 3037 1628
rect 2995 1570 3037 1608
rect 3087 1628 3131 1670
rect 3087 1608 3099 1628
rect 3119 1608 3131 1628
rect 3087 1570 3131 1608
rect 1109 1508 1153 1546
rect 1109 1488 1121 1508
rect 1141 1488 1153 1508
rect 1109 1446 1153 1488
rect 1203 1508 1245 1546
rect 1203 1488 1217 1508
rect 1237 1488 1245 1508
rect 1203 1446 1245 1488
rect 1327 1508 1371 1546
rect 1327 1488 1339 1508
rect 1359 1488 1371 1508
rect 1327 1446 1371 1488
rect 1421 1508 1463 1546
rect 1421 1488 1435 1508
rect 1455 1488 1463 1508
rect 1421 1446 1463 1488
rect 1537 1508 1579 1546
rect 1537 1488 1545 1508
rect 1565 1488 1579 1508
rect 1537 1446 1579 1488
rect 1629 1515 1674 1546
rect 1629 1508 1673 1515
rect 1629 1488 1641 1508
rect 1661 1488 1673 1508
rect 1629 1446 1673 1488
rect 3365 1444 3409 1486
rect 3365 1424 3377 1444
rect 3397 1424 3409 1444
rect 3365 1417 3409 1424
rect 3364 1386 3409 1417
rect 3459 1444 3501 1486
rect 3459 1424 3473 1444
rect 3493 1424 3501 1444
rect 3459 1386 3501 1424
rect 3575 1444 3617 1486
rect 3575 1424 3583 1444
rect 3603 1424 3617 1444
rect 3575 1386 3617 1424
rect 3667 1444 3711 1486
rect 3667 1424 3679 1444
rect 3699 1424 3711 1444
rect 3667 1386 3711 1424
rect 3793 1444 3835 1486
rect 3793 1424 3801 1444
rect 3821 1424 3835 1444
rect 3793 1386 3835 1424
rect 3885 1444 3929 1486
rect 3885 1424 3897 1444
rect 3917 1424 3929 1444
rect 3885 1386 3929 1424
rect 312 1280 356 1318
rect 312 1260 324 1280
rect 344 1260 356 1280
rect 312 1218 356 1260
rect 406 1280 448 1318
rect 406 1260 420 1280
rect 440 1260 448 1280
rect 406 1218 448 1260
rect 530 1280 574 1318
rect 530 1260 542 1280
rect 562 1260 574 1280
rect 530 1218 574 1260
rect 624 1280 666 1318
rect 624 1260 638 1280
rect 658 1260 666 1280
rect 624 1218 666 1260
rect 740 1280 782 1318
rect 740 1260 748 1280
rect 768 1260 782 1280
rect 740 1218 782 1260
rect 832 1287 877 1318
rect 832 1280 876 1287
rect 832 1260 844 1280
rect 864 1260 876 1280
rect 832 1218 876 1260
rect 2468 1218 2512 1260
rect 2468 1198 2480 1218
rect 2500 1198 2512 1218
rect 2468 1191 2512 1198
rect 2467 1160 2512 1191
rect 2562 1218 2604 1260
rect 2562 1198 2576 1218
rect 2596 1198 2604 1218
rect 2562 1160 2604 1198
rect 2678 1218 2720 1260
rect 2678 1198 2686 1218
rect 2706 1198 2720 1218
rect 2678 1160 2720 1198
rect 2770 1218 2814 1260
rect 2770 1198 2782 1218
rect 2802 1198 2814 1218
rect 2770 1160 2814 1198
rect 2896 1218 2938 1260
rect 2896 1198 2904 1218
rect 2924 1198 2938 1218
rect 2896 1160 2938 1198
rect 2988 1218 3032 1260
rect 2988 1198 3000 1218
rect 3020 1198 3032 1218
rect 2988 1160 3032 1198
rect 1191 900 1235 938
rect 1191 880 1203 900
rect 1223 880 1235 900
rect 1191 838 1235 880
rect 1285 900 1327 938
rect 1285 880 1299 900
rect 1319 880 1327 900
rect 1285 838 1327 880
rect 1409 900 1453 938
rect 1409 880 1421 900
rect 1441 880 1453 900
rect 1409 838 1453 880
rect 1503 900 1545 938
rect 1503 880 1517 900
rect 1537 880 1545 900
rect 1503 838 1545 880
rect 1619 900 1661 938
rect 1619 880 1627 900
rect 1647 880 1661 900
rect 1619 838 1661 880
rect 1711 907 1756 938
rect 1711 900 1755 907
rect 1711 880 1723 900
rect 1743 880 1755 900
rect 1711 838 1755 880
rect 3347 838 3391 880
rect 3347 818 3359 838
rect 3379 818 3391 838
rect 3347 811 3391 818
rect 3346 780 3391 811
rect 3441 838 3483 880
rect 3441 818 3455 838
rect 3475 818 3483 838
rect 3441 780 3483 818
rect 3557 838 3599 880
rect 3557 818 3565 838
rect 3585 818 3599 838
rect 3557 780 3599 818
rect 3649 838 3693 880
rect 3649 818 3661 838
rect 3681 818 3693 838
rect 3649 780 3693 818
rect 3775 838 3817 880
rect 3775 818 3783 838
rect 3803 818 3817 838
rect 3775 780 3817 818
rect 3867 838 3911 880
rect 3867 818 3879 838
rect 3899 818 3911 838
rect 3867 780 3911 818
rect 294 674 338 712
rect 294 654 306 674
rect 326 654 338 674
rect 294 612 338 654
rect 388 674 430 712
rect 388 654 402 674
rect 422 654 430 674
rect 388 612 430 654
rect 512 674 556 712
rect 512 654 524 674
rect 544 654 556 674
rect 512 612 556 654
rect 606 674 648 712
rect 606 654 620 674
rect 640 654 648 674
rect 606 612 648 654
rect 722 674 764 712
rect 722 654 730 674
rect 750 654 764 674
rect 722 612 764 654
rect 814 681 859 712
rect 814 674 858 681
rect 814 654 826 674
rect 846 654 858 674
rect 814 612 858 654
rect 2550 610 2594 652
rect 2550 590 2562 610
rect 2582 590 2594 610
rect 2550 583 2594 590
rect 2549 552 2594 583
rect 2644 610 2686 652
rect 2644 590 2658 610
rect 2678 590 2686 610
rect 2644 552 2686 590
rect 2760 610 2802 652
rect 2760 590 2768 610
rect 2788 590 2802 610
rect 2760 552 2802 590
rect 2852 610 2896 652
rect 2852 590 2864 610
rect 2884 590 2896 610
rect 2852 552 2896 590
rect 2978 610 3020 652
rect 2978 590 2986 610
rect 3006 590 3020 610
rect 2978 552 3020 590
rect 3070 610 3114 652
rect 3070 590 3082 610
rect 3102 590 3114 610
rect 3070 552 3114 590
rect 1092 490 1136 528
rect 1092 470 1104 490
rect 1124 470 1136 490
rect 1092 428 1136 470
rect 1186 490 1228 528
rect 1186 470 1200 490
rect 1220 470 1228 490
rect 1186 428 1228 470
rect 1310 490 1354 528
rect 1310 470 1322 490
rect 1342 470 1354 490
rect 1310 428 1354 470
rect 1404 490 1446 528
rect 1404 470 1418 490
rect 1438 470 1446 490
rect 1404 428 1446 470
rect 1520 490 1562 528
rect 1520 470 1528 490
rect 1548 470 1562 490
rect 1520 428 1562 470
rect 1612 497 1657 528
rect 1612 490 1656 497
rect 1612 470 1624 490
rect 1644 470 1656 490
rect 1612 428 1656 470
rect 3348 426 3392 468
rect 3348 406 3360 426
rect 3380 406 3392 426
rect 3348 399 3392 406
rect 3347 368 3392 399
rect 3442 426 3484 468
rect 3442 406 3456 426
rect 3476 406 3484 426
rect 3442 368 3484 406
rect 3558 426 3600 468
rect 3558 406 3566 426
rect 3586 406 3600 426
rect 3558 368 3600 406
rect 3650 426 3694 468
rect 3650 406 3662 426
rect 3682 406 3694 426
rect 3650 368 3694 406
rect 3776 426 3818 468
rect 3776 406 3784 426
rect 3804 406 3818 426
rect 3776 368 3818 406
rect 3868 426 3912 468
rect 3868 406 3880 426
rect 3900 406 3912 426
rect 3868 368 3912 406
rect 295 262 339 300
rect 295 242 307 262
rect 327 242 339 262
rect 295 200 339 242
rect 389 262 431 300
rect 389 242 403 262
rect 423 242 431 262
rect 389 200 431 242
rect 513 262 557 300
rect 513 242 525 262
rect 545 242 557 262
rect 513 200 557 242
rect 607 262 649 300
rect 607 242 621 262
rect 641 242 649 262
rect 607 200 649 242
rect 723 262 765 300
rect 723 242 731 262
rect 751 242 765 262
rect 723 200 765 242
rect 815 269 860 300
rect 815 262 859 269
rect 815 242 827 262
rect 847 242 859 262
rect 815 200 859 242
rect 1508 -314 1552 -276
rect 1508 -334 1520 -314
rect 1540 -334 1552 -314
rect 1508 -376 1552 -334
rect 1602 -314 1644 -276
rect 1602 -334 1616 -314
rect 1636 -334 1644 -314
rect 1602 -376 1644 -334
rect 1726 -314 1770 -276
rect 1726 -334 1738 -314
rect 1758 -334 1770 -314
rect 1726 -376 1770 -334
rect 1820 -314 1862 -276
rect 1820 -334 1834 -314
rect 1854 -334 1862 -314
rect 1820 -376 1862 -334
rect 1936 -314 1978 -276
rect 1936 -334 1944 -314
rect 1964 -334 1978 -314
rect 1936 -376 1978 -334
rect 2028 -307 2073 -276
rect 2028 -314 2072 -307
rect 2028 -334 2040 -314
rect 2060 -334 2072 -314
rect 2028 -376 2072 -334
<< ndiffc >>
rect 3480 8093 3500 8113
rect 3583 8089 3603 8109
rect 3691 8089 3711 8109
rect 3794 8093 3814 8113
rect 3909 8089 3929 8109
rect 4012 8093 4032 8113
rect 4199 8100 4217 8118
rect 263 8038 281 8056
rect 261 7939 279 7957
rect 4197 8001 4215 8019
rect 2683 7865 2703 7885
rect 2786 7861 2806 7881
rect 2894 7861 2914 7881
rect 2997 7865 3017 7885
rect 3112 7861 3132 7881
rect 3215 7865 3235 7885
rect 4192 7882 4210 7900
rect 4190 7783 4208 7801
rect 258 7714 276 7732
rect 3481 7681 3501 7701
rect 256 7615 274 7633
rect 427 7631 447 7651
rect 530 7635 550 7655
rect 645 7631 665 7651
rect 748 7635 768 7655
rect 856 7635 876 7655
rect 3584 7677 3604 7697
rect 3692 7677 3712 7697
rect 3795 7681 3815 7701
rect 3910 7677 3930 7697
rect 4013 7681 4033 7701
rect 4186 7699 4204 7717
rect 959 7631 979 7651
rect 4184 7600 4202 7618
rect 252 7531 270 7549
rect 250 7432 268 7450
rect 1225 7447 1245 7467
rect 1328 7451 1348 7471
rect 1443 7447 1463 7467
rect 1546 7451 1566 7471
rect 1654 7451 1674 7471
rect 1757 7447 1777 7467
rect 2584 7455 2604 7475
rect 2687 7451 2707 7471
rect 2795 7451 2815 7471
rect 2898 7455 2918 7475
rect 3013 7451 3033 7471
rect 3116 7455 3136 7475
rect 245 7313 263 7331
rect 4181 7375 4199 7393
rect 4179 7276 4197 7294
rect 243 7214 261 7232
rect 428 7219 448 7239
rect 531 7223 551 7243
rect 646 7219 666 7239
rect 749 7223 769 7243
rect 857 7223 877 7243
rect 960 7219 980 7239
rect 3463 7075 3483 7095
rect 3566 7071 3586 7091
rect 3674 7071 3694 7091
rect 3777 7075 3797 7095
rect 3892 7071 3912 7091
rect 3995 7075 4015 7095
rect 4182 7082 4200 7100
rect 246 7020 264 7038
rect 244 6921 262 6939
rect 4180 6983 4198 7001
rect 1307 6839 1327 6859
rect 1410 6843 1430 6863
rect 1525 6839 1545 6859
rect 1628 6843 1648 6863
rect 1736 6843 1756 6863
rect 1839 6839 1859 6859
rect 2666 6847 2686 6867
rect 2769 6843 2789 6863
rect 2877 6843 2897 6863
rect 2980 6847 3000 6867
rect 3095 6843 3115 6863
rect 3198 6847 3218 6867
rect 4175 6864 4193 6882
rect 4173 6765 4191 6783
rect 241 6696 259 6714
rect 3464 6663 3484 6683
rect 239 6597 257 6615
rect 410 6613 430 6633
rect 513 6617 533 6637
rect 628 6613 648 6633
rect 731 6617 751 6637
rect 839 6617 859 6637
rect 3567 6659 3587 6679
rect 3675 6659 3695 6679
rect 3778 6663 3798 6683
rect 3893 6659 3913 6679
rect 3996 6663 4016 6683
rect 4169 6681 4187 6699
rect 942 6613 962 6633
rect 4167 6582 4185 6600
rect 235 6513 253 6531
rect 233 6414 251 6432
rect 1208 6429 1228 6449
rect 1311 6433 1331 6453
rect 1426 6429 1446 6449
rect 1529 6433 1549 6453
rect 1637 6433 1657 6453
rect 1740 6429 1760 6449
rect 2501 6439 2521 6459
rect 2604 6435 2624 6455
rect 2712 6435 2732 6455
rect 2815 6439 2835 6459
rect 2930 6435 2950 6455
rect 3033 6439 3053 6459
rect 228 6295 246 6313
rect 4164 6357 4182 6375
rect 4162 6258 4180 6276
rect 226 6196 244 6214
rect 411 6201 431 6221
rect 514 6205 534 6225
rect 629 6201 649 6221
rect 732 6205 752 6225
rect 840 6205 860 6225
rect 943 6201 963 6221
rect 3443 6057 3463 6077
rect 3546 6053 3566 6073
rect 3654 6053 3674 6073
rect 3757 6057 3777 6077
rect 3872 6053 3892 6073
rect 3975 6057 3995 6077
rect 4162 6064 4180 6082
rect 226 6002 244 6020
rect 224 5903 242 5921
rect 4160 5965 4178 5983
rect 1353 5819 1373 5839
rect 1456 5823 1476 5843
rect 1571 5819 1591 5839
rect 1674 5823 1694 5843
rect 1782 5823 1802 5843
rect 1885 5819 1905 5839
rect 2646 5829 2666 5849
rect 2749 5825 2769 5845
rect 2857 5825 2877 5845
rect 2960 5829 2980 5849
rect 3075 5825 3095 5845
rect 3178 5829 3198 5849
rect 4155 5846 4173 5864
rect 4153 5747 4171 5765
rect 221 5678 239 5696
rect 3444 5645 3464 5665
rect 219 5579 237 5597
rect 390 5595 410 5615
rect 493 5599 513 5619
rect 608 5595 628 5615
rect 711 5599 731 5619
rect 819 5599 839 5619
rect 3547 5641 3567 5661
rect 3655 5641 3675 5661
rect 3758 5645 3778 5665
rect 3873 5641 3893 5661
rect 3976 5645 3996 5665
rect 4149 5663 4167 5681
rect 922 5595 942 5615
rect 4147 5564 4165 5582
rect 215 5495 233 5513
rect 213 5396 231 5414
rect 1188 5411 1208 5431
rect 1291 5415 1311 5435
rect 1406 5411 1426 5431
rect 1509 5415 1529 5435
rect 1617 5415 1637 5435
rect 1720 5411 1740 5431
rect 2547 5419 2567 5439
rect 2650 5415 2670 5435
rect 2758 5415 2778 5435
rect 2861 5419 2881 5439
rect 2976 5415 2996 5435
rect 3079 5419 3099 5439
rect 208 5277 226 5295
rect 4144 5339 4162 5357
rect 4142 5240 4160 5258
rect 206 5178 224 5196
rect 391 5183 411 5203
rect 494 5187 514 5207
rect 609 5183 629 5203
rect 712 5187 732 5207
rect 820 5187 840 5207
rect 923 5183 943 5203
rect 3426 5039 3446 5059
rect 3529 5035 3549 5055
rect 3637 5035 3657 5055
rect 3740 5039 3760 5059
rect 3855 5035 3875 5055
rect 3958 5039 3978 5059
rect 4145 5046 4163 5064
rect 209 4984 227 5002
rect 207 4885 225 4903
rect 4143 4947 4161 4965
rect 1270 4803 1290 4823
rect 1373 4807 1393 4827
rect 1488 4803 1508 4823
rect 1591 4807 1611 4827
rect 1699 4807 1719 4827
rect 1802 4803 1822 4823
rect 2629 4811 2649 4831
rect 2732 4807 2752 4827
rect 2840 4807 2860 4827
rect 2943 4811 2963 4831
rect 3058 4807 3078 4827
rect 3161 4811 3181 4831
rect 4138 4828 4156 4846
rect 4136 4729 4154 4747
rect 204 4660 222 4678
rect 3427 4627 3447 4647
rect 202 4561 220 4579
rect 373 4577 393 4597
rect 476 4581 496 4601
rect 591 4577 611 4597
rect 694 4581 714 4601
rect 802 4581 822 4601
rect 3530 4623 3550 4643
rect 3638 4623 3658 4643
rect 3741 4627 3761 4647
rect 3856 4623 3876 4643
rect 3959 4627 3979 4647
rect 4132 4645 4150 4663
rect 905 4577 925 4597
rect 4130 4546 4148 4564
rect 198 4477 216 4495
rect 196 4378 214 4396
rect 1171 4393 1191 4413
rect 1274 4397 1294 4417
rect 1389 4393 1409 4413
rect 1492 4397 1512 4417
rect 1600 4397 1620 4417
rect 1703 4393 1723 4413
rect 2325 4405 2345 4425
rect 2428 4401 2448 4421
rect 2536 4401 2556 4421
rect 2639 4405 2659 4425
rect 2754 4401 2774 4421
rect 2857 4405 2877 4425
rect 191 4259 209 4277
rect 4127 4321 4145 4339
rect 4125 4222 4143 4240
rect 189 4160 207 4178
rect 374 4165 394 4185
rect 477 4169 497 4189
rect 592 4165 612 4185
rect 695 4169 715 4189
rect 803 4169 823 4189
rect 906 4165 926 4185
rect 3407 4021 3427 4041
rect 3510 4017 3530 4037
rect 3618 4017 3638 4037
rect 3721 4021 3741 4041
rect 3836 4017 3856 4037
rect 3939 4021 3959 4041
rect 4126 4028 4144 4046
rect 190 3966 208 3984
rect 188 3867 206 3885
rect 4124 3929 4142 3947
rect 1456 3781 1476 3801
rect 1559 3785 1579 3805
rect 1674 3781 1694 3801
rect 1777 3785 1797 3805
rect 1885 3785 1905 3805
rect 1988 3781 2008 3801
rect 2610 3793 2630 3813
rect 2713 3789 2733 3809
rect 2821 3789 2841 3809
rect 2924 3793 2944 3813
rect 3039 3789 3059 3809
rect 3142 3793 3162 3813
rect 4119 3810 4137 3828
rect 4117 3711 4135 3729
rect 185 3642 203 3660
rect 3408 3609 3428 3629
rect 183 3543 201 3561
rect 354 3559 374 3579
rect 457 3563 477 3583
rect 572 3559 592 3579
rect 675 3563 695 3583
rect 783 3563 803 3583
rect 3511 3605 3531 3625
rect 3619 3605 3639 3625
rect 3722 3609 3742 3629
rect 3837 3605 3857 3625
rect 3940 3609 3960 3629
rect 4113 3627 4131 3645
rect 886 3559 906 3579
rect 4111 3528 4129 3546
rect 179 3459 197 3477
rect 177 3360 195 3378
rect 1152 3375 1172 3395
rect 1255 3379 1275 3399
rect 1370 3375 1390 3395
rect 1473 3379 1493 3399
rect 1581 3379 1601 3399
rect 1684 3375 1704 3395
rect 2511 3383 2531 3403
rect 2614 3379 2634 3399
rect 2722 3379 2742 3399
rect 2825 3383 2845 3403
rect 2940 3379 2960 3399
rect 3043 3383 3063 3403
rect 172 3241 190 3259
rect 4108 3303 4126 3321
rect 4106 3204 4124 3222
rect 170 3142 188 3160
rect 355 3147 375 3167
rect 458 3151 478 3171
rect 573 3147 593 3167
rect 676 3151 696 3171
rect 784 3151 804 3171
rect 887 3147 907 3167
rect 3390 3003 3410 3023
rect 3493 2999 3513 3019
rect 3601 2999 3621 3019
rect 3704 3003 3724 3023
rect 3819 2999 3839 3019
rect 3922 3003 3942 3023
rect 4109 3010 4127 3028
rect 173 2948 191 2966
rect 171 2849 189 2867
rect 4107 2911 4125 2929
rect 1234 2767 1254 2787
rect 1337 2771 1357 2791
rect 1452 2767 1472 2787
rect 1555 2771 1575 2791
rect 1663 2771 1683 2791
rect 1766 2767 1786 2787
rect 2593 2775 2613 2795
rect 2696 2771 2716 2791
rect 2804 2771 2824 2791
rect 2907 2775 2927 2795
rect 3022 2771 3042 2791
rect 3125 2775 3145 2795
rect 4102 2792 4120 2810
rect 4100 2693 4118 2711
rect 168 2624 186 2642
rect 3391 2591 3411 2611
rect 166 2525 184 2543
rect 337 2541 357 2561
rect 440 2545 460 2565
rect 555 2541 575 2561
rect 658 2545 678 2565
rect 766 2545 786 2565
rect 3494 2587 3514 2607
rect 3602 2587 3622 2607
rect 3705 2591 3725 2611
rect 3820 2587 3840 2607
rect 3923 2591 3943 2611
rect 4096 2609 4114 2627
rect 869 2541 889 2561
rect 4094 2510 4112 2528
rect 162 2441 180 2459
rect 160 2342 178 2360
rect 1135 2357 1155 2377
rect 1238 2361 1258 2381
rect 1353 2357 1373 2377
rect 1456 2361 1476 2381
rect 1564 2361 1584 2381
rect 1667 2357 1687 2377
rect 2428 2367 2448 2387
rect 2531 2363 2551 2383
rect 2639 2363 2659 2383
rect 2742 2367 2762 2387
rect 2857 2363 2877 2383
rect 2960 2367 2980 2387
rect 155 2223 173 2241
rect 4091 2285 4109 2303
rect 4089 2186 4107 2204
rect 153 2124 171 2142
rect 338 2129 358 2149
rect 441 2133 461 2153
rect 556 2129 576 2149
rect 659 2133 679 2153
rect 767 2133 787 2153
rect 870 2129 890 2149
rect 3370 1985 3390 2005
rect 3473 1981 3493 2001
rect 3581 1981 3601 2001
rect 3684 1985 3704 2005
rect 3799 1981 3819 2001
rect 3902 1985 3922 2005
rect 4089 1992 4107 2010
rect 153 1930 171 1948
rect 151 1831 169 1849
rect 4087 1893 4105 1911
rect 1280 1747 1300 1767
rect 1383 1751 1403 1771
rect 1498 1747 1518 1767
rect 1601 1751 1621 1771
rect 1709 1751 1729 1771
rect 1812 1747 1832 1767
rect 2573 1757 2593 1777
rect 2676 1753 2696 1773
rect 2784 1753 2804 1773
rect 2887 1757 2907 1777
rect 3002 1753 3022 1773
rect 3105 1757 3125 1777
rect 4082 1774 4100 1792
rect 4080 1675 4098 1693
rect 148 1606 166 1624
rect 3371 1573 3391 1593
rect 146 1507 164 1525
rect 317 1523 337 1543
rect 420 1527 440 1547
rect 535 1523 555 1543
rect 638 1527 658 1547
rect 746 1527 766 1547
rect 3474 1569 3494 1589
rect 3582 1569 3602 1589
rect 3685 1573 3705 1593
rect 3800 1569 3820 1589
rect 3903 1573 3923 1593
rect 4076 1591 4094 1609
rect 849 1523 869 1543
rect 4074 1492 4092 1510
rect 142 1423 160 1441
rect 140 1324 158 1342
rect 1115 1339 1135 1359
rect 1218 1343 1238 1363
rect 1333 1339 1353 1359
rect 1436 1343 1456 1363
rect 1544 1343 1564 1363
rect 1647 1339 1667 1359
rect 2474 1347 2494 1367
rect 2577 1343 2597 1363
rect 2685 1343 2705 1363
rect 2788 1347 2808 1367
rect 2903 1343 2923 1363
rect 3006 1347 3026 1367
rect 135 1205 153 1223
rect 4071 1267 4089 1285
rect 4069 1168 4087 1186
rect 133 1106 151 1124
rect 318 1111 338 1131
rect 421 1115 441 1135
rect 536 1111 556 1131
rect 639 1115 659 1135
rect 747 1115 767 1135
rect 850 1111 870 1131
rect 3353 967 3373 987
rect 3456 963 3476 983
rect 3564 963 3584 983
rect 3667 967 3687 987
rect 3782 963 3802 983
rect 3885 967 3905 987
rect 4072 974 4090 992
rect 136 912 154 930
rect 134 813 152 831
rect 4070 875 4088 893
rect 1197 731 1217 751
rect 1300 735 1320 755
rect 1415 731 1435 751
rect 1518 735 1538 755
rect 1626 735 1646 755
rect 1729 731 1749 751
rect 2556 739 2576 759
rect 2659 735 2679 755
rect 2767 735 2787 755
rect 2870 739 2890 759
rect 2985 735 3005 755
rect 3088 739 3108 759
rect 4065 756 4083 774
rect 4063 657 4081 675
rect 131 588 149 606
rect 3354 555 3374 575
rect 129 489 147 507
rect 300 505 320 525
rect 403 509 423 529
rect 518 505 538 525
rect 621 509 641 529
rect 729 509 749 529
rect 3457 551 3477 571
rect 3565 551 3585 571
rect 3668 555 3688 575
rect 3783 551 3803 571
rect 3886 555 3906 575
rect 4059 573 4077 591
rect 832 505 852 525
rect 4057 474 4075 492
rect 125 405 143 423
rect 123 306 141 324
rect 1098 321 1118 341
rect 1201 325 1221 345
rect 1316 321 1336 341
rect 1419 325 1439 345
rect 1527 325 1547 345
rect 1630 321 1650 341
rect 118 187 136 205
rect 4054 249 4072 267
rect 4052 150 4070 168
rect 116 88 134 106
rect 301 93 321 113
rect 404 97 424 117
rect 519 93 539 113
rect 622 97 642 117
rect 730 97 750 117
rect 833 93 853 113
rect 1514 -483 1534 -463
rect 1617 -479 1637 -459
rect 1732 -483 1752 -463
rect 1835 -479 1855 -459
rect 1943 -479 1963 -459
rect 2046 -483 2066 -463
<< pdiffc >>
rect 3486 7944 3506 7964
rect 3582 7944 3602 7964
rect 3692 7944 3712 7964
rect 3788 7944 3808 7964
rect 3910 7944 3930 7964
rect 4006 7944 4026 7964
rect 433 7780 453 7800
rect 529 7780 549 7800
rect 651 7780 671 7800
rect 747 7780 767 7800
rect 857 7780 877 7800
rect 953 7780 973 7800
rect 2689 7716 2709 7736
rect 2785 7716 2805 7736
rect 2895 7716 2915 7736
rect 2991 7716 3011 7736
rect 3113 7716 3133 7736
rect 3209 7716 3229 7736
rect 1231 7596 1251 7616
rect 1327 7596 1347 7616
rect 1449 7596 1469 7616
rect 1545 7596 1565 7616
rect 1655 7596 1675 7616
rect 1751 7596 1771 7616
rect 3487 7532 3507 7552
rect 3583 7532 3603 7552
rect 3693 7532 3713 7552
rect 3789 7532 3809 7552
rect 3911 7532 3931 7552
rect 4007 7532 4027 7552
rect 434 7368 454 7388
rect 530 7368 550 7388
rect 652 7368 672 7388
rect 748 7368 768 7388
rect 858 7368 878 7388
rect 954 7368 974 7388
rect 2590 7306 2610 7326
rect 2686 7306 2706 7326
rect 2796 7306 2816 7326
rect 2892 7306 2912 7326
rect 3014 7306 3034 7326
rect 3110 7306 3130 7326
rect 1313 6988 1333 7008
rect 1409 6988 1429 7008
rect 1531 6988 1551 7008
rect 1627 6988 1647 7008
rect 1737 6988 1757 7008
rect 1833 6988 1853 7008
rect 3469 6926 3489 6946
rect 3565 6926 3585 6946
rect 3675 6926 3695 6946
rect 3771 6926 3791 6946
rect 3893 6926 3913 6946
rect 3989 6926 4009 6946
rect 416 6762 436 6782
rect 512 6762 532 6782
rect 634 6762 654 6782
rect 730 6762 750 6782
rect 840 6762 860 6782
rect 936 6762 956 6782
rect 2672 6698 2692 6718
rect 2768 6698 2788 6718
rect 2878 6698 2898 6718
rect 2974 6698 2994 6718
rect 3096 6698 3116 6718
rect 3192 6698 3212 6718
rect 1214 6578 1234 6598
rect 1310 6578 1330 6598
rect 1432 6578 1452 6598
rect 1528 6578 1548 6598
rect 1638 6578 1658 6598
rect 1734 6578 1754 6598
rect 3470 6514 3490 6534
rect 3566 6514 3586 6534
rect 3676 6514 3696 6534
rect 3772 6514 3792 6534
rect 3894 6514 3914 6534
rect 3990 6514 4010 6534
rect 417 6350 437 6370
rect 513 6350 533 6370
rect 635 6350 655 6370
rect 731 6350 751 6370
rect 841 6350 861 6370
rect 937 6350 957 6370
rect 2507 6290 2527 6310
rect 2603 6290 2623 6310
rect 2713 6290 2733 6310
rect 2809 6290 2829 6310
rect 2931 6290 2951 6310
rect 3027 6290 3047 6310
rect 1359 5968 1379 5988
rect 1455 5968 1475 5988
rect 1577 5968 1597 5988
rect 1673 5968 1693 5988
rect 1783 5968 1803 5988
rect 1879 5968 1899 5988
rect 3449 5908 3469 5928
rect 3545 5908 3565 5928
rect 3655 5908 3675 5928
rect 3751 5908 3771 5928
rect 3873 5908 3893 5928
rect 3969 5908 3989 5928
rect 396 5744 416 5764
rect 492 5744 512 5764
rect 614 5744 634 5764
rect 710 5744 730 5764
rect 820 5744 840 5764
rect 916 5744 936 5764
rect 2652 5680 2672 5700
rect 2748 5680 2768 5700
rect 2858 5680 2878 5700
rect 2954 5680 2974 5700
rect 3076 5680 3096 5700
rect 3172 5680 3192 5700
rect 1194 5560 1214 5580
rect 1290 5560 1310 5580
rect 1412 5560 1432 5580
rect 1508 5560 1528 5580
rect 1618 5560 1638 5580
rect 1714 5560 1734 5580
rect 3450 5496 3470 5516
rect 3546 5496 3566 5516
rect 3656 5496 3676 5516
rect 3752 5496 3772 5516
rect 3874 5496 3894 5516
rect 3970 5496 3990 5516
rect 397 5332 417 5352
rect 493 5332 513 5352
rect 615 5332 635 5352
rect 711 5332 731 5352
rect 821 5332 841 5352
rect 917 5332 937 5352
rect 2553 5270 2573 5290
rect 2649 5270 2669 5290
rect 2759 5270 2779 5290
rect 2855 5270 2875 5290
rect 2977 5270 2997 5290
rect 3073 5270 3093 5290
rect 1276 4952 1296 4972
rect 1372 4952 1392 4972
rect 1494 4952 1514 4972
rect 1590 4952 1610 4972
rect 1700 4952 1720 4972
rect 1796 4952 1816 4972
rect 3432 4890 3452 4910
rect 3528 4890 3548 4910
rect 3638 4890 3658 4910
rect 3734 4890 3754 4910
rect 3856 4890 3876 4910
rect 3952 4890 3972 4910
rect 379 4726 399 4746
rect 475 4726 495 4746
rect 597 4726 617 4746
rect 693 4726 713 4746
rect 803 4726 823 4746
rect 899 4726 919 4746
rect 2635 4662 2655 4682
rect 2731 4662 2751 4682
rect 2841 4662 2861 4682
rect 2937 4662 2957 4682
rect 3059 4662 3079 4682
rect 3155 4662 3175 4682
rect 1177 4542 1197 4562
rect 1273 4542 1293 4562
rect 1395 4542 1415 4562
rect 1491 4542 1511 4562
rect 1601 4542 1621 4562
rect 1697 4542 1717 4562
rect 3433 4478 3453 4498
rect 3529 4478 3549 4498
rect 3639 4478 3659 4498
rect 3735 4478 3755 4498
rect 3857 4478 3877 4498
rect 3953 4478 3973 4498
rect 380 4314 400 4334
rect 476 4314 496 4334
rect 598 4314 618 4334
rect 694 4314 714 4334
rect 804 4314 824 4334
rect 900 4314 920 4334
rect 2331 4256 2351 4276
rect 2427 4256 2447 4276
rect 2537 4256 2557 4276
rect 2633 4256 2653 4276
rect 2755 4256 2775 4276
rect 2851 4256 2871 4276
rect 1462 3930 1482 3950
rect 1558 3930 1578 3950
rect 1680 3930 1700 3950
rect 1776 3930 1796 3950
rect 1886 3930 1906 3950
rect 1982 3930 2002 3950
rect 3413 3872 3433 3892
rect 3509 3872 3529 3892
rect 3619 3872 3639 3892
rect 3715 3872 3735 3892
rect 3837 3872 3857 3892
rect 3933 3872 3953 3892
rect 360 3708 380 3728
rect 456 3708 476 3728
rect 578 3708 598 3728
rect 674 3708 694 3728
rect 784 3708 804 3728
rect 880 3708 900 3728
rect 2616 3644 2636 3664
rect 2712 3644 2732 3664
rect 2822 3644 2842 3664
rect 2918 3644 2938 3664
rect 3040 3644 3060 3664
rect 3136 3644 3156 3664
rect 1158 3524 1178 3544
rect 1254 3524 1274 3544
rect 1376 3524 1396 3544
rect 1472 3524 1492 3544
rect 1582 3524 1602 3544
rect 1678 3524 1698 3544
rect 3414 3460 3434 3480
rect 3510 3460 3530 3480
rect 3620 3460 3640 3480
rect 3716 3460 3736 3480
rect 3838 3460 3858 3480
rect 3934 3460 3954 3480
rect 361 3296 381 3316
rect 457 3296 477 3316
rect 579 3296 599 3316
rect 675 3296 695 3316
rect 785 3296 805 3316
rect 881 3296 901 3316
rect 2517 3234 2537 3254
rect 2613 3234 2633 3254
rect 2723 3234 2743 3254
rect 2819 3234 2839 3254
rect 2941 3234 2961 3254
rect 3037 3234 3057 3254
rect 1240 2916 1260 2936
rect 1336 2916 1356 2936
rect 1458 2916 1478 2936
rect 1554 2916 1574 2936
rect 1664 2916 1684 2936
rect 1760 2916 1780 2936
rect 3396 2854 3416 2874
rect 3492 2854 3512 2874
rect 3602 2854 3622 2874
rect 3698 2854 3718 2874
rect 3820 2854 3840 2874
rect 3916 2854 3936 2874
rect 343 2690 363 2710
rect 439 2690 459 2710
rect 561 2690 581 2710
rect 657 2690 677 2710
rect 767 2690 787 2710
rect 863 2690 883 2710
rect 2599 2626 2619 2646
rect 2695 2626 2715 2646
rect 2805 2626 2825 2646
rect 2901 2626 2921 2646
rect 3023 2626 3043 2646
rect 3119 2626 3139 2646
rect 1141 2506 1161 2526
rect 1237 2506 1257 2526
rect 1359 2506 1379 2526
rect 1455 2506 1475 2526
rect 1565 2506 1585 2526
rect 1661 2506 1681 2526
rect 3397 2442 3417 2462
rect 3493 2442 3513 2462
rect 3603 2442 3623 2462
rect 3699 2442 3719 2462
rect 3821 2442 3841 2462
rect 3917 2442 3937 2462
rect 344 2278 364 2298
rect 440 2278 460 2298
rect 562 2278 582 2298
rect 658 2278 678 2298
rect 768 2278 788 2298
rect 864 2278 884 2298
rect 2434 2218 2454 2238
rect 2530 2218 2550 2238
rect 2640 2218 2660 2238
rect 2736 2218 2756 2238
rect 2858 2218 2878 2238
rect 2954 2218 2974 2238
rect 1286 1896 1306 1916
rect 1382 1896 1402 1916
rect 1504 1896 1524 1916
rect 1600 1896 1620 1916
rect 1710 1896 1730 1916
rect 1806 1896 1826 1916
rect 3376 1836 3396 1856
rect 3472 1836 3492 1856
rect 3582 1836 3602 1856
rect 3678 1836 3698 1856
rect 3800 1836 3820 1856
rect 3896 1836 3916 1856
rect 323 1672 343 1692
rect 419 1672 439 1692
rect 541 1672 561 1692
rect 637 1672 657 1692
rect 747 1672 767 1692
rect 843 1672 863 1692
rect 2579 1608 2599 1628
rect 2675 1608 2695 1628
rect 2785 1608 2805 1628
rect 2881 1608 2901 1628
rect 3003 1608 3023 1628
rect 3099 1608 3119 1628
rect 1121 1488 1141 1508
rect 1217 1488 1237 1508
rect 1339 1488 1359 1508
rect 1435 1488 1455 1508
rect 1545 1488 1565 1508
rect 1641 1488 1661 1508
rect 3377 1424 3397 1444
rect 3473 1424 3493 1444
rect 3583 1424 3603 1444
rect 3679 1424 3699 1444
rect 3801 1424 3821 1444
rect 3897 1424 3917 1444
rect 324 1260 344 1280
rect 420 1260 440 1280
rect 542 1260 562 1280
rect 638 1260 658 1280
rect 748 1260 768 1280
rect 844 1260 864 1280
rect 2480 1198 2500 1218
rect 2576 1198 2596 1218
rect 2686 1198 2706 1218
rect 2782 1198 2802 1218
rect 2904 1198 2924 1218
rect 3000 1198 3020 1218
rect 1203 880 1223 900
rect 1299 880 1319 900
rect 1421 880 1441 900
rect 1517 880 1537 900
rect 1627 880 1647 900
rect 1723 880 1743 900
rect 3359 818 3379 838
rect 3455 818 3475 838
rect 3565 818 3585 838
rect 3661 818 3681 838
rect 3783 818 3803 838
rect 3879 818 3899 838
rect 306 654 326 674
rect 402 654 422 674
rect 524 654 544 674
rect 620 654 640 674
rect 730 654 750 674
rect 826 654 846 674
rect 2562 590 2582 610
rect 2658 590 2678 610
rect 2768 590 2788 610
rect 2864 590 2884 610
rect 2986 590 3006 610
rect 3082 590 3102 610
rect 1104 470 1124 490
rect 1200 470 1220 490
rect 1322 470 1342 490
rect 1418 470 1438 490
rect 1528 470 1548 490
rect 1624 470 1644 490
rect 3360 406 3380 426
rect 3456 406 3476 426
rect 3566 406 3586 426
rect 3662 406 3682 426
rect 3784 406 3804 426
rect 3880 406 3900 426
rect 307 242 327 262
rect 403 242 423 262
rect 525 242 545 262
rect 621 242 641 262
rect 731 242 751 262
rect 827 242 847 262
rect 1520 -334 1540 -314
rect 1616 -334 1636 -314
rect 1738 -334 1758 -314
rect 1834 -334 1854 -314
rect 1944 -334 1964 -314
rect 2040 -334 2060 -314
<< poly >>
rect 3518 8125 3568 8141
rect 3726 8125 3776 8141
rect 3944 8125 3994 8141
rect 3518 8053 3568 8083
rect 3518 8033 3525 8053
rect 3545 8033 3568 8053
rect 3518 8006 3568 8033
rect 3726 8051 3776 8083
rect 3726 8031 3743 8051
rect 3763 8031 3776 8051
rect 3726 8006 3776 8031
rect 3944 8054 3994 8083
rect 3944 8034 3961 8054
rect 3981 8034 3994 8054
rect 3944 8006 3994 8034
rect 2721 7897 2771 7913
rect 2929 7897 2979 7913
rect 3147 7897 3197 7913
rect 3518 7893 3568 7906
rect 3726 7893 3776 7906
rect 3944 7893 3994 7906
rect 465 7838 515 7851
rect 683 7838 733 7851
rect 891 7838 941 7851
rect 2721 7825 2771 7855
rect 2721 7805 2728 7825
rect 2748 7805 2771 7825
rect 2721 7778 2771 7805
rect 2929 7823 2979 7855
rect 2929 7803 2946 7823
rect 2966 7803 2979 7823
rect 2929 7778 2979 7803
rect 3147 7826 3197 7855
rect 3147 7806 3164 7826
rect 3184 7806 3197 7826
rect 3147 7778 3197 7806
rect 465 7710 515 7738
rect 465 7690 478 7710
rect 498 7690 515 7710
rect 465 7661 515 7690
rect 683 7713 733 7738
rect 683 7693 696 7713
rect 716 7693 733 7713
rect 683 7661 733 7693
rect 891 7711 941 7738
rect 891 7691 914 7711
rect 934 7691 941 7711
rect 891 7661 941 7691
rect 3519 7713 3569 7729
rect 3727 7713 3777 7729
rect 3945 7713 3995 7729
rect 1263 7654 1313 7667
rect 1481 7654 1531 7667
rect 1689 7654 1739 7667
rect 2721 7665 2771 7678
rect 2929 7665 2979 7678
rect 3147 7665 3197 7678
rect 465 7603 515 7619
rect 683 7603 733 7619
rect 891 7603 941 7619
rect 3519 7641 3569 7671
rect 3519 7621 3526 7641
rect 3546 7621 3569 7641
rect 3519 7594 3569 7621
rect 3727 7639 3777 7671
rect 3727 7619 3744 7639
rect 3764 7619 3777 7639
rect 3727 7594 3777 7619
rect 3945 7642 3995 7671
rect 3945 7622 3962 7642
rect 3982 7622 3995 7642
rect 3945 7594 3995 7622
rect 1263 7526 1313 7554
rect 1263 7506 1276 7526
rect 1296 7506 1313 7526
rect 1263 7477 1313 7506
rect 1481 7529 1531 7554
rect 1481 7509 1494 7529
rect 1514 7509 1531 7529
rect 1481 7477 1531 7509
rect 1689 7527 1739 7554
rect 1689 7507 1712 7527
rect 1732 7507 1739 7527
rect 1689 7477 1739 7507
rect 2622 7487 2672 7503
rect 2830 7487 2880 7503
rect 3048 7487 3098 7503
rect 466 7426 516 7439
rect 684 7426 734 7439
rect 892 7426 942 7439
rect 3519 7481 3569 7494
rect 3727 7481 3777 7494
rect 3945 7481 3995 7494
rect 1263 7419 1313 7435
rect 1481 7419 1531 7435
rect 1689 7419 1739 7435
rect 2622 7415 2672 7445
rect 2622 7395 2629 7415
rect 2649 7395 2672 7415
rect 2622 7368 2672 7395
rect 2830 7413 2880 7445
rect 2830 7393 2847 7413
rect 2867 7393 2880 7413
rect 2830 7368 2880 7393
rect 3048 7416 3098 7445
rect 3048 7396 3065 7416
rect 3085 7396 3098 7416
rect 3048 7368 3098 7396
rect 466 7298 516 7326
rect 466 7278 479 7298
rect 499 7278 516 7298
rect 466 7249 516 7278
rect 684 7301 734 7326
rect 684 7281 697 7301
rect 717 7281 734 7301
rect 684 7249 734 7281
rect 892 7299 942 7326
rect 892 7279 915 7299
rect 935 7279 942 7299
rect 892 7249 942 7279
rect 2622 7255 2672 7268
rect 2830 7255 2880 7268
rect 3048 7255 3098 7268
rect 466 7191 516 7207
rect 684 7191 734 7207
rect 892 7191 942 7207
rect 3501 7107 3551 7123
rect 3709 7107 3759 7123
rect 3927 7107 3977 7123
rect 1345 7046 1395 7059
rect 1563 7046 1613 7059
rect 1771 7046 1821 7059
rect 3501 7035 3551 7065
rect 3501 7015 3508 7035
rect 3528 7015 3551 7035
rect 3501 6988 3551 7015
rect 3709 7033 3759 7065
rect 3709 7013 3726 7033
rect 3746 7013 3759 7033
rect 3709 6988 3759 7013
rect 3927 7036 3977 7065
rect 3927 7016 3944 7036
rect 3964 7016 3977 7036
rect 3927 6988 3977 7016
rect 1345 6918 1395 6946
rect 1345 6898 1358 6918
rect 1378 6898 1395 6918
rect 1345 6869 1395 6898
rect 1563 6921 1613 6946
rect 1563 6901 1576 6921
rect 1596 6901 1613 6921
rect 1563 6869 1613 6901
rect 1771 6919 1821 6946
rect 1771 6899 1794 6919
rect 1814 6899 1821 6919
rect 1771 6869 1821 6899
rect 2704 6879 2754 6895
rect 2912 6879 2962 6895
rect 3130 6879 3180 6895
rect 448 6820 498 6833
rect 666 6820 716 6833
rect 874 6820 924 6833
rect 3501 6875 3551 6888
rect 3709 6875 3759 6888
rect 3927 6875 3977 6888
rect 1345 6811 1395 6827
rect 1563 6811 1613 6827
rect 1771 6811 1821 6827
rect 2704 6807 2754 6837
rect 2704 6787 2711 6807
rect 2731 6787 2754 6807
rect 2704 6760 2754 6787
rect 2912 6805 2962 6837
rect 2912 6785 2929 6805
rect 2949 6785 2962 6805
rect 2912 6760 2962 6785
rect 3130 6808 3180 6837
rect 3130 6788 3147 6808
rect 3167 6788 3180 6808
rect 3130 6760 3180 6788
rect 448 6692 498 6720
rect 448 6672 461 6692
rect 481 6672 498 6692
rect 448 6643 498 6672
rect 666 6695 716 6720
rect 666 6675 679 6695
rect 699 6675 716 6695
rect 666 6643 716 6675
rect 874 6693 924 6720
rect 874 6673 897 6693
rect 917 6673 924 6693
rect 874 6643 924 6673
rect 3502 6695 3552 6711
rect 3710 6695 3760 6711
rect 3928 6695 3978 6711
rect 1246 6636 1296 6649
rect 1464 6636 1514 6649
rect 1672 6636 1722 6649
rect 2704 6647 2754 6660
rect 2912 6647 2962 6660
rect 3130 6647 3180 6660
rect 448 6585 498 6601
rect 666 6585 716 6601
rect 874 6585 924 6601
rect 3502 6623 3552 6653
rect 3502 6603 3509 6623
rect 3529 6603 3552 6623
rect 3502 6576 3552 6603
rect 3710 6621 3760 6653
rect 3710 6601 3727 6621
rect 3747 6601 3760 6621
rect 3710 6576 3760 6601
rect 3928 6624 3978 6653
rect 3928 6604 3945 6624
rect 3965 6604 3978 6624
rect 3928 6576 3978 6604
rect 1246 6508 1296 6536
rect 1246 6488 1259 6508
rect 1279 6488 1296 6508
rect 1246 6459 1296 6488
rect 1464 6511 1514 6536
rect 1464 6491 1477 6511
rect 1497 6491 1514 6511
rect 1464 6459 1514 6491
rect 1672 6509 1722 6536
rect 1672 6489 1695 6509
rect 1715 6489 1722 6509
rect 1672 6459 1722 6489
rect 2539 6471 2589 6487
rect 2747 6471 2797 6487
rect 2965 6471 3015 6487
rect 449 6408 499 6421
rect 667 6408 717 6421
rect 875 6408 925 6421
rect 3502 6463 3552 6476
rect 3710 6463 3760 6476
rect 3928 6463 3978 6476
rect 1246 6401 1296 6417
rect 1464 6401 1514 6417
rect 1672 6401 1722 6417
rect 2539 6399 2589 6429
rect 2539 6379 2546 6399
rect 2566 6379 2589 6399
rect 2539 6352 2589 6379
rect 2747 6397 2797 6429
rect 2747 6377 2764 6397
rect 2784 6377 2797 6397
rect 2747 6352 2797 6377
rect 2965 6400 3015 6429
rect 2965 6380 2982 6400
rect 3002 6380 3015 6400
rect 2965 6352 3015 6380
rect 449 6280 499 6308
rect 449 6260 462 6280
rect 482 6260 499 6280
rect 449 6231 499 6260
rect 667 6283 717 6308
rect 667 6263 680 6283
rect 700 6263 717 6283
rect 667 6231 717 6263
rect 875 6281 925 6308
rect 875 6261 898 6281
rect 918 6261 925 6281
rect 875 6231 925 6261
rect 2539 6239 2589 6252
rect 2747 6239 2797 6252
rect 2965 6239 3015 6252
rect 449 6173 499 6189
rect 667 6173 717 6189
rect 875 6173 925 6189
rect 3481 6089 3531 6105
rect 3689 6089 3739 6105
rect 3907 6089 3957 6105
rect 1391 6026 1441 6039
rect 1609 6026 1659 6039
rect 1817 6026 1867 6039
rect 3481 6017 3531 6047
rect 3481 5997 3488 6017
rect 3508 5997 3531 6017
rect 3481 5970 3531 5997
rect 3689 6015 3739 6047
rect 3689 5995 3706 6015
rect 3726 5995 3739 6015
rect 3689 5970 3739 5995
rect 3907 6018 3957 6047
rect 3907 5998 3924 6018
rect 3944 5998 3957 6018
rect 3907 5970 3957 5998
rect 1391 5898 1441 5926
rect 1391 5878 1404 5898
rect 1424 5878 1441 5898
rect 1391 5849 1441 5878
rect 1609 5901 1659 5926
rect 1609 5881 1622 5901
rect 1642 5881 1659 5901
rect 1609 5849 1659 5881
rect 1817 5899 1867 5926
rect 1817 5879 1840 5899
rect 1860 5879 1867 5899
rect 1817 5849 1867 5879
rect 2684 5861 2734 5877
rect 2892 5861 2942 5877
rect 3110 5861 3160 5877
rect 428 5802 478 5815
rect 646 5802 696 5815
rect 854 5802 904 5815
rect 3481 5857 3531 5870
rect 3689 5857 3739 5870
rect 3907 5857 3957 5870
rect 1391 5791 1441 5807
rect 1609 5791 1659 5807
rect 1817 5791 1867 5807
rect 2684 5789 2734 5819
rect 2684 5769 2691 5789
rect 2711 5769 2734 5789
rect 2684 5742 2734 5769
rect 2892 5787 2942 5819
rect 2892 5767 2909 5787
rect 2929 5767 2942 5787
rect 2892 5742 2942 5767
rect 3110 5790 3160 5819
rect 3110 5770 3127 5790
rect 3147 5770 3160 5790
rect 3110 5742 3160 5770
rect 428 5674 478 5702
rect 428 5654 441 5674
rect 461 5654 478 5674
rect 428 5625 478 5654
rect 646 5677 696 5702
rect 646 5657 659 5677
rect 679 5657 696 5677
rect 646 5625 696 5657
rect 854 5675 904 5702
rect 854 5655 877 5675
rect 897 5655 904 5675
rect 854 5625 904 5655
rect 3482 5677 3532 5693
rect 3690 5677 3740 5693
rect 3908 5677 3958 5693
rect 1226 5618 1276 5631
rect 1444 5618 1494 5631
rect 1652 5618 1702 5631
rect 2684 5629 2734 5642
rect 2892 5629 2942 5642
rect 3110 5629 3160 5642
rect 428 5567 478 5583
rect 646 5567 696 5583
rect 854 5567 904 5583
rect 3482 5605 3532 5635
rect 3482 5585 3489 5605
rect 3509 5585 3532 5605
rect 3482 5558 3532 5585
rect 3690 5603 3740 5635
rect 3690 5583 3707 5603
rect 3727 5583 3740 5603
rect 3690 5558 3740 5583
rect 3908 5606 3958 5635
rect 3908 5586 3925 5606
rect 3945 5586 3958 5606
rect 3908 5558 3958 5586
rect 1226 5490 1276 5518
rect 1226 5470 1239 5490
rect 1259 5470 1276 5490
rect 1226 5441 1276 5470
rect 1444 5493 1494 5518
rect 1444 5473 1457 5493
rect 1477 5473 1494 5493
rect 1444 5441 1494 5473
rect 1652 5491 1702 5518
rect 1652 5471 1675 5491
rect 1695 5471 1702 5491
rect 1652 5441 1702 5471
rect 2585 5451 2635 5467
rect 2793 5451 2843 5467
rect 3011 5451 3061 5467
rect 429 5390 479 5403
rect 647 5390 697 5403
rect 855 5390 905 5403
rect 3482 5445 3532 5458
rect 3690 5445 3740 5458
rect 3908 5445 3958 5458
rect 1226 5383 1276 5399
rect 1444 5383 1494 5399
rect 1652 5383 1702 5399
rect 2585 5379 2635 5409
rect 2585 5359 2592 5379
rect 2612 5359 2635 5379
rect 2585 5332 2635 5359
rect 2793 5377 2843 5409
rect 2793 5357 2810 5377
rect 2830 5357 2843 5377
rect 2793 5332 2843 5357
rect 3011 5380 3061 5409
rect 3011 5360 3028 5380
rect 3048 5360 3061 5380
rect 3011 5332 3061 5360
rect 429 5262 479 5290
rect 429 5242 442 5262
rect 462 5242 479 5262
rect 429 5213 479 5242
rect 647 5265 697 5290
rect 647 5245 660 5265
rect 680 5245 697 5265
rect 647 5213 697 5245
rect 855 5263 905 5290
rect 855 5243 878 5263
rect 898 5243 905 5263
rect 855 5213 905 5243
rect 2585 5219 2635 5232
rect 2793 5219 2843 5232
rect 3011 5219 3061 5232
rect 429 5155 479 5171
rect 647 5155 697 5171
rect 855 5155 905 5171
rect 3464 5071 3514 5087
rect 3672 5071 3722 5087
rect 3890 5071 3940 5087
rect 1308 5010 1358 5023
rect 1526 5010 1576 5023
rect 1734 5010 1784 5023
rect 3464 4999 3514 5029
rect 3464 4979 3471 4999
rect 3491 4979 3514 4999
rect 3464 4952 3514 4979
rect 3672 4997 3722 5029
rect 3672 4977 3689 4997
rect 3709 4977 3722 4997
rect 3672 4952 3722 4977
rect 3890 5000 3940 5029
rect 3890 4980 3907 5000
rect 3927 4980 3940 5000
rect 3890 4952 3940 4980
rect 1308 4882 1358 4910
rect 1308 4862 1321 4882
rect 1341 4862 1358 4882
rect 1308 4833 1358 4862
rect 1526 4885 1576 4910
rect 1526 4865 1539 4885
rect 1559 4865 1576 4885
rect 1526 4833 1576 4865
rect 1734 4883 1784 4910
rect 1734 4863 1757 4883
rect 1777 4863 1784 4883
rect 1734 4833 1784 4863
rect 2667 4843 2717 4859
rect 2875 4843 2925 4859
rect 3093 4843 3143 4859
rect 411 4784 461 4797
rect 629 4784 679 4797
rect 837 4784 887 4797
rect 3464 4839 3514 4852
rect 3672 4839 3722 4852
rect 3890 4839 3940 4852
rect 1308 4775 1358 4791
rect 1526 4775 1576 4791
rect 1734 4775 1784 4791
rect 2667 4771 2717 4801
rect 2667 4751 2674 4771
rect 2694 4751 2717 4771
rect 2667 4724 2717 4751
rect 2875 4769 2925 4801
rect 2875 4749 2892 4769
rect 2912 4749 2925 4769
rect 2875 4724 2925 4749
rect 3093 4772 3143 4801
rect 3093 4752 3110 4772
rect 3130 4752 3143 4772
rect 3093 4724 3143 4752
rect 411 4656 461 4684
rect 411 4636 424 4656
rect 444 4636 461 4656
rect 411 4607 461 4636
rect 629 4659 679 4684
rect 629 4639 642 4659
rect 662 4639 679 4659
rect 629 4607 679 4639
rect 837 4657 887 4684
rect 837 4637 860 4657
rect 880 4637 887 4657
rect 837 4607 887 4637
rect 3465 4659 3515 4675
rect 3673 4659 3723 4675
rect 3891 4659 3941 4675
rect 1209 4600 1259 4613
rect 1427 4600 1477 4613
rect 1635 4600 1685 4613
rect 2667 4611 2717 4624
rect 2875 4611 2925 4624
rect 3093 4611 3143 4624
rect 411 4549 461 4565
rect 629 4549 679 4565
rect 837 4549 887 4565
rect 3465 4587 3515 4617
rect 3465 4567 3472 4587
rect 3492 4567 3515 4587
rect 3465 4540 3515 4567
rect 3673 4585 3723 4617
rect 3673 4565 3690 4585
rect 3710 4565 3723 4585
rect 3673 4540 3723 4565
rect 3891 4588 3941 4617
rect 3891 4568 3908 4588
rect 3928 4568 3941 4588
rect 3891 4540 3941 4568
rect 1209 4472 1259 4500
rect 1209 4452 1222 4472
rect 1242 4452 1259 4472
rect 1209 4423 1259 4452
rect 1427 4475 1477 4500
rect 1427 4455 1440 4475
rect 1460 4455 1477 4475
rect 1427 4423 1477 4455
rect 1635 4473 1685 4500
rect 1635 4453 1658 4473
rect 1678 4453 1685 4473
rect 1635 4423 1685 4453
rect 2363 4437 2413 4453
rect 2571 4437 2621 4453
rect 2789 4437 2839 4453
rect 412 4372 462 4385
rect 630 4372 680 4385
rect 838 4372 888 4385
rect 3465 4427 3515 4440
rect 3673 4427 3723 4440
rect 3891 4427 3941 4440
rect 1209 4365 1259 4381
rect 1427 4365 1477 4381
rect 1635 4365 1685 4381
rect 2363 4365 2413 4395
rect 2363 4345 2370 4365
rect 2390 4345 2413 4365
rect 2363 4318 2413 4345
rect 2571 4363 2621 4395
rect 2571 4343 2588 4363
rect 2608 4343 2621 4363
rect 2571 4318 2621 4343
rect 2789 4366 2839 4395
rect 2789 4346 2806 4366
rect 2826 4346 2839 4366
rect 2789 4318 2839 4346
rect 412 4244 462 4272
rect 412 4224 425 4244
rect 445 4224 462 4244
rect 412 4195 462 4224
rect 630 4247 680 4272
rect 630 4227 643 4247
rect 663 4227 680 4247
rect 630 4195 680 4227
rect 838 4245 888 4272
rect 838 4225 861 4245
rect 881 4225 888 4245
rect 838 4195 888 4225
rect 2363 4205 2413 4218
rect 2571 4205 2621 4218
rect 2789 4205 2839 4218
rect 412 4137 462 4153
rect 630 4137 680 4153
rect 838 4137 888 4153
rect 3445 4053 3495 4069
rect 3653 4053 3703 4069
rect 3871 4053 3921 4069
rect 1494 3988 1544 4001
rect 1712 3988 1762 4001
rect 1920 3988 1970 4001
rect 3445 3981 3495 4011
rect 3445 3961 3452 3981
rect 3472 3961 3495 3981
rect 3445 3934 3495 3961
rect 3653 3979 3703 4011
rect 3653 3959 3670 3979
rect 3690 3959 3703 3979
rect 3653 3934 3703 3959
rect 3871 3982 3921 4011
rect 3871 3962 3888 3982
rect 3908 3962 3921 3982
rect 3871 3934 3921 3962
rect 1494 3860 1544 3888
rect 1494 3840 1507 3860
rect 1527 3840 1544 3860
rect 1494 3811 1544 3840
rect 1712 3863 1762 3888
rect 1712 3843 1725 3863
rect 1745 3843 1762 3863
rect 1712 3811 1762 3843
rect 1920 3861 1970 3888
rect 1920 3841 1943 3861
rect 1963 3841 1970 3861
rect 1920 3811 1970 3841
rect 2648 3825 2698 3841
rect 2856 3825 2906 3841
rect 3074 3825 3124 3841
rect 392 3766 442 3779
rect 610 3766 660 3779
rect 818 3766 868 3779
rect 3445 3821 3495 3834
rect 3653 3821 3703 3834
rect 3871 3821 3921 3834
rect 1494 3753 1544 3769
rect 1712 3753 1762 3769
rect 1920 3753 1970 3769
rect 2648 3753 2698 3783
rect 2648 3733 2655 3753
rect 2675 3733 2698 3753
rect 2648 3706 2698 3733
rect 2856 3751 2906 3783
rect 2856 3731 2873 3751
rect 2893 3731 2906 3751
rect 2856 3706 2906 3731
rect 3074 3754 3124 3783
rect 3074 3734 3091 3754
rect 3111 3734 3124 3754
rect 3074 3706 3124 3734
rect 392 3638 442 3666
rect 392 3618 405 3638
rect 425 3618 442 3638
rect 392 3589 442 3618
rect 610 3641 660 3666
rect 610 3621 623 3641
rect 643 3621 660 3641
rect 610 3589 660 3621
rect 818 3639 868 3666
rect 818 3619 841 3639
rect 861 3619 868 3639
rect 818 3589 868 3619
rect 3446 3641 3496 3657
rect 3654 3641 3704 3657
rect 3872 3641 3922 3657
rect 1190 3582 1240 3595
rect 1408 3582 1458 3595
rect 1616 3582 1666 3595
rect 2648 3593 2698 3606
rect 2856 3593 2906 3606
rect 3074 3593 3124 3606
rect 392 3531 442 3547
rect 610 3531 660 3547
rect 818 3531 868 3547
rect 3446 3569 3496 3599
rect 3446 3549 3453 3569
rect 3473 3549 3496 3569
rect 3446 3522 3496 3549
rect 3654 3567 3704 3599
rect 3654 3547 3671 3567
rect 3691 3547 3704 3567
rect 3654 3522 3704 3547
rect 3872 3570 3922 3599
rect 3872 3550 3889 3570
rect 3909 3550 3922 3570
rect 3872 3522 3922 3550
rect 1190 3454 1240 3482
rect 1190 3434 1203 3454
rect 1223 3434 1240 3454
rect 1190 3405 1240 3434
rect 1408 3457 1458 3482
rect 1408 3437 1421 3457
rect 1441 3437 1458 3457
rect 1408 3405 1458 3437
rect 1616 3455 1666 3482
rect 1616 3435 1639 3455
rect 1659 3435 1666 3455
rect 1616 3405 1666 3435
rect 2549 3415 2599 3431
rect 2757 3415 2807 3431
rect 2975 3415 3025 3431
rect 393 3354 443 3367
rect 611 3354 661 3367
rect 819 3354 869 3367
rect 3446 3409 3496 3422
rect 3654 3409 3704 3422
rect 3872 3409 3922 3422
rect 1190 3347 1240 3363
rect 1408 3347 1458 3363
rect 1616 3347 1666 3363
rect 2549 3343 2599 3373
rect 2549 3323 2556 3343
rect 2576 3323 2599 3343
rect 2549 3296 2599 3323
rect 2757 3341 2807 3373
rect 2757 3321 2774 3341
rect 2794 3321 2807 3341
rect 2757 3296 2807 3321
rect 2975 3344 3025 3373
rect 2975 3324 2992 3344
rect 3012 3324 3025 3344
rect 2975 3296 3025 3324
rect 393 3226 443 3254
rect 393 3206 406 3226
rect 426 3206 443 3226
rect 393 3177 443 3206
rect 611 3229 661 3254
rect 611 3209 624 3229
rect 644 3209 661 3229
rect 611 3177 661 3209
rect 819 3227 869 3254
rect 819 3207 842 3227
rect 862 3207 869 3227
rect 819 3177 869 3207
rect 2549 3183 2599 3196
rect 2757 3183 2807 3196
rect 2975 3183 3025 3196
rect 393 3119 443 3135
rect 611 3119 661 3135
rect 819 3119 869 3135
rect 3428 3035 3478 3051
rect 3636 3035 3686 3051
rect 3854 3035 3904 3051
rect 1272 2974 1322 2987
rect 1490 2974 1540 2987
rect 1698 2974 1748 2987
rect 3428 2963 3478 2993
rect 3428 2943 3435 2963
rect 3455 2943 3478 2963
rect 3428 2916 3478 2943
rect 3636 2961 3686 2993
rect 3636 2941 3653 2961
rect 3673 2941 3686 2961
rect 3636 2916 3686 2941
rect 3854 2964 3904 2993
rect 3854 2944 3871 2964
rect 3891 2944 3904 2964
rect 3854 2916 3904 2944
rect 1272 2846 1322 2874
rect 1272 2826 1285 2846
rect 1305 2826 1322 2846
rect 1272 2797 1322 2826
rect 1490 2849 1540 2874
rect 1490 2829 1503 2849
rect 1523 2829 1540 2849
rect 1490 2797 1540 2829
rect 1698 2847 1748 2874
rect 1698 2827 1721 2847
rect 1741 2827 1748 2847
rect 1698 2797 1748 2827
rect 2631 2807 2681 2823
rect 2839 2807 2889 2823
rect 3057 2807 3107 2823
rect 375 2748 425 2761
rect 593 2748 643 2761
rect 801 2748 851 2761
rect 3428 2803 3478 2816
rect 3636 2803 3686 2816
rect 3854 2803 3904 2816
rect 1272 2739 1322 2755
rect 1490 2739 1540 2755
rect 1698 2739 1748 2755
rect 2631 2735 2681 2765
rect 2631 2715 2638 2735
rect 2658 2715 2681 2735
rect 2631 2688 2681 2715
rect 2839 2733 2889 2765
rect 2839 2713 2856 2733
rect 2876 2713 2889 2733
rect 2839 2688 2889 2713
rect 3057 2736 3107 2765
rect 3057 2716 3074 2736
rect 3094 2716 3107 2736
rect 3057 2688 3107 2716
rect 375 2620 425 2648
rect 375 2600 388 2620
rect 408 2600 425 2620
rect 375 2571 425 2600
rect 593 2623 643 2648
rect 593 2603 606 2623
rect 626 2603 643 2623
rect 593 2571 643 2603
rect 801 2621 851 2648
rect 801 2601 824 2621
rect 844 2601 851 2621
rect 801 2571 851 2601
rect 3429 2623 3479 2639
rect 3637 2623 3687 2639
rect 3855 2623 3905 2639
rect 1173 2564 1223 2577
rect 1391 2564 1441 2577
rect 1599 2564 1649 2577
rect 2631 2575 2681 2588
rect 2839 2575 2889 2588
rect 3057 2575 3107 2588
rect 375 2513 425 2529
rect 593 2513 643 2529
rect 801 2513 851 2529
rect 3429 2551 3479 2581
rect 3429 2531 3436 2551
rect 3456 2531 3479 2551
rect 3429 2504 3479 2531
rect 3637 2549 3687 2581
rect 3637 2529 3654 2549
rect 3674 2529 3687 2549
rect 3637 2504 3687 2529
rect 3855 2552 3905 2581
rect 3855 2532 3872 2552
rect 3892 2532 3905 2552
rect 3855 2504 3905 2532
rect 1173 2436 1223 2464
rect 1173 2416 1186 2436
rect 1206 2416 1223 2436
rect 1173 2387 1223 2416
rect 1391 2439 1441 2464
rect 1391 2419 1404 2439
rect 1424 2419 1441 2439
rect 1391 2387 1441 2419
rect 1599 2437 1649 2464
rect 1599 2417 1622 2437
rect 1642 2417 1649 2437
rect 1599 2387 1649 2417
rect 2466 2399 2516 2415
rect 2674 2399 2724 2415
rect 2892 2399 2942 2415
rect 376 2336 426 2349
rect 594 2336 644 2349
rect 802 2336 852 2349
rect 3429 2391 3479 2404
rect 3637 2391 3687 2404
rect 3855 2391 3905 2404
rect 1173 2329 1223 2345
rect 1391 2329 1441 2345
rect 1599 2329 1649 2345
rect 2466 2327 2516 2357
rect 2466 2307 2473 2327
rect 2493 2307 2516 2327
rect 2466 2280 2516 2307
rect 2674 2325 2724 2357
rect 2674 2305 2691 2325
rect 2711 2305 2724 2325
rect 2674 2280 2724 2305
rect 2892 2328 2942 2357
rect 2892 2308 2909 2328
rect 2929 2308 2942 2328
rect 2892 2280 2942 2308
rect 376 2208 426 2236
rect 376 2188 389 2208
rect 409 2188 426 2208
rect 376 2159 426 2188
rect 594 2211 644 2236
rect 594 2191 607 2211
rect 627 2191 644 2211
rect 594 2159 644 2191
rect 802 2209 852 2236
rect 802 2189 825 2209
rect 845 2189 852 2209
rect 802 2159 852 2189
rect 2466 2167 2516 2180
rect 2674 2167 2724 2180
rect 2892 2167 2942 2180
rect 376 2101 426 2117
rect 594 2101 644 2117
rect 802 2101 852 2117
rect 3408 2017 3458 2033
rect 3616 2017 3666 2033
rect 3834 2017 3884 2033
rect 1318 1954 1368 1967
rect 1536 1954 1586 1967
rect 1744 1954 1794 1967
rect 3408 1945 3458 1975
rect 3408 1925 3415 1945
rect 3435 1925 3458 1945
rect 3408 1898 3458 1925
rect 3616 1943 3666 1975
rect 3616 1923 3633 1943
rect 3653 1923 3666 1943
rect 3616 1898 3666 1923
rect 3834 1946 3884 1975
rect 3834 1926 3851 1946
rect 3871 1926 3884 1946
rect 3834 1898 3884 1926
rect 1318 1826 1368 1854
rect 1318 1806 1331 1826
rect 1351 1806 1368 1826
rect 1318 1777 1368 1806
rect 1536 1829 1586 1854
rect 1536 1809 1549 1829
rect 1569 1809 1586 1829
rect 1536 1777 1586 1809
rect 1744 1827 1794 1854
rect 1744 1807 1767 1827
rect 1787 1807 1794 1827
rect 1744 1777 1794 1807
rect 2611 1789 2661 1805
rect 2819 1789 2869 1805
rect 3037 1789 3087 1805
rect 355 1730 405 1743
rect 573 1730 623 1743
rect 781 1730 831 1743
rect 3408 1785 3458 1798
rect 3616 1785 3666 1798
rect 3834 1785 3884 1798
rect 1318 1719 1368 1735
rect 1536 1719 1586 1735
rect 1744 1719 1794 1735
rect 2611 1717 2661 1747
rect 2611 1697 2618 1717
rect 2638 1697 2661 1717
rect 2611 1670 2661 1697
rect 2819 1715 2869 1747
rect 2819 1695 2836 1715
rect 2856 1695 2869 1715
rect 2819 1670 2869 1695
rect 3037 1718 3087 1747
rect 3037 1698 3054 1718
rect 3074 1698 3087 1718
rect 3037 1670 3087 1698
rect 355 1602 405 1630
rect 355 1582 368 1602
rect 388 1582 405 1602
rect 355 1553 405 1582
rect 573 1605 623 1630
rect 573 1585 586 1605
rect 606 1585 623 1605
rect 573 1553 623 1585
rect 781 1603 831 1630
rect 781 1583 804 1603
rect 824 1583 831 1603
rect 781 1553 831 1583
rect 3409 1605 3459 1621
rect 3617 1605 3667 1621
rect 3835 1605 3885 1621
rect 1153 1546 1203 1559
rect 1371 1546 1421 1559
rect 1579 1546 1629 1559
rect 2611 1557 2661 1570
rect 2819 1557 2869 1570
rect 3037 1557 3087 1570
rect 355 1495 405 1511
rect 573 1495 623 1511
rect 781 1495 831 1511
rect 3409 1533 3459 1563
rect 3409 1513 3416 1533
rect 3436 1513 3459 1533
rect 3409 1486 3459 1513
rect 3617 1531 3667 1563
rect 3617 1511 3634 1531
rect 3654 1511 3667 1531
rect 3617 1486 3667 1511
rect 3835 1534 3885 1563
rect 3835 1514 3852 1534
rect 3872 1514 3885 1534
rect 3835 1486 3885 1514
rect 1153 1418 1203 1446
rect 1153 1398 1166 1418
rect 1186 1398 1203 1418
rect 1153 1369 1203 1398
rect 1371 1421 1421 1446
rect 1371 1401 1384 1421
rect 1404 1401 1421 1421
rect 1371 1369 1421 1401
rect 1579 1419 1629 1446
rect 1579 1399 1602 1419
rect 1622 1399 1629 1419
rect 1579 1369 1629 1399
rect 2512 1379 2562 1395
rect 2720 1379 2770 1395
rect 2938 1379 2988 1395
rect 356 1318 406 1331
rect 574 1318 624 1331
rect 782 1318 832 1331
rect 3409 1373 3459 1386
rect 3617 1373 3667 1386
rect 3835 1373 3885 1386
rect 1153 1311 1203 1327
rect 1371 1311 1421 1327
rect 1579 1311 1629 1327
rect 2512 1307 2562 1337
rect 2512 1287 2519 1307
rect 2539 1287 2562 1307
rect 2512 1260 2562 1287
rect 2720 1305 2770 1337
rect 2720 1285 2737 1305
rect 2757 1285 2770 1305
rect 2720 1260 2770 1285
rect 2938 1308 2988 1337
rect 2938 1288 2955 1308
rect 2975 1288 2988 1308
rect 2938 1260 2988 1288
rect 356 1190 406 1218
rect 356 1170 369 1190
rect 389 1170 406 1190
rect 356 1141 406 1170
rect 574 1193 624 1218
rect 574 1173 587 1193
rect 607 1173 624 1193
rect 574 1141 624 1173
rect 782 1191 832 1218
rect 782 1171 805 1191
rect 825 1171 832 1191
rect 782 1141 832 1171
rect 2512 1147 2562 1160
rect 2720 1147 2770 1160
rect 2938 1147 2988 1160
rect 356 1083 406 1099
rect 574 1083 624 1099
rect 782 1083 832 1099
rect 3391 999 3441 1015
rect 3599 999 3649 1015
rect 3817 999 3867 1015
rect 1235 938 1285 951
rect 1453 938 1503 951
rect 1661 938 1711 951
rect 3391 927 3441 957
rect 3391 907 3398 927
rect 3418 907 3441 927
rect 3391 880 3441 907
rect 3599 925 3649 957
rect 3599 905 3616 925
rect 3636 905 3649 925
rect 3599 880 3649 905
rect 3817 928 3867 957
rect 3817 908 3834 928
rect 3854 908 3867 928
rect 3817 880 3867 908
rect 1235 810 1285 838
rect 1235 790 1248 810
rect 1268 790 1285 810
rect 1235 761 1285 790
rect 1453 813 1503 838
rect 1453 793 1466 813
rect 1486 793 1503 813
rect 1453 761 1503 793
rect 1661 811 1711 838
rect 1661 791 1684 811
rect 1704 791 1711 811
rect 1661 761 1711 791
rect 2594 771 2644 787
rect 2802 771 2852 787
rect 3020 771 3070 787
rect 338 712 388 725
rect 556 712 606 725
rect 764 712 814 725
rect 3391 767 3441 780
rect 3599 767 3649 780
rect 3817 767 3867 780
rect 1235 703 1285 719
rect 1453 703 1503 719
rect 1661 703 1711 719
rect 2594 699 2644 729
rect 2594 679 2601 699
rect 2621 679 2644 699
rect 2594 652 2644 679
rect 2802 697 2852 729
rect 2802 677 2819 697
rect 2839 677 2852 697
rect 2802 652 2852 677
rect 3020 700 3070 729
rect 3020 680 3037 700
rect 3057 680 3070 700
rect 3020 652 3070 680
rect 338 584 388 612
rect 338 564 351 584
rect 371 564 388 584
rect 338 535 388 564
rect 556 587 606 612
rect 556 567 569 587
rect 589 567 606 587
rect 556 535 606 567
rect 764 585 814 612
rect 764 565 787 585
rect 807 565 814 585
rect 764 535 814 565
rect 3392 587 3442 603
rect 3600 587 3650 603
rect 3818 587 3868 603
rect 1136 528 1186 541
rect 1354 528 1404 541
rect 1562 528 1612 541
rect 2594 539 2644 552
rect 2802 539 2852 552
rect 3020 539 3070 552
rect 338 477 388 493
rect 556 477 606 493
rect 764 477 814 493
rect 3392 515 3442 545
rect 3392 495 3399 515
rect 3419 495 3442 515
rect 3392 468 3442 495
rect 3600 513 3650 545
rect 3600 493 3617 513
rect 3637 493 3650 513
rect 3600 468 3650 493
rect 3818 516 3868 545
rect 3818 496 3835 516
rect 3855 496 3868 516
rect 3818 468 3868 496
rect 1136 400 1186 428
rect 1136 380 1149 400
rect 1169 380 1186 400
rect 1136 351 1186 380
rect 1354 403 1404 428
rect 1354 383 1367 403
rect 1387 383 1404 403
rect 1354 351 1404 383
rect 1562 401 1612 428
rect 1562 381 1585 401
rect 1605 381 1612 401
rect 1562 351 1612 381
rect 3392 355 3442 368
rect 3600 355 3650 368
rect 3818 355 3868 368
rect 339 300 389 313
rect 557 300 607 313
rect 765 300 815 313
rect 1136 293 1186 309
rect 1354 293 1404 309
rect 1562 293 1612 309
rect 339 172 389 200
rect 339 152 352 172
rect 372 152 389 172
rect 339 123 389 152
rect 557 175 607 200
rect 557 155 570 175
rect 590 155 607 175
rect 557 123 607 155
rect 765 173 815 200
rect 765 153 788 173
rect 808 153 815 173
rect 765 123 815 153
rect 339 65 389 81
rect 557 65 607 81
rect 765 65 815 81
rect 1552 -276 1602 -263
rect 1770 -276 1820 -263
rect 1978 -276 2028 -263
rect 1552 -404 1602 -376
rect 1552 -424 1565 -404
rect 1585 -424 1602 -404
rect 1552 -453 1602 -424
rect 1770 -401 1820 -376
rect 1770 -421 1783 -401
rect 1803 -421 1820 -401
rect 1770 -453 1820 -421
rect 1978 -403 2028 -376
rect 1978 -423 2001 -403
rect 2021 -423 2028 -403
rect 1978 -453 2028 -423
rect 1552 -511 1602 -495
rect 1770 -511 1820 -495
rect 1978 -511 2028 -495
<< polycont >>
rect 3525 8033 3545 8053
rect 3743 8031 3763 8051
rect 3961 8034 3981 8054
rect 2728 7805 2748 7825
rect 2946 7803 2966 7823
rect 3164 7806 3184 7826
rect 478 7690 498 7710
rect 696 7693 716 7713
rect 914 7691 934 7711
rect 3526 7621 3546 7641
rect 3744 7619 3764 7639
rect 3962 7622 3982 7642
rect 1276 7506 1296 7526
rect 1494 7509 1514 7529
rect 1712 7507 1732 7527
rect 2629 7395 2649 7415
rect 2847 7393 2867 7413
rect 3065 7396 3085 7416
rect 479 7278 499 7298
rect 697 7281 717 7301
rect 915 7279 935 7299
rect 3508 7015 3528 7035
rect 3726 7013 3746 7033
rect 3944 7016 3964 7036
rect 1358 6898 1378 6918
rect 1576 6901 1596 6921
rect 1794 6899 1814 6919
rect 2711 6787 2731 6807
rect 2929 6785 2949 6805
rect 3147 6788 3167 6808
rect 461 6672 481 6692
rect 679 6675 699 6695
rect 897 6673 917 6693
rect 3509 6603 3529 6623
rect 3727 6601 3747 6621
rect 3945 6604 3965 6624
rect 1259 6488 1279 6508
rect 1477 6491 1497 6511
rect 1695 6489 1715 6509
rect 2546 6379 2566 6399
rect 2764 6377 2784 6397
rect 2982 6380 3002 6400
rect 462 6260 482 6280
rect 680 6263 700 6283
rect 898 6261 918 6281
rect 3488 5997 3508 6017
rect 3706 5995 3726 6015
rect 3924 5998 3944 6018
rect 1404 5878 1424 5898
rect 1622 5881 1642 5901
rect 1840 5879 1860 5899
rect 2691 5769 2711 5789
rect 2909 5767 2929 5787
rect 3127 5770 3147 5790
rect 441 5654 461 5674
rect 659 5657 679 5677
rect 877 5655 897 5675
rect 3489 5585 3509 5605
rect 3707 5583 3727 5603
rect 3925 5586 3945 5606
rect 1239 5470 1259 5490
rect 1457 5473 1477 5493
rect 1675 5471 1695 5491
rect 2592 5359 2612 5379
rect 2810 5357 2830 5377
rect 3028 5360 3048 5380
rect 442 5242 462 5262
rect 660 5245 680 5265
rect 878 5243 898 5263
rect 3471 4979 3491 4999
rect 3689 4977 3709 4997
rect 3907 4980 3927 5000
rect 1321 4862 1341 4882
rect 1539 4865 1559 4885
rect 1757 4863 1777 4883
rect 2674 4751 2694 4771
rect 2892 4749 2912 4769
rect 3110 4752 3130 4772
rect 424 4636 444 4656
rect 642 4639 662 4659
rect 860 4637 880 4657
rect 3472 4567 3492 4587
rect 3690 4565 3710 4585
rect 3908 4568 3928 4588
rect 1222 4452 1242 4472
rect 1440 4455 1460 4475
rect 1658 4453 1678 4473
rect 2370 4345 2390 4365
rect 2588 4343 2608 4363
rect 2806 4346 2826 4366
rect 425 4224 445 4244
rect 643 4227 663 4247
rect 861 4225 881 4245
rect 3452 3961 3472 3981
rect 3670 3959 3690 3979
rect 3888 3962 3908 3982
rect 1507 3840 1527 3860
rect 1725 3843 1745 3863
rect 1943 3841 1963 3861
rect 2655 3733 2675 3753
rect 2873 3731 2893 3751
rect 3091 3734 3111 3754
rect 405 3618 425 3638
rect 623 3621 643 3641
rect 841 3619 861 3639
rect 3453 3549 3473 3569
rect 3671 3547 3691 3567
rect 3889 3550 3909 3570
rect 1203 3434 1223 3454
rect 1421 3437 1441 3457
rect 1639 3435 1659 3455
rect 2556 3323 2576 3343
rect 2774 3321 2794 3341
rect 2992 3324 3012 3344
rect 406 3206 426 3226
rect 624 3209 644 3229
rect 842 3207 862 3227
rect 3435 2943 3455 2963
rect 3653 2941 3673 2961
rect 3871 2944 3891 2964
rect 1285 2826 1305 2846
rect 1503 2829 1523 2849
rect 1721 2827 1741 2847
rect 2638 2715 2658 2735
rect 2856 2713 2876 2733
rect 3074 2716 3094 2736
rect 388 2600 408 2620
rect 606 2603 626 2623
rect 824 2601 844 2621
rect 3436 2531 3456 2551
rect 3654 2529 3674 2549
rect 3872 2532 3892 2552
rect 1186 2416 1206 2436
rect 1404 2419 1424 2439
rect 1622 2417 1642 2437
rect 2473 2307 2493 2327
rect 2691 2305 2711 2325
rect 2909 2308 2929 2328
rect 389 2188 409 2208
rect 607 2191 627 2211
rect 825 2189 845 2209
rect 3415 1925 3435 1945
rect 3633 1923 3653 1943
rect 3851 1926 3871 1946
rect 1331 1806 1351 1826
rect 1549 1809 1569 1829
rect 1767 1807 1787 1827
rect 2618 1697 2638 1717
rect 2836 1695 2856 1715
rect 3054 1698 3074 1718
rect 368 1582 388 1602
rect 586 1585 606 1605
rect 804 1583 824 1603
rect 3416 1513 3436 1533
rect 3634 1511 3654 1531
rect 3852 1514 3872 1534
rect 1166 1398 1186 1418
rect 1384 1401 1404 1421
rect 1602 1399 1622 1419
rect 2519 1287 2539 1307
rect 2737 1285 2757 1305
rect 2955 1288 2975 1308
rect 369 1170 389 1190
rect 587 1173 607 1193
rect 805 1171 825 1191
rect 3398 907 3418 927
rect 3616 905 3636 925
rect 3834 908 3854 928
rect 1248 790 1268 810
rect 1466 793 1486 813
rect 1684 791 1704 811
rect 2601 679 2621 699
rect 2819 677 2839 697
rect 3037 680 3057 700
rect 351 564 371 584
rect 569 567 589 587
rect 787 565 807 585
rect 3399 495 3419 515
rect 3617 493 3637 513
rect 3835 496 3855 516
rect 1149 380 1169 400
rect 1367 383 1387 403
rect 1585 381 1605 401
rect 352 152 372 172
rect 570 155 590 175
rect 788 153 808 173
rect 1565 -424 1585 -404
rect 1783 -421 1803 -401
rect 2001 -423 2021 -403
<< ndiffres >>
rect 4181 8118 4238 8137
rect 4181 8100 4199 8118
rect 4217 8115 4238 8118
rect 4217 8100 4332 8115
rect 240 8060 301 8076
rect 145 8056 301 8060
rect 145 8038 263 8056
rect 281 8038 301 8056
rect 145 8017 301 8038
rect 145 8016 245 8017
rect 146 7980 188 8016
rect 4181 8077 4332 8100
rect 4290 8041 4332 8077
rect 4233 8040 4333 8041
rect 4177 8019 4333 8040
rect 146 7957 297 7980
rect 146 7942 261 7957
rect 240 7939 261 7942
rect 279 7939 297 7957
rect 240 7920 297 7939
rect 4177 8001 4197 8019
rect 4215 8001 4333 8019
rect 4177 7997 4333 8001
rect 4177 7981 4238 7997
rect 4174 7900 4231 7919
rect 4174 7882 4192 7900
rect 4210 7897 4231 7900
rect 4210 7882 4325 7897
rect 4174 7859 4325 7882
rect 235 7736 296 7752
rect 4283 7823 4325 7859
rect 4226 7822 4326 7823
rect 4170 7801 4326 7822
rect 4170 7783 4190 7801
rect 4208 7783 4326 7801
rect 4170 7779 4326 7783
rect 140 7732 296 7736
rect 140 7714 258 7732
rect 276 7714 296 7732
rect 140 7693 296 7714
rect 140 7692 240 7693
rect 141 7656 183 7692
rect 4170 7763 4231 7779
rect 4168 7717 4225 7736
rect 141 7633 292 7656
rect 141 7618 256 7633
rect 235 7615 256 7618
rect 274 7615 292 7633
rect 4168 7699 4186 7717
rect 4204 7714 4225 7717
rect 4204 7699 4319 7714
rect 4168 7676 4319 7699
rect 235 7596 292 7615
rect 229 7553 290 7569
rect 4277 7640 4319 7676
rect 4220 7639 4320 7640
rect 4164 7618 4320 7639
rect 4164 7600 4184 7618
rect 4202 7600 4320 7618
rect 4164 7596 4320 7600
rect 134 7549 290 7553
rect 134 7531 252 7549
rect 270 7531 290 7549
rect 134 7510 290 7531
rect 134 7509 234 7510
rect 135 7473 177 7509
rect 4164 7580 4225 7596
rect 135 7450 286 7473
rect 135 7435 250 7450
rect 229 7432 250 7435
rect 268 7432 286 7450
rect 229 7413 286 7432
rect 222 7335 283 7351
rect 127 7331 283 7335
rect 127 7313 245 7331
rect 263 7313 283 7331
rect 4163 7393 4220 7412
rect 4163 7375 4181 7393
rect 4199 7390 4220 7393
rect 4199 7375 4314 7390
rect 127 7292 283 7313
rect 127 7291 227 7292
rect 128 7255 170 7291
rect 128 7232 279 7255
rect 4163 7352 4314 7375
rect 4272 7316 4314 7352
rect 4215 7315 4315 7316
rect 4159 7294 4315 7315
rect 4159 7276 4179 7294
rect 4197 7276 4315 7294
rect 4159 7272 4315 7276
rect 4159 7256 4220 7272
rect 128 7217 243 7232
rect 222 7214 243 7217
rect 261 7214 279 7232
rect 222 7195 279 7214
rect 4164 7100 4221 7119
rect 4164 7082 4182 7100
rect 4200 7097 4221 7100
rect 4200 7082 4315 7097
rect 223 7042 284 7058
rect 128 7038 284 7042
rect 128 7020 246 7038
rect 264 7020 284 7038
rect 128 6999 284 7020
rect 128 6998 228 6999
rect 129 6962 171 6998
rect 129 6939 280 6962
rect 4164 7059 4315 7082
rect 4273 7023 4315 7059
rect 4216 7022 4316 7023
rect 4160 7001 4316 7022
rect 129 6924 244 6939
rect 223 6921 244 6924
rect 262 6921 280 6939
rect 223 6902 280 6921
rect 4160 6983 4180 7001
rect 4198 6983 4316 7001
rect 4160 6979 4316 6983
rect 4160 6963 4221 6979
rect 4157 6882 4214 6901
rect 4157 6864 4175 6882
rect 4193 6879 4214 6882
rect 4193 6864 4308 6879
rect 4157 6841 4308 6864
rect 218 6718 279 6734
rect 4266 6805 4308 6841
rect 4209 6804 4309 6805
rect 4153 6783 4309 6804
rect 4153 6765 4173 6783
rect 4191 6765 4309 6783
rect 4153 6761 4309 6765
rect 123 6714 279 6718
rect 123 6696 241 6714
rect 259 6696 279 6714
rect 123 6675 279 6696
rect 123 6674 223 6675
rect 124 6638 166 6674
rect 4153 6745 4214 6761
rect 4151 6699 4208 6718
rect 124 6615 275 6638
rect 124 6600 239 6615
rect 218 6597 239 6600
rect 257 6597 275 6615
rect 4151 6681 4169 6699
rect 4187 6696 4208 6699
rect 4187 6681 4302 6696
rect 4151 6658 4302 6681
rect 218 6578 275 6597
rect 212 6535 273 6551
rect 4260 6622 4302 6658
rect 4203 6621 4303 6622
rect 4147 6600 4303 6621
rect 4147 6582 4167 6600
rect 4185 6582 4303 6600
rect 4147 6578 4303 6582
rect 117 6531 273 6535
rect 117 6513 235 6531
rect 253 6513 273 6531
rect 117 6492 273 6513
rect 117 6491 217 6492
rect 118 6455 160 6491
rect 4147 6562 4208 6578
rect 118 6432 269 6455
rect 118 6417 233 6432
rect 212 6414 233 6417
rect 251 6414 269 6432
rect 212 6395 269 6414
rect 205 6317 266 6333
rect 110 6313 266 6317
rect 110 6295 228 6313
rect 246 6295 266 6313
rect 4146 6375 4203 6394
rect 4146 6357 4164 6375
rect 4182 6372 4203 6375
rect 4182 6357 4297 6372
rect 110 6274 266 6295
rect 110 6273 210 6274
rect 111 6237 153 6273
rect 111 6214 262 6237
rect 4146 6334 4297 6357
rect 4255 6298 4297 6334
rect 4198 6297 4298 6298
rect 4142 6276 4298 6297
rect 4142 6258 4162 6276
rect 4180 6258 4298 6276
rect 4142 6254 4298 6258
rect 4142 6238 4203 6254
rect 111 6199 226 6214
rect 205 6196 226 6199
rect 244 6196 262 6214
rect 205 6177 262 6196
rect 4144 6082 4201 6101
rect 4144 6064 4162 6082
rect 4180 6079 4201 6082
rect 4180 6064 4295 6079
rect 203 6024 264 6040
rect 108 6020 264 6024
rect 108 6002 226 6020
rect 244 6002 264 6020
rect 108 5981 264 6002
rect 108 5980 208 5981
rect 109 5944 151 5980
rect 109 5921 260 5944
rect 4144 6041 4295 6064
rect 4253 6005 4295 6041
rect 4196 6004 4296 6005
rect 4140 5983 4296 6004
rect 109 5906 224 5921
rect 203 5903 224 5906
rect 242 5903 260 5921
rect 203 5884 260 5903
rect 4140 5965 4160 5983
rect 4178 5965 4296 5983
rect 4140 5961 4296 5965
rect 4140 5945 4201 5961
rect 4137 5864 4194 5883
rect 4137 5846 4155 5864
rect 4173 5861 4194 5864
rect 4173 5846 4288 5861
rect 4137 5823 4288 5846
rect 198 5700 259 5716
rect 4246 5787 4288 5823
rect 4189 5786 4289 5787
rect 4133 5765 4289 5786
rect 4133 5747 4153 5765
rect 4171 5747 4289 5765
rect 4133 5743 4289 5747
rect 103 5696 259 5700
rect 103 5678 221 5696
rect 239 5678 259 5696
rect 103 5657 259 5678
rect 103 5656 203 5657
rect 104 5620 146 5656
rect 4133 5727 4194 5743
rect 4131 5681 4188 5700
rect 104 5597 255 5620
rect 104 5582 219 5597
rect 198 5579 219 5582
rect 237 5579 255 5597
rect 4131 5663 4149 5681
rect 4167 5678 4188 5681
rect 4167 5663 4282 5678
rect 4131 5640 4282 5663
rect 198 5560 255 5579
rect 192 5517 253 5533
rect 4240 5604 4282 5640
rect 4183 5603 4283 5604
rect 4127 5582 4283 5603
rect 4127 5564 4147 5582
rect 4165 5564 4283 5582
rect 4127 5560 4283 5564
rect 97 5513 253 5517
rect 97 5495 215 5513
rect 233 5495 253 5513
rect 97 5474 253 5495
rect 97 5473 197 5474
rect 98 5437 140 5473
rect 4127 5544 4188 5560
rect 98 5414 249 5437
rect 98 5399 213 5414
rect 192 5396 213 5399
rect 231 5396 249 5414
rect 192 5377 249 5396
rect 185 5299 246 5315
rect 90 5295 246 5299
rect 90 5277 208 5295
rect 226 5277 246 5295
rect 4126 5357 4183 5376
rect 4126 5339 4144 5357
rect 4162 5354 4183 5357
rect 4162 5339 4277 5354
rect 90 5256 246 5277
rect 90 5255 190 5256
rect 91 5219 133 5255
rect 91 5196 242 5219
rect 4126 5316 4277 5339
rect 4235 5280 4277 5316
rect 4178 5279 4278 5280
rect 4122 5258 4278 5279
rect 4122 5240 4142 5258
rect 4160 5240 4278 5258
rect 4122 5236 4278 5240
rect 4122 5220 4183 5236
rect 91 5181 206 5196
rect 185 5178 206 5181
rect 224 5178 242 5196
rect 185 5159 242 5178
rect 4127 5064 4184 5083
rect 4127 5046 4145 5064
rect 4163 5061 4184 5064
rect 4163 5046 4278 5061
rect 186 5006 247 5022
rect 91 5002 247 5006
rect 91 4984 209 5002
rect 227 4984 247 5002
rect 91 4963 247 4984
rect 91 4962 191 4963
rect 92 4926 134 4962
rect 92 4903 243 4926
rect 4127 5023 4278 5046
rect 4236 4987 4278 5023
rect 4179 4986 4279 4987
rect 4123 4965 4279 4986
rect 92 4888 207 4903
rect 186 4885 207 4888
rect 225 4885 243 4903
rect 186 4866 243 4885
rect 4123 4947 4143 4965
rect 4161 4947 4279 4965
rect 4123 4943 4279 4947
rect 4123 4927 4184 4943
rect 4120 4846 4177 4865
rect 4120 4828 4138 4846
rect 4156 4843 4177 4846
rect 4156 4828 4271 4843
rect 4120 4805 4271 4828
rect 181 4682 242 4698
rect 4229 4769 4271 4805
rect 4172 4768 4272 4769
rect 4116 4747 4272 4768
rect 4116 4729 4136 4747
rect 4154 4729 4272 4747
rect 4116 4725 4272 4729
rect 86 4678 242 4682
rect 86 4660 204 4678
rect 222 4660 242 4678
rect 86 4639 242 4660
rect 86 4638 186 4639
rect 87 4602 129 4638
rect 4116 4709 4177 4725
rect 4114 4663 4171 4682
rect 87 4579 238 4602
rect 87 4564 202 4579
rect 181 4561 202 4564
rect 220 4561 238 4579
rect 4114 4645 4132 4663
rect 4150 4660 4171 4663
rect 4150 4645 4265 4660
rect 4114 4622 4265 4645
rect 181 4542 238 4561
rect 175 4499 236 4515
rect 4223 4586 4265 4622
rect 4166 4585 4266 4586
rect 4110 4564 4266 4585
rect 4110 4546 4130 4564
rect 4148 4546 4266 4564
rect 4110 4542 4266 4546
rect 80 4495 236 4499
rect 80 4477 198 4495
rect 216 4477 236 4495
rect 80 4456 236 4477
rect 80 4455 180 4456
rect 81 4419 123 4455
rect 4110 4526 4171 4542
rect 81 4396 232 4419
rect 81 4381 196 4396
rect 175 4378 196 4381
rect 214 4378 232 4396
rect 175 4359 232 4378
rect 168 4281 229 4297
rect 73 4277 229 4281
rect 73 4259 191 4277
rect 209 4259 229 4277
rect 4109 4339 4166 4358
rect 4109 4321 4127 4339
rect 4145 4336 4166 4339
rect 4145 4321 4260 4336
rect 73 4238 229 4259
rect 73 4237 173 4238
rect 74 4201 116 4237
rect 74 4178 225 4201
rect 4109 4298 4260 4321
rect 4218 4262 4260 4298
rect 4161 4261 4261 4262
rect 4105 4240 4261 4261
rect 4105 4222 4125 4240
rect 4143 4222 4261 4240
rect 4105 4218 4261 4222
rect 4105 4202 4166 4218
rect 74 4163 189 4178
rect 168 4160 189 4163
rect 207 4160 225 4178
rect 168 4141 225 4160
rect 4108 4046 4165 4065
rect 4108 4028 4126 4046
rect 4144 4043 4165 4046
rect 4144 4028 4259 4043
rect 167 3988 228 4004
rect 72 3984 228 3988
rect 72 3966 190 3984
rect 208 3966 228 3984
rect 72 3945 228 3966
rect 72 3944 172 3945
rect 73 3908 115 3944
rect 73 3885 224 3908
rect 4108 4005 4259 4028
rect 4217 3969 4259 4005
rect 4160 3968 4260 3969
rect 4104 3947 4260 3968
rect 73 3870 188 3885
rect 167 3867 188 3870
rect 206 3867 224 3885
rect 167 3848 224 3867
rect 4104 3929 4124 3947
rect 4142 3929 4260 3947
rect 4104 3925 4260 3929
rect 4104 3909 4165 3925
rect 4101 3828 4158 3847
rect 4101 3810 4119 3828
rect 4137 3825 4158 3828
rect 4137 3810 4252 3825
rect 4101 3787 4252 3810
rect 162 3664 223 3680
rect 4210 3751 4252 3787
rect 4153 3750 4253 3751
rect 4097 3729 4253 3750
rect 4097 3711 4117 3729
rect 4135 3711 4253 3729
rect 4097 3707 4253 3711
rect 67 3660 223 3664
rect 67 3642 185 3660
rect 203 3642 223 3660
rect 67 3621 223 3642
rect 67 3620 167 3621
rect 68 3584 110 3620
rect 4097 3691 4158 3707
rect 4095 3645 4152 3664
rect 68 3561 219 3584
rect 68 3546 183 3561
rect 162 3543 183 3546
rect 201 3543 219 3561
rect 4095 3627 4113 3645
rect 4131 3642 4152 3645
rect 4131 3627 4246 3642
rect 4095 3604 4246 3627
rect 162 3524 219 3543
rect 156 3481 217 3497
rect 4204 3568 4246 3604
rect 4147 3567 4247 3568
rect 4091 3546 4247 3567
rect 4091 3528 4111 3546
rect 4129 3528 4247 3546
rect 4091 3524 4247 3528
rect 61 3477 217 3481
rect 61 3459 179 3477
rect 197 3459 217 3477
rect 61 3438 217 3459
rect 61 3437 161 3438
rect 62 3401 104 3437
rect 4091 3508 4152 3524
rect 62 3378 213 3401
rect 62 3363 177 3378
rect 156 3360 177 3363
rect 195 3360 213 3378
rect 156 3341 213 3360
rect 149 3263 210 3279
rect 54 3259 210 3263
rect 54 3241 172 3259
rect 190 3241 210 3259
rect 4090 3321 4147 3340
rect 4090 3303 4108 3321
rect 4126 3318 4147 3321
rect 4126 3303 4241 3318
rect 54 3220 210 3241
rect 54 3219 154 3220
rect 55 3183 97 3219
rect 55 3160 206 3183
rect 4090 3280 4241 3303
rect 4199 3244 4241 3280
rect 4142 3243 4242 3244
rect 4086 3222 4242 3243
rect 4086 3204 4106 3222
rect 4124 3204 4242 3222
rect 4086 3200 4242 3204
rect 4086 3184 4147 3200
rect 55 3145 170 3160
rect 149 3142 170 3145
rect 188 3142 206 3160
rect 149 3123 206 3142
rect 4091 3028 4148 3047
rect 4091 3010 4109 3028
rect 4127 3025 4148 3028
rect 4127 3010 4242 3025
rect 150 2970 211 2986
rect 55 2966 211 2970
rect 55 2948 173 2966
rect 191 2948 211 2966
rect 55 2927 211 2948
rect 55 2926 155 2927
rect 56 2890 98 2926
rect 56 2867 207 2890
rect 4091 2987 4242 3010
rect 4200 2951 4242 2987
rect 4143 2950 4243 2951
rect 4087 2929 4243 2950
rect 56 2852 171 2867
rect 150 2849 171 2852
rect 189 2849 207 2867
rect 150 2830 207 2849
rect 4087 2911 4107 2929
rect 4125 2911 4243 2929
rect 4087 2907 4243 2911
rect 4087 2891 4148 2907
rect 4084 2810 4141 2829
rect 4084 2792 4102 2810
rect 4120 2807 4141 2810
rect 4120 2792 4235 2807
rect 4084 2769 4235 2792
rect 145 2646 206 2662
rect 4193 2733 4235 2769
rect 4136 2732 4236 2733
rect 4080 2711 4236 2732
rect 4080 2693 4100 2711
rect 4118 2693 4236 2711
rect 4080 2689 4236 2693
rect 50 2642 206 2646
rect 50 2624 168 2642
rect 186 2624 206 2642
rect 50 2603 206 2624
rect 50 2602 150 2603
rect 51 2566 93 2602
rect 4080 2673 4141 2689
rect 4078 2627 4135 2646
rect 51 2543 202 2566
rect 51 2528 166 2543
rect 145 2525 166 2528
rect 184 2525 202 2543
rect 4078 2609 4096 2627
rect 4114 2624 4135 2627
rect 4114 2609 4229 2624
rect 4078 2586 4229 2609
rect 145 2506 202 2525
rect 139 2463 200 2479
rect 4187 2550 4229 2586
rect 4130 2549 4230 2550
rect 4074 2528 4230 2549
rect 4074 2510 4094 2528
rect 4112 2510 4230 2528
rect 4074 2506 4230 2510
rect 44 2459 200 2463
rect 44 2441 162 2459
rect 180 2441 200 2459
rect 44 2420 200 2441
rect 44 2419 144 2420
rect 45 2383 87 2419
rect 4074 2490 4135 2506
rect 45 2360 196 2383
rect 45 2345 160 2360
rect 139 2342 160 2345
rect 178 2342 196 2360
rect 139 2323 196 2342
rect 132 2245 193 2261
rect 37 2241 193 2245
rect 37 2223 155 2241
rect 173 2223 193 2241
rect 4073 2303 4130 2322
rect 4073 2285 4091 2303
rect 4109 2300 4130 2303
rect 4109 2285 4224 2300
rect 37 2202 193 2223
rect 37 2201 137 2202
rect 38 2165 80 2201
rect 38 2142 189 2165
rect 4073 2262 4224 2285
rect 4182 2226 4224 2262
rect 4125 2225 4225 2226
rect 4069 2204 4225 2225
rect 4069 2186 4089 2204
rect 4107 2186 4225 2204
rect 4069 2182 4225 2186
rect 4069 2166 4130 2182
rect 38 2127 153 2142
rect 132 2124 153 2127
rect 171 2124 189 2142
rect 132 2105 189 2124
rect 4071 2010 4128 2029
rect 4071 1992 4089 2010
rect 4107 2007 4128 2010
rect 4107 1992 4222 2007
rect 130 1952 191 1968
rect 35 1948 191 1952
rect 35 1930 153 1948
rect 171 1930 191 1948
rect 35 1909 191 1930
rect 35 1908 135 1909
rect 36 1872 78 1908
rect 36 1849 187 1872
rect 4071 1969 4222 1992
rect 4180 1933 4222 1969
rect 4123 1932 4223 1933
rect 4067 1911 4223 1932
rect 36 1834 151 1849
rect 130 1831 151 1834
rect 169 1831 187 1849
rect 130 1812 187 1831
rect 4067 1893 4087 1911
rect 4105 1893 4223 1911
rect 4067 1889 4223 1893
rect 4067 1873 4128 1889
rect 4064 1792 4121 1811
rect 4064 1774 4082 1792
rect 4100 1789 4121 1792
rect 4100 1774 4215 1789
rect 4064 1751 4215 1774
rect 125 1628 186 1644
rect 4173 1715 4215 1751
rect 4116 1714 4216 1715
rect 4060 1693 4216 1714
rect 4060 1675 4080 1693
rect 4098 1675 4216 1693
rect 4060 1671 4216 1675
rect 30 1624 186 1628
rect 30 1606 148 1624
rect 166 1606 186 1624
rect 30 1585 186 1606
rect 30 1584 130 1585
rect 31 1548 73 1584
rect 4060 1655 4121 1671
rect 4058 1609 4115 1628
rect 31 1525 182 1548
rect 31 1510 146 1525
rect 125 1507 146 1510
rect 164 1507 182 1525
rect 4058 1591 4076 1609
rect 4094 1606 4115 1609
rect 4094 1591 4209 1606
rect 4058 1568 4209 1591
rect 125 1488 182 1507
rect 119 1445 180 1461
rect 4167 1532 4209 1568
rect 4110 1531 4210 1532
rect 4054 1510 4210 1531
rect 4054 1492 4074 1510
rect 4092 1492 4210 1510
rect 4054 1488 4210 1492
rect 24 1441 180 1445
rect 24 1423 142 1441
rect 160 1423 180 1441
rect 24 1402 180 1423
rect 24 1401 124 1402
rect 25 1365 67 1401
rect 4054 1472 4115 1488
rect 25 1342 176 1365
rect 25 1327 140 1342
rect 119 1324 140 1327
rect 158 1324 176 1342
rect 119 1305 176 1324
rect 112 1227 173 1243
rect 17 1223 173 1227
rect 17 1205 135 1223
rect 153 1205 173 1223
rect 4053 1285 4110 1304
rect 4053 1267 4071 1285
rect 4089 1282 4110 1285
rect 4089 1267 4204 1282
rect 17 1184 173 1205
rect 17 1183 117 1184
rect 18 1147 60 1183
rect 18 1124 169 1147
rect 4053 1244 4204 1267
rect 4162 1208 4204 1244
rect 4105 1207 4205 1208
rect 4049 1186 4205 1207
rect 4049 1168 4069 1186
rect 4087 1168 4205 1186
rect 4049 1164 4205 1168
rect 4049 1148 4110 1164
rect 18 1109 133 1124
rect 112 1106 133 1109
rect 151 1106 169 1124
rect 112 1087 169 1106
rect 4054 992 4111 1011
rect 4054 974 4072 992
rect 4090 989 4111 992
rect 4090 974 4205 989
rect 113 934 174 950
rect 18 930 174 934
rect 18 912 136 930
rect 154 912 174 930
rect 18 891 174 912
rect 18 890 118 891
rect 19 854 61 890
rect 19 831 170 854
rect 4054 951 4205 974
rect 4163 915 4205 951
rect 4106 914 4206 915
rect 4050 893 4206 914
rect 19 816 134 831
rect 113 813 134 816
rect 152 813 170 831
rect 113 794 170 813
rect 4050 875 4070 893
rect 4088 875 4206 893
rect 4050 871 4206 875
rect 4050 855 4111 871
rect 4047 774 4104 793
rect 4047 756 4065 774
rect 4083 771 4104 774
rect 4083 756 4198 771
rect 4047 733 4198 756
rect 108 610 169 626
rect 4156 697 4198 733
rect 4099 696 4199 697
rect 4043 675 4199 696
rect 4043 657 4063 675
rect 4081 657 4199 675
rect 4043 653 4199 657
rect 13 606 169 610
rect 13 588 131 606
rect 149 588 169 606
rect 13 567 169 588
rect 13 566 113 567
rect 14 530 56 566
rect 4043 637 4104 653
rect 4041 591 4098 610
rect 14 507 165 530
rect 14 492 129 507
rect 108 489 129 492
rect 147 489 165 507
rect 4041 573 4059 591
rect 4077 588 4098 591
rect 4077 573 4192 588
rect 4041 550 4192 573
rect 108 470 165 489
rect 102 427 163 443
rect 4150 514 4192 550
rect 4093 513 4193 514
rect 4037 492 4193 513
rect 4037 474 4057 492
rect 4075 474 4193 492
rect 4037 470 4193 474
rect 7 423 163 427
rect 7 405 125 423
rect 143 405 163 423
rect 7 384 163 405
rect 7 383 107 384
rect 8 347 50 383
rect 4037 454 4098 470
rect 8 324 159 347
rect 8 309 123 324
rect 102 306 123 309
rect 141 306 159 324
rect 102 287 159 306
rect 95 209 156 225
rect 0 205 156 209
rect 0 187 118 205
rect 136 187 156 205
rect 4036 267 4093 286
rect 4036 249 4054 267
rect 4072 264 4093 267
rect 4072 249 4187 264
rect 4036 226 4187 249
rect 0 166 156 187
rect 0 165 100 166
rect 1 129 43 165
rect 1 106 152 129
rect 4145 190 4187 226
rect 4088 189 4188 190
rect 4032 168 4188 189
rect 4032 150 4052 168
rect 4070 150 4188 168
rect 4032 146 4188 150
rect 4032 130 4093 146
rect 1 91 116 106
rect 95 88 116 91
rect 134 88 152 106
rect 95 69 152 88
<< locali >>
rect 2875 8197 2915 8205
rect 2875 8175 2883 8197
rect 2907 8175 2915 8197
rect 253 8056 300 8172
rect 253 8038 263 8056
rect 281 8038 300 8056
rect 253 8034 300 8038
rect 254 8029 291 8034
rect 242 7967 294 7969
rect 240 7963 673 7967
rect 240 7957 679 7963
rect 240 7939 261 7957
rect 279 7939 679 7957
rect 240 7921 679 7939
rect 242 7732 294 7921
rect 640 7896 679 7921
rect 2480 7946 2517 7952
rect 2480 7927 2488 7946
rect 2509 7927 2517 7946
rect 2480 7919 2517 7927
rect 424 7871 611 7895
rect 640 7876 1035 7896
rect 1055 7876 1058 7896
rect 640 7871 1058 7876
rect 424 7800 461 7871
rect 640 7870 983 7871
rect 640 7867 679 7870
rect 945 7869 982 7870
rect 576 7810 607 7811
rect 424 7780 433 7800
rect 453 7780 461 7800
rect 424 7770 461 7780
rect 520 7800 607 7810
rect 520 7780 529 7800
rect 549 7780 607 7800
rect 520 7771 607 7780
rect 520 7770 557 7771
rect 242 7714 258 7732
rect 276 7714 294 7732
rect 576 7720 607 7771
rect 642 7800 679 7867
rect 794 7810 830 7811
rect 642 7780 651 7800
rect 671 7780 679 7800
rect 642 7770 679 7780
rect 738 7800 886 7810
rect 986 7807 1082 7809
rect 738 7780 747 7800
rect 767 7780 857 7800
rect 877 7780 886 7800
rect 738 7771 886 7780
rect 944 7800 1082 7807
rect 944 7780 953 7800
rect 973 7780 1082 7800
rect 944 7771 1082 7780
rect 738 7770 775 7771
rect 468 7717 509 7718
rect 242 7696 294 7714
rect 360 7710 509 7717
rect 360 7690 419 7710
rect 439 7690 478 7710
rect 498 7690 509 7710
rect 360 7682 509 7690
rect 576 7713 733 7720
rect 576 7693 696 7713
rect 716 7693 733 7713
rect 576 7683 733 7693
rect 576 7682 611 7683
rect 576 7661 607 7682
rect 794 7661 830 7771
rect 849 7770 886 7771
rect 945 7770 982 7771
rect 905 7711 995 7717
rect 905 7691 914 7711
rect 934 7709 995 7711
rect 934 7691 959 7709
rect 905 7689 959 7691
rect 979 7689 995 7709
rect 905 7683 995 7689
rect 419 7660 456 7661
rect 418 7651 456 7660
rect 246 7633 286 7643
rect 246 7615 256 7633
rect 274 7615 286 7633
rect 418 7631 427 7651
rect 447 7631 456 7651
rect 418 7623 456 7631
rect 522 7655 607 7661
rect 637 7660 674 7661
rect 522 7635 530 7655
rect 550 7635 607 7655
rect 522 7627 607 7635
rect 636 7651 674 7660
rect 636 7631 645 7651
rect 665 7631 674 7651
rect 522 7626 558 7627
rect 636 7623 674 7631
rect 740 7655 884 7661
rect 740 7635 748 7655
rect 768 7635 801 7655
rect 821 7635 856 7655
rect 876 7635 884 7655
rect 740 7627 884 7635
rect 740 7626 776 7627
rect 848 7626 884 7627
rect 950 7660 987 7661
rect 950 7659 988 7660
rect 950 7651 1014 7659
rect 950 7631 959 7651
rect 979 7637 1014 7651
rect 1034 7637 1037 7657
rect 979 7632 1037 7637
rect 979 7631 1014 7632
rect 246 7559 286 7615
rect 419 7594 456 7623
rect 420 7592 456 7594
rect 420 7570 611 7592
rect 637 7591 674 7623
rect 950 7619 1014 7631
rect 1054 7593 1081 7771
rect 913 7591 1081 7593
rect 637 7581 1081 7591
rect 1222 7687 1409 7711
rect 1440 7692 1833 7712
rect 1853 7692 1856 7712
rect 1440 7687 1856 7692
rect 1222 7616 1259 7687
rect 1440 7686 1781 7687
rect 1374 7626 1405 7627
rect 1222 7596 1231 7616
rect 1251 7596 1259 7616
rect 1222 7586 1259 7596
rect 1318 7616 1405 7626
rect 1318 7596 1327 7616
rect 1347 7596 1405 7616
rect 1318 7587 1405 7596
rect 1318 7586 1355 7587
rect 243 7554 286 7559
rect 634 7565 1081 7581
rect 634 7559 662 7565
rect 913 7564 1081 7565
rect 243 7551 393 7554
rect 634 7551 661 7559
rect 243 7549 661 7551
rect 243 7531 252 7549
rect 270 7531 661 7549
rect 1374 7536 1405 7587
rect 1440 7616 1477 7686
rect 1743 7685 1780 7686
rect 1592 7626 1628 7627
rect 1440 7596 1449 7616
rect 1469 7596 1477 7616
rect 1440 7586 1477 7596
rect 1536 7616 1684 7626
rect 1784 7623 1880 7625
rect 1536 7596 1545 7616
rect 1565 7596 1655 7616
rect 1675 7596 1684 7616
rect 1536 7587 1684 7596
rect 1742 7616 1880 7623
rect 1742 7596 1751 7616
rect 1771 7596 1880 7616
rect 1742 7587 1880 7596
rect 1536 7586 1573 7587
rect 1266 7533 1307 7534
rect 243 7528 661 7531
rect 243 7522 286 7528
rect 246 7519 286 7522
rect 1158 7526 1307 7533
rect 643 7510 683 7511
rect 354 7493 683 7510
rect 1158 7506 1217 7526
rect 1237 7506 1276 7526
rect 1296 7506 1307 7526
rect 1158 7498 1307 7506
rect 1374 7529 1531 7536
rect 1374 7509 1494 7529
rect 1514 7509 1531 7529
rect 1374 7499 1531 7509
rect 1374 7498 1409 7499
rect 238 7450 281 7461
rect 238 7432 250 7450
rect 268 7432 281 7450
rect 238 7406 281 7432
rect 354 7406 381 7493
rect 643 7484 683 7493
rect 238 7385 381 7406
rect 425 7458 459 7474
rect 643 7464 1036 7484
rect 1056 7464 1059 7484
rect 1374 7477 1405 7498
rect 1592 7477 1628 7587
rect 1647 7586 1684 7587
rect 1743 7586 1780 7587
rect 1703 7527 1793 7533
rect 1703 7507 1712 7527
rect 1732 7525 1793 7527
rect 1732 7507 1757 7525
rect 1703 7505 1757 7507
rect 1777 7505 1793 7525
rect 1703 7499 1793 7505
rect 1217 7476 1254 7477
rect 643 7459 1059 7464
rect 1216 7467 1254 7476
rect 643 7458 984 7459
rect 425 7388 462 7458
rect 577 7398 608 7399
rect 238 7383 375 7385
rect 238 7341 281 7383
rect 425 7368 434 7388
rect 454 7368 462 7388
rect 425 7358 462 7368
rect 521 7388 608 7398
rect 521 7368 530 7388
rect 550 7368 608 7388
rect 521 7359 608 7368
rect 521 7358 558 7359
rect 236 7331 281 7341
rect 236 7313 245 7331
rect 263 7313 281 7331
rect 236 7307 281 7313
rect 577 7308 608 7359
rect 643 7388 680 7458
rect 946 7457 983 7458
rect 1216 7447 1225 7467
rect 1245 7447 1254 7467
rect 1216 7439 1254 7447
rect 1320 7471 1405 7477
rect 1435 7476 1472 7477
rect 1320 7451 1328 7471
rect 1348 7451 1405 7471
rect 1320 7443 1405 7451
rect 1434 7467 1472 7476
rect 1434 7447 1443 7467
rect 1463 7447 1472 7467
rect 1320 7442 1356 7443
rect 1434 7439 1472 7447
rect 1538 7471 1682 7477
rect 1538 7451 1546 7471
rect 1566 7452 1598 7471
rect 1619 7452 1654 7471
rect 1566 7451 1654 7452
rect 1674 7451 1682 7471
rect 1538 7443 1682 7451
rect 1538 7442 1574 7443
rect 1646 7442 1682 7443
rect 1748 7476 1785 7477
rect 1748 7475 1786 7476
rect 1748 7467 1812 7475
rect 1748 7447 1757 7467
rect 1777 7453 1812 7467
rect 1832 7453 1835 7473
rect 1777 7448 1835 7453
rect 1777 7447 1812 7448
rect 1217 7410 1254 7439
rect 1218 7408 1254 7410
rect 795 7398 831 7399
rect 643 7368 652 7388
rect 672 7368 680 7388
rect 643 7358 680 7368
rect 739 7388 887 7398
rect 987 7395 1083 7397
rect 739 7368 748 7388
rect 768 7368 858 7388
rect 878 7368 887 7388
rect 739 7359 887 7368
rect 945 7388 1083 7395
rect 945 7368 954 7388
rect 974 7368 1083 7388
rect 1218 7386 1409 7408
rect 1435 7407 1472 7439
rect 1748 7435 1812 7447
rect 1852 7409 1879 7587
rect 2484 7586 2517 7919
rect 2581 7951 2749 7952
rect 2875 7951 2915 8175
rect 3378 8179 3546 8180
rect 3378 8178 3822 8179
rect 4185 8178 4226 8179
rect 3378 8153 4226 8178
rect 3378 8151 3546 8153
rect 3742 8152 4226 8153
rect 3378 7973 3405 8151
rect 3445 8113 3509 8125
rect 3785 8121 3822 8152
rect 4003 8121 4040 8152
rect 4185 8127 4226 8152
rect 3445 8112 3480 8113
rect 3422 8107 3480 8112
rect 3422 8087 3425 8107
rect 3445 8093 3480 8107
rect 3500 8093 3509 8113
rect 3445 8085 3509 8093
rect 3471 8084 3509 8085
rect 3472 8083 3509 8084
rect 3575 8117 3611 8118
rect 3683 8117 3719 8118
rect 3575 8109 3719 8117
rect 3575 8089 3583 8109
rect 3603 8105 3691 8109
rect 3603 8089 3647 8105
rect 3575 8085 3647 8089
rect 3667 8089 3691 8105
rect 3711 8089 3719 8109
rect 3667 8085 3719 8089
rect 3575 8083 3719 8085
rect 3785 8113 3823 8121
rect 3901 8117 3937 8118
rect 3785 8093 3794 8113
rect 3814 8093 3823 8113
rect 3785 8084 3823 8093
rect 3852 8109 3937 8117
rect 3852 8089 3909 8109
rect 3929 8089 3937 8109
rect 3785 8083 3822 8084
rect 3852 8083 3937 8089
rect 4003 8113 4041 8121
rect 4003 8093 4012 8113
rect 4032 8093 4041 8113
rect 4003 8084 4041 8093
rect 4185 8118 4227 8127
rect 4185 8100 4199 8118
rect 4217 8100 4227 8118
rect 4185 8092 4227 8100
rect 4190 8090 4227 8092
rect 4003 8083 4040 8084
rect 3464 8055 3554 8061
rect 3464 8035 3480 8055
rect 3500 8053 3554 8055
rect 3500 8035 3525 8053
rect 3464 8033 3525 8035
rect 3545 8033 3554 8053
rect 3464 8027 3554 8033
rect 3477 7973 3514 7974
rect 3573 7973 3610 7974
rect 3629 7973 3665 8083
rect 3852 8062 3883 8083
rect 3848 8061 3883 8062
rect 3726 8051 3883 8061
rect 3726 8031 3743 8051
rect 3763 8031 3883 8051
rect 3726 8024 3883 8031
rect 3950 8054 4099 8062
rect 3950 8034 3961 8054
rect 3981 8034 4020 8054
rect 4040 8034 4099 8054
rect 3950 8027 4099 8034
rect 3950 8026 3991 8027
rect 4187 8025 4224 8028
rect 3684 7973 3721 7974
rect 3377 7964 3515 7973
rect 2581 7925 3025 7951
rect 2581 7923 2749 7925
rect 2581 7745 2608 7923
rect 2648 7885 2712 7897
rect 2988 7893 3025 7925
rect 3051 7924 3242 7946
rect 3377 7944 3486 7964
rect 3506 7944 3515 7964
rect 3377 7937 3515 7944
rect 3573 7964 3721 7973
rect 3573 7944 3582 7964
rect 3602 7944 3692 7964
rect 3712 7944 3721 7964
rect 3377 7935 3473 7937
rect 3573 7934 3721 7944
rect 3780 7964 3817 7974
rect 3780 7944 3788 7964
rect 3808 7944 3817 7964
rect 3629 7933 3665 7934
rect 3206 7922 3242 7924
rect 3206 7893 3243 7922
rect 2648 7884 2683 7885
rect 2625 7879 2683 7884
rect 2625 7859 2628 7879
rect 2648 7865 2683 7879
rect 2703 7865 2712 7885
rect 2648 7859 2712 7865
rect 2625 7857 2712 7859
rect 2625 7853 2652 7857
rect 2674 7856 2712 7857
rect 2675 7855 2712 7856
rect 2778 7889 2814 7890
rect 2886 7889 2922 7890
rect 2778 7882 2922 7889
rect 2778 7881 2840 7882
rect 2778 7861 2786 7881
rect 2806 7864 2840 7881
rect 2859 7881 2922 7882
rect 2859 7864 2894 7881
rect 2806 7861 2894 7864
rect 2914 7861 2922 7881
rect 2778 7855 2922 7861
rect 2988 7885 3026 7893
rect 3104 7889 3140 7890
rect 2988 7865 2997 7885
rect 3017 7865 3026 7885
rect 2988 7856 3026 7865
rect 3055 7881 3140 7889
rect 3055 7861 3112 7881
rect 3132 7861 3140 7881
rect 2988 7855 3025 7856
rect 3055 7855 3140 7861
rect 3206 7885 3244 7893
rect 3206 7865 3215 7885
rect 3235 7865 3244 7885
rect 3477 7874 3514 7875
rect 3780 7874 3817 7944
rect 3852 7973 3883 8024
rect 4179 8019 4224 8025
rect 4179 8001 4197 8019
rect 4215 8001 4224 8019
rect 4179 7991 4224 8001
rect 3902 7973 3939 7974
rect 3852 7964 3939 7973
rect 3852 7944 3910 7964
rect 3930 7944 3939 7964
rect 3852 7934 3939 7944
rect 3998 7964 4035 7974
rect 3998 7944 4006 7964
rect 4026 7944 4035 7964
rect 4179 7949 4222 7991
rect 4085 7947 4222 7949
rect 3852 7933 3883 7934
rect 3998 7874 4035 7944
rect 3476 7873 3817 7874
rect 3206 7856 3244 7865
rect 3401 7868 3817 7873
rect 3206 7855 3243 7856
rect 2667 7827 2757 7833
rect 2667 7807 2683 7827
rect 2703 7825 2757 7827
rect 2703 7807 2728 7825
rect 2667 7805 2728 7807
rect 2748 7805 2757 7825
rect 2667 7799 2757 7805
rect 2680 7745 2717 7746
rect 2776 7745 2813 7746
rect 2832 7745 2868 7855
rect 3055 7834 3086 7855
rect 3401 7848 3404 7868
rect 3424 7848 3817 7868
rect 4001 7858 4035 7874
rect 4079 7926 4222 7947
rect 3777 7839 3817 7848
rect 4079 7839 4106 7926
rect 4179 7900 4222 7926
rect 4179 7882 4192 7900
rect 4210 7882 4222 7900
rect 4179 7871 4222 7882
rect 3051 7833 3086 7834
rect 2929 7823 3086 7833
rect 2929 7803 2946 7823
rect 2966 7803 3086 7823
rect 2929 7796 3086 7803
rect 3153 7826 3299 7834
rect 3153 7806 3164 7826
rect 3184 7806 3223 7826
rect 3243 7806 3299 7826
rect 3777 7822 4106 7839
rect 3777 7821 3817 7822
rect 3153 7799 3299 7806
rect 4174 7810 4214 7813
rect 4174 7804 4217 7810
rect 3799 7801 4217 7804
rect 3153 7798 3194 7799
rect 2887 7745 2924 7746
rect 2580 7736 2718 7745
rect 2580 7716 2689 7736
rect 2709 7716 2718 7736
rect 2580 7709 2718 7716
rect 2776 7736 2924 7745
rect 2776 7716 2785 7736
rect 2805 7716 2895 7736
rect 2915 7716 2924 7736
rect 2580 7707 2676 7709
rect 2776 7706 2924 7716
rect 2983 7736 3020 7746
rect 2983 7716 2991 7736
rect 3011 7716 3020 7736
rect 2832 7705 2868 7706
rect 2680 7646 2717 7647
rect 2983 7646 3020 7716
rect 3055 7745 3086 7796
rect 3799 7783 4190 7801
rect 4208 7783 4217 7801
rect 3799 7781 4217 7783
rect 3799 7773 3826 7781
rect 4067 7778 4217 7781
rect 3379 7767 3547 7768
rect 3798 7767 3826 7773
rect 3379 7751 3826 7767
rect 4174 7773 4217 7778
rect 3105 7745 3142 7746
rect 3055 7736 3142 7745
rect 3055 7716 3113 7736
rect 3133 7716 3142 7736
rect 3055 7706 3142 7716
rect 3201 7736 3238 7746
rect 3201 7716 3209 7736
rect 3229 7716 3238 7736
rect 3055 7705 3086 7706
rect 2679 7645 3020 7646
rect 3201 7645 3238 7716
rect 2604 7640 3020 7645
rect 2604 7620 2607 7640
rect 2627 7620 3020 7640
rect 3051 7621 3238 7645
rect 3379 7741 3823 7751
rect 3379 7739 3547 7741
rect 2479 7541 2521 7586
rect 3379 7561 3406 7739
rect 3446 7701 3510 7713
rect 3786 7709 3823 7741
rect 3849 7740 4040 7762
rect 4004 7738 4040 7740
rect 4004 7709 4041 7738
rect 4174 7717 4214 7773
rect 3446 7700 3481 7701
rect 3423 7695 3481 7700
rect 3423 7675 3426 7695
rect 3446 7681 3481 7695
rect 3501 7681 3510 7701
rect 3446 7673 3510 7681
rect 3472 7672 3510 7673
rect 3473 7671 3510 7672
rect 3576 7705 3612 7706
rect 3684 7705 3720 7706
rect 3576 7697 3720 7705
rect 3576 7677 3584 7697
rect 3604 7677 3639 7697
rect 3659 7677 3692 7697
rect 3712 7677 3720 7697
rect 3576 7671 3720 7677
rect 3786 7701 3824 7709
rect 3902 7705 3938 7706
rect 3786 7681 3795 7701
rect 3815 7681 3824 7701
rect 3786 7672 3824 7681
rect 3853 7697 3938 7705
rect 3853 7677 3910 7697
rect 3930 7677 3938 7697
rect 3786 7671 3823 7672
rect 3853 7671 3938 7677
rect 4004 7701 4042 7709
rect 4004 7681 4013 7701
rect 4033 7681 4042 7701
rect 4174 7699 4186 7717
rect 4204 7699 4214 7717
rect 4174 7689 4214 7699
rect 4004 7672 4042 7681
rect 4004 7671 4041 7672
rect 3465 7643 3555 7649
rect 3465 7623 3481 7643
rect 3501 7641 3555 7643
rect 3501 7623 3526 7641
rect 3465 7621 3526 7623
rect 3546 7621 3555 7641
rect 3465 7615 3555 7621
rect 3478 7561 3515 7562
rect 3574 7561 3611 7562
rect 3630 7561 3666 7671
rect 3853 7650 3884 7671
rect 3849 7649 3884 7650
rect 3727 7639 3884 7649
rect 3727 7619 3744 7639
rect 3764 7619 3884 7639
rect 3727 7612 3884 7619
rect 3951 7642 4100 7650
rect 3951 7622 3962 7642
rect 3982 7622 4021 7642
rect 4041 7622 4100 7642
rect 3951 7615 4100 7622
rect 4166 7618 4218 7636
rect 3951 7614 3992 7615
rect 3685 7561 3722 7562
rect 3378 7552 3516 7561
rect 2850 7541 2883 7543
rect 2479 7529 2926 7541
rect 1711 7407 1879 7409
rect 1435 7381 1879 7407
rect 945 7359 1083 7368
rect 739 7358 776 7359
rect 236 7304 273 7307
rect 469 7305 510 7306
rect 361 7298 510 7305
rect 361 7278 420 7298
rect 440 7278 479 7298
rect 499 7278 510 7298
rect 361 7270 510 7278
rect 577 7301 734 7308
rect 577 7281 697 7301
rect 717 7281 734 7301
rect 577 7271 734 7281
rect 577 7270 612 7271
rect 577 7249 608 7270
rect 795 7249 831 7359
rect 850 7358 887 7359
rect 946 7358 983 7359
rect 906 7299 996 7305
rect 906 7279 915 7299
rect 935 7297 996 7299
rect 935 7279 960 7297
rect 906 7277 960 7279
rect 980 7277 996 7297
rect 906 7271 996 7277
rect 420 7248 457 7249
rect 233 7240 270 7242
rect 233 7232 275 7240
rect 233 7214 243 7232
rect 261 7214 275 7232
rect 233 7205 275 7214
rect 419 7239 457 7248
rect 419 7219 428 7239
rect 448 7219 457 7239
rect 419 7211 457 7219
rect 523 7243 608 7249
rect 638 7248 675 7249
rect 523 7223 531 7243
rect 551 7223 608 7243
rect 523 7215 608 7223
rect 637 7239 675 7248
rect 637 7219 646 7239
rect 666 7219 675 7239
rect 523 7214 559 7215
rect 637 7211 675 7219
rect 741 7247 885 7249
rect 741 7243 793 7247
rect 741 7223 749 7243
rect 769 7227 793 7243
rect 813 7243 885 7247
rect 813 7227 857 7243
rect 769 7223 857 7227
rect 877 7223 885 7243
rect 741 7215 885 7223
rect 741 7214 777 7215
rect 849 7214 885 7215
rect 951 7248 988 7249
rect 951 7247 989 7248
rect 951 7239 1015 7247
rect 951 7219 960 7239
rect 980 7225 1015 7239
rect 1035 7225 1038 7245
rect 980 7220 1038 7225
rect 980 7219 1015 7220
rect 234 7180 275 7205
rect 420 7180 457 7211
rect 638 7180 675 7211
rect 951 7207 1015 7219
rect 1055 7181 1082 7359
rect 234 7153 283 7180
rect 419 7154 468 7180
rect 637 7179 718 7180
rect 914 7179 1082 7181
rect 637 7154 1082 7179
rect 638 7153 1082 7154
rect 236 7120 283 7153
rect 639 7120 679 7153
rect 914 7152 1082 7153
rect 1545 7157 1585 7381
rect 1711 7380 1879 7381
rect 2482 7515 2926 7529
rect 2482 7513 2650 7515
rect 2482 7335 2509 7513
rect 2549 7475 2613 7487
rect 2889 7483 2926 7515
rect 2952 7514 3143 7536
rect 3378 7532 3487 7552
rect 3507 7532 3516 7552
rect 3378 7525 3516 7532
rect 3574 7552 3722 7561
rect 3574 7532 3583 7552
rect 3603 7532 3693 7552
rect 3713 7532 3722 7552
rect 3378 7523 3474 7525
rect 3574 7522 3722 7532
rect 3781 7552 3818 7562
rect 3781 7532 3789 7552
rect 3809 7532 3818 7552
rect 3630 7521 3666 7522
rect 3107 7512 3143 7514
rect 3107 7483 3144 7512
rect 2549 7474 2584 7475
rect 2526 7469 2584 7474
rect 2526 7449 2529 7469
rect 2549 7455 2584 7469
rect 2604 7455 2613 7475
rect 2549 7447 2613 7455
rect 2575 7446 2613 7447
rect 2576 7445 2613 7446
rect 2679 7479 2715 7480
rect 2787 7479 2823 7480
rect 2679 7473 2823 7479
rect 2679 7471 2740 7473
rect 2679 7451 2687 7471
rect 2707 7456 2740 7471
rect 2759 7471 2823 7473
rect 2759 7456 2795 7471
rect 2707 7451 2795 7456
rect 2815 7451 2823 7471
rect 2679 7445 2823 7451
rect 2889 7475 2927 7483
rect 3005 7479 3041 7480
rect 2889 7455 2898 7475
rect 2918 7455 2927 7475
rect 2889 7446 2927 7455
rect 2956 7471 3041 7479
rect 2956 7451 3013 7471
rect 3033 7451 3041 7471
rect 2889 7445 2926 7446
rect 2956 7445 3041 7451
rect 3107 7475 3145 7483
rect 3107 7455 3116 7475
rect 3136 7455 3145 7475
rect 3781 7465 3818 7532
rect 3853 7561 3884 7612
rect 4166 7600 4184 7618
rect 4202 7600 4218 7618
rect 3903 7561 3940 7562
rect 3853 7552 3940 7561
rect 3853 7532 3911 7552
rect 3931 7532 3940 7552
rect 3853 7522 3940 7532
rect 3999 7552 4036 7562
rect 3999 7532 4007 7552
rect 4027 7532 4036 7552
rect 3853 7521 3884 7522
rect 3478 7462 3515 7463
rect 3781 7462 3820 7465
rect 3477 7461 3820 7462
rect 3999 7461 4036 7532
rect 3107 7446 3145 7455
rect 3402 7456 3820 7461
rect 3107 7445 3144 7446
rect 2568 7417 2658 7423
rect 2568 7397 2584 7417
rect 2604 7415 2658 7417
rect 2604 7397 2629 7415
rect 2568 7395 2629 7397
rect 2649 7395 2658 7415
rect 2568 7389 2658 7395
rect 2581 7335 2618 7336
rect 2677 7335 2714 7336
rect 2733 7335 2769 7445
rect 2956 7424 2987 7445
rect 3402 7436 3405 7456
rect 3425 7436 3820 7456
rect 3849 7437 4036 7461
rect 2952 7423 2987 7424
rect 2830 7413 2987 7423
rect 2830 7393 2847 7413
rect 2867 7393 2987 7413
rect 2830 7386 2987 7393
rect 3054 7416 3203 7424
rect 3054 7396 3065 7416
rect 3085 7396 3124 7416
rect 3144 7396 3203 7416
rect 3054 7389 3203 7396
rect 3781 7411 3820 7436
rect 4166 7411 4218 7600
rect 3781 7393 4220 7411
rect 3054 7388 3095 7389
rect 2788 7335 2825 7336
rect 2481 7326 2619 7335
rect 2481 7306 2590 7326
rect 2610 7306 2619 7326
rect 2481 7299 2619 7306
rect 2677 7326 2825 7335
rect 2677 7306 2686 7326
rect 2706 7306 2796 7326
rect 2816 7306 2825 7326
rect 2481 7297 2577 7299
rect 2677 7296 2825 7306
rect 2884 7326 2921 7336
rect 2884 7306 2892 7326
rect 2912 7306 2921 7326
rect 2733 7295 2769 7296
rect 2581 7236 2618 7237
rect 2884 7236 2921 7306
rect 2956 7335 2987 7386
rect 3781 7375 4181 7393
rect 4199 7375 4220 7393
rect 3781 7369 4220 7375
rect 3787 7365 4220 7369
rect 4166 7363 4218 7365
rect 3006 7335 3043 7336
rect 2956 7326 3043 7335
rect 2956 7306 3014 7326
rect 3034 7306 3043 7326
rect 2956 7296 3043 7306
rect 3102 7326 3139 7336
rect 3102 7306 3110 7326
rect 3130 7306 3139 7326
rect 2956 7295 2987 7296
rect 2580 7235 2921 7236
rect 3102 7235 3139 7306
rect 4169 7298 4206 7303
rect 4160 7294 4207 7298
rect 4160 7276 4179 7294
rect 4197 7276 4207 7294
rect 2505 7230 2921 7235
rect 2505 7210 2508 7230
rect 2528 7210 2921 7230
rect 2952 7211 3139 7235
rect 3764 7233 3804 7238
rect 4160 7233 4207 7276
rect 3764 7194 4207 7233
rect 1545 7135 1553 7157
rect 1577 7135 1585 7157
rect 1545 7127 1585 7135
rect 2858 7179 2898 7187
rect 2858 7157 2866 7179
rect 2890 7157 2898 7179
rect 236 7081 679 7120
rect 236 7038 283 7081
rect 639 7076 679 7081
rect 1304 7079 1491 7103
rect 1522 7084 1915 7104
rect 1935 7084 1938 7104
rect 1522 7079 1938 7084
rect 236 7020 246 7038
rect 264 7020 283 7038
rect 236 7016 283 7020
rect 237 7011 274 7016
rect 1304 7008 1341 7079
rect 1522 7078 1863 7079
rect 1456 7018 1487 7019
rect 1304 6988 1313 7008
rect 1333 6988 1341 7008
rect 1304 6978 1341 6988
rect 1400 7008 1487 7018
rect 1400 6988 1409 7008
rect 1429 6988 1487 7008
rect 1400 6979 1487 6988
rect 1400 6978 1437 6979
rect 225 6949 277 6951
rect 223 6945 656 6949
rect 223 6939 662 6945
rect 223 6921 244 6939
rect 262 6921 662 6939
rect 1456 6928 1487 6979
rect 1522 7008 1559 7078
rect 1825 7077 1862 7078
rect 1674 7018 1710 7019
rect 1522 6988 1531 7008
rect 1551 6988 1559 7008
rect 1522 6978 1559 6988
rect 1618 7008 1766 7018
rect 1866 7015 1962 7017
rect 1618 6988 1627 7008
rect 1647 6988 1737 7008
rect 1757 6988 1766 7008
rect 1618 6979 1766 6988
rect 1824 7008 1962 7015
rect 1824 6988 1833 7008
rect 1853 6988 1962 7008
rect 1824 6979 1962 6988
rect 1618 6978 1655 6979
rect 1348 6925 1389 6926
rect 223 6903 662 6921
rect 225 6714 277 6903
rect 623 6878 662 6903
rect 1240 6918 1389 6925
rect 1240 6898 1299 6918
rect 1319 6898 1358 6918
rect 1378 6898 1389 6918
rect 1240 6890 1389 6898
rect 1456 6921 1613 6928
rect 1456 6901 1576 6921
rect 1596 6901 1613 6921
rect 1456 6891 1613 6901
rect 1456 6890 1491 6891
rect 407 6853 594 6877
rect 623 6858 1018 6878
rect 1038 6858 1041 6878
rect 1456 6869 1487 6890
rect 1674 6869 1710 6979
rect 1729 6978 1766 6979
rect 1825 6978 1862 6979
rect 1785 6919 1875 6925
rect 1785 6899 1794 6919
rect 1814 6917 1875 6919
rect 1814 6899 1839 6917
rect 1785 6897 1839 6899
rect 1859 6897 1875 6917
rect 1785 6891 1875 6897
rect 1299 6868 1336 6869
rect 623 6853 1041 6858
rect 1298 6859 1336 6868
rect 407 6782 444 6853
rect 623 6852 966 6853
rect 623 6849 662 6852
rect 928 6851 965 6852
rect 559 6792 590 6793
rect 407 6762 416 6782
rect 436 6762 444 6782
rect 407 6752 444 6762
rect 503 6782 590 6792
rect 503 6762 512 6782
rect 532 6762 590 6782
rect 503 6753 590 6762
rect 503 6752 540 6753
rect 225 6696 241 6714
rect 259 6696 277 6714
rect 559 6702 590 6753
rect 625 6782 662 6849
rect 1298 6839 1307 6859
rect 1327 6839 1336 6859
rect 1298 6831 1336 6839
rect 1402 6863 1487 6869
rect 1517 6868 1554 6869
rect 1402 6843 1410 6863
rect 1430 6843 1487 6863
rect 1402 6835 1487 6843
rect 1516 6859 1554 6868
rect 1516 6839 1525 6859
rect 1545 6839 1554 6859
rect 1402 6834 1438 6835
rect 1516 6831 1554 6839
rect 1620 6864 1764 6869
rect 1620 6863 1682 6864
rect 1620 6843 1628 6863
rect 1648 6845 1682 6863
rect 1703 6863 1764 6864
rect 1703 6845 1736 6863
rect 1648 6843 1736 6845
rect 1756 6843 1764 6863
rect 1620 6835 1764 6843
rect 1620 6834 1656 6835
rect 1728 6834 1764 6835
rect 1830 6868 1867 6869
rect 1830 6867 1868 6868
rect 1830 6859 1894 6867
rect 1830 6839 1839 6859
rect 1859 6845 1894 6859
rect 1914 6845 1917 6865
rect 1859 6840 1917 6845
rect 1859 6839 1894 6840
rect 1299 6802 1336 6831
rect 1300 6800 1336 6802
rect 777 6792 813 6793
rect 625 6762 634 6782
rect 654 6762 662 6782
rect 625 6752 662 6762
rect 721 6782 869 6792
rect 969 6789 1065 6791
rect 721 6762 730 6782
rect 750 6762 840 6782
rect 860 6762 869 6782
rect 721 6753 869 6762
rect 927 6782 1065 6789
rect 927 6762 936 6782
rect 956 6762 1065 6782
rect 1300 6778 1491 6800
rect 1517 6799 1554 6831
rect 1830 6827 1894 6839
rect 1934 6801 1961 6979
rect 1793 6799 1961 6801
rect 1517 6785 1961 6799
rect 2564 6933 2732 6934
rect 2858 6933 2898 7157
rect 3361 7161 3529 7162
rect 3764 7161 3804 7194
rect 4160 7161 4207 7194
rect 3361 7160 3805 7161
rect 3361 7135 3806 7160
rect 3361 7133 3529 7135
rect 3725 7134 3806 7135
rect 3975 7134 4024 7160
rect 4160 7134 4209 7161
rect 3361 6955 3388 7133
rect 3428 7095 3492 7107
rect 3768 7103 3805 7134
rect 3986 7103 4023 7134
rect 4168 7109 4209 7134
rect 3428 7094 3463 7095
rect 3405 7089 3463 7094
rect 3405 7069 3408 7089
rect 3428 7075 3463 7089
rect 3483 7075 3492 7095
rect 3428 7067 3492 7075
rect 3454 7066 3492 7067
rect 3455 7065 3492 7066
rect 3558 7099 3594 7100
rect 3666 7099 3702 7100
rect 3558 7091 3702 7099
rect 3558 7071 3566 7091
rect 3586 7087 3674 7091
rect 3586 7071 3630 7087
rect 3558 7067 3630 7071
rect 3650 7071 3674 7087
rect 3694 7071 3702 7091
rect 3650 7067 3702 7071
rect 3558 7065 3702 7067
rect 3768 7095 3806 7103
rect 3884 7099 3920 7100
rect 3768 7075 3777 7095
rect 3797 7075 3806 7095
rect 3768 7066 3806 7075
rect 3835 7091 3920 7099
rect 3835 7071 3892 7091
rect 3912 7071 3920 7091
rect 3768 7065 3805 7066
rect 3835 7065 3920 7071
rect 3986 7095 4024 7103
rect 3986 7075 3995 7095
rect 4015 7075 4024 7095
rect 3986 7066 4024 7075
rect 4168 7100 4210 7109
rect 4168 7082 4182 7100
rect 4200 7082 4210 7100
rect 4168 7074 4210 7082
rect 4173 7072 4210 7074
rect 3986 7065 4023 7066
rect 3447 7037 3537 7043
rect 3447 7017 3463 7037
rect 3483 7035 3537 7037
rect 3483 7017 3508 7035
rect 3447 7015 3508 7017
rect 3528 7015 3537 7035
rect 3447 7009 3537 7015
rect 3460 6955 3497 6956
rect 3556 6955 3593 6956
rect 3612 6955 3648 7065
rect 3835 7044 3866 7065
rect 3831 7043 3866 7044
rect 3709 7033 3866 7043
rect 3709 7013 3726 7033
rect 3746 7013 3866 7033
rect 3709 7006 3866 7013
rect 3933 7036 4082 7044
rect 3933 7016 3944 7036
rect 3964 7016 4003 7036
rect 4023 7016 4082 7036
rect 3933 7009 4082 7016
rect 3933 7008 3974 7009
rect 4170 7007 4207 7010
rect 3667 6955 3704 6956
rect 3360 6946 3498 6955
rect 2564 6907 3008 6933
rect 2564 6905 2732 6907
rect 1517 6773 1964 6785
rect 1560 6771 1593 6773
rect 927 6753 1065 6762
rect 721 6752 758 6753
rect 451 6699 492 6700
rect 225 6678 277 6696
rect 343 6692 492 6699
rect 343 6672 402 6692
rect 422 6672 461 6692
rect 481 6672 492 6692
rect 343 6664 492 6672
rect 559 6695 716 6702
rect 559 6675 679 6695
rect 699 6675 716 6695
rect 559 6665 716 6675
rect 559 6664 594 6665
rect 559 6643 590 6664
rect 777 6643 813 6753
rect 832 6752 869 6753
rect 928 6752 965 6753
rect 888 6693 978 6699
rect 888 6673 897 6693
rect 917 6691 978 6693
rect 917 6673 942 6691
rect 888 6671 942 6673
rect 962 6671 978 6691
rect 888 6665 978 6671
rect 402 6642 439 6643
rect 401 6633 439 6642
rect 229 6615 269 6625
rect 229 6597 239 6615
rect 257 6597 269 6615
rect 401 6613 410 6633
rect 430 6613 439 6633
rect 401 6605 439 6613
rect 505 6637 590 6643
rect 620 6642 657 6643
rect 505 6617 513 6637
rect 533 6617 590 6637
rect 505 6609 590 6617
rect 619 6633 657 6642
rect 619 6613 628 6633
rect 648 6613 657 6633
rect 505 6608 541 6609
rect 619 6605 657 6613
rect 723 6637 867 6643
rect 723 6617 731 6637
rect 751 6617 784 6637
rect 804 6617 839 6637
rect 859 6617 867 6637
rect 723 6609 867 6617
rect 723 6608 759 6609
rect 831 6608 867 6609
rect 933 6642 970 6643
rect 933 6641 971 6642
rect 933 6633 997 6641
rect 933 6613 942 6633
rect 962 6619 997 6633
rect 1017 6619 1020 6639
rect 962 6614 1020 6619
rect 962 6613 997 6614
rect 229 6541 269 6597
rect 402 6576 439 6605
rect 403 6574 439 6576
rect 403 6552 594 6574
rect 620 6573 657 6605
rect 933 6601 997 6613
rect 1037 6575 1064 6753
rect 1922 6728 1964 6773
rect 896 6573 1064 6575
rect 620 6563 1064 6573
rect 1205 6669 1392 6693
rect 1423 6674 1816 6694
rect 1836 6674 1839 6694
rect 1423 6669 1839 6674
rect 1205 6598 1242 6669
rect 1423 6668 1764 6669
rect 1357 6608 1388 6609
rect 1205 6578 1214 6598
rect 1234 6578 1242 6598
rect 1205 6568 1242 6578
rect 1301 6598 1388 6608
rect 1301 6578 1310 6598
rect 1330 6578 1388 6598
rect 1301 6569 1388 6578
rect 1301 6568 1338 6569
rect 226 6536 269 6541
rect 617 6547 1064 6563
rect 617 6541 645 6547
rect 896 6546 1064 6547
rect 226 6533 376 6536
rect 617 6533 644 6541
rect 226 6531 644 6533
rect 226 6513 235 6531
rect 253 6513 644 6531
rect 1357 6518 1388 6569
rect 1423 6598 1460 6668
rect 1726 6667 1763 6668
rect 1575 6608 1611 6609
rect 1423 6578 1432 6598
rect 1452 6578 1460 6598
rect 1423 6568 1460 6578
rect 1519 6598 1667 6608
rect 1767 6605 1863 6607
rect 1519 6578 1528 6598
rect 1548 6578 1638 6598
rect 1658 6578 1667 6598
rect 1519 6569 1667 6578
rect 1725 6598 1863 6605
rect 1725 6578 1734 6598
rect 1754 6578 1863 6598
rect 1725 6569 1863 6578
rect 1519 6568 1556 6569
rect 1249 6515 1290 6516
rect 226 6510 644 6513
rect 226 6504 269 6510
rect 229 6501 269 6504
rect 1144 6508 1290 6515
rect 626 6492 666 6493
rect 337 6475 666 6492
rect 1144 6488 1200 6508
rect 1220 6488 1259 6508
rect 1279 6488 1290 6508
rect 1144 6480 1290 6488
rect 1357 6511 1514 6518
rect 1357 6491 1477 6511
rect 1497 6491 1514 6511
rect 1357 6481 1514 6491
rect 1357 6480 1392 6481
rect 221 6432 264 6443
rect 221 6414 233 6432
rect 251 6414 264 6432
rect 221 6388 264 6414
rect 337 6388 364 6475
rect 626 6466 666 6475
rect 221 6367 364 6388
rect 408 6440 442 6456
rect 626 6446 1019 6466
rect 1039 6446 1042 6466
rect 1357 6459 1388 6480
rect 1575 6459 1611 6569
rect 1630 6568 1667 6569
rect 1726 6568 1763 6569
rect 1686 6509 1776 6515
rect 1686 6489 1695 6509
rect 1715 6507 1776 6509
rect 1715 6489 1740 6507
rect 1686 6487 1740 6489
rect 1760 6487 1776 6507
rect 1686 6481 1776 6487
rect 1200 6458 1237 6459
rect 626 6441 1042 6446
rect 1199 6449 1237 6458
rect 626 6440 967 6441
rect 408 6370 445 6440
rect 560 6380 591 6381
rect 221 6365 358 6367
rect 221 6323 264 6365
rect 408 6350 417 6370
rect 437 6350 445 6370
rect 408 6340 445 6350
rect 504 6370 591 6380
rect 504 6350 513 6370
rect 533 6350 591 6370
rect 504 6341 591 6350
rect 504 6340 541 6341
rect 219 6313 264 6323
rect 219 6295 228 6313
rect 246 6295 264 6313
rect 219 6289 264 6295
rect 560 6290 591 6341
rect 626 6370 663 6440
rect 929 6439 966 6440
rect 1199 6429 1208 6449
rect 1228 6429 1237 6449
rect 1199 6421 1237 6429
rect 1303 6453 1388 6459
rect 1418 6458 1455 6459
rect 1303 6433 1311 6453
rect 1331 6433 1388 6453
rect 1303 6425 1388 6433
rect 1417 6449 1455 6458
rect 1417 6429 1426 6449
rect 1446 6429 1455 6449
rect 1303 6424 1339 6425
rect 1417 6421 1455 6429
rect 1521 6453 1665 6459
rect 1521 6433 1529 6453
rect 1549 6450 1637 6453
rect 1549 6433 1584 6450
rect 1521 6432 1584 6433
rect 1603 6433 1637 6450
rect 1657 6433 1665 6453
rect 1603 6432 1665 6433
rect 1521 6425 1665 6432
rect 1521 6424 1557 6425
rect 1629 6424 1665 6425
rect 1731 6458 1768 6459
rect 1731 6457 1769 6458
rect 1791 6457 1818 6461
rect 1731 6455 1818 6457
rect 1731 6449 1795 6455
rect 1731 6429 1740 6449
rect 1760 6435 1795 6449
rect 1815 6435 1818 6455
rect 1760 6430 1818 6435
rect 1760 6429 1795 6430
rect 1200 6392 1237 6421
rect 1201 6390 1237 6392
rect 778 6380 814 6381
rect 626 6350 635 6370
rect 655 6350 663 6370
rect 626 6340 663 6350
rect 722 6370 870 6380
rect 970 6377 1066 6379
rect 722 6350 731 6370
rect 751 6350 841 6370
rect 861 6350 870 6370
rect 722 6341 870 6350
rect 928 6370 1066 6377
rect 928 6350 937 6370
rect 957 6350 1066 6370
rect 1201 6368 1392 6390
rect 1418 6389 1455 6421
rect 1731 6417 1795 6429
rect 1835 6391 1862 6569
rect 1694 6389 1862 6391
rect 1418 6363 1862 6389
rect 928 6341 1066 6350
rect 722 6340 759 6341
rect 219 6286 256 6289
rect 452 6287 493 6288
rect 344 6280 493 6287
rect 344 6260 403 6280
rect 423 6260 462 6280
rect 482 6260 493 6280
rect 344 6252 493 6260
rect 560 6283 717 6290
rect 560 6263 680 6283
rect 700 6263 717 6283
rect 560 6253 717 6263
rect 560 6252 595 6253
rect 560 6231 591 6252
rect 778 6231 814 6341
rect 833 6340 870 6341
rect 929 6340 966 6341
rect 889 6281 979 6287
rect 889 6261 898 6281
rect 918 6279 979 6281
rect 918 6261 943 6279
rect 889 6259 943 6261
rect 963 6259 979 6279
rect 889 6253 979 6259
rect 403 6230 440 6231
rect 215 6222 253 6224
rect 215 6214 258 6222
rect 215 6196 226 6214
rect 244 6196 258 6214
rect 215 6169 258 6196
rect 402 6221 440 6230
rect 402 6201 411 6221
rect 431 6201 440 6221
rect 402 6193 440 6201
rect 506 6225 591 6231
rect 621 6230 658 6231
rect 506 6205 514 6225
rect 534 6205 591 6225
rect 506 6197 591 6205
rect 620 6221 658 6230
rect 620 6201 629 6221
rect 649 6201 658 6221
rect 506 6196 542 6197
rect 620 6193 658 6201
rect 724 6229 868 6231
rect 724 6225 776 6229
rect 724 6205 732 6225
rect 752 6209 776 6225
rect 796 6225 868 6229
rect 796 6209 840 6225
rect 752 6205 840 6209
rect 860 6205 868 6225
rect 724 6197 868 6205
rect 724 6196 760 6197
rect 832 6196 868 6197
rect 934 6230 971 6231
rect 934 6229 972 6230
rect 934 6221 998 6229
rect 934 6201 943 6221
rect 963 6207 998 6221
rect 1018 6207 1021 6227
rect 963 6202 1021 6207
rect 963 6201 998 6202
rect 216 6162 258 6169
rect 403 6162 440 6193
rect 621 6162 658 6193
rect 934 6189 998 6201
rect 1038 6163 1065 6341
rect 216 6122 261 6162
rect 403 6137 548 6162
rect 621 6161 701 6162
rect 897 6161 1065 6163
rect 621 6145 1065 6161
rect 405 6136 548 6137
rect 620 6135 1065 6145
rect 216 6101 263 6122
rect 620 6101 661 6135
rect 897 6134 1065 6135
rect 1528 6139 1568 6363
rect 1694 6362 1862 6363
rect 1926 6395 1959 6728
rect 2564 6727 2591 6905
rect 2631 6867 2695 6879
rect 2971 6875 3008 6907
rect 3034 6906 3225 6928
rect 3360 6926 3469 6946
rect 3489 6926 3498 6946
rect 3360 6919 3498 6926
rect 3556 6946 3704 6955
rect 3556 6926 3565 6946
rect 3585 6926 3675 6946
rect 3695 6926 3704 6946
rect 3360 6917 3456 6919
rect 3556 6916 3704 6926
rect 3763 6946 3800 6956
rect 3763 6926 3771 6946
rect 3791 6926 3800 6946
rect 3612 6915 3648 6916
rect 3189 6904 3225 6906
rect 3189 6875 3226 6904
rect 2631 6866 2666 6867
rect 2608 6861 2666 6866
rect 2608 6841 2611 6861
rect 2631 6847 2666 6861
rect 2686 6847 2695 6867
rect 2631 6839 2695 6847
rect 2657 6838 2695 6839
rect 2658 6837 2695 6838
rect 2761 6871 2797 6872
rect 2869 6871 2905 6872
rect 2761 6863 2905 6871
rect 2761 6843 2769 6863
rect 2789 6862 2877 6863
rect 2789 6843 2824 6862
rect 2845 6843 2877 6862
rect 2897 6843 2905 6863
rect 2761 6837 2905 6843
rect 2971 6867 3009 6875
rect 3087 6871 3123 6872
rect 2971 6847 2980 6867
rect 3000 6847 3009 6867
rect 2971 6838 3009 6847
rect 3038 6863 3123 6871
rect 3038 6843 3095 6863
rect 3115 6843 3123 6863
rect 2971 6837 3008 6838
rect 3038 6837 3123 6843
rect 3189 6867 3227 6875
rect 3189 6847 3198 6867
rect 3218 6847 3227 6867
rect 3460 6856 3497 6857
rect 3763 6856 3800 6926
rect 3835 6955 3866 7006
rect 4162 7001 4207 7007
rect 4162 6983 4180 7001
rect 4198 6983 4207 7001
rect 4162 6973 4207 6983
rect 3885 6955 3922 6956
rect 3835 6946 3922 6955
rect 3835 6926 3893 6946
rect 3913 6926 3922 6946
rect 3835 6916 3922 6926
rect 3981 6946 4018 6956
rect 3981 6926 3989 6946
rect 4009 6926 4018 6946
rect 4162 6931 4205 6973
rect 4068 6929 4205 6931
rect 3835 6915 3866 6916
rect 3981 6856 4018 6926
rect 3459 6855 3800 6856
rect 3189 6838 3227 6847
rect 3384 6850 3800 6855
rect 3189 6837 3226 6838
rect 2650 6809 2740 6815
rect 2650 6789 2666 6809
rect 2686 6807 2740 6809
rect 2686 6789 2711 6807
rect 2650 6787 2711 6789
rect 2731 6787 2740 6807
rect 2650 6781 2740 6787
rect 2663 6727 2700 6728
rect 2759 6727 2796 6728
rect 2815 6727 2851 6837
rect 3038 6816 3069 6837
rect 3384 6830 3387 6850
rect 3407 6830 3800 6850
rect 3984 6840 4018 6856
rect 4062 6908 4205 6929
rect 3760 6821 3800 6830
rect 4062 6821 4089 6908
rect 4162 6882 4205 6908
rect 4162 6864 4175 6882
rect 4193 6864 4205 6882
rect 4162 6853 4205 6864
rect 3034 6815 3069 6816
rect 2912 6805 3069 6815
rect 2912 6785 2929 6805
rect 2949 6785 3069 6805
rect 2912 6778 3069 6785
rect 3136 6808 3285 6816
rect 3136 6788 3147 6808
rect 3167 6788 3206 6808
rect 3226 6788 3285 6808
rect 3760 6804 4089 6821
rect 3760 6803 3800 6804
rect 3136 6781 3285 6788
rect 4157 6792 4197 6795
rect 4157 6786 4200 6792
rect 3782 6783 4200 6786
rect 3136 6780 3177 6781
rect 2870 6727 2907 6728
rect 2563 6718 2701 6727
rect 2426 6708 2462 6714
rect 2426 6690 2431 6708
rect 2453 6690 2462 6708
rect 2426 6686 2462 6690
rect 2563 6698 2672 6718
rect 2692 6698 2701 6718
rect 2563 6691 2701 6698
rect 2759 6718 2907 6727
rect 2759 6698 2768 6718
rect 2788 6698 2878 6718
rect 2898 6698 2907 6718
rect 2563 6689 2659 6691
rect 2759 6688 2907 6698
rect 2966 6718 3003 6728
rect 2966 6698 2974 6718
rect 2994 6698 3003 6718
rect 2815 6687 2851 6688
rect 2429 6527 2462 6686
rect 2663 6628 2700 6629
rect 2966 6628 3003 6698
rect 3038 6727 3069 6778
rect 3782 6765 4173 6783
rect 4191 6765 4200 6783
rect 3782 6763 4200 6765
rect 3782 6755 3809 6763
rect 4050 6760 4200 6763
rect 3362 6749 3530 6750
rect 3781 6749 3809 6755
rect 3362 6733 3809 6749
rect 4157 6755 4200 6760
rect 3088 6727 3125 6728
rect 3038 6718 3125 6727
rect 3038 6698 3096 6718
rect 3116 6698 3125 6718
rect 3038 6688 3125 6698
rect 3184 6718 3221 6728
rect 3184 6698 3192 6718
rect 3212 6698 3221 6718
rect 3038 6687 3069 6688
rect 2662 6627 3003 6628
rect 3184 6627 3221 6698
rect 2587 6622 3003 6627
rect 2587 6602 2590 6622
rect 2610 6602 3003 6622
rect 3034 6603 3221 6627
rect 3362 6723 3806 6733
rect 3362 6721 3530 6723
rect 3362 6543 3389 6721
rect 3429 6683 3493 6695
rect 3769 6691 3806 6723
rect 3832 6722 4023 6744
rect 3987 6720 4023 6722
rect 3987 6691 4024 6720
rect 4157 6699 4197 6755
rect 3429 6682 3464 6683
rect 3406 6677 3464 6682
rect 3406 6657 3409 6677
rect 3429 6663 3464 6677
rect 3484 6663 3493 6683
rect 3429 6655 3493 6663
rect 3455 6654 3493 6655
rect 3456 6653 3493 6654
rect 3559 6687 3595 6688
rect 3667 6687 3703 6688
rect 3559 6679 3703 6687
rect 3559 6659 3567 6679
rect 3587 6659 3622 6679
rect 3642 6659 3675 6679
rect 3695 6659 3703 6679
rect 3559 6653 3703 6659
rect 3769 6683 3807 6691
rect 3885 6687 3921 6688
rect 3769 6663 3778 6683
rect 3798 6663 3807 6683
rect 3769 6654 3807 6663
rect 3836 6679 3921 6687
rect 3836 6659 3893 6679
rect 3913 6659 3921 6679
rect 3769 6653 3806 6654
rect 3836 6653 3921 6659
rect 3987 6683 4025 6691
rect 3987 6663 3996 6683
rect 4016 6663 4025 6683
rect 4157 6681 4169 6699
rect 4187 6681 4197 6699
rect 4157 6671 4197 6681
rect 3987 6654 4025 6663
rect 3987 6653 4024 6654
rect 3448 6625 3538 6631
rect 3448 6605 3464 6625
rect 3484 6623 3538 6625
rect 3484 6605 3509 6623
rect 3448 6603 3509 6605
rect 3529 6603 3538 6623
rect 3448 6597 3538 6603
rect 3461 6543 3498 6544
rect 3557 6543 3594 6544
rect 3613 6543 3649 6653
rect 3836 6632 3867 6653
rect 3832 6631 3867 6632
rect 3710 6621 3867 6631
rect 3710 6601 3727 6621
rect 3747 6601 3867 6621
rect 3710 6594 3867 6601
rect 3934 6624 4083 6632
rect 3934 6604 3945 6624
rect 3965 6604 4004 6624
rect 4024 6604 4083 6624
rect 3934 6597 4083 6604
rect 4149 6600 4201 6618
rect 3934 6596 3975 6597
rect 3668 6543 3705 6544
rect 3361 6534 3499 6543
rect 2428 6526 2465 6527
rect 2399 6525 2567 6526
rect 2693 6525 2733 6527
rect 2224 6516 2263 6522
rect 2224 6494 2232 6516
rect 2256 6494 2263 6516
rect 1926 6387 1963 6395
rect 1926 6368 1934 6387
rect 1955 6368 1963 6387
rect 1926 6362 1963 6368
rect 1528 6117 1536 6139
rect 1560 6117 1568 6139
rect 1528 6109 1568 6117
rect 216 6071 661 6101
rect 1699 6084 1764 6085
rect 216 6068 639 6071
rect 216 6020 263 6068
rect 216 6002 226 6020
rect 244 6002 263 6020
rect 216 5998 263 6002
rect 1350 6059 1537 6083
rect 1568 6064 1961 6084
rect 1981 6064 1984 6084
rect 1568 6059 1984 6064
rect 217 5993 254 5998
rect 1350 5988 1387 6059
rect 1568 6058 1909 6059
rect 1502 5998 1533 5999
rect 1350 5968 1359 5988
rect 1379 5968 1387 5988
rect 1350 5958 1387 5968
rect 1446 5988 1533 5998
rect 1446 5968 1455 5988
rect 1475 5968 1533 5988
rect 1446 5959 1533 5968
rect 1446 5958 1483 5959
rect 205 5931 257 5933
rect 203 5927 636 5931
rect 203 5921 642 5927
rect 203 5903 224 5921
rect 242 5903 642 5921
rect 1502 5908 1533 5959
rect 1568 5988 1605 6058
rect 1871 6057 1908 6058
rect 1720 5998 1756 5999
rect 1568 5968 1577 5988
rect 1597 5968 1605 5988
rect 1568 5958 1605 5968
rect 1664 5988 1812 5998
rect 1912 5995 2008 5997
rect 1664 5968 1673 5988
rect 1693 5968 1783 5988
rect 1803 5968 1812 5988
rect 1664 5959 1812 5968
rect 1870 5988 2008 5995
rect 1870 5968 1879 5988
rect 1899 5968 2008 5988
rect 1870 5959 2008 5968
rect 1664 5958 1701 5959
rect 1394 5905 1435 5906
rect 203 5885 642 5903
rect 205 5696 257 5885
rect 603 5860 642 5885
rect 1286 5898 1435 5905
rect 1286 5878 1345 5898
rect 1365 5878 1404 5898
rect 1424 5878 1435 5898
rect 1286 5870 1435 5878
rect 1502 5901 1659 5908
rect 1502 5881 1622 5901
rect 1642 5881 1659 5901
rect 1502 5871 1659 5881
rect 1502 5870 1537 5871
rect 387 5835 574 5859
rect 603 5840 998 5860
rect 1018 5840 1021 5860
rect 1502 5849 1533 5870
rect 1720 5849 1756 5959
rect 1775 5958 1812 5959
rect 1871 5958 1908 5959
rect 1831 5899 1921 5905
rect 1831 5879 1840 5899
rect 1860 5897 1921 5899
rect 1860 5879 1885 5897
rect 1831 5877 1885 5879
rect 1905 5877 1921 5897
rect 1831 5871 1921 5877
rect 1345 5848 1382 5849
rect 603 5835 1021 5840
rect 1344 5839 1382 5848
rect 387 5764 424 5835
rect 603 5834 946 5835
rect 603 5831 642 5834
rect 908 5833 945 5834
rect 539 5774 570 5775
rect 387 5744 396 5764
rect 416 5744 424 5764
rect 387 5734 424 5744
rect 483 5764 570 5774
rect 483 5744 492 5764
rect 512 5744 570 5764
rect 483 5735 570 5744
rect 483 5734 520 5735
rect 205 5678 221 5696
rect 239 5678 257 5696
rect 539 5684 570 5735
rect 605 5764 642 5831
rect 1344 5819 1353 5839
rect 1373 5819 1382 5839
rect 1344 5811 1382 5819
rect 1448 5843 1533 5849
rect 1563 5848 1600 5849
rect 1448 5823 1456 5843
rect 1476 5823 1533 5843
rect 1448 5815 1533 5823
rect 1562 5839 1600 5848
rect 1562 5819 1571 5839
rect 1591 5819 1600 5839
rect 1448 5814 1484 5815
rect 1562 5811 1600 5819
rect 1666 5843 1810 5849
rect 1666 5823 1674 5843
rect 1694 5842 1782 5843
rect 1694 5824 1729 5842
rect 1747 5824 1782 5842
rect 1694 5823 1782 5824
rect 1802 5823 1810 5843
rect 1666 5815 1810 5823
rect 1666 5814 1702 5815
rect 1774 5814 1810 5815
rect 1876 5848 1913 5849
rect 1876 5847 1914 5848
rect 1876 5839 1940 5847
rect 1876 5819 1885 5839
rect 1905 5825 1940 5839
rect 1960 5825 1963 5845
rect 1905 5820 1963 5825
rect 1905 5819 1940 5820
rect 1345 5782 1382 5811
rect 1346 5780 1382 5782
rect 757 5774 793 5775
rect 605 5744 614 5764
rect 634 5744 642 5764
rect 605 5734 642 5744
rect 701 5764 849 5774
rect 949 5771 1045 5773
rect 701 5744 710 5764
rect 730 5744 820 5764
rect 840 5744 849 5764
rect 701 5735 849 5744
rect 907 5764 1045 5771
rect 907 5744 916 5764
rect 936 5744 1045 5764
rect 1346 5758 1537 5780
rect 1563 5779 1600 5811
rect 1876 5807 1940 5819
rect 1980 5783 2007 5959
rect 1926 5781 2007 5783
rect 1839 5779 2007 5781
rect 1563 5753 2007 5779
rect 1673 5751 1713 5753
rect 1839 5752 2007 5753
rect 907 5735 1045 5744
rect 1948 5750 2007 5752
rect 701 5734 738 5735
rect 431 5681 472 5682
rect 205 5660 257 5678
rect 323 5674 472 5681
rect 323 5654 382 5674
rect 402 5654 441 5674
rect 461 5654 472 5674
rect 323 5646 472 5654
rect 539 5677 696 5684
rect 539 5657 659 5677
rect 679 5657 696 5677
rect 539 5647 696 5657
rect 539 5646 574 5647
rect 539 5625 570 5646
rect 757 5625 793 5735
rect 812 5734 849 5735
rect 908 5734 945 5735
rect 868 5675 958 5681
rect 868 5655 877 5675
rect 897 5673 958 5675
rect 897 5655 922 5673
rect 868 5653 922 5655
rect 942 5653 958 5673
rect 868 5647 958 5653
rect 382 5624 419 5625
rect 381 5615 419 5624
rect 209 5597 249 5607
rect 209 5579 219 5597
rect 237 5579 249 5597
rect 381 5595 390 5615
rect 410 5595 419 5615
rect 381 5587 419 5595
rect 485 5619 570 5625
rect 600 5624 637 5625
rect 485 5599 493 5619
rect 513 5599 570 5619
rect 485 5591 570 5599
rect 599 5615 637 5624
rect 599 5595 608 5615
rect 628 5595 637 5615
rect 485 5590 521 5591
rect 599 5587 637 5595
rect 703 5619 847 5625
rect 703 5599 711 5619
rect 731 5599 764 5619
rect 784 5599 819 5619
rect 839 5599 847 5619
rect 703 5591 847 5599
rect 703 5590 739 5591
rect 811 5590 847 5591
rect 913 5624 950 5625
rect 913 5623 951 5624
rect 913 5615 977 5623
rect 913 5595 922 5615
rect 942 5601 977 5615
rect 997 5601 1000 5621
rect 942 5596 1000 5601
rect 942 5595 977 5596
rect 209 5523 249 5579
rect 382 5558 419 5587
rect 383 5556 419 5558
rect 383 5534 574 5556
rect 600 5555 637 5587
rect 913 5583 977 5595
rect 1017 5557 1044 5735
rect 1948 5732 1977 5750
rect 876 5555 1044 5557
rect 600 5545 1044 5555
rect 1185 5651 1372 5675
rect 1403 5656 1796 5676
rect 1816 5656 1819 5676
rect 1403 5651 1819 5656
rect 1185 5580 1222 5651
rect 1403 5650 1744 5651
rect 1337 5590 1368 5591
rect 1185 5560 1194 5580
rect 1214 5560 1222 5580
rect 1185 5550 1222 5560
rect 1281 5580 1368 5590
rect 1281 5560 1290 5580
rect 1310 5560 1368 5580
rect 1281 5551 1368 5560
rect 1281 5550 1318 5551
rect 206 5518 249 5523
rect 597 5529 1044 5545
rect 597 5523 625 5529
rect 876 5528 1044 5529
rect 206 5515 356 5518
rect 597 5515 624 5523
rect 206 5513 624 5515
rect 206 5495 215 5513
rect 233 5495 624 5513
rect 1337 5500 1368 5551
rect 1403 5580 1440 5650
rect 1706 5649 1743 5650
rect 1555 5590 1591 5591
rect 1403 5560 1412 5580
rect 1432 5560 1440 5580
rect 1403 5550 1440 5560
rect 1499 5580 1647 5590
rect 1747 5587 1843 5589
rect 1499 5560 1508 5580
rect 1528 5560 1618 5580
rect 1638 5560 1647 5580
rect 1499 5551 1647 5560
rect 1705 5580 1843 5587
rect 1705 5560 1714 5580
rect 1734 5560 1843 5580
rect 1705 5551 1843 5560
rect 1499 5550 1536 5551
rect 1229 5497 1270 5498
rect 206 5492 624 5495
rect 206 5486 249 5492
rect 209 5483 249 5486
rect 1121 5490 1270 5497
rect 606 5474 646 5475
rect 317 5457 646 5474
rect 1121 5470 1180 5490
rect 1200 5470 1239 5490
rect 1259 5470 1270 5490
rect 1121 5462 1270 5470
rect 1337 5493 1494 5500
rect 1337 5473 1457 5493
rect 1477 5473 1494 5493
rect 1337 5463 1494 5473
rect 1337 5462 1372 5463
rect 201 5414 244 5425
rect 201 5396 213 5414
rect 231 5396 244 5414
rect 201 5370 244 5396
rect 317 5370 344 5457
rect 606 5448 646 5457
rect 201 5349 344 5370
rect 388 5422 422 5438
rect 606 5428 999 5448
rect 1019 5428 1022 5448
rect 1337 5441 1368 5462
rect 1555 5441 1591 5551
rect 1610 5550 1647 5551
rect 1706 5550 1743 5551
rect 1666 5491 1756 5497
rect 1666 5471 1675 5491
rect 1695 5489 1756 5491
rect 1695 5471 1720 5489
rect 1666 5469 1720 5471
rect 1740 5469 1756 5489
rect 1666 5463 1756 5469
rect 1180 5440 1217 5441
rect 606 5423 1022 5428
rect 1179 5431 1217 5440
rect 606 5422 947 5423
rect 388 5352 425 5422
rect 540 5362 571 5363
rect 201 5347 338 5349
rect 201 5305 244 5347
rect 388 5332 397 5352
rect 417 5332 425 5352
rect 388 5322 425 5332
rect 484 5352 571 5362
rect 484 5332 493 5352
rect 513 5332 571 5352
rect 484 5323 571 5332
rect 484 5322 521 5323
rect 199 5295 244 5305
rect 199 5277 208 5295
rect 226 5277 244 5295
rect 199 5271 244 5277
rect 540 5272 571 5323
rect 606 5352 643 5422
rect 909 5421 946 5422
rect 1179 5411 1188 5431
rect 1208 5411 1217 5431
rect 1179 5403 1217 5411
rect 1283 5435 1368 5441
rect 1398 5440 1435 5441
rect 1283 5415 1291 5435
rect 1311 5415 1368 5435
rect 1283 5407 1368 5415
rect 1397 5431 1435 5440
rect 1397 5411 1406 5431
rect 1426 5411 1435 5431
rect 1283 5406 1319 5407
rect 1397 5403 1435 5411
rect 1501 5435 1645 5441
rect 1501 5415 1509 5435
rect 1529 5416 1561 5435
rect 1582 5416 1617 5435
rect 1529 5415 1617 5416
rect 1637 5415 1645 5435
rect 1501 5407 1645 5415
rect 1501 5406 1537 5407
rect 1609 5406 1645 5407
rect 1711 5440 1748 5441
rect 1711 5439 1749 5440
rect 1711 5431 1775 5439
rect 1711 5411 1720 5431
rect 1740 5417 1775 5431
rect 1795 5417 1798 5437
rect 1740 5412 1798 5417
rect 1740 5411 1775 5412
rect 1180 5374 1217 5403
rect 1181 5372 1217 5374
rect 758 5362 794 5363
rect 606 5332 615 5352
rect 635 5332 643 5352
rect 606 5322 643 5332
rect 702 5352 850 5362
rect 950 5359 1046 5361
rect 702 5332 711 5352
rect 731 5332 821 5352
rect 841 5332 850 5352
rect 702 5323 850 5332
rect 908 5352 1046 5359
rect 908 5332 917 5352
rect 937 5332 1046 5352
rect 1181 5350 1372 5372
rect 1398 5371 1435 5403
rect 1711 5399 1775 5411
rect 1815 5373 1842 5551
rect 1674 5371 1842 5373
rect 1398 5345 1842 5371
rect 908 5323 1046 5332
rect 702 5322 739 5323
rect 199 5268 236 5271
rect 432 5269 473 5270
rect 324 5262 473 5269
rect 324 5242 383 5262
rect 403 5242 442 5262
rect 462 5242 473 5262
rect 324 5234 473 5242
rect 540 5265 697 5272
rect 540 5245 660 5265
rect 680 5245 697 5265
rect 540 5235 697 5245
rect 540 5234 575 5235
rect 540 5213 571 5234
rect 758 5213 794 5323
rect 813 5322 850 5323
rect 909 5322 946 5323
rect 869 5263 959 5269
rect 869 5243 878 5263
rect 898 5261 959 5263
rect 898 5243 923 5261
rect 869 5241 923 5243
rect 943 5241 959 5261
rect 869 5235 959 5241
rect 383 5212 420 5213
rect 196 5204 233 5206
rect 196 5196 238 5204
rect 196 5178 206 5196
rect 224 5178 238 5196
rect 196 5169 238 5178
rect 382 5203 420 5212
rect 382 5183 391 5203
rect 411 5183 420 5203
rect 382 5175 420 5183
rect 486 5207 571 5213
rect 601 5212 638 5213
rect 486 5187 494 5207
rect 514 5187 571 5207
rect 486 5179 571 5187
rect 600 5203 638 5212
rect 600 5183 609 5203
rect 629 5183 638 5203
rect 486 5178 522 5179
rect 600 5175 638 5183
rect 704 5211 848 5213
rect 704 5207 756 5211
rect 704 5187 712 5207
rect 732 5191 756 5207
rect 776 5207 848 5211
rect 776 5191 820 5207
rect 732 5187 820 5191
rect 840 5187 848 5207
rect 704 5179 848 5187
rect 704 5178 740 5179
rect 812 5178 848 5179
rect 914 5212 951 5213
rect 914 5211 952 5212
rect 914 5203 978 5211
rect 914 5183 923 5203
rect 943 5189 978 5203
rect 998 5189 1001 5209
rect 943 5184 1001 5189
rect 943 5183 978 5184
rect 197 5144 238 5169
rect 383 5144 420 5175
rect 601 5144 638 5175
rect 914 5171 978 5183
rect 1018 5145 1045 5323
rect 197 5117 246 5144
rect 382 5118 431 5144
rect 600 5143 681 5144
rect 877 5143 1045 5145
rect 600 5118 1045 5143
rect 601 5117 1045 5118
rect 199 5084 246 5117
rect 602 5084 642 5117
rect 877 5116 1045 5117
rect 1508 5121 1548 5345
rect 1674 5344 1842 5345
rect 1508 5099 1516 5121
rect 1540 5099 1548 5121
rect 1508 5091 1548 5099
rect 199 5045 642 5084
rect 199 5002 246 5045
rect 602 5040 642 5045
rect 1267 5043 1454 5067
rect 1485 5048 1878 5068
rect 1898 5048 1901 5068
rect 1485 5043 1901 5048
rect 199 4984 209 5002
rect 227 4984 246 5002
rect 199 4980 246 4984
rect 200 4975 237 4980
rect 1267 4972 1304 5043
rect 1485 5042 1826 5043
rect 1419 4982 1450 4983
rect 1267 4952 1276 4972
rect 1296 4952 1304 4972
rect 1267 4942 1304 4952
rect 1363 4972 1450 4982
rect 1363 4952 1372 4972
rect 1392 4952 1450 4972
rect 1363 4943 1450 4952
rect 1363 4942 1400 4943
rect 188 4913 240 4915
rect 186 4909 619 4913
rect 186 4903 625 4909
rect 186 4885 207 4903
rect 225 4885 625 4903
rect 1419 4892 1450 4943
rect 1485 4972 1522 5042
rect 1788 5041 1825 5042
rect 1637 4982 1673 4983
rect 1485 4952 1494 4972
rect 1514 4952 1522 4972
rect 1485 4942 1522 4952
rect 1581 4972 1729 4982
rect 1829 4979 1925 4981
rect 1581 4952 1590 4972
rect 1610 4952 1700 4972
rect 1720 4952 1729 4972
rect 1581 4943 1729 4952
rect 1787 4972 1925 4979
rect 1787 4952 1796 4972
rect 1816 4952 1925 4972
rect 1787 4943 1925 4952
rect 1581 4942 1618 4943
rect 1311 4889 1352 4890
rect 186 4867 625 4885
rect 188 4678 240 4867
rect 586 4842 625 4867
rect 1203 4882 1352 4889
rect 1203 4862 1262 4882
rect 1282 4862 1321 4882
rect 1341 4862 1352 4882
rect 1203 4854 1352 4862
rect 1419 4885 1576 4892
rect 1419 4865 1539 4885
rect 1559 4865 1576 4885
rect 1419 4855 1576 4865
rect 1419 4854 1454 4855
rect 370 4817 557 4841
rect 586 4822 981 4842
rect 1001 4822 1004 4842
rect 1419 4833 1450 4854
rect 1637 4833 1673 4943
rect 1692 4942 1729 4943
rect 1788 4942 1825 4943
rect 1748 4883 1838 4889
rect 1748 4863 1757 4883
rect 1777 4881 1838 4883
rect 1777 4863 1802 4881
rect 1748 4861 1802 4863
rect 1822 4861 1838 4881
rect 1748 4855 1838 4861
rect 1262 4832 1299 4833
rect 586 4817 1004 4822
rect 1261 4823 1299 4832
rect 370 4746 407 4817
rect 586 4816 929 4817
rect 586 4813 625 4816
rect 891 4815 928 4816
rect 522 4756 553 4757
rect 370 4726 379 4746
rect 399 4726 407 4746
rect 370 4716 407 4726
rect 466 4746 553 4756
rect 466 4726 475 4746
rect 495 4726 553 4746
rect 466 4717 553 4726
rect 466 4716 503 4717
rect 188 4660 204 4678
rect 222 4660 240 4678
rect 522 4666 553 4717
rect 588 4746 625 4813
rect 1261 4803 1270 4823
rect 1290 4803 1299 4823
rect 1261 4795 1299 4803
rect 1365 4827 1450 4833
rect 1480 4832 1517 4833
rect 1365 4807 1373 4827
rect 1393 4807 1450 4827
rect 1365 4799 1450 4807
rect 1479 4823 1517 4832
rect 1479 4803 1488 4823
rect 1508 4803 1517 4823
rect 1365 4798 1401 4799
rect 1479 4795 1517 4803
rect 1583 4827 1727 4833
rect 1583 4807 1591 4827
rect 1611 4822 1699 4827
rect 1611 4807 1647 4822
rect 1583 4805 1647 4807
rect 1666 4807 1699 4822
rect 1719 4807 1727 4827
rect 1666 4805 1727 4807
rect 1583 4799 1727 4805
rect 1583 4798 1619 4799
rect 1691 4798 1727 4799
rect 1793 4832 1830 4833
rect 1793 4831 1831 4832
rect 1793 4823 1857 4831
rect 1793 4803 1802 4823
rect 1822 4809 1857 4823
rect 1877 4809 1880 4829
rect 1822 4804 1880 4809
rect 1822 4803 1857 4804
rect 1262 4766 1299 4795
rect 1263 4764 1299 4766
rect 740 4756 776 4757
rect 588 4726 597 4746
rect 617 4726 625 4746
rect 588 4716 625 4726
rect 684 4746 832 4756
rect 932 4753 1028 4755
rect 684 4726 693 4746
rect 713 4726 803 4746
rect 823 4726 832 4746
rect 684 4717 832 4726
rect 890 4746 1028 4753
rect 890 4726 899 4746
rect 919 4726 1028 4746
rect 1263 4742 1454 4764
rect 1480 4763 1517 4795
rect 1793 4791 1857 4803
rect 1897 4765 1924 4943
rect 1756 4763 1924 4765
rect 1480 4749 1924 4763
rect 1948 4786 1976 5732
rect 1948 4756 1993 4786
rect 1480 4737 1927 4749
rect 1523 4735 1556 4737
rect 890 4717 1028 4726
rect 684 4716 721 4717
rect 414 4663 455 4664
rect 188 4642 240 4660
rect 306 4656 455 4663
rect 306 4636 365 4656
rect 385 4636 424 4656
rect 444 4636 455 4656
rect 306 4628 455 4636
rect 522 4659 679 4666
rect 522 4639 642 4659
rect 662 4639 679 4659
rect 522 4629 679 4639
rect 522 4628 557 4629
rect 522 4607 553 4628
rect 740 4607 776 4717
rect 795 4716 832 4717
rect 891 4716 928 4717
rect 851 4657 941 4663
rect 851 4637 860 4657
rect 880 4655 941 4657
rect 880 4637 905 4655
rect 851 4635 905 4637
rect 925 4635 941 4655
rect 851 4629 941 4635
rect 365 4606 402 4607
rect 364 4597 402 4606
rect 192 4579 232 4589
rect 192 4561 202 4579
rect 220 4561 232 4579
rect 364 4577 373 4597
rect 393 4577 402 4597
rect 364 4569 402 4577
rect 468 4601 553 4607
rect 583 4606 620 4607
rect 468 4581 476 4601
rect 496 4581 553 4601
rect 468 4573 553 4581
rect 582 4597 620 4606
rect 582 4577 591 4597
rect 611 4577 620 4597
rect 468 4572 504 4573
rect 582 4569 620 4577
rect 686 4601 830 4607
rect 686 4581 694 4601
rect 714 4581 747 4601
rect 767 4581 802 4601
rect 822 4581 830 4601
rect 686 4573 830 4581
rect 686 4572 722 4573
rect 794 4572 830 4573
rect 896 4606 933 4607
rect 896 4605 934 4606
rect 896 4597 960 4605
rect 896 4577 905 4597
rect 925 4583 960 4597
rect 980 4583 983 4603
rect 925 4578 983 4583
rect 925 4577 960 4578
rect 192 4505 232 4561
rect 365 4540 402 4569
rect 366 4538 402 4540
rect 366 4516 557 4538
rect 583 4537 620 4569
rect 896 4565 960 4577
rect 1000 4539 1027 4717
rect 1885 4692 1927 4737
rect 1948 4738 1959 4756
rect 1981 4738 1993 4756
rect 1948 4732 1993 4738
rect 1949 4731 1993 4732
rect 859 4537 1027 4539
rect 583 4527 1027 4537
rect 1168 4633 1355 4657
rect 1386 4638 1779 4658
rect 1799 4638 1802 4658
rect 1386 4633 1802 4638
rect 1168 4562 1205 4633
rect 1386 4632 1727 4633
rect 1320 4572 1351 4573
rect 1168 4542 1177 4562
rect 1197 4542 1205 4562
rect 1168 4532 1205 4542
rect 1264 4562 1351 4572
rect 1264 4542 1273 4562
rect 1293 4542 1351 4562
rect 1264 4533 1351 4542
rect 1264 4532 1301 4533
rect 189 4500 232 4505
rect 580 4511 1027 4527
rect 580 4505 608 4511
rect 859 4510 1027 4511
rect 189 4497 339 4500
rect 580 4497 607 4505
rect 189 4495 607 4497
rect 189 4477 198 4495
rect 216 4477 607 4495
rect 1320 4482 1351 4533
rect 1386 4562 1423 4632
rect 1689 4631 1726 4632
rect 1538 4572 1574 4573
rect 1386 4542 1395 4562
rect 1415 4542 1423 4562
rect 1386 4532 1423 4542
rect 1482 4562 1630 4572
rect 1730 4569 1826 4571
rect 1482 4542 1491 4562
rect 1511 4542 1601 4562
rect 1621 4542 1630 4562
rect 1482 4533 1630 4542
rect 1688 4562 1826 4569
rect 1688 4542 1697 4562
rect 1717 4542 1826 4562
rect 1688 4533 1826 4542
rect 1482 4532 1519 4533
rect 1212 4479 1253 4480
rect 189 4474 607 4477
rect 189 4468 232 4474
rect 192 4465 232 4468
rect 1107 4472 1253 4479
rect 589 4456 629 4457
rect 300 4439 629 4456
rect 1107 4452 1163 4472
rect 1183 4452 1222 4472
rect 1242 4452 1253 4472
rect 1107 4444 1253 4452
rect 1320 4475 1477 4482
rect 1320 4455 1440 4475
rect 1460 4455 1477 4475
rect 1320 4445 1477 4455
rect 1320 4444 1355 4445
rect 184 4396 227 4407
rect 184 4378 196 4396
rect 214 4378 227 4396
rect 184 4352 227 4378
rect 300 4352 327 4439
rect 589 4430 629 4439
rect 184 4331 327 4352
rect 371 4404 405 4420
rect 589 4410 982 4430
rect 1002 4410 1005 4430
rect 1320 4423 1351 4444
rect 1538 4423 1574 4533
rect 1593 4532 1630 4533
rect 1689 4532 1726 4533
rect 1649 4473 1739 4479
rect 1649 4453 1658 4473
rect 1678 4471 1739 4473
rect 1678 4453 1703 4471
rect 1649 4451 1703 4453
rect 1723 4451 1739 4471
rect 1649 4445 1739 4451
rect 1163 4422 1200 4423
rect 589 4405 1005 4410
rect 1162 4413 1200 4422
rect 589 4404 930 4405
rect 371 4334 408 4404
rect 523 4344 554 4345
rect 184 4329 321 4331
rect 184 4287 227 4329
rect 371 4314 380 4334
rect 400 4314 408 4334
rect 371 4304 408 4314
rect 467 4334 554 4344
rect 467 4314 476 4334
rect 496 4314 554 4334
rect 467 4305 554 4314
rect 467 4304 504 4305
rect 182 4277 227 4287
rect 182 4259 191 4277
rect 209 4259 227 4277
rect 182 4253 227 4259
rect 523 4254 554 4305
rect 589 4334 626 4404
rect 892 4403 929 4404
rect 1162 4393 1171 4413
rect 1191 4393 1200 4413
rect 1162 4385 1200 4393
rect 1266 4417 1351 4423
rect 1381 4422 1418 4423
rect 1266 4397 1274 4417
rect 1294 4397 1351 4417
rect 1266 4389 1351 4397
rect 1380 4413 1418 4422
rect 1380 4393 1389 4413
rect 1409 4393 1418 4413
rect 1266 4388 1302 4389
rect 1380 4385 1418 4393
rect 1484 4417 1628 4423
rect 1484 4397 1492 4417
rect 1512 4414 1600 4417
rect 1512 4397 1547 4414
rect 1484 4396 1547 4397
rect 1566 4397 1600 4414
rect 1620 4397 1628 4417
rect 1566 4396 1628 4397
rect 1484 4389 1628 4396
rect 1484 4388 1520 4389
rect 1592 4388 1628 4389
rect 1694 4422 1731 4423
rect 1694 4421 1732 4422
rect 1754 4421 1781 4425
rect 1694 4419 1781 4421
rect 1694 4413 1758 4419
rect 1694 4393 1703 4413
rect 1723 4399 1758 4413
rect 1778 4399 1781 4419
rect 1723 4394 1781 4399
rect 1723 4393 1758 4394
rect 1163 4356 1200 4385
rect 1164 4354 1200 4356
rect 741 4344 777 4345
rect 589 4314 598 4334
rect 618 4314 626 4334
rect 589 4304 626 4314
rect 685 4334 833 4344
rect 933 4341 1029 4343
rect 685 4314 694 4334
rect 714 4314 804 4334
rect 824 4314 833 4334
rect 685 4305 833 4314
rect 891 4334 1029 4341
rect 891 4314 900 4334
rect 920 4314 1029 4334
rect 1164 4332 1355 4354
rect 1381 4353 1418 4385
rect 1694 4381 1758 4393
rect 1798 4355 1825 4533
rect 1657 4353 1825 4355
rect 1381 4327 1825 4353
rect 891 4305 1029 4314
rect 685 4304 722 4305
rect 182 4250 219 4253
rect 415 4251 456 4252
rect 307 4244 456 4251
rect 307 4224 366 4244
rect 386 4224 425 4244
rect 445 4224 456 4244
rect 307 4216 456 4224
rect 523 4247 680 4254
rect 523 4227 643 4247
rect 663 4227 680 4247
rect 523 4217 680 4227
rect 523 4216 558 4217
rect 523 4195 554 4216
rect 741 4195 777 4305
rect 796 4304 833 4305
rect 892 4304 929 4305
rect 852 4245 942 4251
rect 852 4225 861 4245
rect 881 4243 942 4245
rect 881 4225 906 4243
rect 852 4223 906 4225
rect 926 4223 942 4243
rect 852 4217 942 4223
rect 366 4194 403 4195
rect 179 4186 216 4188
rect 179 4178 221 4186
rect 179 4160 189 4178
rect 207 4160 221 4178
rect 179 4151 221 4160
rect 365 4185 403 4194
rect 365 4165 374 4185
rect 394 4165 403 4185
rect 365 4157 403 4165
rect 469 4189 554 4195
rect 584 4194 621 4195
rect 469 4169 477 4189
rect 497 4169 554 4189
rect 469 4161 554 4169
rect 583 4185 621 4194
rect 583 4165 592 4185
rect 612 4165 621 4185
rect 469 4160 505 4161
rect 583 4157 621 4165
rect 687 4193 831 4195
rect 687 4189 739 4193
rect 687 4169 695 4189
rect 715 4173 739 4189
rect 759 4189 831 4193
rect 759 4173 803 4189
rect 715 4169 803 4173
rect 823 4169 831 4189
rect 687 4161 831 4169
rect 687 4160 723 4161
rect 795 4160 831 4161
rect 897 4194 934 4195
rect 897 4193 935 4194
rect 897 4185 961 4193
rect 897 4165 906 4185
rect 926 4171 961 4185
rect 981 4171 984 4191
rect 926 4166 984 4171
rect 926 4165 961 4166
rect 180 4126 221 4151
rect 366 4126 403 4157
rect 584 4126 621 4157
rect 897 4153 961 4165
rect 1001 4127 1028 4305
rect 180 4092 223 4126
rect 362 4100 429 4126
rect 584 4125 664 4126
rect 860 4125 1028 4127
rect 584 4099 1028 4125
rect 180 4081 227 4092
rect 584 4082 619 4099
rect 860 4098 1028 4099
rect 1491 4103 1531 4327
rect 1657 4326 1825 4327
rect 1889 4359 1922 4692
rect 2224 4679 2263 6494
rect 2399 6500 2843 6525
rect 2399 6319 2426 6500
rect 2568 6499 2843 6500
rect 2466 6459 2530 6471
rect 2806 6467 2843 6499
rect 2869 6498 3060 6520
rect 3361 6514 3470 6534
rect 3490 6514 3499 6534
rect 3361 6507 3499 6514
rect 3557 6534 3705 6543
rect 3557 6514 3566 6534
rect 3586 6514 3676 6534
rect 3696 6514 3705 6534
rect 3361 6505 3457 6507
rect 3557 6504 3705 6514
rect 3764 6534 3801 6544
rect 3764 6514 3772 6534
rect 3792 6514 3801 6534
rect 3613 6503 3649 6504
rect 3024 6496 3060 6498
rect 3024 6467 3061 6496
rect 2466 6458 2501 6459
rect 2443 6453 2501 6458
rect 2443 6433 2446 6453
rect 2466 6439 2501 6453
rect 2521 6439 2530 6459
rect 2466 6431 2530 6439
rect 2492 6430 2530 6431
rect 2493 6429 2530 6430
rect 2596 6463 2632 6464
rect 2704 6463 2740 6464
rect 2596 6455 2740 6463
rect 2596 6435 2604 6455
rect 2624 6453 2712 6455
rect 2624 6435 2657 6453
rect 2596 6431 2657 6435
rect 2680 6435 2712 6453
rect 2732 6435 2740 6455
rect 2680 6431 2740 6435
rect 2596 6429 2740 6431
rect 2806 6459 2844 6467
rect 2922 6463 2958 6464
rect 2806 6439 2815 6459
rect 2835 6439 2844 6459
rect 2806 6430 2844 6439
rect 2873 6455 2958 6463
rect 2873 6435 2930 6455
rect 2950 6435 2958 6455
rect 2806 6429 2843 6430
rect 2873 6429 2958 6435
rect 3024 6459 3062 6467
rect 3024 6439 3033 6459
rect 3053 6439 3062 6459
rect 3764 6447 3801 6514
rect 3836 6543 3867 6594
rect 4149 6582 4167 6600
rect 4185 6582 4201 6600
rect 3886 6543 3923 6544
rect 3836 6534 3923 6543
rect 3836 6514 3894 6534
rect 3914 6514 3923 6534
rect 3836 6504 3923 6514
rect 3982 6534 4019 6544
rect 3982 6514 3990 6534
rect 4010 6514 4019 6534
rect 3836 6503 3867 6504
rect 3461 6444 3498 6445
rect 3764 6444 3803 6447
rect 3460 6443 3803 6444
rect 3982 6443 4019 6514
rect 3024 6430 3062 6439
rect 3385 6438 3803 6443
rect 3024 6429 3061 6430
rect 2485 6401 2575 6407
rect 2485 6381 2501 6401
rect 2521 6399 2575 6401
rect 2521 6381 2546 6399
rect 2485 6379 2546 6381
rect 2566 6379 2575 6399
rect 2485 6373 2575 6379
rect 2498 6319 2535 6320
rect 2594 6319 2631 6320
rect 2650 6319 2686 6429
rect 2873 6408 2904 6429
rect 3385 6418 3388 6438
rect 3408 6418 3803 6438
rect 3832 6419 4019 6443
rect 2869 6407 2904 6408
rect 2747 6397 2904 6407
rect 2747 6377 2764 6397
rect 2784 6377 2904 6397
rect 2747 6370 2904 6377
rect 2971 6400 3120 6408
rect 2971 6380 2982 6400
rect 3002 6380 3041 6400
rect 3061 6380 3120 6400
rect 2971 6373 3120 6380
rect 3764 6393 3803 6418
rect 4149 6393 4201 6582
rect 3764 6375 4203 6393
rect 2971 6372 3012 6373
rect 2705 6319 2742 6320
rect 2398 6310 2536 6319
rect 2398 6290 2507 6310
rect 2527 6290 2536 6310
rect 2398 6283 2536 6290
rect 2594 6310 2742 6319
rect 2594 6290 2603 6310
rect 2623 6290 2713 6310
rect 2733 6290 2742 6310
rect 2398 6281 2494 6283
rect 2594 6280 2742 6290
rect 2801 6310 2838 6320
rect 2801 6290 2809 6310
rect 2829 6290 2838 6310
rect 2650 6279 2686 6280
rect 2498 6220 2535 6221
rect 2801 6220 2838 6290
rect 2873 6319 2904 6370
rect 3764 6357 4164 6375
rect 4182 6357 4203 6375
rect 3764 6351 4203 6357
rect 3770 6347 4203 6351
rect 4149 6345 4201 6347
rect 2923 6319 2960 6320
rect 2873 6310 2960 6319
rect 2873 6290 2931 6310
rect 2951 6290 2960 6310
rect 2873 6280 2960 6290
rect 3019 6310 3056 6320
rect 3019 6290 3027 6310
rect 3047 6290 3056 6310
rect 2873 6279 2904 6280
rect 2497 6219 2838 6220
rect 3019 6219 3056 6290
rect 4152 6280 4189 6285
rect 2422 6214 2838 6219
rect 2422 6194 2425 6214
rect 2445 6194 2838 6214
rect 2869 6195 3056 6219
rect 4143 6276 4190 6280
rect 4143 6258 4162 6276
rect 4180 6258 4190 6276
rect 4143 6210 4190 6258
rect 3767 6207 4190 6210
rect 2642 6193 2707 6194
rect 3745 6177 4190 6207
rect 2838 6161 2878 6169
rect 2838 6139 2846 6161
rect 2870 6139 2878 6161
rect 2443 5910 2480 5916
rect 2443 5891 2451 5910
rect 2472 5891 2480 5910
rect 2443 5883 2480 5891
rect 2447 5550 2480 5883
rect 2544 5915 2712 5916
rect 2838 5915 2878 6139
rect 3341 6143 3509 6144
rect 3745 6143 3786 6177
rect 4143 6156 4190 6177
rect 3341 6133 3786 6143
rect 3858 6141 4001 6142
rect 3341 6117 3785 6133
rect 3341 6115 3509 6117
rect 3705 6116 3785 6117
rect 3858 6116 4003 6141
rect 4145 6116 4190 6156
rect 3341 5937 3368 6115
rect 3408 6077 3472 6089
rect 3748 6085 3785 6116
rect 3966 6085 4003 6116
rect 4148 6109 4190 6116
rect 3408 6076 3443 6077
rect 3385 6071 3443 6076
rect 3385 6051 3388 6071
rect 3408 6057 3443 6071
rect 3463 6057 3472 6077
rect 3408 6049 3472 6057
rect 3434 6048 3472 6049
rect 3435 6047 3472 6048
rect 3538 6081 3574 6082
rect 3646 6081 3682 6082
rect 3538 6073 3682 6081
rect 3538 6053 3546 6073
rect 3566 6069 3654 6073
rect 3566 6053 3610 6069
rect 3538 6049 3610 6053
rect 3630 6053 3654 6069
rect 3674 6053 3682 6073
rect 3630 6049 3682 6053
rect 3538 6047 3682 6049
rect 3748 6077 3786 6085
rect 3864 6081 3900 6082
rect 3748 6057 3757 6077
rect 3777 6057 3786 6077
rect 3748 6048 3786 6057
rect 3815 6073 3900 6081
rect 3815 6053 3872 6073
rect 3892 6053 3900 6073
rect 3748 6047 3785 6048
rect 3815 6047 3900 6053
rect 3966 6077 4004 6085
rect 3966 6057 3975 6077
rect 3995 6057 4004 6077
rect 3966 6048 4004 6057
rect 4148 6082 4191 6109
rect 4148 6064 4162 6082
rect 4180 6064 4191 6082
rect 4148 6056 4191 6064
rect 4153 6054 4191 6056
rect 3966 6047 4003 6048
rect 3427 6019 3517 6025
rect 3427 5999 3443 6019
rect 3463 6017 3517 6019
rect 3463 5999 3488 6017
rect 3427 5997 3488 5999
rect 3508 5997 3517 6017
rect 3427 5991 3517 5997
rect 3440 5937 3477 5938
rect 3536 5937 3573 5938
rect 3592 5937 3628 6047
rect 3815 6026 3846 6047
rect 3811 6025 3846 6026
rect 3689 6015 3846 6025
rect 3689 5995 3706 6015
rect 3726 5995 3846 6015
rect 3689 5988 3846 5995
rect 3913 6018 4062 6026
rect 3913 5998 3924 6018
rect 3944 5998 3983 6018
rect 4003 5998 4062 6018
rect 3913 5991 4062 5998
rect 3913 5990 3954 5991
rect 4150 5989 4187 5992
rect 3647 5937 3684 5938
rect 3340 5928 3478 5937
rect 2544 5889 2988 5915
rect 2544 5887 2712 5889
rect 2544 5709 2571 5887
rect 2611 5849 2675 5861
rect 2951 5857 2988 5889
rect 3014 5888 3205 5910
rect 3340 5908 3449 5928
rect 3469 5908 3478 5928
rect 3340 5901 3478 5908
rect 3536 5928 3684 5937
rect 3536 5908 3545 5928
rect 3565 5908 3655 5928
rect 3675 5908 3684 5928
rect 3340 5899 3436 5901
rect 3536 5898 3684 5908
rect 3743 5928 3780 5938
rect 3743 5908 3751 5928
rect 3771 5908 3780 5928
rect 3592 5897 3628 5898
rect 3169 5886 3205 5888
rect 3169 5857 3206 5886
rect 2611 5848 2646 5849
rect 2588 5843 2646 5848
rect 2588 5823 2591 5843
rect 2611 5829 2646 5843
rect 2666 5829 2675 5849
rect 2611 5823 2675 5829
rect 2588 5821 2675 5823
rect 2588 5817 2615 5821
rect 2637 5820 2675 5821
rect 2638 5819 2675 5820
rect 2741 5853 2777 5854
rect 2849 5853 2885 5854
rect 2741 5846 2885 5853
rect 2741 5845 2803 5846
rect 2741 5825 2749 5845
rect 2769 5828 2803 5845
rect 2822 5845 2885 5846
rect 2822 5828 2857 5845
rect 2769 5825 2857 5828
rect 2877 5825 2885 5845
rect 2741 5819 2885 5825
rect 2951 5849 2989 5857
rect 3067 5853 3103 5854
rect 2951 5829 2960 5849
rect 2980 5829 2989 5849
rect 2951 5820 2989 5829
rect 3018 5845 3103 5853
rect 3018 5825 3075 5845
rect 3095 5825 3103 5845
rect 2951 5819 2988 5820
rect 3018 5819 3103 5825
rect 3169 5849 3207 5857
rect 3169 5829 3178 5849
rect 3198 5829 3207 5849
rect 3440 5838 3477 5839
rect 3743 5838 3780 5908
rect 3815 5937 3846 5988
rect 4142 5983 4187 5989
rect 4142 5965 4160 5983
rect 4178 5965 4187 5983
rect 4142 5955 4187 5965
rect 3865 5937 3902 5938
rect 3815 5928 3902 5937
rect 3815 5908 3873 5928
rect 3893 5908 3902 5928
rect 3815 5898 3902 5908
rect 3961 5928 3998 5938
rect 3961 5908 3969 5928
rect 3989 5908 3998 5928
rect 4142 5913 4185 5955
rect 4048 5911 4185 5913
rect 3815 5897 3846 5898
rect 3961 5838 3998 5908
rect 3439 5837 3780 5838
rect 3169 5820 3207 5829
rect 3364 5832 3780 5837
rect 3169 5819 3206 5820
rect 2630 5791 2720 5797
rect 2630 5771 2646 5791
rect 2666 5789 2720 5791
rect 2666 5771 2691 5789
rect 2630 5769 2691 5771
rect 2711 5769 2720 5789
rect 2630 5763 2720 5769
rect 2643 5709 2680 5710
rect 2739 5709 2776 5710
rect 2795 5709 2831 5819
rect 3018 5798 3049 5819
rect 3364 5812 3367 5832
rect 3387 5812 3780 5832
rect 3964 5822 3998 5838
rect 4042 5890 4185 5911
rect 3740 5803 3780 5812
rect 4042 5803 4069 5890
rect 4142 5864 4185 5890
rect 4142 5846 4155 5864
rect 4173 5846 4185 5864
rect 4142 5835 4185 5846
rect 3014 5797 3049 5798
rect 2892 5787 3049 5797
rect 2892 5767 2909 5787
rect 2929 5767 3049 5787
rect 2892 5760 3049 5767
rect 3116 5790 3262 5798
rect 3116 5770 3127 5790
rect 3147 5770 3186 5790
rect 3206 5770 3262 5790
rect 3740 5786 4069 5803
rect 3740 5785 3780 5786
rect 3116 5763 3262 5770
rect 4137 5774 4177 5777
rect 4137 5768 4180 5774
rect 3762 5765 4180 5768
rect 3116 5762 3157 5763
rect 2850 5709 2887 5710
rect 2543 5700 2681 5709
rect 2543 5680 2652 5700
rect 2672 5680 2681 5700
rect 2543 5673 2681 5680
rect 2739 5700 2887 5709
rect 2739 5680 2748 5700
rect 2768 5680 2858 5700
rect 2878 5680 2887 5700
rect 2543 5671 2639 5673
rect 2739 5670 2887 5680
rect 2946 5700 2983 5710
rect 2946 5680 2954 5700
rect 2974 5680 2983 5700
rect 2795 5669 2831 5670
rect 2643 5610 2680 5611
rect 2946 5610 2983 5680
rect 3018 5709 3049 5760
rect 3762 5747 4153 5765
rect 4171 5747 4180 5765
rect 3762 5745 4180 5747
rect 3762 5737 3789 5745
rect 4030 5742 4180 5745
rect 3342 5731 3510 5732
rect 3761 5731 3789 5737
rect 3342 5715 3789 5731
rect 4137 5737 4180 5742
rect 3068 5709 3105 5710
rect 3018 5700 3105 5709
rect 3018 5680 3076 5700
rect 3096 5680 3105 5700
rect 3018 5670 3105 5680
rect 3164 5700 3201 5710
rect 3164 5680 3172 5700
rect 3192 5680 3201 5700
rect 3018 5669 3049 5670
rect 2642 5609 2983 5610
rect 3164 5609 3201 5680
rect 2567 5604 2983 5609
rect 2567 5584 2570 5604
rect 2590 5584 2983 5604
rect 3014 5585 3201 5609
rect 3342 5705 3786 5715
rect 3342 5703 3510 5705
rect 2442 5505 2484 5550
rect 3342 5525 3369 5703
rect 3409 5665 3473 5677
rect 3749 5673 3786 5705
rect 3812 5704 4003 5726
rect 3967 5702 4003 5704
rect 3967 5673 4004 5702
rect 4137 5681 4177 5737
rect 3409 5664 3444 5665
rect 3386 5659 3444 5664
rect 3386 5639 3389 5659
rect 3409 5645 3444 5659
rect 3464 5645 3473 5665
rect 3409 5637 3473 5645
rect 3435 5636 3473 5637
rect 3436 5635 3473 5636
rect 3539 5669 3575 5670
rect 3647 5669 3683 5670
rect 3539 5661 3683 5669
rect 3539 5641 3547 5661
rect 3567 5641 3602 5661
rect 3622 5641 3655 5661
rect 3675 5641 3683 5661
rect 3539 5635 3683 5641
rect 3749 5665 3787 5673
rect 3865 5669 3901 5670
rect 3749 5645 3758 5665
rect 3778 5645 3787 5665
rect 3749 5636 3787 5645
rect 3816 5661 3901 5669
rect 3816 5641 3873 5661
rect 3893 5641 3901 5661
rect 3749 5635 3786 5636
rect 3816 5635 3901 5641
rect 3967 5665 4005 5673
rect 3967 5645 3976 5665
rect 3996 5645 4005 5665
rect 4137 5663 4149 5681
rect 4167 5663 4177 5681
rect 4137 5653 4177 5663
rect 3967 5636 4005 5645
rect 3967 5635 4004 5636
rect 3428 5607 3518 5613
rect 3428 5587 3444 5607
rect 3464 5605 3518 5607
rect 3464 5587 3489 5605
rect 3428 5585 3489 5587
rect 3509 5585 3518 5605
rect 3428 5579 3518 5585
rect 3441 5525 3478 5526
rect 3537 5525 3574 5526
rect 3593 5525 3629 5635
rect 3816 5614 3847 5635
rect 3812 5613 3847 5614
rect 3690 5603 3847 5613
rect 3690 5583 3707 5603
rect 3727 5583 3847 5603
rect 3690 5576 3847 5583
rect 3914 5606 4063 5614
rect 3914 5586 3925 5606
rect 3945 5586 3984 5606
rect 4004 5586 4063 5606
rect 3914 5579 4063 5586
rect 4129 5582 4181 5600
rect 3914 5578 3955 5579
rect 3648 5525 3685 5526
rect 3341 5516 3479 5525
rect 2813 5505 2846 5507
rect 2442 5493 2889 5505
rect 2445 5479 2889 5493
rect 2445 5477 2613 5479
rect 2445 5299 2472 5477
rect 2512 5439 2576 5451
rect 2852 5447 2889 5479
rect 2915 5478 3106 5500
rect 3341 5496 3450 5516
rect 3470 5496 3479 5516
rect 3341 5489 3479 5496
rect 3537 5516 3685 5525
rect 3537 5496 3546 5516
rect 3566 5496 3656 5516
rect 3676 5496 3685 5516
rect 3341 5487 3437 5489
rect 3537 5486 3685 5496
rect 3744 5516 3781 5526
rect 3744 5496 3752 5516
rect 3772 5496 3781 5516
rect 3593 5485 3629 5486
rect 3070 5476 3106 5478
rect 3070 5447 3107 5476
rect 2512 5438 2547 5439
rect 2489 5433 2547 5438
rect 2489 5413 2492 5433
rect 2512 5419 2547 5433
rect 2567 5419 2576 5439
rect 2512 5411 2576 5419
rect 2538 5410 2576 5411
rect 2539 5409 2576 5410
rect 2642 5443 2678 5444
rect 2750 5443 2786 5444
rect 2642 5435 2786 5443
rect 2642 5415 2650 5435
rect 2670 5433 2758 5435
rect 2670 5415 2703 5433
rect 2642 5414 2703 5415
rect 2724 5415 2758 5433
rect 2778 5415 2786 5435
rect 2724 5414 2786 5415
rect 2642 5409 2786 5414
rect 2852 5439 2890 5447
rect 2968 5443 3004 5444
rect 2852 5419 2861 5439
rect 2881 5419 2890 5439
rect 2852 5410 2890 5419
rect 2919 5435 3004 5443
rect 2919 5415 2976 5435
rect 2996 5415 3004 5435
rect 2852 5409 2889 5410
rect 2919 5409 3004 5415
rect 3070 5439 3108 5447
rect 3070 5419 3079 5439
rect 3099 5419 3108 5439
rect 3744 5429 3781 5496
rect 3816 5525 3847 5576
rect 4129 5564 4147 5582
rect 4165 5564 4181 5582
rect 3866 5525 3903 5526
rect 3816 5516 3903 5525
rect 3816 5496 3874 5516
rect 3894 5496 3903 5516
rect 3816 5486 3903 5496
rect 3962 5516 3999 5526
rect 3962 5496 3970 5516
rect 3990 5496 3999 5516
rect 3816 5485 3847 5486
rect 3441 5426 3478 5427
rect 3744 5426 3783 5429
rect 3440 5425 3783 5426
rect 3962 5425 3999 5496
rect 3070 5410 3108 5419
rect 3365 5420 3783 5425
rect 3070 5409 3107 5410
rect 2531 5381 2621 5387
rect 2531 5361 2547 5381
rect 2567 5379 2621 5381
rect 2567 5361 2592 5379
rect 2531 5359 2592 5361
rect 2612 5359 2621 5379
rect 2531 5353 2621 5359
rect 2544 5299 2581 5300
rect 2640 5299 2677 5300
rect 2696 5299 2732 5409
rect 2919 5388 2950 5409
rect 3365 5400 3368 5420
rect 3388 5400 3783 5420
rect 3812 5401 3999 5425
rect 2915 5387 2950 5388
rect 2793 5377 2950 5387
rect 2793 5357 2810 5377
rect 2830 5357 2950 5377
rect 2793 5350 2950 5357
rect 3017 5380 3166 5388
rect 3017 5360 3028 5380
rect 3048 5360 3087 5380
rect 3107 5360 3166 5380
rect 3017 5353 3166 5360
rect 3744 5375 3783 5400
rect 4129 5375 4181 5564
rect 3744 5357 4183 5375
rect 3017 5352 3058 5353
rect 2751 5299 2788 5300
rect 2444 5290 2582 5299
rect 2444 5270 2553 5290
rect 2573 5270 2582 5290
rect 2444 5263 2582 5270
rect 2640 5290 2788 5299
rect 2640 5270 2649 5290
rect 2669 5270 2759 5290
rect 2779 5270 2788 5290
rect 2444 5261 2540 5263
rect 2640 5260 2788 5270
rect 2847 5290 2884 5300
rect 2847 5270 2855 5290
rect 2875 5270 2884 5290
rect 2696 5259 2732 5260
rect 2544 5200 2581 5201
rect 2847 5200 2884 5270
rect 2919 5299 2950 5350
rect 3744 5339 4144 5357
rect 4162 5339 4183 5357
rect 3744 5333 4183 5339
rect 3750 5329 4183 5333
rect 4129 5327 4181 5329
rect 2969 5299 3006 5300
rect 2919 5290 3006 5299
rect 2919 5270 2977 5290
rect 2997 5270 3006 5290
rect 2919 5260 3006 5270
rect 3065 5290 3102 5300
rect 3065 5270 3073 5290
rect 3093 5270 3102 5290
rect 2919 5259 2950 5260
rect 2543 5199 2884 5200
rect 3065 5199 3102 5270
rect 4132 5262 4169 5267
rect 4123 5258 4170 5262
rect 4123 5240 4142 5258
rect 4160 5240 4170 5258
rect 2468 5194 2884 5199
rect 2468 5174 2471 5194
rect 2491 5174 2884 5194
rect 2915 5175 3102 5199
rect 3727 5197 3767 5202
rect 4123 5197 4170 5240
rect 3727 5158 4170 5197
rect 2821 5143 2861 5151
rect 2821 5121 2829 5143
rect 2853 5121 2861 5143
rect 2527 4897 2695 4898
rect 2821 4897 2861 5121
rect 3324 5125 3492 5126
rect 3727 5125 3767 5158
rect 4123 5125 4170 5158
rect 3324 5124 3768 5125
rect 3324 5099 3769 5124
rect 3324 5097 3492 5099
rect 3688 5098 3769 5099
rect 3938 5098 3987 5124
rect 4123 5098 4172 5125
rect 3324 4919 3351 5097
rect 3391 5059 3455 5071
rect 3731 5067 3768 5098
rect 3949 5067 3986 5098
rect 4131 5073 4172 5098
rect 3391 5058 3426 5059
rect 3368 5053 3426 5058
rect 3368 5033 3371 5053
rect 3391 5039 3426 5053
rect 3446 5039 3455 5059
rect 3391 5031 3455 5039
rect 3417 5030 3455 5031
rect 3418 5029 3455 5030
rect 3521 5063 3557 5064
rect 3629 5063 3665 5064
rect 3521 5055 3665 5063
rect 3521 5035 3529 5055
rect 3549 5051 3637 5055
rect 3549 5035 3593 5051
rect 3521 5031 3593 5035
rect 3613 5035 3637 5051
rect 3657 5035 3665 5055
rect 3613 5031 3665 5035
rect 3521 5029 3665 5031
rect 3731 5059 3769 5067
rect 3847 5063 3883 5064
rect 3731 5039 3740 5059
rect 3760 5039 3769 5059
rect 3731 5030 3769 5039
rect 3798 5055 3883 5063
rect 3798 5035 3855 5055
rect 3875 5035 3883 5055
rect 3731 5029 3768 5030
rect 3798 5029 3883 5035
rect 3949 5059 3987 5067
rect 3949 5039 3958 5059
rect 3978 5039 3987 5059
rect 3949 5030 3987 5039
rect 4131 5064 4173 5073
rect 4131 5046 4145 5064
rect 4163 5046 4173 5064
rect 4131 5038 4173 5046
rect 4136 5036 4173 5038
rect 3949 5029 3986 5030
rect 3410 5001 3500 5007
rect 3410 4981 3426 5001
rect 3446 4999 3500 5001
rect 3446 4981 3471 4999
rect 3410 4979 3471 4981
rect 3491 4979 3500 4999
rect 3410 4973 3500 4979
rect 3423 4919 3460 4920
rect 3519 4919 3556 4920
rect 3575 4919 3611 5029
rect 3798 5008 3829 5029
rect 3794 5007 3829 5008
rect 3672 4997 3829 5007
rect 3672 4977 3689 4997
rect 3709 4977 3829 4997
rect 3672 4970 3829 4977
rect 3896 5000 4045 5008
rect 3896 4980 3907 5000
rect 3927 4980 3966 5000
rect 3986 4980 4045 5000
rect 3896 4973 4045 4980
rect 3896 4972 3937 4973
rect 4133 4971 4170 4974
rect 3630 4919 3667 4920
rect 3323 4910 3461 4919
rect 2527 4871 2971 4897
rect 2527 4869 2695 4871
rect 2527 4691 2554 4869
rect 2594 4831 2658 4843
rect 2934 4839 2971 4871
rect 2997 4870 3188 4892
rect 3323 4890 3432 4910
rect 3452 4890 3461 4910
rect 3323 4883 3461 4890
rect 3519 4910 3667 4919
rect 3519 4890 3528 4910
rect 3548 4890 3638 4910
rect 3658 4890 3667 4910
rect 3323 4881 3419 4883
rect 3519 4880 3667 4890
rect 3726 4910 3763 4920
rect 3726 4890 3734 4910
rect 3754 4890 3763 4910
rect 3575 4879 3611 4880
rect 3152 4868 3188 4870
rect 3152 4839 3189 4868
rect 2594 4830 2629 4831
rect 2571 4825 2629 4830
rect 2571 4805 2574 4825
rect 2594 4811 2629 4825
rect 2649 4811 2658 4831
rect 2594 4803 2658 4811
rect 2620 4802 2658 4803
rect 2621 4801 2658 4802
rect 2724 4835 2760 4836
rect 2832 4835 2868 4836
rect 2724 4827 2868 4835
rect 2724 4807 2732 4827
rect 2752 4826 2840 4827
rect 2752 4807 2787 4826
rect 2808 4807 2840 4826
rect 2860 4807 2868 4827
rect 2724 4801 2868 4807
rect 2934 4831 2972 4839
rect 3050 4835 3086 4836
rect 2934 4811 2943 4831
rect 2963 4811 2972 4831
rect 2934 4802 2972 4811
rect 3001 4827 3086 4835
rect 3001 4807 3058 4827
rect 3078 4807 3086 4827
rect 2934 4801 2971 4802
rect 3001 4801 3086 4807
rect 3152 4831 3190 4839
rect 3152 4811 3161 4831
rect 3181 4811 3190 4831
rect 3423 4820 3460 4821
rect 3726 4820 3763 4890
rect 3798 4919 3829 4970
rect 4125 4965 4170 4971
rect 4125 4947 4143 4965
rect 4161 4947 4170 4965
rect 4125 4937 4170 4947
rect 3848 4919 3885 4920
rect 3798 4910 3885 4919
rect 3798 4890 3856 4910
rect 3876 4890 3885 4910
rect 3798 4880 3885 4890
rect 3944 4910 3981 4920
rect 3944 4890 3952 4910
rect 3972 4890 3981 4910
rect 4125 4895 4168 4937
rect 4031 4893 4168 4895
rect 3798 4879 3829 4880
rect 3944 4820 3981 4890
rect 3422 4819 3763 4820
rect 3152 4802 3190 4811
rect 3347 4814 3763 4819
rect 3152 4801 3189 4802
rect 2613 4773 2703 4779
rect 2613 4753 2629 4773
rect 2649 4771 2703 4773
rect 2649 4753 2674 4771
rect 2613 4751 2674 4753
rect 2694 4751 2703 4771
rect 2613 4745 2703 4751
rect 2626 4691 2663 4692
rect 2722 4691 2759 4692
rect 2778 4691 2814 4801
rect 3001 4780 3032 4801
rect 3347 4794 3350 4814
rect 3370 4794 3763 4814
rect 3947 4804 3981 4820
rect 4025 4872 4168 4893
rect 3723 4785 3763 4794
rect 4025 4785 4052 4872
rect 4125 4846 4168 4872
rect 4125 4828 4138 4846
rect 4156 4828 4168 4846
rect 4125 4817 4168 4828
rect 2997 4779 3032 4780
rect 2875 4769 3032 4779
rect 2875 4749 2892 4769
rect 2912 4749 3032 4769
rect 2875 4742 3032 4749
rect 3099 4772 3248 4780
rect 3099 4752 3110 4772
rect 3130 4752 3169 4772
rect 3189 4752 3248 4772
rect 3723 4768 4052 4785
rect 3723 4767 3763 4768
rect 3099 4745 3248 4752
rect 4120 4756 4160 4759
rect 4120 4750 4163 4756
rect 3745 4747 4163 4750
rect 3099 4744 3140 4745
rect 2833 4691 2870 4692
rect 2526 4682 2664 4691
rect 2224 4507 2264 4679
rect 2526 4662 2635 4682
rect 2655 4662 2664 4682
rect 2526 4655 2664 4662
rect 2722 4682 2870 4691
rect 2722 4662 2731 4682
rect 2751 4662 2841 4682
rect 2861 4662 2870 4682
rect 2526 4653 2622 4655
rect 2722 4652 2870 4662
rect 2929 4682 2966 4692
rect 2929 4662 2937 4682
rect 2957 4662 2966 4682
rect 2778 4651 2814 4652
rect 2626 4592 2663 4593
rect 2929 4592 2966 4662
rect 3001 4691 3032 4742
rect 3745 4729 4136 4747
rect 4154 4729 4163 4747
rect 3745 4727 4163 4729
rect 3745 4719 3772 4727
rect 4013 4724 4163 4727
rect 3325 4713 3493 4714
rect 3744 4713 3772 4719
rect 3325 4697 3772 4713
rect 4120 4719 4163 4724
rect 3051 4691 3088 4692
rect 3001 4682 3088 4691
rect 3001 4662 3059 4682
rect 3079 4662 3088 4682
rect 3001 4652 3088 4662
rect 3147 4682 3184 4692
rect 3147 4662 3155 4682
rect 3175 4662 3184 4682
rect 3001 4651 3032 4652
rect 2625 4591 2966 4592
rect 3147 4591 3184 4662
rect 2550 4586 2966 4591
rect 2550 4566 2553 4586
rect 2573 4566 2966 4586
rect 2997 4567 3184 4591
rect 3325 4687 3769 4697
rect 3325 4685 3493 4687
rect 3325 4507 3352 4685
rect 3392 4647 3456 4659
rect 3732 4655 3769 4687
rect 3795 4686 3986 4708
rect 3950 4684 3986 4686
rect 3950 4655 3987 4684
rect 4120 4663 4160 4719
rect 3392 4646 3427 4647
rect 3369 4641 3427 4646
rect 3369 4621 3372 4641
rect 3392 4627 3427 4641
rect 3447 4627 3456 4647
rect 3392 4619 3456 4627
rect 3418 4618 3456 4619
rect 3419 4617 3456 4618
rect 3522 4651 3558 4652
rect 3630 4651 3666 4652
rect 3522 4643 3666 4651
rect 3522 4623 3530 4643
rect 3550 4623 3585 4643
rect 3605 4623 3638 4643
rect 3658 4623 3666 4643
rect 3522 4617 3666 4623
rect 3732 4647 3770 4655
rect 3848 4651 3884 4652
rect 3732 4627 3741 4647
rect 3761 4627 3770 4647
rect 3732 4618 3770 4627
rect 3799 4643 3884 4651
rect 3799 4623 3856 4643
rect 3876 4623 3884 4643
rect 3732 4617 3769 4618
rect 3799 4617 3884 4623
rect 3950 4647 3988 4655
rect 3950 4627 3959 4647
rect 3979 4627 3988 4647
rect 4120 4645 4132 4663
rect 4150 4645 4160 4663
rect 4120 4635 4160 4645
rect 3950 4618 3988 4627
rect 3950 4617 3987 4618
rect 3411 4589 3501 4595
rect 3411 4569 3427 4589
rect 3447 4587 3501 4589
rect 3447 4569 3472 4587
rect 3411 4567 3472 4569
rect 3492 4567 3501 4587
rect 3411 4561 3501 4567
rect 3424 4507 3461 4508
rect 3520 4507 3557 4508
rect 3576 4507 3612 4617
rect 3799 4596 3830 4617
rect 3795 4595 3830 4596
rect 3673 4585 3830 4595
rect 3673 4565 3690 4585
rect 3710 4565 3830 4585
rect 3673 4558 3830 4565
rect 3897 4588 4046 4596
rect 3897 4568 3908 4588
rect 3928 4568 3967 4588
rect 3987 4568 4046 4588
rect 3897 4561 4046 4568
rect 4112 4564 4164 4582
rect 3897 4560 3938 4561
rect 3631 4507 3668 4508
rect 2225 4492 2264 4507
rect 3324 4498 3462 4507
rect 2225 4491 2391 4492
rect 2517 4491 2557 4493
rect 2225 4465 2667 4491
rect 2225 4463 2391 4465
rect 1889 4351 1926 4359
rect 1889 4332 1897 4351
rect 1918 4332 1926 4351
rect 1889 4326 1926 4332
rect 2225 4285 2250 4463
rect 2290 4425 2354 4437
rect 2630 4433 2667 4465
rect 2693 4464 2884 4486
rect 3324 4478 3433 4498
rect 3453 4478 3462 4498
rect 3324 4471 3462 4478
rect 3520 4498 3668 4507
rect 3520 4478 3529 4498
rect 3549 4478 3639 4498
rect 3659 4478 3668 4498
rect 3324 4469 3420 4471
rect 3520 4468 3668 4478
rect 3727 4498 3764 4508
rect 3727 4478 3735 4498
rect 3755 4478 3764 4498
rect 3576 4467 3612 4468
rect 2848 4462 2884 4464
rect 2848 4433 2885 4462
rect 2290 4424 2325 4425
rect 2267 4419 2325 4424
rect 2267 4399 2270 4419
rect 2290 4405 2325 4419
rect 2345 4405 2354 4425
rect 2290 4397 2354 4405
rect 2316 4396 2354 4397
rect 2317 4395 2354 4396
rect 2420 4429 2456 4430
rect 2528 4429 2564 4430
rect 2420 4424 2564 4429
rect 2420 4421 2482 4424
rect 2420 4401 2428 4421
rect 2448 4401 2482 4421
rect 2420 4398 2482 4401
rect 2508 4421 2564 4424
rect 2508 4401 2536 4421
rect 2556 4401 2564 4421
rect 2508 4398 2564 4401
rect 2420 4395 2564 4398
rect 2630 4425 2668 4433
rect 2746 4429 2782 4430
rect 2630 4405 2639 4425
rect 2659 4405 2668 4425
rect 2630 4396 2668 4405
rect 2697 4421 2782 4429
rect 2697 4401 2754 4421
rect 2774 4401 2782 4421
rect 2630 4395 2667 4396
rect 2697 4395 2782 4401
rect 2848 4425 2886 4433
rect 2848 4405 2857 4425
rect 2877 4405 2886 4425
rect 3727 4411 3764 4478
rect 3799 4507 3830 4558
rect 4112 4546 4130 4564
rect 4148 4546 4164 4564
rect 3849 4507 3886 4508
rect 3799 4498 3886 4507
rect 3799 4478 3857 4498
rect 3877 4478 3886 4498
rect 3799 4468 3886 4478
rect 3945 4498 3982 4508
rect 3945 4478 3953 4498
rect 3973 4478 3982 4498
rect 3799 4467 3830 4468
rect 3424 4408 3461 4409
rect 3727 4408 3766 4411
rect 3423 4407 3766 4408
rect 3945 4407 3982 4478
rect 2848 4396 2886 4405
rect 3348 4402 3766 4407
rect 2848 4395 2885 4396
rect 2309 4367 2399 4373
rect 2309 4347 2325 4367
rect 2345 4365 2399 4367
rect 2345 4347 2370 4365
rect 2309 4345 2370 4347
rect 2390 4345 2399 4365
rect 2309 4339 2399 4345
rect 2322 4285 2359 4286
rect 2418 4285 2455 4286
rect 2474 4285 2510 4395
rect 2697 4374 2728 4395
rect 3348 4382 3351 4402
rect 3371 4382 3766 4402
rect 3795 4383 3982 4407
rect 2693 4373 2728 4374
rect 2571 4363 2728 4373
rect 2571 4343 2588 4363
rect 2608 4343 2728 4363
rect 2571 4336 2728 4343
rect 2795 4366 2944 4374
rect 2795 4346 2806 4366
rect 2826 4346 2865 4366
rect 2885 4346 2944 4366
rect 2795 4339 2944 4346
rect 3727 4357 3766 4382
rect 4112 4357 4164 4546
rect 3727 4339 4166 4357
rect 2795 4338 2836 4339
rect 2529 4285 2566 4286
rect 2225 4276 2360 4285
rect 2225 4256 2331 4276
rect 2351 4256 2360 4276
rect 2225 4249 2360 4256
rect 2418 4276 2566 4285
rect 2418 4256 2427 4276
rect 2447 4256 2537 4276
rect 2557 4256 2566 4276
rect 2225 4247 2318 4249
rect 2418 4246 2566 4256
rect 2625 4276 2662 4286
rect 2625 4256 2633 4276
rect 2653 4256 2662 4276
rect 2474 4245 2510 4246
rect 2322 4186 2359 4187
rect 2625 4186 2662 4256
rect 2697 4285 2728 4336
rect 3727 4321 4127 4339
rect 4145 4321 4166 4339
rect 3727 4315 4166 4321
rect 3733 4311 4166 4315
rect 4112 4309 4164 4311
rect 2747 4285 2784 4286
rect 2697 4276 2784 4285
rect 2697 4256 2755 4276
rect 2775 4256 2784 4276
rect 2697 4246 2784 4256
rect 2843 4276 2880 4286
rect 2843 4256 2851 4276
rect 2871 4256 2880 4276
rect 2697 4245 2728 4246
rect 2321 4185 2662 4186
rect 2843 4185 2880 4256
rect 4115 4244 4152 4249
rect 2246 4180 2662 4185
rect 2246 4160 2249 4180
rect 2269 4160 2662 4180
rect 2693 4161 2880 4185
rect 4106 4240 4153 4244
rect 4106 4222 4125 4240
rect 4143 4222 4153 4240
rect 3714 4163 3752 4164
rect 4106 4163 4153 4222
rect 2466 4159 2531 4160
rect 581 4081 619 4082
rect 180 4043 619 4081
rect 1491 4081 1499 4103
rect 1523 4081 1531 4103
rect 1491 4073 1531 4081
rect 2802 4125 2842 4133
rect 2802 4103 2810 4125
rect 2834 4103 2842 4125
rect 3714 4125 4153 4163
rect 3714 4124 3752 4125
rect 1802 4046 1867 4047
rect 180 3984 227 4043
rect 581 4042 619 4043
rect 180 3966 190 3984
rect 208 3966 227 3984
rect 180 3962 227 3966
rect 1453 4021 1640 4045
rect 1671 4026 2064 4046
rect 2084 4026 2087 4046
rect 1671 4021 2087 4026
rect 181 3957 218 3962
rect 1453 3950 1490 4021
rect 1671 4020 2012 4021
rect 1605 3960 1636 3961
rect 1453 3930 1462 3950
rect 1482 3930 1490 3950
rect 1453 3920 1490 3930
rect 1549 3950 1636 3960
rect 1549 3930 1558 3950
rect 1578 3930 1636 3950
rect 1549 3921 1636 3930
rect 1549 3920 1586 3921
rect 169 3895 221 3897
rect 167 3891 600 3895
rect 167 3885 606 3891
rect 167 3867 188 3885
rect 206 3867 606 3885
rect 1605 3870 1636 3921
rect 1671 3950 1708 4020
rect 1974 4019 2011 4020
rect 1823 3960 1859 3961
rect 1671 3930 1680 3950
rect 1700 3930 1708 3950
rect 1671 3920 1708 3930
rect 1767 3950 1915 3960
rect 2015 3957 2111 3959
rect 1767 3930 1776 3950
rect 1796 3930 1886 3950
rect 1906 3930 1915 3950
rect 1767 3921 1915 3930
rect 1973 3950 2111 3957
rect 1973 3930 1982 3950
rect 2002 3930 2111 3950
rect 1973 3921 2111 3930
rect 1767 3920 1804 3921
rect 1497 3867 1538 3868
rect 167 3849 606 3867
rect 169 3660 221 3849
rect 567 3824 606 3849
rect 1389 3860 1538 3867
rect 1389 3840 1448 3860
rect 1468 3840 1507 3860
rect 1527 3840 1538 3860
rect 1389 3832 1538 3840
rect 1605 3863 1762 3870
rect 1605 3843 1725 3863
rect 1745 3843 1762 3863
rect 1605 3833 1762 3843
rect 1605 3832 1640 3833
rect 351 3799 538 3823
rect 567 3804 962 3824
rect 982 3804 985 3824
rect 1605 3811 1636 3832
rect 1823 3811 1859 3921
rect 1878 3920 1915 3921
rect 1974 3920 2011 3921
rect 1934 3861 2024 3867
rect 1934 3841 1943 3861
rect 1963 3859 2024 3861
rect 1963 3841 1988 3859
rect 1934 3839 1988 3841
rect 2008 3839 2024 3859
rect 1934 3833 2024 3839
rect 1448 3810 1485 3811
rect 567 3799 985 3804
rect 1447 3801 1485 3810
rect 351 3728 388 3799
rect 567 3798 910 3799
rect 567 3795 606 3798
rect 872 3797 909 3798
rect 503 3738 534 3739
rect 351 3708 360 3728
rect 380 3708 388 3728
rect 351 3698 388 3708
rect 447 3728 534 3738
rect 447 3708 456 3728
rect 476 3708 534 3728
rect 447 3699 534 3708
rect 447 3698 484 3699
rect 169 3642 185 3660
rect 203 3642 221 3660
rect 503 3648 534 3699
rect 569 3728 606 3795
rect 1447 3781 1456 3801
rect 1476 3781 1485 3801
rect 1447 3773 1485 3781
rect 1551 3805 1636 3811
rect 1666 3810 1703 3811
rect 1551 3785 1559 3805
rect 1579 3785 1636 3805
rect 1551 3777 1636 3785
rect 1665 3801 1703 3810
rect 1665 3781 1674 3801
rect 1694 3781 1703 3801
rect 1551 3776 1587 3777
rect 1665 3773 1703 3781
rect 1769 3805 1913 3811
rect 1769 3785 1777 3805
rect 1797 3799 1885 3805
rect 1797 3785 1826 3799
rect 1769 3777 1826 3785
rect 1769 3776 1805 3777
rect 1849 3785 1885 3799
rect 1905 3785 1913 3805
rect 1849 3777 1913 3785
rect 1877 3776 1913 3777
rect 1979 3810 2016 3811
rect 1979 3809 2017 3810
rect 1979 3801 2043 3809
rect 1979 3781 1988 3801
rect 2008 3787 2043 3801
rect 2063 3787 2066 3807
rect 2008 3782 2066 3787
rect 2008 3781 2043 3782
rect 1448 3744 1485 3773
rect 1449 3742 1485 3744
rect 721 3738 757 3739
rect 569 3708 578 3728
rect 598 3708 606 3728
rect 569 3698 606 3708
rect 665 3728 813 3738
rect 913 3735 1009 3737
rect 665 3708 674 3728
rect 694 3708 784 3728
rect 804 3708 813 3728
rect 665 3699 813 3708
rect 871 3728 1009 3735
rect 871 3708 880 3728
rect 900 3708 1009 3728
rect 1449 3720 1640 3742
rect 1666 3741 1703 3773
rect 1979 3769 2043 3781
rect 2083 3743 2110 3921
rect 2407 3874 2444 3880
rect 2407 3855 2415 3874
rect 2436 3855 2444 3874
rect 2407 3847 2444 3855
rect 1942 3741 2110 3743
rect 1666 3715 2110 3741
rect 1776 3713 1816 3715
rect 1942 3714 2110 3715
rect 871 3699 1009 3708
rect 2069 3709 2110 3714
rect 665 3698 702 3699
rect 395 3645 436 3646
rect 169 3624 221 3642
rect 287 3638 436 3645
rect 287 3618 346 3638
rect 366 3618 405 3638
rect 425 3618 436 3638
rect 287 3610 436 3618
rect 503 3641 660 3648
rect 503 3621 623 3641
rect 643 3621 660 3641
rect 503 3611 660 3621
rect 503 3610 538 3611
rect 503 3589 534 3610
rect 721 3589 757 3699
rect 776 3698 813 3699
rect 872 3698 909 3699
rect 832 3639 922 3645
rect 832 3619 841 3639
rect 861 3637 922 3639
rect 861 3619 886 3637
rect 832 3617 886 3619
rect 906 3617 922 3637
rect 832 3611 922 3617
rect 346 3588 383 3589
rect 345 3579 383 3588
rect 173 3561 213 3571
rect 173 3543 183 3561
rect 201 3543 213 3561
rect 345 3559 354 3579
rect 374 3559 383 3579
rect 345 3551 383 3559
rect 449 3583 534 3589
rect 564 3588 601 3589
rect 449 3563 457 3583
rect 477 3563 534 3583
rect 449 3555 534 3563
rect 563 3579 601 3588
rect 563 3559 572 3579
rect 592 3559 601 3579
rect 449 3554 485 3555
rect 563 3551 601 3559
rect 667 3583 811 3589
rect 667 3563 675 3583
rect 695 3563 728 3583
rect 748 3563 783 3583
rect 803 3563 811 3583
rect 667 3555 811 3563
rect 667 3554 703 3555
rect 775 3554 811 3555
rect 877 3588 914 3589
rect 877 3587 915 3588
rect 877 3579 941 3587
rect 877 3559 886 3579
rect 906 3565 941 3579
rect 961 3565 964 3585
rect 906 3560 964 3565
rect 906 3559 941 3560
rect 173 3487 213 3543
rect 346 3522 383 3551
rect 347 3520 383 3522
rect 347 3498 538 3520
rect 564 3519 601 3551
rect 877 3547 941 3559
rect 981 3521 1008 3699
rect 840 3519 1008 3521
rect 564 3509 1008 3519
rect 1149 3615 1336 3639
rect 1367 3620 1760 3640
rect 1780 3620 1783 3640
rect 1367 3615 1783 3620
rect 1149 3544 1186 3615
rect 1367 3614 1708 3615
rect 1301 3554 1332 3555
rect 1149 3524 1158 3544
rect 1178 3524 1186 3544
rect 1149 3514 1186 3524
rect 1245 3544 1332 3554
rect 1245 3524 1254 3544
rect 1274 3524 1332 3544
rect 1245 3515 1332 3524
rect 1245 3514 1282 3515
rect 170 3482 213 3487
rect 561 3493 1008 3509
rect 561 3487 589 3493
rect 840 3492 1008 3493
rect 170 3479 320 3482
rect 561 3479 588 3487
rect 170 3477 588 3479
rect 170 3459 179 3477
rect 197 3459 588 3477
rect 1301 3464 1332 3515
rect 1367 3544 1404 3614
rect 1670 3613 1707 3614
rect 1519 3554 1555 3555
rect 1367 3524 1376 3544
rect 1396 3524 1404 3544
rect 1367 3514 1404 3524
rect 1463 3544 1611 3554
rect 1711 3551 1807 3553
rect 1463 3524 1472 3544
rect 1492 3524 1582 3544
rect 1602 3524 1611 3544
rect 1463 3515 1611 3524
rect 1669 3544 1807 3551
rect 1669 3524 1678 3544
rect 1698 3524 1807 3544
rect 2069 3527 2109 3709
rect 1669 3515 1807 3524
rect 1463 3514 1500 3515
rect 1193 3461 1234 3462
rect 170 3456 588 3459
rect 170 3450 213 3456
rect 173 3447 213 3450
rect 1085 3454 1234 3461
rect 570 3438 610 3439
rect 281 3421 610 3438
rect 1085 3434 1144 3454
rect 1164 3434 1203 3454
rect 1223 3434 1234 3454
rect 1085 3426 1234 3434
rect 1301 3457 1458 3464
rect 1301 3437 1421 3457
rect 1441 3437 1458 3457
rect 1301 3427 1458 3437
rect 1301 3426 1336 3427
rect 165 3378 208 3389
rect 165 3360 177 3378
rect 195 3360 208 3378
rect 165 3334 208 3360
rect 281 3334 308 3421
rect 570 3412 610 3421
rect 165 3313 308 3334
rect 352 3386 386 3402
rect 570 3392 963 3412
rect 983 3392 986 3412
rect 1301 3405 1332 3426
rect 1519 3405 1555 3515
rect 1574 3514 1611 3515
rect 1670 3514 1707 3515
rect 1630 3455 1720 3461
rect 1630 3435 1639 3455
rect 1659 3453 1720 3455
rect 1659 3435 1684 3453
rect 1630 3433 1684 3435
rect 1704 3433 1720 3453
rect 1630 3427 1720 3433
rect 1144 3404 1181 3405
rect 570 3387 986 3392
rect 1143 3395 1181 3404
rect 570 3386 911 3387
rect 352 3316 389 3386
rect 504 3326 535 3327
rect 165 3311 302 3313
rect 165 3269 208 3311
rect 352 3296 361 3316
rect 381 3296 389 3316
rect 352 3286 389 3296
rect 448 3316 535 3326
rect 448 3296 457 3316
rect 477 3296 535 3316
rect 448 3287 535 3296
rect 448 3286 485 3287
rect 163 3259 208 3269
rect 163 3241 172 3259
rect 190 3241 208 3259
rect 163 3235 208 3241
rect 504 3236 535 3287
rect 570 3316 607 3386
rect 873 3385 910 3386
rect 1143 3375 1152 3395
rect 1172 3375 1181 3395
rect 1143 3367 1181 3375
rect 1247 3399 1332 3405
rect 1362 3404 1399 3405
rect 1247 3379 1255 3399
rect 1275 3379 1332 3399
rect 1247 3371 1332 3379
rect 1361 3395 1399 3404
rect 1361 3375 1370 3395
rect 1390 3375 1399 3395
rect 1247 3370 1283 3371
rect 1361 3367 1399 3375
rect 1465 3399 1609 3405
rect 1465 3379 1473 3399
rect 1493 3380 1525 3399
rect 1546 3380 1581 3399
rect 1493 3379 1581 3380
rect 1601 3379 1609 3399
rect 1465 3371 1609 3379
rect 1465 3370 1501 3371
rect 1573 3370 1609 3371
rect 1675 3404 1712 3405
rect 1675 3403 1713 3404
rect 1675 3395 1739 3403
rect 1675 3375 1684 3395
rect 1704 3381 1739 3395
rect 1759 3381 1762 3401
rect 1704 3376 1762 3381
rect 1704 3375 1739 3376
rect 1144 3338 1181 3367
rect 1145 3336 1181 3338
rect 722 3326 758 3327
rect 570 3296 579 3316
rect 599 3296 607 3316
rect 570 3286 607 3296
rect 666 3316 814 3326
rect 914 3323 1010 3325
rect 666 3296 675 3316
rect 695 3296 785 3316
rect 805 3296 814 3316
rect 666 3287 814 3296
rect 872 3316 1010 3323
rect 872 3296 881 3316
rect 901 3296 1010 3316
rect 1145 3314 1336 3336
rect 1362 3335 1399 3367
rect 1675 3363 1739 3375
rect 1779 3337 1806 3515
rect 1638 3335 1806 3337
rect 1362 3309 1806 3335
rect 872 3287 1010 3296
rect 666 3286 703 3287
rect 163 3232 200 3235
rect 396 3233 437 3234
rect 288 3226 437 3233
rect 288 3206 347 3226
rect 367 3206 406 3226
rect 426 3206 437 3226
rect 288 3198 437 3206
rect 504 3229 661 3236
rect 504 3209 624 3229
rect 644 3209 661 3229
rect 504 3199 661 3209
rect 504 3198 539 3199
rect 504 3177 535 3198
rect 722 3177 758 3287
rect 777 3286 814 3287
rect 873 3286 910 3287
rect 833 3227 923 3233
rect 833 3207 842 3227
rect 862 3225 923 3227
rect 862 3207 887 3225
rect 833 3205 887 3207
rect 907 3205 923 3225
rect 833 3199 923 3205
rect 347 3176 384 3177
rect 160 3168 197 3170
rect 160 3160 202 3168
rect 160 3142 170 3160
rect 188 3142 202 3160
rect 160 3133 202 3142
rect 346 3167 384 3176
rect 346 3147 355 3167
rect 375 3147 384 3167
rect 346 3139 384 3147
rect 450 3171 535 3177
rect 565 3176 602 3177
rect 450 3151 458 3171
rect 478 3151 535 3171
rect 450 3143 535 3151
rect 564 3167 602 3176
rect 564 3147 573 3167
rect 593 3147 602 3167
rect 450 3142 486 3143
rect 564 3139 602 3147
rect 668 3175 812 3177
rect 668 3171 720 3175
rect 668 3151 676 3171
rect 696 3155 720 3171
rect 740 3171 812 3175
rect 740 3155 784 3171
rect 696 3151 784 3155
rect 804 3151 812 3171
rect 668 3143 812 3151
rect 668 3142 704 3143
rect 776 3142 812 3143
rect 878 3176 915 3177
rect 878 3175 916 3176
rect 878 3167 942 3175
rect 878 3147 887 3167
rect 907 3153 942 3167
rect 962 3153 965 3173
rect 907 3148 965 3153
rect 907 3147 942 3148
rect 161 3108 202 3133
rect 347 3108 384 3139
rect 565 3108 602 3139
rect 878 3135 942 3147
rect 982 3109 1009 3287
rect 161 3081 210 3108
rect 346 3082 395 3108
rect 564 3107 645 3108
rect 841 3107 1009 3109
rect 564 3082 1009 3107
rect 565 3081 1009 3082
rect 163 3048 210 3081
rect 566 3048 606 3081
rect 841 3080 1009 3081
rect 1472 3085 1512 3309
rect 1638 3308 1806 3309
rect 1472 3063 1480 3085
rect 1504 3063 1512 3085
rect 1472 3055 1512 3063
rect 163 3009 606 3048
rect 163 2966 210 3009
rect 566 3004 606 3009
rect 1231 3007 1418 3031
rect 1449 3012 1842 3032
rect 1862 3012 1865 3032
rect 1449 3007 1865 3012
rect 163 2948 173 2966
rect 191 2948 210 2966
rect 163 2944 210 2948
rect 164 2939 201 2944
rect 1231 2936 1268 3007
rect 1449 3006 1790 3007
rect 1383 2946 1414 2947
rect 1231 2916 1240 2936
rect 1260 2916 1268 2936
rect 1231 2906 1268 2916
rect 1327 2936 1414 2946
rect 1327 2916 1336 2936
rect 1356 2916 1414 2936
rect 1327 2907 1414 2916
rect 1327 2906 1364 2907
rect 152 2877 204 2879
rect 150 2873 583 2877
rect 150 2867 589 2873
rect 150 2849 171 2867
rect 189 2849 589 2867
rect 1383 2856 1414 2907
rect 1449 2936 1486 3006
rect 1752 3005 1789 3006
rect 1601 2946 1637 2947
rect 1449 2916 1458 2936
rect 1478 2916 1486 2936
rect 1449 2906 1486 2916
rect 1545 2936 1693 2946
rect 1793 2943 1889 2945
rect 1545 2916 1554 2936
rect 1574 2916 1664 2936
rect 1684 2916 1693 2936
rect 1545 2907 1693 2916
rect 1751 2936 1889 2943
rect 1751 2916 1760 2936
rect 1780 2916 1889 2936
rect 1751 2907 1889 2916
rect 1545 2906 1582 2907
rect 1275 2853 1316 2854
rect 150 2831 589 2849
rect 152 2642 204 2831
rect 550 2806 589 2831
rect 1167 2846 1316 2853
rect 1167 2826 1226 2846
rect 1246 2826 1285 2846
rect 1305 2826 1316 2846
rect 1167 2818 1316 2826
rect 1383 2849 1540 2856
rect 1383 2829 1503 2849
rect 1523 2829 1540 2849
rect 1383 2819 1540 2829
rect 1383 2818 1418 2819
rect 334 2781 521 2805
rect 550 2786 945 2806
rect 965 2786 968 2806
rect 1383 2797 1414 2818
rect 1601 2797 1637 2907
rect 1656 2906 1693 2907
rect 1752 2906 1789 2907
rect 1712 2847 1802 2853
rect 1712 2827 1721 2847
rect 1741 2845 1802 2847
rect 1741 2827 1766 2845
rect 1712 2825 1766 2827
rect 1786 2825 1802 2845
rect 1712 2819 1802 2825
rect 1226 2796 1263 2797
rect 550 2781 968 2786
rect 1225 2787 1263 2796
rect 334 2710 371 2781
rect 550 2780 893 2781
rect 550 2777 589 2780
rect 855 2779 892 2780
rect 486 2720 517 2721
rect 334 2690 343 2710
rect 363 2690 371 2710
rect 334 2680 371 2690
rect 430 2710 517 2720
rect 430 2690 439 2710
rect 459 2690 517 2710
rect 430 2681 517 2690
rect 430 2680 467 2681
rect 152 2624 168 2642
rect 186 2624 204 2642
rect 486 2630 517 2681
rect 552 2710 589 2777
rect 1225 2767 1234 2787
rect 1254 2767 1263 2787
rect 1225 2759 1263 2767
rect 1329 2791 1414 2797
rect 1444 2796 1481 2797
rect 1329 2771 1337 2791
rect 1357 2771 1414 2791
rect 1329 2763 1414 2771
rect 1443 2787 1481 2796
rect 1443 2767 1452 2787
rect 1472 2767 1481 2787
rect 1329 2762 1365 2763
rect 1443 2759 1481 2767
rect 1547 2792 1691 2797
rect 1547 2791 1609 2792
rect 1547 2771 1555 2791
rect 1575 2773 1609 2791
rect 1630 2791 1691 2792
rect 1630 2773 1663 2791
rect 1575 2771 1663 2773
rect 1683 2771 1691 2791
rect 1547 2763 1691 2771
rect 1547 2762 1583 2763
rect 1655 2762 1691 2763
rect 1757 2796 1794 2797
rect 1757 2795 1795 2796
rect 1757 2787 1821 2795
rect 1757 2767 1766 2787
rect 1786 2773 1821 2787
rect 1841 2773 1844 2793
rect 1786 2768 1844 2773
rect 1786 2767 1821 2768
rect 1226 2730 1263 2759
rect 1227 2728 1263 2730
rect 704 2720 740 2721
rect 552 2690 561 2710
rect 581 2690 589 2710
rect 552 2680 589 2690
rect 648 2710 796 2720
rect 896 2717 992 2719
rect 648 2690 657 2710
rect 677 2690 767 2710
rect 787 2690 796 2710
rect 648 2681 796 2690
rect 854 2710 992 2717
rect 854 2690 863 2710
rect 883 2690 992 2710
rect 1227 2706 1418 2728
rect 1444 2727 1481 2759
rect 1757 2755 1821 2767
rect 1861 2729 1888 2907
rect 1720 2727 1888 2729
rect 1444 2713 1888 2727
rect 1444 2701 1891 2713
rect 1487 2699 1520 2701
rect 854 2681 992 2690
rect 648 2680 685 2681
rect 378 2627 419 2628
rect 152 2606 204 2624
rect 270 2620 419 2627
rect 270 2600 329 2620
rect 349 2600 388 2620
rect 408 2600 419 2620
rect 270 2592 419 2600
rect 486 2623 643 2630
rect 486 2603 606 2623
rect 626 2603 643 2623
rect 486 2593 643 2603
rect 486 2592 521 2593
rect 486 2571 517 2592
rect 704 2571 740 2681
rect 759 2680 796 2681
rect 855 2680 892 2681
rect 815 2621 905 2627
rect 815 2601 824 2621
rect 844 2619 905 2621
rect 844 2601 869 2619
rect 815 2599 869 2601
rect 889 2599 905 2619
rect 815 2593 905 2599
rect 329 2570 366 2571
rect 328 2561 366 2570
rect 156 2543 196 2553
rect 156 2525 166 2543
rect 184 2525 196 2543
rect 328 2541 337 2561
rect 357 2541 366 2561
rect 328 2533 366 2541
rect 432 2565 517 2571
rect 547 2570 584 2571
rect 432 2545 440 2565
rect 460 2545 517 2565
rect 432 2537 517 2545
rect 546 2561 584 2570
rect 546 2541 555 2561
rect 575 2541 584 2561
rect 432 2536 468 2537
rect 546 2533 584 2541
rect 650 2565 794 2571
rect 650 2545 658 2565
rect 678 2545 711 2565
rect 731 2545 766 2565
rect 786 2545 794 2565
rect 650 2537 794 2545
rect 650 2536 686 2537
rect 758 2536 794 2537
rect 860 2570 897 2571
rect 860 2569 898 2570
rect 860 2561 924 2569
rect 860 2541 869 2561
rect 889 2547 924 2561
rect 944 2547 947 2567
rect 889 2542 947 2547
rect 889 2541 924 2542
rect 156 2469 196 2525
rect 329 2504 366 2533
rect 330 2502 366 2504
rect 330 2480 521 2502
rect 547 2501 584 2533
rect 860 2529 924 2541
rect 964 2503 991 2681
rect 1849 2656 1891 2701
rect 823 2501 991 2503
rect 547 2491 991 2501
rect 1132 2597 1319 2621
rect 1350 2602 1743 2622
rect 1763 2602 1766 2622
rect 1350 2597 1766 2602
rect 1132 2526 1169 2597
rect 1350 2596 1691 2597
rect 1284 2536 1315 2537
rect 1132 2506 1141 2526
rect 1161 2506 1169 2526
rect 1132 2496 1169 2506
rect 1228 2526 1315 2536
rect 1228 2506 1237 2526
rect 1257 2506 1315 2526
rect 1228 2497 1315 2506
rect 1228 2496 1265 2497
rect 153 2464 196 2469
rect 544 2475 991 2491
rect 544 2469 572 2475
rect 823 2474 991 2475
rect 153 2461 303 2464
rect 544 2461 571 2469
rect 153 2459 571 2461
rect 153 2441 162 2459
rect 180 2441 571 2459
rect 1284 2446 1315 2497
rect 1350 2526 1387 2596
rect 1653 2595 1690 2596
rect 1502 2536 1538 2537
rect 1350 2506 1359 2526
rect 1379 2506 1387 2526
rect 1350 2496 1387 2506
rect 1446 2526 1594 2536
rect 1694 2533 1790 2535
rect 1446 2506 1455 2526
rect 1475 2506 1565 2526
rect 1585 2506 1594 2526
rect 1446 2497 1594 2506
rect 1652 2526 1790 2533
rect 1652 2506 1661 2526
rect 1681 2506 1790 2526
rect 1652 2497 1790 2506
rect 1446 2496 1483 2497
rect 1176 2443 1217 2444
rect 153 2438 571 2441
rect 153 2432 196 2438
rect 156 2429 196 2432
rect 1071 2436 1217 2443
rect 553 2420 593 2421
rect 264 2403 593 2420
rect 1071 2416 1127 2436
rect 1147 2416 1186 2436
rect 1206 2416 1217 2436
rect 1071 2408 1217 2416
rect 1284 2439 1441 2446
rect 1284 2419 1404 2439
rect 1424 2419 1441 2439
rect 1284 2409 1441 2419
rect 1284 2408 1319 2409
rect 148 2360 191 2371
rect 148 2342 160 2360
rect 178 2342 191 2360
rect 148 2316 191 2342
rect 264 2316 291 2403
rect 553 2394 593 2403
rect 148 2295 291 2316
rect 335 2368 369 2384
rect 553 2374 946 2394
rect 966 2374 969 2394
rect 1284 2387 1315 2408
rect 1502 2387 1538 2497
rect 1557 2496 1594 2497
rect 1653 2496 1690 2497
rect 1613 2437 1703 2443
rect 1613 2417 1622 2437
rect 1642 2435 1703 2437
rect 1642 2417 1667 2435
rect 1613 2415 1667 2417
rect 1687 2415 1703 2435
rect 1613 2409 1703 2415
rect 1127 2386 1164 2387
rect 553 2369 969 2374
rect 1126 2377 1164 2386
rect 553 2368 894 2369
rect 335 2298 372 2368
rect 487 2308 518 2309
rect 148 2293 285 2295
rect 148 2251 191 2293
rect 335 2278 344 2298
rect 364 2278 372 2298
rect 335 2268 372 2278
rect 431 2298 518 2308
rect 431 2278 440 2298
rect 460 2278 518 2298
rect 431 2269 518 2278
rect 431 2268 468 2269
rect 146 2241 191 2251
rect 146 2223 155 2241
rect 173 2223 191 2241
rect 146 2217 191 2223
rect 487 2218 518 2269
rect 553 2298 590 2368
rect 856 2367 893 2368
rect 1126 2357 1135 2377
rect 1155 2357 1164 2377
rect 1126 2349 1164 2357
rect 1230 2381 1315 2387
rect 1345 2386 1382 2387
rect 1230 2361 1238 2381
rect 1258 2361 1315 2381
rect 1230 2353 1315 2361
rect 1344 2377 1382 2386
rect 1344 2357 1353 2377
rect 1373 2357 1382 2377
rect 1230 2352 1266 2353
rect 1344 2349 1382 2357
rect 1448 2381 1592 2387
rect 1448 2361 1456 2381
rect 1476 2378 1564 2381
rect 1476 2361 1511 2378
rect 1448 2360 1511 2361
rect 1530 2361 1564 2378
rect 1584 2361 1592 2381
rect 1530 2360 1592 2361
rect 1448 2353 1592 2360
rect 1448 2352 1484 2353
rect 1556 2352 1592 2353
rect 1658 2386 1695 2387
rect 1658 2385 1696 2386
rect 1718 2385 1745 2389
rect 1658 2383 1745 2385
rect 1658 2377 1722 2383
rect 1658 2357 1667 2377
rect 1687 2363 1722 2377
rect 1742 2363 1745 2383
rect 1687 2358 1745 2363
rect 1687 2357 1722 2358
rect 1127 2320 1164 2349
rect 1128 2318 1164 2320
rect 705 2308 741 2309
rect 553 2278 562 2298
rect 582 2278 590 2298
rect 553 2268 590 2278
rect 649 2298 797 2308
rect 897 2305 993 2307
rect 649 2278 658 2298
rect 678 2278 768 2298
rect 788 2278 797 2298
rect 649 2269 797 2278
rect 855 2298 993 2305
rect 855 2278 864 2298
rect 884 2278 993 2298
rect 1128 2296 1319 2318
rect 1345 2317 1382 2349
rect 1658 2345 1722 2357
rect 1762 2319 1789 2497
rect 1621 2317 1789 2319
rect 1345 2291 1789 2317
rect 855 2269 993 2278
rect 649 2268 686 2269
rect 146 2214 183 2217
rect 379 2215 420 2216
rect 271 2208 420 2215
rect 271 2188 330 2208
rect 350 2188 389 2208
rect 409 2188 420 2208
rect 271 2180 420 2188
rect 487 2211 644 2218
rect 487 2191 607 2211
rect 627 2191 644 2211
rect 487 2181 644 2191
rect 487 2180 522 2181
rect 487 2159 518 2180
rect 705 2159 741 2269
rect 760 2268 797 2269
rect 856 2268 893 2269
rect 816 2209 906 2215
rect 816 2189 825 2209
rect 845 2207 906 2209
rect 845 2189 870 2207
rect 816 2187 870 2189
rect 890 2187 906 2207
rect 816 2181 906 2187
rect 330 2158 367 2159
rect 142 2150 180 2152
rect 142 2142 185 2150
rect 142 2124 153 2142
rect 171 2124 185 2142
rect 142 2097 185 2124
rect 329 2149 367 2158
rect 329 2129 338 2149
rect 358 2129 367 2149
rect 329 2121 367 2129
rect 433 2153 518 2159
rect 548 2158 585 2159
rect 433 2133 441 2153
rect 461 2133 518 2153
rect 433 2125 518 2133
rect 547 2149 585 2158
rect 547 2129 556 2149
rect 576 2129 585 2149
rect 433 2124 469 2125
rect 547 2121 585 2129
rect 651 2157 795 2159
rect 651 2153 703 2157
rect 651 2133 659 2153
rect 679 2137 703 2153
rect 723 2153 795 2157
rect 723 2137 767 2153
rect 679 2133 767 2137
rect 787 2133 795 2153
rect 651 2125 795 2133
rect 651 2124 687 2125
rect 759 2124 795 2125
rect 861 2158 898 2159
rect 861 2157 899 2158
rect 861 2149 925 2157
rect 861 2129 870 2149
rect 890 2135 925 2149
rect 945 2135 948 2155
rect 890 2130 948 2135
rect 890 2129 925 2130
rect 143 2090 185 2097
rect 330 2090 367 2121
rect 548 2090 585 2121
rect 861 2117 925 2129
rect 965 2091 992 2269
rect 143 2050 188 2090
rect 330 2065 475 2090
rect 548 2089 628 2090
rect 824 2089 992 2091
rect 548 2073 992 2089
rect 332 2064 475 2065
rect 547 2063 992 2073
rect 143 2029 190 2050
rect 547 2029 588 2063
rect 824 2062 992 2063
rect 1455 2067 1495 2291
rect 1621 2290 1789 2291
rect 1853 2323 1886 2656
rect 1853 2315 1890 2323
rect 1853 2296 1861 2315
rect 1882 2296 1890 2315
rect 1853 2290 1890 2296
rect 1455 2045 1463 2067
rect 1487 2045 1495 2067
rect 1455 2037 1495 2045
rect 143 1999 588 2029
rect 1626 2012 1691 2013
rect 143 1996 566 1999
rect 143 1948 190 1996
rect 143 1930 153 1948
rect 171 1930 190 1948
rect 143 1926 190 1930
rect 1277 1987 1464 2011
rect 1495 1992 1888 2012
rect 1908 1992 1911 2012
rect 1495 1987 1911 1992
rect 144 1921 181 1926
rect 1277 1916 1314 1987
rect 1495 1986 1836 1987
rect 1429 1926 1460 1927
rect 1277 1896 1286 1916
rect 1306 1896 1314 1916
rect 1277 1886 1314 1896
rect 1373 1916 1460 1926
rect 1373 1896 1382 1916
rect 1402 1896 1460 1916
rect 1373 1887 1460 1896
rect 1373 1886 1410 1887
rect 132 1859 184 1861
rect 130 1855 563 1859
rect 130 1849 569 1855
rect 130 1831 151 1849
rect 169 1831 569 1849
rect 1429 1836 1460 1887
rect 1495 1916 1532 1986
rect 1798 1985 1835 1986
rect 1647 1926 1683 1927
rect 1495 1896 1504 1916
rect 1524 1896 1532 1916
rect 1495 1886 1532 1896
rect 1591 1916 1739 1926
rect 1839 1923 1935 1925
rect 1591 1896 1600 1916
rect 1620 1896 1710 1916
rect 1730 1896 1739 1916
rect 1591 1887 1739 1896
rect 1797 1916 1935 1923
rect 1797 1896 1806 1916
rect 1826 1896 1935 1916
rect 1797 1887 1935 1896
rect 1591 1886 1628 1887
rect 1321 1833 1362 1834
rect 130 1813 569 1831
rect 132 1624 184 1813
rect 530 1788 569 1813
rect 1213 1826 1362 1833
rect 1213 1806 1272 1826
rect 1292 1806 1331 1826
rect 1351 1806 1362 1826
rect 1213 1798 1362 1806
rect 1429 1829 1586 1836
rect 1429 1809 1549 1829
rect 1569 1809 1586 1829
rect 1429 1799 1586 1809
rect 1429 1798 1464 1799
rect 314 1763 501 1787
rect 530 1768 925 1788
rect 945 1768 948 1788
rect 1429 1777 1460 1798
rect 1647 1777 1683 1887
rect 1702 1886 1739 1887
rect 1798 1886 1835 1887
rect 1758 1827 1848 1833
rect 1758 1807 1767 1827
rect 1787 1825 1848 1827
rect 1787 1807 1812 1825
rect 1758 1805 1812 1807
rect 1832 1805 1848 1825
rect 1758 1799 1848 1805
rect 1272 1776 1309 1777
rect 530 1763 948 1768
rect 1271 1767 1309 1776
rect 314 1692 351 1763
rect 530 1762 873 1763
rect 530 1759 569 1762
rect 835 1761 872 1762
rect 466 1702 497 1703
rect 314 1672 323 1692
rect 343 1672 351 1692
rect 314 1662 351 1672
rect 410 1692 497 1702
rect 410 1672 419 1692
rect 439 1672 497 1692
rect 410 1663 497 1672
rect 410 1662 447 1663
rect 132 1606 148 1624
rect 166 1606 184 1624
rect 466 1612 497 1663
rect 532 1692 569 1759
rect 1271 1747 1280 1767
rect 1300 1747 1309 1767
rect 1271 1739 1309 1747
rect 1375 1771 1460 1777
rect 1490 1776 1527 1777
rect 1375 1751 1383 1771
rect 1403 1751 1460 1771
rect 1375 1743 1460 1751
rect 1489 1767 1527 1776
rect 1489 1747 1498 1767
rect 1518 1747 1527 1767
rect 1375 1742 1411 1743
rect 1489 1739 1527 1747
rect 1593 1775 1737 1777
rect 1593 1771 1653 1775
rect 1593 1751 1601 1771
rect 1621 1753 1653 1771
rect 1676 1771 1737 1775
rect 1676 1753 1709 1771
rect 1621 1751 1709 1753
rect 1729 1751 1737 1771
rect 1593 1743 1737 1751
rect 1593 1742 1629 1743
rect 1701 1742 1737 1743
rect 1803 1776 1840 1777
rect 1803 1775 1841 1776
rect 1803 1767 1867 1775
rect 1803 1747 1812 1767
rect 1832 1753 1867 1767
rect 1887 1753 1890 1773
rect 1832 1748 1890 1753
rect 1832 1747 1867 1748
rect 1272 1710 1309 1739
rect 1273 1708 1309 1710
rect 684 1702 720 1703
rect 532 1672 541 1692
rect 561 1672 569 1692
rect 532 1662 569 1672
rect 628 1692 776 1702
rect 876 1699 972 1701
rect 628 1672 637 1692
rect 657 1672 747 1692
rect 767 1672 776 1692
rect 628 1663 776 1672
rect 834 1692 972 1699
rect 834 1672 843 1692
rect 863 1672 972 1692
rect 1273 1686 1464 1708
rect 1490 1707 1527 1739
rect 1803 1735 1867 1747
rect 1490 1706 1765 1707
rect 1907 1706 1934 1887
rect 1490 1681 1934 1706
rect 2070 1712 2109 3527
rect 2411 3514 2444 3847
rect 2508 3879 2676 3880
rect 2802 3879 2842 4103
rect 3305 4107 3473 4108
rect 3714 4107 3749 4124
rect 4106 4114 4153 4125
rect 3305 4081 3749 4107
rect 3305 4079 3473 4081
rect 3669 4080 3749 4081
rect 3904 4080 3971 4106
rect 4110 4080 4153 4114
rect 3305 3901 3332 4079
rect 3372 4041 3436 4053
rect 3712 4049 3749 4080
rect 3930 4049 3967 4080
rect 4112 4055 4153 4080
rect 3372 4040 3407 4041
rect 3349 4035 3407 4040
rect 3349 4015 3352 4035
rect 3372 4021 3407 4035
rect 3427 4021 3436 4041
rect 3372 4013 3436 4021
rect 3398 4012 3436 4013
rect 3399 4011 3436 4012
rect 3502 4045 3538 4046
rect 3610 4045 3646 4046
rect 3502 4037 3646 4045
rect 3502 4017 3510 4037
rect 3530 4033 3618 4037
rect 3530 4017 3574 4033
rect 3502 4013 3574 4017
rect 3594 4017 3618 4033
rect 3638 4017 3646 4037
rect 3594 4013 3646 4017
rect 3502 4011 3646 4013
rect 3712 4041 3750 4049
rect 3828 4045 3864 4046
rect 3712 4021 3721 4041
rect 3741 4021 3750 4041
rect 3712 4012 3750 4021
rect 3779 4037 3864 4045
rect 3779 4017 3836 4037
rect 3856 4017 3864 4037
rect 3712 4011 3749 4012
rect 3779 4011 3864 4017
rect 3930 4041 3968 4049
rect 3930 4021 3939 4041
rect 3959 4021 3968 4041
rect 3930 4012 3968 4021
rect 4112 4046 4154 4055
rect 4112 4028 4126 4046
rect 4144 4028 4154 4046
rect 4112 4020 4154 4028
rect 4117 4018 4154 4020
rect 3930 4011 3967 4012
rect 3391 3983 3481 3989
rect 3391 3963 3407 3983
rect 3427 3981 3481 3983
rect 3427 3963 3452 3981
rect 3391 3961 3452 3963
rect 3472 3961 3481 3981
rect 3391 3955 3481 3961
rect 3404 3901 3441 3902
rect 3500 3901 3537 3902
rect 3556 3901 3592 4011
rect 3779 3990 3810 4011
rect 3775 3989 3810 3990
rect 3653 3979 3810 3989
rect 3653 3959 3670 3979
rect 3690 3959 3810 3979
rect 3653 3952 3810 3959
rect 3877 3982 4026 3990
rect 3877 3962 3888 3982
rect 3908 3962 3947 3982
rect 3967 3962 4026 3982
rect 3877 3955 4026 3962
rect 3877 3954 3918 3955
rect 4114 3953 4151 3956
rect 3611 3901 3648 3902
rect 3304 3892 3442 3901
rect 2508 3853 2952 3879
rect 2508 3851 2676 3853
rect 2508 3673 2535 3851
rect 2575 3813 2639 3825
rect 2915 3821 2952 3853
rect 2978 3852 3169 3874
rect 3304 3872 3413 3892
rect 3433 3872 3442 3892
rect 3304 3865 3442 3872
rect 3500 3892 3648 3901
rect 3500 3872 3509 3892
rect 3529 3872 3619 3892
rect 3639 3872 3648 3892
rect 3304 3863 3400 3865
rect 3500 3862 3648 3872
rect 3707 3892 3744 3902
rect 3707 3872 3715 3892
rect 3735 3872 3744 3892
rect 3556 3861 3592 3862
rect 3133 3850 3169 3852
rect 3133 3821 3170 3850
rect 2575 3812 2610 3813
rect 2552 3807 2610 3812
rect 2552 3787 2555 3807
rect 2575 3793 2610 3807
rect 2630 3793 2639 3813
rect 2575 3787 2639 3793
rect 2552 3785 2639 3787
rect 2552 3781 2579 3785
rect 2601 3784 2639 3785
rect 2602 3783 2639 3784
rect 2705 3817 2741 3818
rect 2813 3817 2849 3818
rect 2705 3810 2849 3817
rect 2705 3809 2767 3810
rect 2705 3789 2713 3809
rect 2733 3792 2767 3809
rect 2786 3809 2849 3810
rect 2786 3792 2821 3809
rect 2733 3789 2821 3792
rect 2841 3789 2849 3809
rect 2705 3783 2849 3789
rect 2915 3813 2953 3821
rect 3031 3817 3067 3818
rect 2915 3793 2924 3813
rect 2944 3793 2953 3813
rect 2915 3784 2953 3793
rect 2982 3809 3067 3817
rect 2982 3789 3039 3809
rect 3059 3789 3067 3809
rect 2915 3783 2952 3784
rect 2982 3783 3067 3789
rect 3133 3813 3171 3821
rect 3133 3793 3142 3813
rect 3162 3793 3171 3813
rect 3404 3802 3441 3803
rect 3707 3802 3744 3872
rect 3779 3901 3810 3952
rect 4106 3947 4151 3953
rect 4106 3929 4124 3947
rect 4142 3929 4151 3947
rect 4106 3919 4151 3929
rect 3829 3901 3866 3902
rect 3779 3892 3866 3901
rect 3779 3872 3837 3892
rect 3857 3872 3866 3892
rect 3779 3862 3866 3872
rect 3925 3892 3962 3902
rect 3925 3872 3933 3892
rect 3953 3872 3962 3892
rect 4106 3877 4149 3919
rect 4012 3875 4149 3877
rect 3779 3861 3810 3862
rect 3925 3802 3962 3872
rect 3403 3801 3744 3802
rect 3133 3784 3171 3793
rect 3328 3796 3744 3801
rect 3133 3783 3170 3784
rect 2594 3755 2684 3761
rect 2594 3735 2610 3755
rect 2630 3753 2684 3755
rect 2630 3735 2655 3753
rect 2594 3733 2655 3735
rect 2675 3733 2684 3753
rect 2594 3727 2684 3733
rect 2607 3673 2644 3674
rect 2703 3673 2740 3674
rect 2759 3673 2795 3783
rect 2982 3762 3013 3783
rect 3328 3776 3331 3796
rect 3351 3776 3744 3796
rect 3928 3786 3962 3802
rect 4006 3854 4149 3875
rect 3704 3767 3744 3776
rect 4006 3767 4033 3854
rect 4106 3828 4149 3854
rect 4106 3810 4119 3828
rect 4137 3810 4149 3828
rect 4106 3799 4149 3810
rect 2978 3761 3013 3762
rect 2856 3751 3013 3761
rect 2856 3731 2873 3751
rect 2893 3731 3013 3751
rect 2856 3724 3013 3731
rect 3080 3754 3226 3762
rect 3080 3734 3091 3754
rect 3111 3734 3150 3754
rect 3170 3734 3226 3754
rect 3704 3750 4033 3767
rect 3704 3749 3744 3750
rect 3080 3727 3226 3734
rect 4101 3738 4141 3741
rect 4101 3732 4144 3738
rect 3726 3729 4144 3732
rect 3080 3726 3121 3727
rect 2814 3673 2851 3674
rect 2507 3664 2645 3673
rect 2507 3644 2616 3664
rect 2636 3644 2645 3664
rect 2507 3637 2645 3644
rect 2703 3664 2851 3673
rect 2703 3644 2712 3664
rect 2732 3644 2822 3664
rect 2842 3644 2851 3664
rect 2507 3635 2603 3637
rect 2703 3634 2851 3644
rect 2910 3664 2947 3674
rect 2910 3644 2918 3664
rect 2938 3644 2947 3664
rect 2759 3633 2795 3634
rect 2607 3574 2644 3575
rect 2910 3574 2947 3644
rect 2982 3673 3013 3724
rect 3726 3711 4117 3729
rect 4135 3711 4144 3729
rect 3726 3709 4144 3711
rect 3726 3701 3753 3709
rect 3994 3706 4144 3709
rect 3306 3695 3474 3696
rect 3725 3695 3753 3701
rect 3306 3679 3753 3695
rect 4101 3701 4144 3706
rect 3032 3673 3069 3674
rect 2982 3664 3069 3673
rect 2982 3644 3040 3664
rect 3060 3644 3069 3664
rect 2982 3634 3069 3644
rect 3128 3664 3165 3674
rect 3128 3644 3136 3664
rect 3156 3644 3165 3664
rect 2982 3633 3013 3634
rect 2606 3573 2947 3574
rect 3128 3573 3165 3644
rect 2531 3568 2947 3573
rect 2531 3548 2534 3568
rect 2554 3548 2947 3568
rect 2978 3549 3165 3573
rect 3306 3669 3750 3679
rect 3306 3667 3474 3669
rect 2340 3474 2384 3475
rect 2340 3468 2385 3474
rect 2340 3450 2352 3468
rect 2374 3450 2385 3468
rect 2406 3469 2448 3514
rect 3306 3489 3333 3667
rect 3373 3629 3437 3641
rect 3713 3637 3750 3669
rect 3776 3668 3967 3690
rect 3931 3666 3967 3668
rect 3931 3637 3968 3666
rect 4101 3645 4141 3701
rect 3373 3628 3408 3629
rect 3350 3623 3408 3628
rect 3350 3603 3353 3623
rect 3373 3609 3408 3623
rect 3428 3609 3437 3629
rect 3373 3601 3437 3609
rect 3399 3600 3437 3601
rect 3400 3599 3437 3600
rect 3503 3633 3539 3634
rect 3611 3633 3647 3634
rect 3503 3625 3647 3633
rect 3503 3605 3511 3625
rect 3531 3605 3566 3625
rect 3586 3605 3619 3625
rect 3639 3605 3647 3625
rect 3503 3599 3647 3605
rect 3713 3629 3751 3637
rect 3829 3633 3865 3634
rect 3713 3609 3722 3629
rect 3742 3609 3751 3629
rect 3713 3600 3751 3609
rect 3780 3625 3865 3633
rect 3780 3605 3837 3625
rect 3857 3605 3865 3625
rect 3713 3599 3750 3600
rect 3780 3599 3865 3605
rect 3931 3629 3969 3637
rect 3931 3609 3940 3629
rect 3960 3609 3969 3629
rect 4101 3627 4113 3645
rect 4131 3627 4141 3645
rect 4101 3617 4141 3627
rect 3931 3600 3969 3609
rect 3931 3599 3968 3600
rect 3392 3571 3482 3577
rect 3392 3551 3408 3571
rect 3428 3569 3482 3571
rect 3428 3551 3453 3569
rect 3392 3549 3453 3551
rect 3473 3549 3482 3569
rect 3392 3543 3482 3549
rect 3405 3489 3442 3490
rect 3501 3489 3538 3490
rect 3557 3489 3593 3599
rect 3780 3578 3811 3599
rect 3776 3577 3811 3578
rect 3654 3567 3811 3577
rect 3654 3547 3671 3567
rect 3691 3547 3811 3567
rect 3654 3540 3811 3547
rect 3878 3570 4027 3578
rect 3878 3550 3889 3570
rect 3909 3550 3948 3570
rect 3968 3550 4027 3570
rect 3878 3543 4027 3550
rect 4093 3546 4145 3564
rect 3878 3542 3919 3543
rect 3612 3489 3649 3490
rect 3305 3480 3443 3489
rect 2777 3469 2810 3471
rect 2406 3457 2853 3469
rect 2340 3420 2385 3450
rect 2357 2474 2385 3420
rect 2409 3443 2853 3457
rect 2409 3441 2577 3443
rect 2409 3263 2436 3441
rect 2476 3403 2540 3415
rect 2816 3411 2853 3443
rect 2879 3442 3070 3464
rect 3305 3460 3414 3480
rect 3434 3460 3443 3480
rect 3305 3453 3443 3460
rect 3501 3480 3649 3489
rect 3501 3460 3510 3480
rect 3530 3460 3620 3480
rect 3640 3460 3649 3480
rect 3305 3451 3401 3453
rect 3501 3450 3649 3460
rect 3708 3480 3745 3490
rect 3708 3460 3716 3480
rect 3736 3460 3745 3480
rect 3557 3449 3593 3450
rect 3034 3440 3070 3442
rect 3034 3411 3071 3440
rect 2476 3402 2511 3403
rect 2453 3397 2511 3402
rect 2453 3377 2456 3397
rect 2476 3383 2511 3397
rect 2531 3383 2540 3403
rect 2476 3375 2540 3383
rect 2502 3374 2540 3375
rect 2503 3373 2540 3374
rect 2606 3407 2642 3408
rect 2714 3407 2750 3408
rect 2606 3401 2750 3407
rect 2606 3399 2667 3401
rect 2606 3379 2614 3399
rect 2634 3384 2667 3399
rect 2686 3399 2750 3401
rect 2686 3384 2722 3399
rect 2634 3379 2722 3384
rect 2742 3379 2750 3399
rect 2606 3373 2750 3379
rect 2816 3403 2854 3411
rect 2932 3407 2968 3408
rect 2816 3383 2825 3403
rect 2845 3383 2854 3403
rect 2816 3374 2854 3383
rect 2883 3399 2968 3407
rect 2883 3379 2940 3399
rect 2960 3379 2968 3399
rect 2816 3373 2853 3374
rect 2883 3373 2968 3379
rect 3034 3403 3072 3411
rect 3034 3383 3043 3403
rect 3063 3383 3072 3403
rect 3708 3393 3745 3460
rect 3780 3489 3811 3540
rect 4093 3528 4111 3546
rect 4129 3528 4145 3546
rect 3830 3489 3867 3490
rect 3780 3480 3867 3489
rect 3780 3460 3838 3480
rect 3858 3460 3867 3480
rect 3780 3450 3867 3460
rect 3926 3480 3963 3490
rect 3926 3460 3934 3480
rect 3954 3460 3963 3480
rect 3780 3449 3811 3450
rect 3405 3390 3442 3391
rect 3708 3390 3747 3393
rect 3404 3389 3747 3390
rect 3926 3389 3963 3460
rect 3034 3374 3072 3383
rect 3329 3384 3747 3389
rect 3034 3373 3071 3374
rect 2495 3345 2585 3351
rect 2495 3325 2511 3345
rect 2531 3343 2585 3345
rect 2531 3325 2556 3343
rect 2495 3323 2556 3325
rect 2576 3323 2585 3343
rect 2495 3317 2585 3323
rect 2508 3263 2545 3264
rect 2604 3263 2641 3264
rect 2660 3263 2696 3373
rect 2883 3352 2914 3373
rect 3329 3364 3332 3384
rect 3352 3364 3747 3384
rect 3776 3365 3963 3389
rect 2879 3351 2914 3352
rect 2757 3341 2914 3351
rect 2757 3321 2774 3341
rect 2794 3321 2914 3341
rect 2757 3314 2914 3321
rect 2981 3344 3130 3352
rect 2981 3324 2992 3344
rect 3012 3324 3051 3344
rect 3071 3324 3130 3344
rect 2981 3317 3130 3324
rect 3708 3339 3747 3364
rect 4093 3339 4145 3528
rect 3708 3321 4147 3339
rect 2981 3316 3022 3317
rect 2715 3263 2752 3264
rect 2408 3254 2546 3263
rect 2408 3234 2517 3254
rect 2537 3234 2546 3254
rect 2408 3227 2546 3234
rect 2604 3254 2752 3263
rect 2604 3234 2613 3254
rect 2633 3234 2723 3254
rect 2743 3234 2752 3254
rect 2408 3225 2504 3227
rect 2604 3224 2752 3234
rect 2811 3254 2848 3264
rect 2811 3234 2819 3254
rect 2839 3234 2848 3254
rect 2660 3223 2696 3224
rect 2508 3164 2545 3165
rect 2811 3164 2848 3234
rect 2883 3263 2914 3314
rect 3708 3303 4108 3321
rect 4126 3303 4147 3321
rect 3708 3297 4147 3303
rect 3714 3293 4147 3297
rect 4093 3291 4145 3293
rect 2933 3263 2970 3264
rect 2883 3254 2970 3263
rect 2883 3234 2941 3254
rect 2961 3234 2970 3254
rect 2883 3224 2970 3234
rect 3029 3254 3066 3264
rect 3029 3234 3037 3254
rect 3057 3234 3066 3254
rect 2883 3223 2914 3224
rect 2507 3163 2848 3164
rect 3029 3163 3066 3234
rect 4096 3226 4133 3231
rect 4087 3222 4134 3226
rect 4087 3204 4106 3222
rect 4124 3204 4134 3222
rect 2432 3158 2848 3163
rect 2432 3138 2435 3158
rect 2455 3138 2848 3158
rect 2879 3139 3066 3163
rect 3691 3161 3731 3166
rect 4087 3161 4134 3204
rect 3691 3122 4134 3161
rect 2785 3107 2825 3115
rect 2785 3085 2793 3107
rect 2817 3085 2825 3107
rect 2491 2861 2659 2862
rect 2785 2861 2825 3085
rect 3288 3089 3456 3090
rect 3691 3089 3731 3122
rect 4087 3089 4134 3122
rect 3288 3088 3732 3089
rect 3288 3063 3733 3088
rect 3288 3061 3456 3063
rect 3652 3062 3733 3063
rect 3902 3062 3951 3088
rect 4087 3062 4136 3089
rect 3288 2883 3315 3061
rect 3355 3023 3419 3035
rect 3695 3031 3732 3062
rect 3913 3031 3950 3062
rect 4095 3037 4136 3062
rect 3355 3022 3390 3023
rect 3332 3017 3390 3022
rect 3332 2997 3335 3017
rect 3355 3003 3390 3017
rect 3410 3003 3419 3023
rect 3355 2995 3419 3003
rect 3381 2994 3419 2995
rect 3382 2993 3419 2994
rect 3485 3027 3521 3028
rect 3593 3027 3629 3028
rect 3485 3019 3629 3027
rect 3485 2999 3493 3019
rect 3513 3015 3601 3019
rect 3513 2999 3557 3015
rect 3485 2995 3557 2999
rect 3577 2999 3601 3015
rect 3621 2999 3629 3019
rect 3577 2995 3629 2999
rect 3485 2993 3629 2995
rect 3695 3023 3733 3031
rect 3811 3027 3847 3028
rect 3695 3003 3704 3023
rect 3724 3003 3733 3023
rect 3695 2994 3733 3003
rect 3762 3019 3847 3027
rect 3762 2999 3819 3019
rect 3839 2999 3847 3019
rect 3695 2993 3732 2994
rect 3762 2993 3847 2999
rect 3913 3023 3951 3031
rect 3913 3003 3922 3023
rect 3942 3003 3951 3023
rect 3913 2994 3951 3003
rect 4095 3028 4137 3037
rect 4095 3010 4109 3028
rect 4127 3010 4137 3028
rect 4095 3002 4137 3010
rect 4100 3000 4137 3002
rect 3913 2993 3950 2994
rect 3374 2965 3464 2971
rect 3374 2945 3390 2965
rect 3410 2963 3464 2965
rect 3410 2945 3435 2963
rect 3374 2943 3435 2945
rect 3455 2943 3464 2963
rect 3374 2937 3464 2943
rect 3387 2883 3424 2884
rect 3483 2883 3520 2884
rect 3539 2883 3575 2993
rect 3762 2972 3793 2993
rect 3758 2971 3793 2972
rect 3636 2961 3793 2971
rect 3636 2941 3653 2961
rect 3673 2941 3793 2961
rect 3636 2934 3793 2941
rect 3860 2964 4009 2972
rect 3860 2944 3871 2964
rect 3891 2944 3930 2964
rect 3950 2944 4009 2964
rect 3860 2937 4009 2944
rect 3860 2936 3901 2937
rect 4097 2935 4134 2938
rect 3594 2883 3631 2884
rect 3287 2874 3425 2883
rect 2491 2835 2935 2861
rect 2491 2833 2659 2835
rect 2491 2655 2518 2833
rect 2558 2795 2622 2807
rect 2898 2803 2935 2835
rect 2961 2834 3152 2856
rect 3287 2854 3396 2874
rect 3416 2854 3425 2874
rect 3287 2847 3425 2854
rect 3483 2874 3631 2883
rect 3483 2854 3492 2874
rect 3512 2854 3602 2874
rect 3622 2854 3631 2874
rect 3287 2845 3383 2847
rect 3483 2844 3631 2854
rect 3690 2874 3727 2884
rect 3690 2854 3698 2874
rect 3718 2854 3727 2874
rect 3539 2843 3575 2844
rect 3116 2832 3152 2834
rect 3116 2803 3153 2832
rect 2558 2794 2593 2795
rect 2535 2789 2593 2794
rect 2535 2769 2538 2789
rect 2558 2775 2593 2789
rect 2613 2775 2622 2795
rect 2558 2767 2622 2775
rect 2584 2766 2622 2767
rect 2585 2765 2622 2766
rect 2688 2799 2724 2800
rect 2796 2799 2832 2800
rect 2688 2791 2832 2799
rect 2688 2771 2696 2791
rect 2716 2790 2804 2791
rect 2716 2771 2751 2790
rect 2772 2771 2804 2790
rect 2824 2771 2832 2791
rect 2688 2765 2832 2771
rect 2898 2795 2936 2803
rect 3014 2799 3050 2800
rect 2898 2775 2907 2795
rect 2927 2775 2936 2795
rect 2898 2766 2936 2775
rect 2965 2791 3050 2799
rect 2965 2771 3022 2791
rect 3042 2771 3050 2791
rect 2898 2765 2935 2766
rect 2965 2765 3050 2771
rect 3116 2795 3154 2803
rect 3116 2775 3125 2795
rect 3145 2775 3154 2795
rect 3387 2784 3424 2785
rect 3690 2784 3727 2854
rect 3762 2883 3793 2934
rect 4089 2929 4134 2935
rect 4089 2911 4107 2929
rect 4125 2911 4134 2929
rect 4089 2901 4134 2911
rect 3812 2883 3849 2884
rect 3762 2874 3849 2883
rect 3762 2854 3820 2874
rect 3840 2854 3849 2874
rect 3762 2844 3849 2854
rect 3908 2874 3945 2884
rect 3908 2854 3916 2874
rect 3936 2854 3945 2874
rect 4089 2859 4132 2901
rect 3995 2857 4132 2859
rect 3762 2843 3793 2844
rect 3908 2784 3945 2854
rect 3386 2783 3727 2784
rect 3116 2766 3154 2775
rect 3311 2778 3727 2783
rect 3116 2765 3153 2766
rect 2577 2737 2667 2743
rect 2577 2717 2593 2737
rect 2613 2735 2667 2737
rect 2613 2717 2638 2735
rect 2577 2715 2638 2717
rect 2658 2715 2667 2735
rect 2577 2709 2667 2715
rect 2590 2655 2627 2656
rect 2686 2655 2723 2656
rect 2742 2655 2778 2765
rect 2965 2744 2996 2765
rect 3311 2758 3314 2778
rect 3334 2758 3727 2778
rect 3911 2768 3945 2784
rect 3989 2836 4132 2857
rect 3687 2749 3727 2758
rect 3989 2749 4016 2836
rect 4089 2810 4132 2836
rect 4089 2792 4102 2810
rect 4120 2792 4132 2810
rect 4089 2781 4132 2792
rect 2961 2743 2996 2744
rect 2839 2733 2996 2743
rect 2839 2713 2856 2733
rect 2876 2713 2996 2733
rect 2839 2706 2996 2713
rect 3063 2736 3212 2744
rect 3063 2716 3074 2736
rect 3094 2716 3133 2736
rect 3153 2716 3212 2736
rect 3687 2732 4016 2749
rect 3687 2731 3727 2732
rect 3063 2709 3212 2716
rect 4084 2720 4124 2723
rect 4084 2714 4127 2720
rect 3709 2711 4127 2714
rect 3063 2708 3104 2709
rect 2797 2655 2834 2656
rect 2490 2646 2628 2655
rect 2490 2626 2599 2646
rect 2619 2626 2628 2646
rect 2490 2619 2628 2626
rect 2686 2646 2834 2655
rect 2686 2626 2695 2646
rect 2715 2626 2805 2646
rect 2825 2626 2834 2646
rect 2490 2617 2586 2619
rect 2686 2616 2834 2626
rect 2893 2646 2930 2656
rect 2893 2626 2901 2646
rect 2921 2626 2930 2646
rect 2742 2615 2778 2616
rect 2590 2556 2627 2557
rect 2893 2556 2930 2626
rect 2965 2655 2996 2706
rect 3709 2693 4100 2711
rect 4118 2693 4127 2711
rect 3709 2691 4127 2693
rect 3709 2683 3736 2691
rect 3977 2688 4127 2691
rect 3289 2677 3457 2678
rect 3708 2677 3736 2683
rect 3289 2661 3736 2677
rect 4084 2683 4127 2688
rect 3015 2655 3052 2656
rect 2965 2646 3052 2655
rect 2965 2626 3023 2646
rect 3043 2626 3052 2646
rect 2965 2616 3052 2626
rect 3111 2646 3148 2656
rect 3111 2626 3119 2646
rect 3139 2626 3148 2646
rect 2965 2615 2996 2616
rect 2589 2555 2930 2556
rect 3111 2555 3148 2626
rect 2514 2550 2930 2555
rect 2514 2530 2517 2550
rect 2537 2530 2930 2550
rect 2961 2531 3148 2555
rect 3289 2651 3733 2661
rect 3289 2649 3457 2651
rect 2356 2456 2385 2474
rect 3289 2471 3316 2649
rect 3356 2611 3420 2623
rect 3696 2619 3733 2651
rect 3759 2650 3950 2672
rect 3914 2648 3950 2650
rect 3914 2619 3951 2648
rect 4084 2627 4124 2683
rect 3356 2610 3391 2611
rect 3333 2605 3391 2610
rect 3333 2585 3336 2605
rect 3356 2591 3391 2605
rect 3411 2591 3420 2611
rect 3356 2583 3420 2591
rect 3382 2582 3420 2583
rect 3383 2581 3420 2582
rect 3486 2615 3522 2616
rect 3594 2615 3630 2616
rect 3486 2607 3630 2615
rect 3486 2587 3494 2607
rect 3514 2587 3549 2607
rect 3569 2587 3602 2607
rect 3622 2587 3630 2607
rect 3486 2581 3630 2587
rect 3696 2611 3734 2619
rect 3812 2615 3848 2616
rect 3696 2591 3705 2611
rect 3725 2591 3734 2611
rect 3696 2582 3734 2591
rect 3763 2607 3848 2615
rect 3763 2587 3820 2607
rect 3840 2587 3848 2607
rect 3696 2581 3733 2582
rect 3763 2581 3848 2587
rect 3914 2611 3952 2619
rect 3914 2591 3923 2611
rect 3943 2591 3952 2611
rect 4084 2609 4096 2627
rect 4114 2609 4124 2627
rect 4084 2599 4124 2609
rect 3914 2582 3952 2591
rect 3914 2581 3951 2582
rect 3375 2553 3465 2559
rect 3375 2533 3391 2553
rect 3411 2551 3465 2553
rect 3411 2533 3436 2551
rect 3375 2531 3436 2533
rect 3456 2531 3465 2551
rect 3375 2525 3465 2531
rect 3388 2471 3425 2472
rect 3484 2471 3521 2472
rect 3540 2471 3576 2581
rect 3763 2560 3794 2581
rect 3759 2559 3794 2560
rect 3637 2549 3794 2559
rect 3637 2529 3654 2549
rect 3674 2529 3794 2549
rect 3637 2522 3794 2529
rect 3861 2552 4010 2560
rect 3861 2532 3872 2552
rect 3892 2532 3931 2552
rect 3951 2532 4010 2552
rect 3861 2525 4010 2532
rect 4076 2528 4128 2546
rect 3861 2524 3902 2525
rect 3595 2471 3632 2472
rect 2326 2454 2385 2456
rect 3288 2462 3426 2471
rect 2326 2453 2494 2454
rect 2620 2453 2660 2455
rect 2326 2427 2770 2453
rect 2326 2425 2494 2427
rect 2326 2423 2407 2425
rect 2326 2247 2353 2423
rect 2393 2387 2457 2399
rect 2733 2395 2770 2427
rect 2796 2426 2987 2448
rect 3288 2442 3397 2462
rect 3417 2442 3426 2462
rect 3288 2435 3426 2442
rect 3484 2462 3632 2471
rect 3484 2442 3493 2462
rect 3513 2442 3603 2462
rect 3623 2442 3632 2462
rect 3288 2433 3384 2435
rect 3484 2432 3632 2442
rect 3691 2462 3728 2472
rect 3691 2442 3699 2462
rect 3719 2442 3728 2462
rect 3540 2431 3576 2432
rect 2951 2424 2987 2426
rect 2951 2395 2988 2424
rect 2393 2386 2428 2387
rect 2370 2381 2428 2386
rect 2370 2361 2373 2381
rect 2393 2367 2428 2381
rect 2448 2367 2457 2387
rect 2393 2359 2457 2367
rect 2419 2358 2457 2359
rect 2420 2357 2457 2358
rect 2523 2391 2559 2392
rect 2631 2391 2667 2392
rect 2523 2383 2667 2391
rect 2523 2363 2531 2383
rect 2551 2382 2639 2383
rect 2551 2364 2586 2382
rect 2604 2364 2639 2382
rect 2551 2363 2639 2364
rect 2659 2363 2667 2383
rect 2523 2357 2667 2363
rect 2733 2387 2771 2395
rect 2849 2391 2885 2392
rect 2733 2367 2742 2387
rect 2762 2367 2771 2387
rect 2733 2358 2771 2367
rect 2800 2383 2885 2391
rect 2800 2363 2857 2383
rect 2877 2363 2885 2383
rect 2733 2357 2770 2358
rect 2800 2357 2885 2363
rect 2951 2387 2989 2395
rect 2951 2367 2960 2387
rect 2980 2367 2989 2387
rect 3691 2375 3728 2442
rect 3763 2471 3794 2522
rect 4076 2510 4094 2528
rect 4112 2510 4128 2528
rect 3813 2471 3850 2472
rect 3763 2462 3850 2471
rect 3763 2442 3821 2462
rect 3841 2442 3850 2462
rect 3763 2432 3850 2442
rect 3909 2462 3946 2472
rect 3909 2442 3917 2462
rect 3937 2442 3946 2462
rect 3763 2431 3794 2432
rect 3388 2372 3425 2373
rect 3691 2372 3730 2375
rect 3387 2371 3730 2372
rect 3909 2371 3946 2442
rect 2951 2358 2989 2367
rect 3312 2366 3730 2371
rect 2951 2357 2988 2358
rect 2412 2329 2502 2335
rect 2412 2309 2428 2329
rect 2448 2327 2502 2329
rect 2448 2309 2473 2327
rect 2412 2307 2473 2309
rect 2493 2307 2502 2327
rect 2412 2301 2502 2307
rect 2425 2247 2462 2248
rect 2521 2247 2558 2248
rect 2577 2247 2613 2357
rect 2800 2336 2831 2357
rect 3312 2346 3315 2366
rect 3335 2346 3730 2366
rect 3759 2347 3946 2371
rect 2796 2335 2831 2336
rect 2674 2325 2831 2335
rect 2674 2305 2691 2325
rect 2711 2305 2831 2325
rect 2674 2298 2831 2305
rect 2898 2328 3047 2336
rect 2898 2308 2909 2328
rect 2929 2308 2968 2328
rect 2988 2308 3047 2328
rect 2898 2301 3047 2308
rect 3691 2321 3730 2346
rect 4076 2321 4128 2510
rect 3691 2303 4130 2321
rect 2898 2300 2939 2301
rect 2632 2247 2669 2248
rect 2325 2238 2463 2247
rect 2325 2218 2434 2238
rect 2454 2218 2463 2238
rect 2325 2211 2463 2218
rect 2521 2238 2669 2247
rect 2521 2218 2530 2238
rect 2550 2218 2640 2238
rect 2660 2218 2669 2238
rect 2325 2209 2421 2211
rect 2521 2208 2669 2218
rect 2728 2238 2765 2248
rect 2728 2218 2736 2238
rect 2756 2218 2765 2238
rect 2577 2207 2613 2208
rect 2425 2148 2462 2149
rect 2728 2148 2765 2218
rect 2800 2247 2831 2298
rect 3691 2285 4091 2303
rect 4109 2285 4130 2303
rect 3691 2279 4130 2285
rect 3697 2275 4130 2279
rect 4076 2273 4128 2275
rect 2850 2247 2887 2248
rect 2800 2238 2887 2247
rect 2800 2218 2858 2238
rect 2878 2218 2887 2238
rect 2800 2208 2887 2218
rect 2946 2238 2983 2248
rect 2946 2218 2954 2238
rect 2974 2218 2983 2238
rect 2800 2207 2831 2208
rect 2424 2147 2765 2148
rect 2946 2147 2983 2218
rect 4079 2208 4116 2213
rect 2349 2142 2765 2147
rect 2349 2122 2352 2142
rect 2372 2122 2765 2142
rect 2796 2123 2983 2147
rect 4070 2204 4117 2208
rect 4070 2186 4089 2204
rect 4107 2186 4117 2204
rect 4070 2138 4117 2186
rect 3694 2135 4117 2138
rect 2569 2121 2634 2122
rect 3672 2105 4117 2135
rect 2765 2089 2805 2097
rect 2765 2067 2773 2089
rect 2797 2067 2805 2089
rect 2370 1838 2407 1844
rect 2370 1819 2378 1838
rect 2399 1819 2407 1838
rect 2370 1811 2407 1819
rect 2070 1690 2077 1712
rect 2101 1690 2109 1712
rect 2070 1684 2109 1690
rect 1600 1679 1640 1681
rect 1766 1680 1934 1681
rect 1868 1679 1905 1680
rect 834 1663 972 1672
rect 628 1662 665 1663
rect 358 1609 399 1610
rect 132 1588 184 1606
rect 250 1602 399 1609
rect 250 1582 309 1602
rect 329 1582 368 1602
rect 388 1582 399 1602
rect 250 1574 399 1582
rect 466 1605 623 1612
rect 466 1585 586 1605
rect 606 1585 623 1605
rect 466 1575 623 1585
rect 466 1574 501 1575
rect 466 1553 497 1574
rect 684 1553 720 1663
rect 739 1662 776 1663
rect 835 1662 872 1663
rect 795 1603 885 1609
rect 795 1583 804 1603
rect 824 1601 885 1603
rect 824 1583 849 1601
rect 795 1581 849 1583
rect 869 1581 885 1601
rect 795 1575 885 1581
rect 309 1552 346 1553
rect 308 1543 346 1552
rect 136 1525 176 1535
rect 136 1507 146 1525
rect 164 1507 176 1525
rect 308 1523 317 1543
rect 337 1523 346 1543
rect 308 1515 346 1523
rect 412 1547 497 1553
rect 527 1552 564 1553
rect 412 1527 420 1547
rect 440 1527 497 1547
rect 412 1519 497 1527
rect 526 1543 564 1552
rect 526 1523 535 1543
rect 555 1523 564 1543
rect 412 1518 448 1519
rect 526 1515 564 1523
rect 630 1547 774 1553
rect 630 1527 638 1547
rect 658 1527 691 1547
rect 711 1527 746 1547
rect 766 1527 774 1547
rect 630 1519 774 1527
rect 630 1518 666 1519
rect 738 1518 774 1519
rect 840 1552 877 1553
rect 840 1551 878 1552
rect 840 1543 904 1551
rect 840 1523 849 1543
rect 869 1529 904 1543
rect 924 1529 927 1549
rect 869 1524 927 1529
rect 869 1523 904 1524
rect 136 1451 176 1507
rect 309 1486 346 1515
rect 310 1484 346 1486
rect 310 1462 501 1484
rect 527 1483 564 1515
rect 840 1511 904 1523
rect 944 1485 971 1663
rect 803 1483 971 1485
rect 527 1473 971 1483
rect 1112 1579 1299 1603
rect 1330 1584 1723 1604
rect 1743 1584 1746 1604
rect 1330 1579 1746 1584
rect 1112 1508 1149 1579
rect 1330 1578 1671 1579
rect 1264 1518 1295 1519
rect 1112 1488 1121 1508
rect 1141 1488 1149 1508
rect 1112 1478 1149 1488
rect 1208 1508 1295 1518
rect 1208 1488 1217 1508
rect 1237 1488 1295 1508
rect 1208 1479 1295 1488
rect 1208 1478 1245 1479
rect 133 1446 176 1451
rect 524 1457 971 1473
rect 524 1451 552 1457
rect 803 1456 971 1457
rect 133 1443 283 1446
rect 524 1443 551 1451
rect 133 1441 551 1443
rect 133 1423 142 1441
rect 160 1423 551 1441
rect 1264 1428 1295 1479
rect 1330 1508 1367 1578
rect 1633 1577 1670 1578
rect 1871 1520 1904 1679
rect 1482 1518 1518 1519
rect 1330 1488 1339 1508
rect 1359 1488 1367 1508
rect 1330 1478 1367 1488
rect 1426 1508 1574 1518
rect 1674 1515 1770 1517
rect 1426 1488 1435 1508
rect 1455 1488 1545 1508
rect 1565 1488 1574 1508
rect 1426 1479 1574 1488
rect 1632 1508 1770 1515
rect 1632 1488 1641 1508
rect 1661 1488 1770 1508
rect 1871 1516 1907 1520
rect 1871 1498 1880 1516
rect 1902 1498 1907 1516
rect 1871 1492 1907 1498
rect 1632 1479 1770 1488
rect 1426 1478 1463 1479
rect 1156 1425 1197 1426
rect 133 1420 551 1423
rect 133 1414 176 1420
rect 136 1411 176 1414
rect 1048 1418 1197 1425
rect 533 1402 573 1403
rect 244 1385 573 1402
rect 1048 1398 1107 1418
rect 1127 1398 1166 1418
rect 1186 1398 1197 1418
rect 1048 1390 1197 1398
rect 1264 1421 1421 1428
rect 1264 1401 1384 1421
rect 1404 1401 1421 1421
rect 1264 1391 1421 1401
rect 1264 1390 1299 1391
rect 128 1342 171 1353
rect 128 1324 140 1342
rect 158 1324 171 1342
rect 128 1298 171 1324
rect 244 1298 271 1385
rect 533 1376 573 1385
rect 128 1277 271 1298
rect 315 1350 349 1366
rect 533 1356 926 1376
rect 946 1356 949 1376
rect 1264 1369 1295 1390
rect 1482 1369 1518 1479
rect 1537 1478 1574 1479
rect 1633 1478 1670 1479
rect 1593 1419 1683 1425
rect 1593 1399 1602 1419
rect 1622 1417 1683 1419
rect 1622 1399 1647 1417
rect 1593 1397 1647 1399
rect 1667 1397 1683 1417
rect 1593 1391 1683 1397
rect 1107 1368 1144 1369
rect 533 1351 949 1356
rect 1106 1359 1144 1368
rect 533 1350 874 1351
rect 315 1280 352 1350
rect 467 1290 498 1291
rect 128 1275 265 1277
rect 128 1233 171 1275
rect 315 1260 324 1280
rect 344 1260 352 1280
rect 315 1250 352 1260
rect 411 1280 498 1290
rect 411 1260 420 1280
rect 440 1260 498 1280
rect 411 1251 498 1260
rect 411 1250 448 1251
rect 126 1223 171 1233
rect 126 1205 135 1223
rect 153 1205 171 1223
rect 126 1199 171 1205
rect 467 1200 498 1251
rect 533 1280 570 1350
rect 836 1349 873 1350
rect 1106 1339 1115 1359
rect 1135 1339 1144 1359
rect 1106 1331 1144 1339
rect 1210 1363 1295 1369
rect 1325 1368 1362 1369
rect 1210 1343 1218 1363
rect 1238 1343 1295 1363
rect 1210 1335 1295 1343
rect 1324 1359 1362 1368
rect 1324 1339 1333 1359
rect 1353 1339 1362 1359
rect 1210 1334 1246 1335
rect 1324 1331 1362 1339
rect 1428 1363 1572 1369
rect 1428 1343 1436 1363
rect 1456 1344 1488 1363
rect 1509 1344 1544 1363
rect 1456 1343 1544 1344
rect 1564 1343 1572 1363
rect 1428 1335 1572 1343
rect 1428 1334 1464 1335
rect 1536 1334 1572 1335
rect 1638 1368 1675 1369
rect 1638 1367 1676 1368
rect 1638 1359 1702 1367
rect 1638 1339 1647 1359
rect 1667 1345 1702 1359
rect 1722 1345 1725 1365
rect 1667 1340 1725 1345
rect 1667 1339 1702 1340
rect 1107 1302 1144 1331
rect 1108 1300 1144 1302
rect 685 1290 721 1291
rect 533 1260 542 1280
rect 562 1260 570 1280
rect 533 1250 570 1260
rect 629 1280 777 1290
rect 877 1287 973 1289
rect 629 1260 638 1280
rect 658 1260 748 1280
rect 768 1260 777 1280
rect 629 1251 777 1260
rect 835 1280 973 1287
rect 835 1260 844 1280
rect 864 1260 973 1280
rect 1108 1278 1299 1300
rect 1325 1299 1362 1331
rect 1638 1327 1702 1339
rect 1742 1301 1769 1479
rect 2374 1478 2407 1811
rect 2471 1843 2639 1844
rect 2765 1843 2805 2067
rect 3268 2071 3436 2072
rect 3672 2071 3713 2105
rect 4070 2084 4117 2105
rect 3268 2061 3713 2071
rect 3785 2069 3928 2070
rect 3268 2045 3712 2061
rect 3268 2043 3436 2045
rect 3632 2044 3712 2045
rect 3785 2044 3930 2069
rect 4072 2044 4117 2084
rect 3268 1865 3295 2043
rect 3335 2005 3399 2017
rect 3675 2013 3712 2044
rect 3893 2013 3930 2044
rect 4075 2037 4117 2044
rect 3335 2004 3370 2005
rect 3312 1999 3370 2004
rect 3312 1979 3315 1999
rect 3335 1985 3370 1999
rect 3390 1985 3399 2005
rect 3335 1977 3399 1985
rect 3361 1976 3399 1977
rect 3362 1975 3399 1976
rect 3465 2009 3501 2010
rect 3573 2009 3609 2010
rect 3465 2001 3609 2009
rect 3465 1981 3473 2001
rect 3493 1997 3581 2001
rect 3493 1981 3537 1997
rect 3465 1977 3537 1981
rect 3557 1981 3581 1997
rect 3601 1981 3609 2001
rect 3557 1977 3609 1981
rect 3465 1975 3609 1977
rect 3675 2005 3713 2013
rect 3791 2009 3827 2010
rect 3675 1985 3684 2005
rect 3704 1985 3713 2005
rect 3675 1976 3713 1985
rect 3742 2001 3827 2009
rect 3742 1981 3799 2001
rect 3819 1981 3827 2001
rect 3675 1975 3712 1976
rect 3742 1975 3827 1981
rect 3893 2005 3931 2013
rect 3893 1985 3902 2005
rect 3922 1985 3931 2005
rect 3893 1976 3931 1985
rect 4075 2010 4118 2037
rect 4075 1992 4089 2010
rect 4107 1992 4118 2010
rect 4075 1984 4118 1992
rect 4080 1982 4118 1984
rect 3893 1975 3930 1976
rect 3354 1947 3444 1953
rect 3354 1927 3370 1947
rect 3390 1945 3444 1947
rect 3390 1927 3415 1945
rect 3354 1925 3415 1927
rect 3435 1925 3444 1945
rect 3354 1919 3444 1925
rect 3367 1865 3404 1866
rect 3463 1865 3500 1866
rect 3519 1865 3555 1975
rect 3742 1954 3773 1975
rect 3738 1953 3773 1954
rect 3616 1943 3773 1953
rect 3616 1923 3633 1943
rect 3653 1923 3773 1943
rect 3616 1916 3773 1923
rect 3840 1946 3989 1954
rect 3840 1926 3851 1946
rect 3871 1926 3910 1946
rect 3930 1926 3989 1946
rect 3840 1919 3989 1926
rect 3840 1918 3881 1919
rect 4077 1917 4114 1920
rect 3574 1865 3611 1866
rect 3267 1856 3405 1865
rect 2471 1817 2915 1843
rect 2471 1815 2639 1817
rect 2471 1637 2498 1815
rect 2538 1777 2602 1789
rect 2878 1785 2915 1817
rect 2941 1816 3132 1838
rect 3267 1836 3376 1856
rect 3396 1836 3405 1856
rect 3267 1829 3405 1836
rect 3463 1856 3611 1865
rect 3463 1836 3472 1856
rect 3492 1836 3582 1856
rect 3602 1836 3611 1856
rect 3267 1827 3363 1829
rect 3463 1826 3611 1836
rect 3670 1856 3707 1866
rect 3670 1836 3678 1856
rect 3698 1836 3707 1856
rect 3519 1825 3555 1826
rect 3096 1814 3132 1816
rect 3096 1785 3133 1814
rect 2538 1776 2573 1777
rect 2515 1771 2573 1776
rect 2515 1751 2518 1771
rect 2538 1757 2573 1771
rect 2593 1757 2602 1777
rect 2538 1751 2602 1757
rect 2515 1749 2602 1751
rect 2515 1745 2542 1749
rect 2564 1748 2602 1749
rect 2565 1747 2602 1748
rect 2668 1781 2704 1782
rect 2776 1781 2812 1782
rect 2668 1774 2812 1781
rect 2668 1773 2730 1774
rect 2668 1753 2676 1773
rect 2696 1756 2730 1773
rect 2749 1773 2812 1774
rect 2749 1756 2784 1773
rect 2696 1753 2784 1756
rect 2804 1753 2812 1773
rect 2668 1747 2812 1753
rect 2878 1777 2916 1785
rect 2994 1781 3030 1782
rect 2878 1757 2887 1777
rect 2907 1757 2916 1777
rect 2878 1748 2916 1757
rect 2945 1773 3030 1781
rect 2945 1753 3002 1773
rect 3022 1753 3030 1773
rect 2878 1747 2915 1748
rect 2945 1747 3030 1753
rect 3096 1777 3134 1785
rect 3096 1757 3105 1777
rect 3125 1757 3134 1777
rect 3367 1766 3404 1767
rect 3670 1766 3707 1836
rect 3742 1865 3773 1916
rect 4069 1911 4114 1917
rect 4069 1893 4087 1911
rect 4105 1893 4114 1911
rect 4069 1883 4114 1893
rect 3792 1865 3829 1866
rect 3742 1856 3829 1865
rect 3742 1836 3800 1856
rect 3820 1836 3829 1856
rect 3742 1826 3829 1836
rect 3888 1856 3925 1866
rect 3888 1836 3896 1856
rect 3916 1836 3925 1856
rect 4069 1841 4112 1883
rect 3975 1839 4112 1841
rect 3742 1825 3773 1826
rect 3888 1766 3925 1836
rect 3366 1765 3707 1766
rect 3096 1748 3134 1757
rect 3291 1760 3707 1765
rect 3096 1747 3133 1748
rect 2557 1719 2647 1725
rect 2557 1699 2573 1719
rect 2593 1717 2647 1719
rect 2593 1699 2618 1717
rect 2557 1697 2618 1699
rect 2638 1697 2647 1717
rect 2557 1691 2647 1697
rect 2570 1637 2607 1638
rect 2666 1637 2703 1638
rect 2722 1637 2758 1747
rect 2945 1726 2976 1747
rect 3291 1740 3294 1760
rect 3314 1740 3707 1760
rect 3891 1750 3925 1766
rect 3969 1818 4112 1839
rect 3667 1731 3707 1740
rect 3969 1731 3996 1818
rect 4069 1792 4112 1818
rect 4069 1774 4082 1792
rect 4100 1774 4112 1792
rect 4069 1763 4112 1774
rect 2941 1725 2976 1726
rect 2819 1715 2976 1725
rect 2819 1695 2836 1715
rect 2856 1695 2976 1715
rect 2819 1688 2976 1695
rect 3043 1718 3189 1726
rect 3043 1698 3054 1718
rect 3074 1698 3113 1718
rect 3133 1698 3189 1718
rect 3667 1714 3996 1731
rect 3667 1713 3707 1714
rect 3043 1691 3189 1698
rect 4064 1702 4104 1705
rect 4064 1696 4107 1702
rect 3689 1693 4107 1696
rect 3043 1690 3084 1691
rect 2777 1637 2814 1638
rect 2470 1628 2608 1637
rect 2470 1608 2579 1628
rect 2599 1608 2608 1628
rect 2470 1601 2608 1608
rect 2666 1628 2814 1637
rect 2666 1608 2675 1628
rect 2695 1608 2785 1628
rect 2805 1608 2814 1628
rect 2470 1599 2566 1601
rect 2666 1598 2814 1608
rect 2873 1628 2910 1638
rect 2873 1608 2881 1628
rect 2901 1608 2910 1628
rect 2722 1597 2758 1598
rect 2570 1538 2607 1539
rect 2873 1538 2910 1608
rect 2945 1637 2976 1688
rect 3689 1675 4080 1693
rect 4098 1675 4107 1693
rect 3689 1673 4107 1675
rect 3689 1665 3716 1673
rect 3957 1670 4107 1673
rect 3269 1659 3437 1660
rect 3688 1659 3716 1665
rect 3269 1643 3716 1659
rect 4064 1665 4107 1670
rect 2995 1637 3032 1638
rect 2945 1628 3032 1637
rect 2945 1608 3003 1628
rect 3023 1608 3032 1628
rect 2945 1598 3032 1608
rect 3091 1628 3128 1638
rect 3091 1608 3099 1628
rect 3119 1608 3128 1628
rect 2945 1597 2976 1598
rect 2569 1537 2910 1538
rect 3091 1537 3128 1608
rect 2494 1532 2910 1537
rect 2494 1512 2497 1532
rect 2517 1512 2910 1532
rect 2941 1513 3128 1537
rect 3269 1633 3713 1643
rect 3269 1631 3437 1633
rect 2369 1433 2411 1478
rect 3269 1453 3296 1631
rect 3336 1593 3400 1605
rect 3676 1601 3713 1633
rect 3739 1632 3930 1654
rect 3894 1630 3930 1632
rect 3894 1601 3931 1630
rect 4064 1609 4104 1665
rect 3336 1592 3371 1593
rect 3313 1587 3371 1592
rect 3313 1567 3316 1587
rect 3336 1573 3371 1587
rect 3391 1573 3400 1593
rect 3336 1565 3400 1573
rect 3362 1564 3400 1565
rect 3363 1563 3400 1564
rect 3466 1597 3502 1598
rect 3574 1597 3610 1598
rect 3466 1589 3610 1597
rect 3466 1569 3474 1589
rect 3494 1569 3529 1589
rect 3549 1569 3582 1589
rect 3602 1569 3610 1589
rect 3466 1563 3610 1569
rect 3676 1593 3714 1601
rect 3792 1597 3828 1598
rect 3676 1573 3685 1593
rect 3705 1573 3714 1593
rect 3676 1564 3714 1573
rect 3743 1589 3828 1597
rect 3743 1569 3800 1589
rect 3820 1569 3828 1589
rect 3676 1563 3713 1564
rect 3743 1563 3828 1569
rect 3894 1593 3932 1601
rect 3894 1573 3903 1593
rect 3923 1573 3932 1593
rect 4064 1591 4076 1609
rect 4094 1591 4104 1609
rect 4064 1581 4104 1591
rect 3894 1564 3932 1573
rect 3894 1563 3931 1564
rect 3355 1535 3445 1541
rect 3355 1515 3371 1535
rect 3391 1533 3445 1535
rect 3391 1515 3416 1533
rect 3355 1513 3416 1515
rect 3436 1513 3445 1533
rect 3355 1507 3445 1513
rect 3368 1453 3405 1454
rect 3464 1453 3501 1454
rect 3520 1453 3556 1563
rect 3743 1542 3774 1563
rect 3739 1541 3774 1542
rect 3617 1531 3774 1541
rect 3617 1511 3634 1531
rect 3654 1511 3774 1531
rect 3617 1504 3774 1511
rect 3841 1534 3990 1542
rect 3841 1514 3852 1534
rect 3872 1514 3911 1534
rect 3931 1514 3990 1534
rect 3841 1507 3990 1514
rect 4056 1510 4108 1528
rect 3841 1506 3882 1507
rect 3575 1453 3612 1454
rect 3268 1444 3406 1453
rect 2740 1433 2773 1435
rect 2369 1421 2816 1433
rect 1601 1299 1769 1301
rect 1325 1273 1769 1299
rect 835 1251 973 1260
rect 629 1250 666 1251
rect 126 1196 163 1199
rect 359 1197 400 1198
rect 251 1190 400 1197
rect 251 1170 310 1190
rect 330 1170 369 1190
rect 389 1170 400 1190
rect 251 1162 400 1170
rect 467 1193 624 1200
rect 467 1173 587 1193
rect 607 1173 624 1193
rect 467 1163 624 1173
rect 467 1162 502 1163
rect 467 1141 498 1162
rect 685 1141 721 1251
rect 740 1250 777 1251
rect 836 1250 873 1251
rect 796 1191 886 1197
rect 796 1171 805 1191
rect 825 1189 886 1191
rect 825 1171 850 1189
rect 796 1169 850 1171
rect 870 1169 886 1189
rect 796 1163 886 1169
rect 310 1140 347 1141
rect 123 1132 160 1134
rect 123 1124 165 1132
rect 123 1106 133 1124
rect 151 1106 165 1124
rect 123 1097 165 1106
rect 309 1131 347 1140
rect 309 1111 318 1131
rect 338 1111 347 1131
rect 309 1103 347 1111
rect 413 1135 498 1141
rect 528 1140 565 1141
rect 413 1115 421 1135
rect 441 1115 498 1135
rect 413 1107 498 1115
rect 527 1131 565 1140
rect 527 1111 536 1131
rect 556 1111 565 1131
rect 413 1106 449 1107
rect 527 1103 565 1111
rect 631 1139 775 1141
rect 631 1135 683 1139
rect 631 1115 639 1135
rect 659 1119 683 1135
rect 703 1135 775 1139
rect 703 1119 747 1135
rect 659 1115 747 1119
rect 767 1115 775 1135
rect 631 1107 775 1115
rect 631 1106 667 1107
rect 739 1106 775 1107
rect 841 1140 878 1141
rect 841 1139 879 1140
rect 841 1131 905 1139
rect 841 1111 850 1131
rect 870 1117 905 1131
rect 925 1117 928 1137
rect 870 1112 928 1117
rect 870 1111 905 1112
rect 124 1072 165 1097
rect 310 1072 347 1103
rect 528 1072 565 1103
rect 841 1099 905 1111
rect 945 1073 972 1251
rect 124 1045 173 1072
rect 309 1046 358 1072
rect 527 1071 608 1072
rect 804 1071 972 1073
rect 527 1046 972 1071
rect 528 1045 972 1046
rect 126 1012 173 1045
rect 529 1012 569 1045
rect 804 1044 972 1045
rect 1435 1049 1475 1273
rect 1601 1272 1769 1273
rect 2372 1407 2816 1421
rect 2372 1405 2540 1407
rect 2372 1227 2399 1405
rect 2439 1367 2503 1379
rect 2779 1375 2816 1407
rect 2842 1406 3033 1428
rect 3268 1424 3377 1444
rect 3397 1424 3406 1444
rect 3268 1417 3406 1424
rect 3464 1444 3612 1453
rect 3464 1424 3473 1444
rect 3493 1424 3583 1444
rect 3603 1424 3612 1444
rect 3268 1415 3364 1417
rect 3464 1414 3612 1424
rect 3671 1444 3708 1454
rect 3671 1424 3679 1444
rect 3699 1424 3708 1444
rect 3520 1413 3556 1414
rect 2997 1404 3033 1406
rect 2997 1375 3034 1404
rect 2439 1366 2474 1367
rect 2416 1361 2474 1366
rect 2416 1341 2419 1361
rect 2439 1347 2474 1361
rect 2494 1347 2503 1367
rect 2439 1339 2503 1347
rect 2465 1338 2503 1339
rect 2466 1337 2503 1338
rect 2569 1371 2605 1372
rect 2677 1371 2713 1372
rect 2569 1363 2713 1371
rect 2569 1343 2577 1363
rect 2597 1361 2685 1363
rect 2597 1343 2630 1361
rect 2569 1342 2630 1343
rect 2651 1343 2685 1361
rect 2705 1343 2713 1363
rect 2651 1342 2713 1343
rect 2569 1337 2713 1342
rect 2779 1367 2817 1375
rect 2895 1371 2931 1372
rect 2779 1347 2788 1367
rect 2808 1347 2817 1367
rect 2779 1338 2817 1347
rect 2846 1363 2931 1371
rect 2846 1343 2903 1363
rect 2923 1343 2931 1363
rect 2779 1337 2816 1338
rect 2846 1337 2931 1343
rect 2997 1367 3035 1375
rect 2997 1347 3006 1367
rect 3026 1347 3035 1367
rect 3671 1357 3708 1424
rect 3743 1453 3774 1504
rect 4056 1492 4074 1510
rect 4092 1492 4108 1510
rect 3793 1453 3830 1454
rect 3743 1444 3830 1453
rect 3743 1424 3801 1444
rect 3821 1424 3830 1444
rect 3743 1414 3830 1424
rect 3889 1444 3926 1454
rect 3889 1424 3897 1444
rect 3917 1424 3926 1444
rect 3743 1413 3774 1414
rect 3368 1354 3405 1355
rect 3671 1354 3710 1357
rect 3367 1353 3710 1354
rect 3889 1353 3926 1424
rect 2997 1338 3035 1347
rect 3292 1348 3710 1353
rect 2997 1337 3034 1338
rect 2458 1309 2548 1315
rect 2458 1289 2474 1309
rect 2494 1307 2548 1309
rect 2494 1289 2519 1307
rect 2458 1287 2519 1289
rect 2539 1287 2548 1307
rect 2458 1281 2548 1287
rect 2471 1227 2508 1228
rect 2567 1227 2604 1228
rect 2623 1227 2659 1337
rect 2846 1316 2877 1337
rect 3292 1328 3295 1348
rect 3315 1328 3710 1348
rect 3739 1329 3926 1353
rect 2842 1315 2877 1316
rect 2720 1305 2877 1315
rect 2720 1285 2737 1305
rect 2757 1285 2877 1305
rect 2720 1278 2877 1285
rect 2944 1308 3093 1316
rect 2944 1288 2955 1308
rect 2975 1288 3014 1308
rect 3034 1288 3093 1308
rect 2944 1281 3093 1288
rect 3671 1303 3710 1328
rect 4056 1303 4108 1492
rect 3671 1285 4110 1303
rect 2944 1280 2985 1281
rect 2678 1227 2715 1228
rect 2371 1218 2509 1227
rect 2371 1198 2480 1218
rect 2500 1198 2509 1218
rect 2371 1191 2509 1198
rect 2567 1218 2715 1227
rect 2567 1198 2576 1218
rect 2596 1198 2686 1218
rect 2706 1198 2715 1218
rect 2371 1189 2467 1191
rect 2567 1188 2715 1198
rect 2774 1218 2811 1228
rect 2774 1198 2782 1218
rect 2802 1198 2811 1218
rect 2623 1187 2659 1188
rect 2471 1128 2508 1129
rect 2774 1128 2811 1198
rect 2846 1227 2877 1278
rect 3671 1267 4071 1285
rect 4089 1267 4110 1285
rect 3671 1261 4110 1267
rect 3677 1257 4110 1261
rect 4056 1255 4108 1257
rect 2896 1227 2933 1228
rect 2846 1218 2933 1227
rect 2846 1198 2904 1218
rect 2924 1198 2933 1218
rect 2846 1188 2933 1198
rect 2992 1218 3029 1228
rect 2992 1198 3000 1218
rect 3020 1198 3029 1218
rect 2846 1187 2877 1188
rect 2470 1127 2811 1128
rect 2992 1127 3029 1198
rect 4059 1190 4096 1195
rect 4050 1186 4097 1190
rect 4050 1168 4069 1186
rect 4087 1168 4097 1186
rect 2395 1122 2811 1127
rect 2395 1102 2398 1122
rect 2418 1102 2811 1122
rect 2842 1103 3029 1127
rect 3654 1125 3694 1130
rect 4050 1125 4097 1168
rect 3654 1086 4097 1125
rect 1435 1027 1443 1049
rect 1467 1027 1475 1049
rect 1435 1019 1475 1027
rect 2748 1071 2788 1079
rect 2748 1049 2756 1071
rect 2780 1049 2788 1071
rect 126 973 569 1012
rect 126 930 173 973
rect 529 968 569 973
rect 1194 971 1381 995
rect 1412 976 1805 996
rect 1825 976 1828 996
rect 1412 971 1828 976
rect 126 912 136 930
rect 154 912 173 930
rect 126 908 173 912
rect 127 903 164 908
rect 1194 900 1231 971
rect 1412 970 1753 971
rect 1346 910 1377 911
rect 1194 880 1203 900
rect 1223 880 1231 900
rect 1194 870 1231 880
rect 1290 900 1377 910
rect 1290 880 1299 900
rect 1319 880 1377 900
rect 1290 871 1377 880
rect 1290 870 1327 871
rect 115 841 167 843
rect 113 837 546 841
rect 113 831 552 837
rect 113 813 134 831
rect 152 813 552 831
rect 1346 820 1377 871
rect 1412 900 1449 970
rect 1715 969 1752 970
rect 1564 910 1600 911
rect 1412 880 1421 900
rect 1441 880 1449 900
rect 1412 870 1449 880
rect 1508 900 1656 910
rect 1756 907 1852 909
rect 1508 880 1517 900
rect 1537 880 1627 900
rect 1647 880 1656 900
rect 1508 871 1656 880
rect 1714 900 1852 907
rect 1714 880 1723 900
rect 1743 880 1852 900
rect 1714 871 1852 880
rect 1508 870 1545 871
rect 1238 817 1279 818
rect 113 795 552 813
rect 115 606 167 795
rect 513 770 552 795
rect 1130 810 1279 817
rect 1130 790 1189 810
rect 1209 790 1248 810
rect 1268 790 1279 810
rect 1130 782 1279 790
rect 1346 813 1503 820
rect 1346 793 1466 813
rect 1486 793 1503 813
rect 1346 783 1503 793
rect 1346 782 1381 783
rect 297 745 484 769
rect 513 750 908 770
rect 928 750 931 770
rect 1346 761 1377 782
rect 1564 761 1600 871
rect 1619 870 1656 871
rect 1715 870 1752 871
rect 1675 811 1765 817
rect 1675 791 1684 811
rect 1704 809 1765 811
rect 1704 791 1729 809
rect 1675 789 1729 791
rect 1749 789 1765 809
rect 1675 783 1765 789
rect 1189 760 1226 761
rect 513 745 931 750
rect 1188 751 1226 760
rect 297 674 334 745
rect 513 744 856 745
rect 513 741 552 744
rect 818 743 855 744
rect 449 684 480 685
rect 297 654 306 674
rect 326 654 334 674
rect 297 644 334 654
rect 393 674 480 684
rect 393 654 402 674
rect 422 654 480 674
rect 393 645 480 654
rect 393 644 430 645
rect 115 588 131 606
rect 149 588 167 606
rect 449 594 480 645
rect 515 674 552 741
rect 1188 731 1197 751
rect 1217 731 1226 751
rect 1188 723 1226 731
rect 1292 755 1377 761
rect 1407 760 1444 761
rect 1292 735 1300 755
rect 1320 735 1377 755
rect 1292 727 1377 735
rect 1406 751 1444 760
rect 1406 731 1415 751
rect 1435 731 1444 751
rect 1292 726 1328 727
rect 1406 723 1444 731
rect 1510 755 1654 761
rect 1510 735 1518 755
rect 1538 750 1626 755
rect 1538 735 1574 750
rect 1510 733 1574 735
rect 1593 735 1626 750
rect 1646 735 1654 755
rect 1593 733 1654 735
rect 1510 727 1654 733
rect 1510 726 1546 727
rect 1618 726 1654 727
rect 1720 760 1757 761
rect 1720 759 1758 760
rect 1720 751 1784 759
rect 1720 731 1729 751
rect 1749 737 1784 751
rect 1804 737 1807 757
rect 1749 732 1807 737
rect 1749 731 1784 732
rect 1189 694 1226 723
rect 1190 692 1226 694
rect 667 684 703 685
rect 515 654 524 674
rect 544 654 552 674
rect 515 644 552 654
rect 611 674 759 684
rect 859 681 955 683
rect 611 654 620 674
rect 640 654 730 674
rect 750 654 759 674
rect 611 645 759 654
rect 817 674 955 681
rect 817 654 826 674
rect 846 654 955 674
rect 1190 670 1381 692
rect 1407 691 1444 723
rect 1720 719 1784 731
rect 1824 693 1851 871
rect 1683 691 1851 693
rect 1407 677 1851 691
rect 2454 825 2622 826
rect 2748 825 2788 1049
rect 3251 1053 3419 1054
rect 3654 1053 3694 1086
rect 4050 1053 4097 1086
rect 3251 1052 3695 1053
rect 3251 1027 3696 1052
rect 3251 1025 3419 1027
rect 3615 1026 3696 1027
rect 3865 1026 3914 1052
rect 4050 1026 4099 1053
rect 3251 847 3278 1025
rect 3318 987 3382 999
rect 3658 995 3695 1026
rect 3876 995 3913 1026
rect 4058 1001 4099 1026
rect 3318 986 3353 987
rect 3295 981 3353 986
rect 3295 961 3298 981
rect 3318 967 3353 981
rect 3373 967 3382 987
rect 3318 959 3382 967
rect 3344 958 3382 959
rect 3345 957 3382 958
rect 3448 991 3484 992
rect 3556 991 3592 992
rect 3448 983 3592 991
rect 3448 963 3456 983
rect 3476 979 3564 983
rect 3476 963 3520 979
rect 3448 959 3520 963
rect 3540 963 3564 979
rect 3584 963 3592 983
rect 3540 959 3592 963
rect 3448 957 3592 959
rect 3658 987 3696 995
rect 3774 991 3810 992
rect 3658 967 3667 987
rect 3687 967 3696 987
rect 3658 958 3696 967
rect 3725 983 3810 991
rect 3725 963 3782 983
rect 3802 963 3810 983
rect 3658 957 3695 958
rect 3725 957 3810 963
rect 3876 987 3914 995
rect 3876 967 3885 987
rect 3905 967 3914 987
rect 3876 958 3914 967
rect 4058 992 4100 1001
rect 4058 974 4072 992
rect 4090 974 4100 992
rect 4058 966 4100 974
rect 4063 964 4100 966
rect 3876 957 3913 958
rect 3337 929 3427 935
rect 3337 909 3353 929
rect 3373 927 3427 929
rect 3373 909 3398 927
rect 3337 907 3398 909
rect 3418 907 3427 927
rect 3337 901 3427 907
rect 3350 847 3387 848
rect 3446 847 3483 848
rect 3502 847 3538 957
rect 3725 936 3756 957
rect 3721 935 3756 936
rect 3599 925 3756 935
rect 3599 905 3616 925
rect 3636 905 3756 925
rect 3599 898 3756 905
rect 3823 928 3972 936
rect 3823 908 3834 928
rect 3854 908 3893 928
rect 3913 908 3972 928
rect 3823 901 3972 908
rect 3823 900 3864 901
rect 4060 899 4097 902
rect 3557 847 3594 848
rect 3250 838 3388 847
rect 2454 799 2898 825
rect 2454 797 2622 799
rect 1407 665 1854 677
rect 1450 663 1483 665
rect 817 645 955 654
rect 611 644 648 645
rect 341 591 382 592
rect 115 570 167 588
rect 233 584 382 591
rect 233 564 292 584
rect 312 564 351 584
rect 371 564 382 584
rect 233 556 382 564
rect 449 587 606 594
rect 449 567 569 587
rect 589 567 606 587
rect 449 557 606 567
rect 449 556 484 557
rect 449 535 480 556
rect 667 535 703 645
rect 722 644 759 645
rect 818 644 855 645
rect 778 585 868 591
rect 778 565 787 585
rect 807 583 868 585
rect 807 565 832 583
rect 778 563 832 565
rect 852 563 868 583
rect 778 557 868 563
rect 292 534 329 535
rect 291 525 329 534
rect 119 507 159 517
rect 119 489 129 507
rect 147 489 159 507
rect 291 505 300 525
rect 320 505 329 525
rect 291 497 329 505
rect 395 529 480 535
rect 510 534 547 535
rect 395 509 403 529
rect 423 509 480 529
rect 395 501 480 509
rect 509 525 547 534
rect 509 505 518 525
rect 538 505 547 525
rect 395 500 431 501
rect 509 497 547 505
rect 613 529 757 535
rect 613 509 621 529
rect 641 509 674 529
rect 694 509 729 529
rect 749 509 757 529
rect 613 501 757 509
rect 613 500 649 501
rect 721 500 757 501
rect 823 534 860 535
rect 823 533 861 534
rect 823 525 887 533
rect 823 505 832 525
rect 852 511 887 525
rect 907 511 910 531
rect 852 506 910 511
rect 852 505 887 506
rect 119 433 159 489
rect 292 468 329 497
rect 293 466 329 468
rect 293 444 484 466
rect 510 465 547 497
rect 823 493 887 505
rect 927 467 954 645
rect 1812 620 1854 665
rect 786 465 954 467
rect 510 455 954 465
rect 1095 561 1282 585
rect 1313 566 1706 586
rect 1726 566 1729 586
rect 1313 561 1729 566
rect 1095 490 1132 561
rect 1313 560 1654 561
rect 1247 500 1278 501
rect 1095 470 1104 490
rect 1124 470 1132 490
rect 1095 460 1132 470
rect 1191 490 1278 500
rect 1191 470 1200 490
rect 1220 470 1278 490
rect 1191 461 1278 470
rect 1191 460 1228 461
rect 116 428 159 433
rect 507 439 954 455
rect 507 433 535 439
rect 786 438 954 439
rect 116 425 266 428
rect 507 425 534 433
rect 116 423 534 425
rect 116 405 125 423
rect 143 405 534 423
rect 1247 410 1278 461
rect 1313 490 1350 560
rect 1616 559 1653 560
rect 1465 500 1501 501
rect 1313 470 1322 490
rect 1342 470 1350 490
rect 1313 460 1350 470
rect 1409 490 1557 500
rect 1657 497 1753 499
rect 1409 470 1418 490
rect 1438 470 1528 490
rect 1548 470 1557 490
rect 1409 461 1557 470
rect 1615 490 1753 497
rect 1615 470 1624 490
rect 1644 470 1753 490
rect 1615 461 1753 470
rect 1409 460 1446 461
rect 1139 407 1180 408
rect 116 402 534 405
rect 116 396 159 402
rect 119 393 159 396
rect 1034 400 1180 407
rect 516 384 556 385
rect 227 367 556 384
rect 1034 380 1090 400
rect 1110 380 1149 400
rect 1169 380 1180 400
rect 1034 372 1180 380
rect 1247 403 1404 410
rect 1247 383 1367 403
rect 1387 383 1404 403
rect 1247 373 1404 383
rect 1247 372 1282 373
rect 111 324 154 335
rect 111 306 123 324
rect 141 306 154 324
rect 111 280 154 306
rect 227 280 254 367
rect 516 358 556 367
rect 111 259 254 280
rect 298 332 332 348
rect 516 338 909 358
rect 929 338 932 358
rect 1247 351 1278 372
rect 1465 351 1501 461
rect 1520 460 1557 461
rect 1616 460 1653 461
rect 1576 401 1666 407
rect 1576 381 1585 401
rect 1605 399 1666 401
rect 1605 381 1630 399
rect 1576 379 1630 381
rect 1650 379 1666 399
rect 1576 373 1666 379
rect 1090 350 1127 351
rect 516 333 932 338
rect 1089 341 1127 350
rect 516 332 857 333
rect 298 262 335 332
rect 450 272 481 273
rect 111 257 248 259
rect 111 215 154 257
rect 298 242 307 262
rect 327 242 335 262
rect 298 232 335 242
rect 394 262 481 272
rect 394 242 403 262
rect 423 242 481 262
rect 394 233 481 242
rect 394 232 431 233
rect 109 205 154 215
rect 109 187 118 205
rect 136 187 154 205
rect 109 181 154 187
rect 450 182 481 233
rect 516 262 553 332
rect 819 331 856 332
rect 1089 321 1098 341
rect 1118 321 1127 341
rect 1089 313 1127 321
rect 1193 345 1278 351
rect 1308 350 1345 351
rect 1193 325 1201 345
rect 1221 325 1278 345
rect 1193 317 1278 325
rect 1307 341 1345 350
rect 1307 321 1316 341
rect 1336 321 1345 341
rect 1193 316 1229 317
rect 1307 313 1345 321
rect 1411 345 1555 351
rect 1411 325 1419 345
rect 1439 342 1527 345
rect 1439 325 1474 342
rect 1411 324 1474 325
rect 1493 325 1527 342
rect 1547 325 1555 345
rect 1493 324 1555 325
rect 1411 317 1555 324
rect 1411 316 1447 317
rect 1519 316 1555 317
rect 1621 350 1658 351
rect 1621 349 1659 350
rect 1681 349 1708 353
rect 1621 347 1708 349
rect 1621 341 1685 347
rect 1621 321 1630 341
rect 1650 327 1685 341
rect 1705 327 1708 347
rect 1650 322 1708 327
rect 1650 321 1685 322
rect 1090 284 1127 313
rect 1091 282 1127 284
rect 668 272 704 273
rect 516 242 525 262
rect 545 242 553 262
rect 516 232 553 242
rect 612 262 760 272
rect 860 269 956 271
rect 612 242 621 262
rect 641 242 731 262
rect 751 242 760 262
rect 612 233 760 242
rect 818 262 956 269
rect 818 242 827 262
rect 847 242 956 262
rect 1091 260 1282 282
rect 1308 281 1345 313
rect 1621 309 1685 321
rect 1725 283 1752 461
rect 1584 281 1752 283
rect 1308 255 1752 281
rect 818 233 956 242
rect 612 232 649 233
rect 109 178 146 181
rect 342 179 383 180
rect 234 172 383 179
rect 234 152 293 172
rect 313 152 352 172
rect 372 152 383 172
rect 234 144 383 152
rect 450 175 607 182
rect 450 155 570 175
rect 590 155 607 175
rect 450 145 607 155
rect 450 144 485 145
rect 450 123 481 144
rect 668 123 704 233
rect 723 232 760 233
rect 819 232 856 233
rect 779 173 869 179
rect 779 153 788 173
rect 808 171 869 173
rect 808 153 833 171
rect 779 151 833 153
rect 853 151 869 171
rect 779 145 869 151
rect 293 122 330 123
rect 106 114 143 116
rect 106 106 148 114
rect 106 88 116 106
rect 134 88 148 106
rect 106 79 148 88
rect 292 113 330 122
rect 292 93 301 113
rect 321 93 330 113
rect 292 85 330 93
rect 396 117 481 123
rect 511 122 548 123
rect 396 97 404 117
rect 424 97 481 117
rect 396 89 481 97
rect 510 113 548 122
rect 510 93 519 113
rect 539 93 548 113
rect 396 88 432 89
rect 510 85 548 93
rect 614 121 758 123
rect 614 117 666 121
rect 614 97 622 117
rect 642 101 666 117
rect 686 117 758 121
rect 686 101 730 117
rect 642 97 730 101
rect 750 97 758 117
rect 614 89 758 97
rect 614 88 650 89
rect 722 88 758 89
rect 824 122 861 123
rect 824 121 862 122
rect 824 113 888 121
rect 824 93 833 113
rect 853 99 888 113
rect 908 99 911 119
rect 853 94 911 99
rect 853 93 888 94
rect 107 54 148 79
rect 293 54 330 85
rect 511 63 548 85
rect 824 81 888 93
rect 506 54 548 63
rect 928 55 955 233
rect 107 42 152 54
rect 103 -16 152 42
rect 293 28 355 54
rect 506 53 591 54
rect 787 53 955 55
rect 506 27 955 53
rect 506 -16 545 27
rect 787 26 955 27
rect 1418 31 1458 255
rect 1584 254 1752 255
rect 1816 287 1849 620
rect 2454 619 2481 797
rect 2521 759 2585 771
rect 2861 767 2898 799
rect 2924 798 3115 820
rect 3250 818 3359 838
rect 3379 818 3388 838
rect 3250 811 3388 818
rect 3446 838 3594 847
rect 3446 818 3455 838
rect 3475 818 3565 838
rect 3585 818 3594 838
rect 3250 809 3346 811
rect 3446 808 3594 818
rect 3653 838 3690 848
rect 3653 818 3661 838
rect 3681 818 3690 838
rect 3502 807 3538 808
rect 3079 796 3115 798
rect 3079 767 3116 796
rect 2521 758 2556 759
rect 2498 753 2556 758
rect 2498 733 2501 753
rect 2521 739 2556 753
rect 2576 739 2585 759
rect 2521 731 2585 739
rect 2547 730 2585 731
rect 2548 729 2585 730
rect 2651 763 2687 764
rect 2759 763 2795 764
rect 2651 755 2795 763
rect 2651 735 2659 755
rect 2679 754 2767 755
rect 2679 735 2714 754
rect 2735 735 2767 754
rect 2787 735 2795 755
rect 2651 729 2795 735
rect 2861 759 2899 767
rect 2977 763 3013 764
rect 2861 739 2870 759
rect 2890 739 2899 759
rect 2861 730 2899 739
rect 2928 755 3013 763
rect 2928 735 2985 755
rect 3005 735 3013 755
rect 2861 729 2898 730
rect 2928 729 3013 735
rect 3079 759 3117 767
rect 3079 739 3088 759
rect 3108 739 3117 759
rect 3350 748 3387 749
rect 3653 748 3690 818
rect 3725 847 3756 898
rect 4052 893 4097 899
rect 4052 875 4070 893
rect 4088 875 4097 893
rect 4052 865 4097 875
rect 3775 847 3812 848
rect 3725 838 3812 847
rect 3725 818 3783 838
rect 3803 818 3812 838
rect 3725 808 3812 818
rect 3871 838 3908 848
rect 3871 818 3879 838
rect 3899 818 3908 838
rect 4052 823 4095 865
rect 3958 821 4095 823
rect 3725 807 3756 808
rect 3871 748 3908 818
rect 3349 747 3690 748
rect 3079 730 3117 739
rect 3274 742 3690 747
rect 3079 729 3116 730
rect 2540 701 2630 707
rect 2540 681 2556 701
rect 2576 699 2630 701
rect 2576 681 2601 699
rect 2540 679 2601 681
rect 2621 679 2630 699
rect 2540 673 2630 679
rect 2553 619 2590 620
rect 2649 619 2686 620
rect 2705 619 2741 729
rect 2928 708 2959 729
rect 3274 722 3277 742
rect 3297 722 3690 742
rect 3874 732 3908 748
rect 3952 800 4095 821
rect 3650 713 3690 722
rect 3952 713 3979 800
rect 4052 774 4095 800
rect 4052 756 4065 774
rect 4083 756 4095 774
rect 4052 745 4095 756
rect 2924 707 2959 708
rect 2802 697 2959 707
rect 2802 677 2819 697
rect 2839 677 2959 697
rect 2802 670 2959 677
rect 3026 700 3175 708
rect 3026 680 3037 700
rect 3057 680 3096 700
rect 3116 680 3175 700
rect 3650 696 3979 713
rect 3650 695 3690 696
rect 3026 673 3175 680
rect 4047 684 4087 687
rect 4047 678 4090 684
rect 3672 675 4090 678
rect 3026 672 3067 673
rect 2760 619 2797 620
rect 2453 610 2591 619
rect 2453 590 2562 610
rect 2582 590 2591 610
rect 2453 583 2591 590
rect 2649 610 2797 619
rect 2649 590 2658 610
rect 2678 590 2768 610
rect 2788 590 2797 610
rect 2453 581 2549 583
rect 2649 580 2797 590
rect 2856 610 2893 620
rect 2856 590 2864 610
rect 2884 590 2893 610
rect 2705 579 2741 580
rect 2553 520 2590 521
rect 2856 520 2893 590
rect 2928 619 2959 670
rect 3672 657 4063 675
rect 4081 657 4090 675
rect 3672 655 4090 657
rect 3672 647 3699 655
rect 3940 652 4090 655
rect 3252 641 3420 642
rect 3671 641 3699 647
rect 3252 625 3699 641
rect 4047 647 4090 652
rect 2978 619 3015 620
rect 2928 610 3015 619
rect 2928 590 2986 610
rect 3006 590 3015 610
rect 2928 580 3015 590
rect 3074 610 3111 620
rect 3074 590 3082 610
rect 3102 590 3111 610
rect 2928 579 2959 580
rect 2552 519 2893 520
rect 3074 519 3111 590
rect 2477 514 2893 519
rect 2477 494 2480 514
rect 2500 494 2893 514
rect 2924 495 3111 519
rect 3252 615 3696 625
rect 3252 613 3420 615
rect 3252 435 3279 613
rect 3319 575 3383 587
rect 3659 583 3696 615
rect 3722 614 3913 636
rect 3877 612 3913 614
rect 3877 583 3914 612
rect 4047 591 4087 647
rect 3319 574 3354 575
rect 3296 569 3354 574
rect 3296 549 3299 569
rect 3319 555 3354 569
rect 3374 555 3383 575
rect 3319 547 3383 555
rect 3345 546 3383 547
rect 3346 545 3383 546
rect 3449 579 3485 580
rect 3557 579 3593 580
rect 3449 571 3593 579
rect 3449 551 3457 571
rect 3477 551 3512 571
rect 3532 551 3565 571
rect 3585 551 3593 571
rect 3449 545 3593 551
rect 3659 575 3697 583
rect 3775 579 3811 580
rect 3659 555 3668 575
rect 3688 555 3697 575
rect 3659 546 3697 555
rect 3726 571 3811 579
rect 3726 551 3783 571
rect 3803 551 3811 571
rect 3659 545 3696 546
rect 3726 545 3811 551
rect 3877 575 3915 583
rect 3877 555 3886 575
rect 3906 555 3915 575
rect 4047 573 4059 591
rect 4077 573 4087 591
rect 4047 563 4087 573
rect 3877 546 3915 555
rect 3877 545 3914 546
rect 3338 517 3428 523
rect 3338 497 3354 517
rect 3374 515 3428 517
rect 3374 497 3399 515
rect 3338 495 3399 497
rect 3419 495 3428 515
rect 3338 489 3428 495
rect 3351 435 3388 436
rect 3447 435 3484 436
rect 3503 435 3539 545
rect 3726 524 3757 545
rect 3722 523 3757 524
rect 3600 513 3757 523
rect 3600 493 3617 513
rect 3637 493 3757 513
rect 3600 486 3757 493
rect 3824 516 3973 524
rect 3824 496 3835 516
rect 3855 496 3894 516
rect 3914 496 3973 516
rect 3824 489 3973 496
rect 4039 492 4091 510
rect 3824 488 3865 489
rect 3558 435 3595 436
rect 3251 426 3389 435
rect 3251 406 3360 426
rect 3380 406 3389 426
rect 3251 399 3389 406
rect 3447 426 3595 435
rect 3447 406 3456 426
rect 3476 406 3566 426
rect 3586 406 3595 426
rect 3251 397 3347 399
rect 3447 396 3595 406
rect 3654 426 3691 436
rect 3654 406 3662 426
rect 3682 406 3691 426
rect 3503 395 3539 396
rect 3654 339 3691 406
rect 3726 435 3757 486
rect 4039 474 4057 492
rect 4075 474 4091 492
rect 3776 435 3813 436
rect 3726 426 3813 435
rect 3726 406 3784 426
rect 3804 406 3813 426
rect 3726 396 3813 406
rect 3872 426 3909 436
rect 3872 406 3880 426
rect 3900 406 3909 426
rect 3726 395 3757 396
rect 3351 336 3388 337
rect 3654 336 3693 339
rect 3350 335 3693 336
rect 3872 335 3909 406
rect 3275 330 3693 335
rect 3275 310 3278 330
rect 3298 310 3693 330
rect 3722 311 3909 335
rect 1816 279 1853 287
rect 1816 260 1824 279
rect 1845 260 1853 279
rect 1816 254 1853 260
rect 3654 285 3693 310
rect 4039 285 4091 474
rect 3654 267 4093 285
rect 3654 249 4054 267
rect 4072 249 4093 267
rect 3654 243 4093 249
rect 3660 239 4093 243
rect 4039 237 4091 239
rect 4042 172 4079 177
rect 4033 168 4080 172
rect 4033 150 4052 168
rect 4070 150 4080 168
rect 4033 87 4080 150
rect 4033 72 4083 87
rect 4033 47 4047 72
rect 4079 47 4083 72
rect 4033 34 4080 47
rect 1418 9 1426 31
rect 1450 9 1458 31
rect 1418 1 1458 9
rect 101 -43 506 -16
rect 542 -43 545 -16
rect 101 -47 545 -43
rect 101 -48 527 -47
rect 1860 -218 1925 -217
rect 1511 -243 1698 -219
rect 1729 -239 2122 -218
rect 2143 -239 2145 -218
rect 1729 -243 2145 -239
rect 1511 -314 1548 -243
rect 1729 -244 2070 -243
rect 1663 -304 1694 -303
rect 1511 -334 1520 -314
rect 1540 -334 1548 -314
rect 1511 -344 1548 -334
rect 1607 -314 1694 -304
rect 1607 -334 1616 -314
rect 1636 -334 1694 -314
rect 1607 -343 1694 -334
rect 1607 -344 1644 -343
rect 1663 -394 1694 -343
rect 1729 -314 1766 -244
rect 2032 -245 2069 -244
rect 1881 -304 1917 -303
rect 1729 -334 1738 -314
rect 1758 -334 1766 -314
rect 1729 -344 1766 -334
rect 1825 -314 1973 -304
rect 2073 -307 2234 -305
rect 1825 -334 1834 -314
rect 1854 -334 1944 -314
rect 1964 -334 1973 -314
rect 1825 -343 1973 -334
rect 2031 -312 2234 -307
rect 2031 -314 2204 -312
rect 2031 -334 2040 -314
rect 2060 -332 2204 -314
rect 2224 -332 2234 -312
rect 2060 -334 2234 -332
rect 2031 -341 2234 -334
rect 2031 -343 2169 -341
rect 1825 -344 1862 -343
rect 1555 -397 1596 -396
rect 1447 -404 1596 -397
rect 1447 -424 1506 -404
rect 1526 -424 1565 -404
rect 1585 -424 1596 -404
rect 1447 -432 1596 -424
rect 1663 -401 1820 -394
rect 1663 -421 1783 -401
rect 1803 -421 1820 -401
rect 1663 -431 1820 -421
rect 1663 -432 1698 -431
rect 1663 -453 1694 -432
rect 1881 -453 1917 -343
rect 1936 -344 1973 -343
rect 2032 -344 2069 -343
rect 1992 -403 2082 -397
rect 1992 -423 2001 -403
rect 2021 -405 2082 -403
rect 2021 -423 2046 -405
rect 1992 -425 2046 -423
rect 2066 -425 2082 -405
rect 1992 -431 2082 -425
rect 1506 -454 1543 -453
rect 1505 -463 1543 -454
rect 1505 -483 1514 -463
rect 1534 -483 1543 -463
rect 1505 -491 1543 -483
rect 1609 -459 1694 -453
rect 1724 -454 1761 -453
rect 1609 -479 1617 -459
rect 1637 -479 1694 -459
rect 1609 -487 1694 -479
rect 1723 -463 1761 -454
rect 1723 -483 1732 -463
rect 1752 -483 1761 -463
rect 1609 -488 1645 -487
rect 1723 -491 1761 -483
rect 1827 -459 1971 -453
rect 1827 -479 1835 -459
rect 1855 -479 1943 -459
rect 1963 -479 1971 -459
rect 1827 -487 1971 -479
rect 1827 -488 1863 -487
rect 1935 -488 1971 -487
rect 2037 -454 2074 -453
rect 2037 -455 2075 -454
rect 2037 -463 2101 -455
rect 2037 -483 2046 -463
rect 2066 -477 2101 -463
rect 2121 -477 2124 -457
rect 2066 -482 2124 -477
rect 2066 -483 2101 -482
rect 1506 -520 1543 -491
rect 1507 -522 1543 -520
rect 1507 -544 1698 -522
rect 1724 -523 1761 -491
rect 2037 -495 2101 -483
rect 2141 -521 2168 -343
rect 2000 -523 2168 -521
rect 1724 -549 2168 -523
rect 1834 -552 1874 -549
rect 2000 -550 2168 -549
<< viali >>
rect 2883 8175 2907 8197
rect 2488 7927 2509 7946
rect 1035 7876 1055 7896
rect 419 7690 439 7710
rect 959 7689 979 7709
rect 801 7635 821 7655
rect 1014 7637 1034 7657
rect 1833 7692 1853 7712
rect 1217 7506 1237 7526
rect 1036 7464 1056 7484
rect 1757 7505 1777 7525
rect 1598 7452 1619 7471
rect 1812 7453 1832 7473
rect 3425 8087 3445 8107
rect 3647 8085 3667 8105
rect 3480 8035 3500 8055
rect 4020 8034 4040 8054
rect 2628 7859 2648 7879
rect 2840 7864 2859 7882
rect 2683 7807 2703 7827
rect 3404 7848 3424 7868
rect 3223 7806 3243 7826
rect 2607 7620 2627 7640
rect 3426 7675 3446 7695
rect 3639 7677 3659 7697
rect 3481 7623 3501 7643
rect 4021 7622 4041 7642
rect 420 7278 440 7298
rect 960 7277 980 7297
rect 793 7227 813 7247
rect 1015 7225 1035 7245
rect 2529 7449 2549 7469
rect 2740 7456 2759 7473
rect 2584 7397 2604 7417
rect 3405 7436 3425 7456
rect 3124 7396 3144 7416
rect 2508 7210 2528 7230
rect 1553 7135 1577 7157
rect 2866 7157 2890 7179
rect 1915 7084 1935 7104
rect 1299 6898 1319 6918
rect 1018 6858 1038 6878
rect 1839 6897 1859 6917
rect 1682 6845 1703 6864
rect 1894 6845 1914 6865
rect 3408 7069 3428 7089
rect 3630 7067 3650 7087
rect 3463 7017 3483 7037
rect 4003 7016 4023 7036
rect 402 6672 422 6692
rect 942 6671 962 6691
rect 784 6617 804 6637
rect 997 6619 1017 6639
rect 1816 6674 1836 6694
rect 1200 6488 1220 6508
rect 1019 6446 1039 6466
rect 1740 6487 1760 6507
rect 1584 6432 1603 6450
rect 1795 6435 1815 6455
rect 403 6260 423 6280
rect 943 6259 963 6279
rect 776 6209 796 6229
rect 998 6207 1018 6227
rect 2611 6841 2631 6861
rect 2824 6843 2845 6862
rect 2666 6789 2686 6809
rect 3387 6830 3407 6850
rect 3206 6788 3226 6808
rect 2431 6690 2453 6708
rect 2590 6602 2610 6622
rect 3409 6657 3429 6677
rect 3622 6659 3642 6679
rect 3464 6605 3484 6625
rect 4004 6604 4024 6624
rect 2232 6494 2256 6516
rect 1934 6368 1955 6387
rect 1536 6117 1560 6139
rect 1961 6064 1981 6084
rect 1345 5878 1365 5898
rect 998 5840 1018 5860
rect 1885 5877 1905 5897
rect 1729 5824 1747 5842
rect 1940 5825 1960 5845
rect 382 5654 402 5674
rect 922 5653 942 5673
rect 764 5599 784 5619
rect 977 5601 997 5621
rect 1796 5656 1816 5676
rect 1180 5470 1200 5490
rect 999 5428 1019 5448
rect 1720 5469 1740 5489
rect 1561 5416 1582 5435
rect 1775 5417 1795 5437
rect 383 5242 403 5262
rect 923 5241 943 5261
rect 756 5191 776 5211
rect 978 5189 998 5209
rect 1516 5099 1540 5121
rect 1878 5048 1898 5068
rect 1262 4862 1282 4882
rect 981 4822 1001 4842
rect 1802 4861 1822 4881
rect 1647 4805 1666 4822
rect 1857 4809 1877 4829
rect 365 4636 385 4656
rect 905 4635 925 4655
rect 747 4581 767 4601
rect 960 4583 980 4603
rect 1959 4738 1981 4756
rect 1779 4638 1799 4658
rect 1163 4452 1183 4472
rect 982 4410 1002 4430
rect 1703 4451 1723 4471
rect 1547 4396 1566 4414
rect 1758 4399 1778 4419
rect 366 4224 386 4244
rect 906 4223 926 4243
rect 739 4173 759 4193
rect 961 4171 981 4191
rect 2446 6433 2466 6453
rect 2657 6431 2680 6453
rect 2501 6381 2521 6401
rect 3388 6418 3408 6438
rect 3041 6380 3061 6400
rect 2425 6194 2445 6214
rect 2846 6139 2870 6161
rect 2451 5891 2472 5910
rect 3388 6051 3408 6071
rect 3610 6049 3630 6069
rect 3443 5999 3463 6019
rect 3983 5998 4003 6018
rect 2591 5823 2611 5843
rect 2803 5828 2822 5846
rect 2646 5771 2666 5791
rect 3367 5812 3387 5832
rect 3186 5770 3206 5790
rect 2570 5584 2590 5604
rect 3389 5639 3409 5659
rect 3602 5641 3622 5661
rect 3444 5587 3464 5607
rect 3984 5586 4004 5606
rect 2492 5413 2512 5433
rect 2703 5414 2724 5433
rect 2547 5361 2567 5381
rect 3368 5400 3388 5420
rect 3087 5360 3107 5380
rect 2471 5174 2491 5194
rect 2829 5121 2853 5143
rect 3371 5033 3391 5053
rect 3593 5031 3613 5051
rect 3426 4981 3446 5001
rect 3966 4980 3986 5000
rect 2574 4805 2594 4825
rect 2787 4807 2808 4826
rect 2629 4753 2649 4773
rect 3350 4794 3370 4814
rect 3169 4752 3189 4772
rect 2553 4566 2573 4586
rect 3372 4621 3392 4641
rect 3585 4623 3605 4643
rect 3427 4569 3447 4589
rect 3967 4568 3987 4588
rect 1897 4332 1918 4351
rect 2270 4399 2290 4419
rect 2482 4398 2508 4424
rect 2325 4347 2345 4367
rect 3351 4382 3371 4402
rect 2865 4346 2885 4366
rect 2249 4160 2269 4180
rect 1499 4081 1523 4103
rect 2810 4103 2834 4125
rect 2064 4026 2084 4046
rect 1448 3840 1468 3860
rect 962 3804 982 3824
rect 1988 3839 2008 3859
rect 1826 3776 1849 3799
rect 2043 3787 2063 3807
rect 2415 3855 2436 3874
rect 346 3618 366 3638
rect 886 3617 906 3637
rect 728 3563 748 3583
rect 941 3565 961 3585
rect 1760 3620 1780 3640
rect 1144 3434 1164 3454
rect 963 3392 983 3412
rect 1684 3433 1704 3453
rect 1525 3380 1546 3399
rect 1739 3381 1759 3401
rect 347 3206 367 3226
rect 887 3205 907 3225
rect 720 3155 740 3175
rect 942 3153 962 3173
rect 1480 3063 1504 3085
rect 1842 3012 1862 3032
rect 1226 2826 1246 2846
rect 945 2786 965 2806
rect 1766 2825 1786 2845
rect 1609 2773 1630 2792
rect 1821 2773 1841 2793
rect 329 2600 349 2620
rect 869 2599 889 2619
rect 711 2545 731 2565
rect 924 2547 944 2567
rect 1743 2602 1763 2622
rect 1127 2416 1147 2436
rect 946 2374 966 2394
rect 1667 2415 1687 2435
rect 1511 2360 1530 2378
rect 1722 2363 1742 2383
rect 330 2188 350 2208
rect 870 2187 890 2207
rect 703 2137 723 2157
rect 925 2135 945 2155
rect 1861 2296 1882 2315
rect 1463 2045 1487 2067
rect 1888 1992 1908 2012
rect 1272 1806 1292 1826
rect 925 1768 945 1788
rect 1812 1805 1832 1825
rect 1653 1753 1676 1775
rect 1867 1753 1887 1773
rect 3352 4015 3372 4035
rect 3574 4013 3594 4033
rect 3407 3963 3427 3983
rect 3947 3962 3967 3982
rect 2555 3787 2575 3807
rect 2767 3792 2786 3810
rect 2610 3735 2630 3755
rect 3331 3776 3351 3796
rect 3150 3734 3170 3754
rect 2534 3548 2554 3568
rect 2352 3450 2374 3468
rect 3353 3603 3373 3623
rect 3566 3605 3586 3625
rect 3408 3551 3428 3571
rect 3948 3550 3968 3570
rect 2456 3377 2476 3397
rect 2667 3384 2686 3401
rect 2511 3325 2531 3345
rect 3332 3364 3352 3384
rect 3051 3324 3071 3344
rect 2435 3138 2455 3158
rect 2793 3085 2817 3107
rect 3335 2997 3355 3017
rect 3557 2995 3577 3015
rect 3390 2945 3410 2965
rect 3930 2944 3950 2964
rect 2538 2769 2558 2789
rect 2751 2771 2772 2790
rect 2593 2717 2613 2737
rect 3314 2758 3334 2778
rect 3133 2716 3153 2736
rect 2517 2530 2537 2550
rect 3336 2585 3356 2605
rect 3549 2587 3569 2607
rect 3391 2533 3411 2553
rect 3931 2532 3951 2552
rect 2373 2361 2393 2381
rect 2586 2364 2604 2382
rect 2428 2309 2448 2329
rect 3315 2346 3335 2366
rect 2968 2308 2988 2328
rect 2352 2122 2372 2142
rect 2773 2067 2797 2089
rect 2378 1819 2399 1838
rect 2077 1690 2101 1712
rect 309 1582 329 1602
rect 849 1581 869 1601
rect 691 1527 711 1547
rect 904 1529 924 1549
rect 1723 1584 1743 1604
rect 1880 1498 1902 1516
rect 1107 1398 1127 1418
rect 926 1356 946 1376
rect 1647 1397 1667 1417
rect 1488 1344 1509 1363
rect 1702 1345 1722 1365
rect 3315 1979 3335 1999
rect 3537 1977 3557 1997
rect 3370 1927 3390 1947
rect 3910 1926 3930 1946
rect 2518 1751 2538 1771
rect 2730 1756 2749 1774
rect 2573 1699 2593 1719
rect 3294 1740 3314 1760
rect 3113 1698 3133 1718
rect 2497 1512 2517 1532
rect 3316 1567 3336 1587
rect 3529 1569 3549 1589
rect 3371 1515 3391 1535
rect 3911 1514 3931 1534
rect 310 1170 330 1190
rect 850 1169 870 1189
rect 683 1119 703 1139
rect 905 1117 925 1137
rect 2419 1341 2439 1361
rect 2630 1342 2651 1361
rect 2474 1289 2494 1309
rect 3295 1328 3315 1348
rect 3014 1288 3034 1308
rect 2398 1102 2418 1122
rect 1443 1027 1467 1049
rect 2756 1049 2780 1071
rect 1805 976 1825 996
rect 1189 790 1209 810
rect 908 750 928 770
rect 1729 789 1749 809
rect 1574 733 1593 750
rect 1784 737 1804 757
rect 3298 961 3318 981
rect 3520 959 3540 979
rect 3353 909 3373 929
rect 3893 908 3913 928
rect 292 564 312 584
rect 832 563 852 583
rect 674 509 694 529
rect 887 511 907 531
rect 1706 566 1726 586
rect 1090 380 1110 400
rect 909 338 929 358
rect 1630 379 1650 399
rect 1474 324 1493 342
rect 1685 327 1705 347
rect 293 152 313 172
rect 833 151 853 171
rect 666 101 686 121
rect 888 99 908 119
rect 2501 733 2521 753
rect 2714 735 2735 754
rect 2556 681 2576 701
rect 3277 722 3297 742
rect 3096 680 3116 700
rect 2480 494 2500 514
rect 3299 549 3319 569
rect 3512 551 3532 571
rect 3354 497 3374 517
rect 3894 496 3914 516
rect 3278 310 3298 330
rect 1824 260 1845 279
rect 4047 47 4079 72
rect 1426 9 1450 31
rect 506 -43 542 -16
rect 2122 -239 2143 -218
rect 2204 -332 2224 -312
rect 1506 -424 1526 -404
rect 2046 -425 2066 -405
rect 2101 -477 2121 -457
<< metal1 >>
rect 3387 8205 3673 8206
rect 2872 8197 3675 8205
rect 2872 8180 2883 8197
rect 2873 8175 2883 8180
rect 2907 8180 3675 8197
rect 2907 8175 2912 8180
rect 2873 8162 2912 8175
rect 3417 8114 3452 8115
rect 3396 8107 3452 8114
rect 3396 8087 3425 8107
rect 3445 8087 3452 8107
rect 3396 8082 3452 8087
rect 3636 8105 3675 8180
rect 3636 8085 3647 8105
rect 3667 8085 3675 8105
rect 2480 7946 2862 7951
rect 2480 7927 2488 7946
rect 2509 7927 2862 7946
rect 2480 7919 2862 7927
rect 1031 7901 1063 7902
rect 1028 7896 1063 7901
rect 1028 7876 1035 7896
rect 1055 7876 1063 7896
rect 2833 7889 2862 7919
rect 2620 7886 2655 7887
rect 1028 7868 1063 7876
rect 410 7710 995 7718
rect 410 7690 419 7710
rect 439 7709 995 7710
rect 439 7690 959 7709
rect 410 7689 959 7690
rect 979 7689 995 7709
rect 410 7683 995 7689
rect 1029 7662 1063 7868
rect 2599 7879 2655 7886
rect 2599 7859 2628 7879
rect 2648 7859 2655 7879
rect 2599 7854 2655 7859
rect 2832 7882 2866 7889
rect 2832 7864 2840 7882
rect 2859 7864 2866 7882
rect 2832 7856 2866 7864
rect 3396 7876 3430 8082
rect 3636 8081 3675 8085
rect 3464 8055 4049 8061
rect 3464 8035 3480 8055
rect 3500 8054 4049 8055
rect 3500 8035 4020 8054
rect 3464 8034 4020 8035
rect 4040 8034 4049 8054
rect 3464 8026 4049 8034
rect 3396 7868 3431 7876
rect 793 7655 828 7662
rect 793 7635 801 7655
rect 821 7635 828 7655
rect 793 7562 828 7635
rect 1007 7657 1063 7662
rect 1007 7637 1014 7657
rect 1034 7637 1063 7657
rect 1007 7630 1063 7637
rect 1098 7764 1128 7766
rect 1827 7764 1860 7765
rect 1098 7738 1861 7764
rect 1007 7629 1042 7630
rect 1098 7563 1128 7738
rect 1827 7717 1861 7738
rect 1826 7712 1861 7717
rect 1826 7692 1833 7712
rect 1853 7692 1861 7712
rect 1826 7684 1861 7692
rect 1093 7562 1128 7563
rect 792 7535 1128 7562
rect 1098 7534 1128 7535
rect 1208 7526 1793 7534
rect 1208 7506 1217 7526
rect 1237 7525 1793 7526
rect 1237 7506 1757 7525
rect 1208 7505 1757 7506
rect 1777 7505 1793 7525
rect 1208 7499 1793 7505
rect 1032 7489 1064 7490
rect 1029 7484 1064 7489
rect 1029 7464 1036 7484
rect 1056 7464 1064 7484
rect 1827 7478 1861 7684
rect 2599 7648 2633 7854
rect 3396 7848 3404 7868
rect 3424 7848 3431 7868
rect 3396 7843 3431 7848
rect 3396 7842 3428 7843
rect 2667 7827 3252 7833
rect 2667 7807 2683 7827
rect 2703 7826 3252 7827
rect 2703 7807 3223 7826
rect 2667 7806 3223 7807
rect 3243 7806 3252 7826
rect 2667 7798 3252 7806
rect 3332 7797 3362 7798
rect 3332 7770 3668 7797
rect 3332 7769 3367 7770
rect 2599 7640 2634 7648
rect 2599 7620 2607 7640
rect 2627 7620 2634 7640
rect 2599 7615 2634 7620
rect 2599 7594 2633 7615
rect 3332 7594 3362 7769
rect 3418 7702 3453 7703
rect 2599 7568 3362 7594
rect 2600 7567 2633 7568
rect 3332 7566 3362 7568
rect 3397 7695 3453 7702
rect 3397 7675 3426 7695
rect 3446 7675 3453 7695
rect 3397 7670 3453 7675
rect 3632 7697 3667 7770
rect 3632 7677 3639 7697
rect 3659 7677 3667 7697
rect 3632 7670 3667 7677
rect 1029 7456 1064 7464
rect 411 7298 996 7306
rect 411 7278 420 7298
rect 440 7297 996 7298
rect 440 7278 960 7297
rect 411 7277 960 7278
rect 980 7277 996 7297
rect 411 7271 996 7277
rect 785 7247 824 7251
rect 1030 7250 1064 7456
rect 1593 7471 1628 7477
rect 1593 7452 1598 7471
rect 1619 7452 1628 7471
rect 1593 7443 1628 7452
rect 1805 7473 1861 7478
rect 1805 7453 1812 7473
rect 1832 7453 1861 7473
rect 1805 7446 1861 7453
rect 2428 7517 2762 7545
rect 1805 7445 1840 7446
rect 1597 7375 1626 7443
rect 1597 7341 1943 7375
rect 785 7227 793 7247
rect 813 7227 824 7247
rect 785 7152 824 7227
rect 1008 7245 1064 7250
rect 1008 7225 1015 7245
rect 1035 7225 1064 7245
rect 1008 7218 1064 7225
rect 1008 7217 1043 7218
rect 1548 7157 1587 7170
rect 1548 7152 1553 7157
rect 785 7135 1553 7152
rect 1577 7152 1587 7157
rect 1577 7135 1588 7152
rect 785 7127 1588 7135
rect 787 7126 1073 7127
rect 1904 7104 1943 7341
rect 1904 7092 1915 7104
rect 1908 7084 1915 7092
rect 1935 7084 1943 7104
rect 1908 7076 1943 7084
rect 1290 6918 1875 6926
rect 1290 6898 1299 6918
rect 1319 6917 1875 6918
rect 1319 6898 1839 6917
rect 1290 6897 1839 6898
rect 1859 6897 1875 6917
rect 1290 6891 1875 6897
rect 1014 6883 1046 6884
rect 1011 6878 1046 6883
rect 1011 6858 1018 6878
rect 1038 6858 1046 6878
rect 1909 6870 1943 7076
rect 1011 6850 1046 6858
rect 393 6692 978 6700
rect 393 6672 402 6692
rect 422 6691 978 6692
rect 422 6672 942 6691
rect 393 6671 942 6672
rect 962 6671 978 6691
rect 393 6665 978 6671
rect 1012 6644 1046 6850
rect 1677 6864 1708 6870
rect 1677 6845 1682 6864
rect 1703 6845 1708 6864
rect 1677 6803 1708 6845
rect 1887 6865 1943 6870
rect 1887 6845 1894 6865
rect 1914 6845 1943 6865
rect 1887 6838 1943 6845
rect 1887 6837 1922 6838
rect 1677 6775 2016 6803
rect 776 6637 811 6644
rect 776 6617 784 6637
rect 804 6617 811 6637
rect 776 6544 811 6617
rect 990 6639 1046 6644
rect 990 6619 997 6639
rect 1017 6619 1046 6639
rect 990 6612 1046 6619
rect 1081 6746 1111 6748
rect 1810 6746 1843 6747
rect 1081 6720 1844 6746
rect 990 6611 1025 6612
rect 1081 6545 1111 6720
rect 1810 6699 1844 6720
rect 1809 6694 1844 6699
rect 1809 6674 1816 6694
rect 1836 6674 1844 6694
rect 1809 6666 1844 6674
rect 1076 6544 1111 6545
rect 775 6517 1111 6544
rect 1081 6516 1111 6517
rect 1191 6508 1776 6516
rect 1191 6488 1200 6508
rect 1220 6507 1776 6508
rect 1220 6488 1740 6507
rect 1191 6487 1740 6488
rect 1760 6487 1776 6507
rect 1191 6481 1776 6487
rect 1015 6471 1047 6472
rect 1012 6466 1047 6471
rect 1012 6446 1019 6466
rect 1039 6446 1047 6466
rect 1810 6460 1844 6666
rect 1012 6438 1047 6446
rect 394 6280 979 6288
rect 394 6260 403 6280
rect 423 6279 979 6280
rect 423 6260 943 6279
rect 394 6259 943 6260
rect 963 6259 979 6279
rect 394 6253 979 6259
rect 768 6229 807 6233
rect 1013 6232 1047 6438
rect 1577 6450 1611 6458
rect 1577 6432 1584 6450
rect 1603 6432 1611 6450
rect 1577 6425 1611 6432
rect 1788 6455 1844 6460
rect 1788 6435 1795 6455
rect 1815 6435 1844 6455
rect 1788 6428 1844 6435
rect 1788 6427 1823 6428
rect 1581 6395 1610 6425
rect 1581 6387 1963 6395
rect 1581 6368 1934 6387
rect 1955 6368 1963 6387
rect 1581 6363 1963 6368
rect 768 6209 776 6229
rect 796 6209 807 6229
rect 768 6134 807 6209
rect 991 6227 1047 6232
rect 991 6207 998 6227
rect 1018 6207 1047 6227
rect 991 6200 1047 6207
rect 991 6199 1026 6200
rect 1531 6139 1570 6152
rect 1531 6134 1536 6139
rect 768 6117 1536 6134
rect 1560 6134 1570 6139
rect 1560 6117 1571 6134
rect 768 6109 1571 6117
rect 770 6108 1056 6109
rect 1987 6090 2016 6775
rect 2428 6708 2460 7517
rect 2736 7482 2762 7517
rect 2521 7476 2556 7477
rect 2500 7469 2556 7476
rect 2500 7449 2529 7469
rect 2549 7449 2556 7469
rect 2500 7444 2556 7449
rect 2732 7473 2768 7482
rect 2732 7456 2740 7473
rect 2759 7456 2768 7473
rect 2732 7447 2768 7456
rect 3397 7464 3431 7670
rect 3465 7643 4050 7649
rect 3465 7623 3481 7643
rect 3501 7642 4050 7643
rect 3501 7623 4021 7642
rect 3465 7622 4021 7623
rect 4041 7622 4050 7642
rect 3465 7614 4050 7622
rect 3397 7456 3432 7464
rect 2500 7238 2534 7444
rect 3397 7436 3405 7456
rect 3425 7436 3432 7456
rect 3397 7431 3432 7436
rect 3397 7430 3429 7431
rect 2568 7417 3153 7423
rect 2568 7397 2584 7417
rect 2604 7416 3153 7417
rect 2604 7397 3124 7416
rect 2568 7396 3124 7397
rect 3144 7396 3153 7416
rect 2568 7388 3153 7396
rect 2500 7230 2535 7238
rect 2500 7210 2508 7230
rect 2528 7222 2535 7230
rect 2528 7210 2539 7222
rect 2500 6973 2539 7210
rect 3370 7187 3656 7188
rect 2855 7179 3658 7187
rect 2855 7162 2866 7179
rect 2856 7157 2866 7162
rect 2890 7162 3658 7179
rect 2890 7157 2895 7162
rect 2856 7144 2895 7157
rect 3400 7096 3435 7097
rect 3379 7089 3435 7096
rect 3379 7069 3408 7089
rect 3428 7069 3435 7089
rect 3379 7064 3435 7069
rect 3619 7087 3658 7162
rect 3619 7067 3630 7087
rect 3650 7067 3658 7087
rect 2500 6939 2846 6973
rect 2817 6871 2846 6939
rect 2603 6868 2638 6869
rect 2428 6690 2431 6708
rect 2453 6690 2460 6708
rect 2428 6678 2460 6690
rect 2582 6861 2638 6868
rect 2582 6841 2611 6861
rect 2631 6841 2638 6861
rect 2582 6836 2638 6841
rect 2815 6862 2850 6871
rect 2815 6843 2824 6862
rect 2845 6843 2850 6862
rect 2815 6837 2850 6843
rect 3379 6858 3413 7064
rect 3619 7063 3658 7067
rect 3447 7037 4032 7043
rect 3447 7017 3463 7037
rect 3483 7036 4032 7037
rect 3483 7017 4003 7036
rect 3447 7016 4003 7017
rect 4023 7016 4032 7036
rect 3447 7008 4032 7016
rect 3379 6850 3414 6858
rect 2582 6630 2616 6836
rect 3379 6830 3387 6850
rect 3407 6830 3414 6850
rect 3379 6825 3414 6830
rect 3379 6824 3411 6825
rect 2650 6809 3235 6815
rect 2650 6789 2666 6809
rect 2686 6808 3235 6809
rect 2686 6789 3206 6808
rect 2650 6788 3206 6789
rect 3226 6788 3235 6808
rect 2650 6780 3235 6788
rect 3315 6779 3345 6780
rect 3315 6752 3651 6779
rect 3315 6751 3350 6752
rect 2582 6622 2617 6630
rect 2582 6602 2590 6622
rect 2610 6602 2617 6622
rect 2582 6597 2617 6602
rect 2582 6576 2616 6597
rect 3315 6576 3345 6751
rect 3401 6684 3436 6685
rect 2582 6550 3345 6576
rect 2583 6549 2616 6550
rect 3315 6548 3345 6550
rect 3380 6677 3436 6684
rect 3380 6657 3409 6677
rect 3429 6657 3436 6677
rect 3380 6652 3436 6657
rect 3615 6679 3650 6752
rect 3615 6659 3622 6679
rect 3642 6659 3650 6679
rect 3615 6652 3650 6659
rect 2220 6516 2683 6524
rect 2220 6494 2232 6516
rect 2256 6494 2683 6516
rect 2220 6493 2683 6494
rect 2222 6481 2261 6493
rect 2656 6462 2683 6493
rect 2438 6460 2473 6461
rect 2417 6453 2473 6460
rect 2417 6433 2446 6453
rect 2466 6433 2473 6453
rect 2417 6428 2473 6433
rect 2652 6453 2685 6462
rect 2652 6431 2657 6453
rect 2680 6431 2685 6453
rect 2417 6222 2451 6428
rect 2652 6425 2685 6431
rect 3380 6446 3414 6652
rect 3448 6625 4033 6631
rect 3448 6605 3464 6625
rect 3484 6624 4033 6625
rect 3484 6605 4004 6624
rect 3448 6604 4004 6605
rect 4024 6604 4033 6624
rect 3448 6596 4033 6604
rect 3380 6438 3415 6446
rect 3380 6418 3388 6438
rect 3408 6418 3415 6438
rect 3380 6413 3415 6418
rect 3380 6412 3412 6413
rect 2485 6401 3070 6407
rect 2485 6381 2501 6401
rect 2521 6400 3070 6401
rect 2521 6381 3041 6400
rect 2485 6380 3041 6381
rect 3061 6380 3070 6400
rect 2485 6372 3070 6380
rect 2417 6221 2452 6222
rect 2385 6214 2452 6221
rect 2385 6194 2425 6214
rect 2445 6194 2452 6214
rect 2385 6191 2452 6194
rect 2385 6188 2450 6191
rect 1956 6087 2021 6090
rect 1954 6084 2021 6087
rect 1954 6064 1961 6084
rect 1981 6064 2021 6084
rect 1954 6057 2021 6064
rect 1954 6056 1989 6057
rect 1336 5898 1921 5906
rect 1336 5878 1345 5898
rect 1365 5897 1921 5898
rect 1365 5878 1885 5897
rect 1336 5877 1885 5878
rect 1905 5877 1921 5897
rect 1336 5871 1921 5877
rect 994 5865 1026 5866
rect 991 5860 1026 5865
rect 991 5840 998 5860
rect 1018 5840 1026 5860
rect 991 5832 1026 5840
rect 373 5674 958 5682
rect 373 5654 382 5674
rect 402 5673 958 5674
rect 402 5654 922 5673
rect 373 5653 922 5654
rect 942 5653 958 5673
rect 373 5647 958 5653
rect 992 5626 1026 5832
rect 1719 5842 1760 5853
rect 1955 5850 1989 6056
rect 1719 5824 1729 5842
rect 1747 5824 1760 5842
rect 1719 5816 1760 5824
rect 1933 5845 1989 5850
rect 1933 5825 1940 5845
rect 1960 5825 1989 5845
rect 1933 5818 1989 5825
rect 1933 5817 1968 5818
rect 1728 5786 1754 5816
rect 1728 5785 2066 5786
rect 1728 5749 2082 5785
rect 756 5619 791 5626
rect 756 5599 764 5619
rect 784 5599 791 5619
rect 756 5526 791 5599
rect 970 5621 1026 5626
rect 970 5601 977 5621
rect 997 5601 1026 5621
rect 970 5594 1026 5601
rect 1061 5728 1091 5730
rect 1790 5728 1823 5729
rect 1061 5702 1824 5728
rect 970 5593 1005 5594
rect 1061 5527 1091 5702
rect 1790 5681 1824 5702
rect 1789 5676 1824 5681
rect 1789 5656 1796 5676
rect 1816 5656 1824 5676
rect 1789 5648 1824 5656
rect 1056 5526 1091 5527
rect 755 5499 1091 5526
rect 1061 5498 1091 5499
rect 1171 5490 1756 5498
rect 1171 5470 1180 5490
rect 1200 5489 1756 5490
rect 1200 5470 1720 5489
rect 1171 5469 1720 5470
rect 1740 5469 1756 5489
rect 1171 5463 1756 5469
rect 995 5453 1027 5454
rect 992 5448 1027 5453
rect 992 5428 999 5448
rect 1019 5428 1027 5448
rect 1790 5442 1824 5648
rect 992 5420 1027 5428
rect 374 5262 959 5270
rect 374 5242 383 5262
rect 403 5261 959 5262
rect 403 5242 923 5261
rect 374 5241 923 5242
rect 943 5241 959 5261
rect 374 5235 959 5241
rect 748 5211 787 5215
rect 993 5214 1027 5420
rect 1556 5435 1591 5441
rect 1556 5416 1561 5435
rect 1582 5416 1591 5435
rect 1556 5407 1591 5416
rect 1768 5437 1824 5442
rect 1768 5417 1775 5437
rect 1795 5417 1824 5437
rect 1768 5410 1824 5417
rect 1768 5409 1803 5410
rect 1560 5339 1589 5407
rect 1560 5305 1906 5339
rect 748 5191 756 5211
rect 776 5191 787 5211
rect 748 5116 787 5191
rect 971 5209 1027 5214
rect 971 5189 978 5209
rect 998 5189 1027 5209
rect 971 5182 1027 5189
rect 971 5181 1006 5182
rect 1511 5121 1550 5134
rect 1511 5116 1516 5121
rect 748 5099 1516 5116
rect 1540 5116 1550 5121
rect 1540 5099 1551 5116
rect 748 5091 1551 5099
rect 750 5090 1036 5091
rect 1867 5068 1906 5305
rect 1867 5056 1878 5068
rect 1871 5048 1878 5056
rect 1898 5048 1906 5068
rect 1871 5040 1906 5048
rect 1253 4882 1838 4890
rect 1253 4862 1262 4882
rect 1282 4881 1838 4882
rect 1282 4862 1802 4881
rect 1253 4861 1802 4862
rect 1822 4861 1838 4881
rect 1253 4855 1838 4861
rect 977 4847 1009 4848
rect 974 4842 1009 4847
rect 974 4822 981 4842
rect 1001 4822 1009 4842
rect 1872 4834 1906 5040
rect 974 4814 1009 4822
rect 356 4656 941 4664
rect 356 4636 365 4656
rect 385 4655 941 4656
rect 385 4636 905 4655
rect 356 4635 905 4636
rect 925 4635 941 4655
rect 356 4629 941 4635
rect 975 4608 1009 4814
rect 1638 4822 1674 4831
rect 1638 4805 1647 4822
rect 1666 4805 1674 4822
rect 1638 4796 1674 4805
rect 1850 4829 1906 4834
rect 1850 4809 1857 4829
rect 1877 4809 1906 4829
rect 1850 4802 1906 4809
rect 1850 4801 1885 4802
rect 1644 4761 1670 4796
rect 1952 4761 1984 4762
rect 1644 4756 1984 4761
rect 1644 4738 1959 4756
rect 1981 4738 1984 4756
rect 1644 4733 1984 4738
rect 1952 4732 1984 4733
rect 739 4601 774 4608
rect 739 4581 747 4601
rect 767 4581 774 4601
rect 739 4508 774 4581
rect 953 4603 1009 4608
rect 953 4583 960 4603
rect 980 4583 1009 4603
rect 953 4576 1009 4583
rect 1044 4710 1074 4712
rect 1773 4710 1806 4711
rect 1044 4684 1807 4710
rect 953 4575 988 4576
rect 1044 4509 1074 4684
rect 1773 4663 1807 4684
rect 1772 4658 1807 4663
rect 1772 4638 1779 4658
rect 1799 4638 1807 4658
rect 1772 4630 1807 4638
rect 1039 4508 1074 4509
rect 738 4481 1074 4508
rect 1044 4480 1074 4481
rect 1154 4472 1739 4480
rect 1154 4452 1163 4472
rect 1183 4471 1739 4472
rect 1183 4452 1703 4471
rect 1154 4451 1703 4452
rect 1723 4451 1739 4471
rect 1154 4445 1739 4451
rect 978 4435 1010 4436
rect 975 4430 1010 4435
rect 975 4410 982 4430
rect 1002 4410 1010 4430
rect 1773 4424 1807 4630
rect 975 4402 1010 4410
rect 357 4244 942 4252
rect 357 4224 366 4244
rect 386 4243 942 4244
rect 386 4224 906 4243
rect 357 4223 906 4224
rect 926 4223 942 4243
rect 357 4217 942 4223
rect 731 4193 770 4197
rect 976 4196 1010 4402
rect 1540 4414 1574 4422
rect 1540 4396 1547 4414
rect 1566 4396 1574 4414
rect 1540 4389 1574 4396
rect 1751 4419 1807 4424
rect 1751 4399 1758 4419
rect 1778 4399 1807 4419
rect 1751 4392 1807 4399
rect 1751 4391 1786 4392
rect 1544 4359 1573 4389
rect 1544 4351 1926 4359
rect 1544 4332 1897 4351
rect 1918 4332 1926 4351
rect 1544 4327 1926 4332
rect 731 4173 739 4193
rect 759 4173 770 4193
rect 731 4098 770 4173
rect 954 4191 1010 4196
rect 954 4171 961 4191
rect 981 4171 1010 4191
rect 954 4164 1010 4171
rect 954 4163 989 4164
rect 1494 4103 1533 4116
rect 1494 4098 1499 4103
rect 731 4081 1499 4098
rect 1523 4098 1533 4103
rect 1523 4081 1534 4098
rect 731 4073 1534 4081
rect 733 4072 1019 4073
rect 2055 4049 2082 5749
rect 2390 5503 2419 6188
rect 3350 6169 3636 6170
rect 2835 6161 3638 6169
rect 2835 6144 2846 6161
rect 2836 6139 2846 6144
rect 2870 6144 3638 6161
rect 2870 6139 2875 6144
rect 2836 6126 2875 6139
rect 3380 6078 3415 6079
rect 3359 6071 3415 6078
rect 3359 6051 3388 6071
rect 3408 6051 3415 6071
rect 3359 6046 3415 6051
rect 3599 6069 3638 6144
rect 3599 6049 3610 6069
rect 3630 6049 3638 6069
rect 2443 5910 2825 5915
rect 2443 5891 2451 5910
rect 2472 5891 2825 5910
rect 2443 5883 2825 5891
rect 2796 5853 2825 5883
rect 2583 5850 2618 5851
rect 2562 5843 2618 5850
rect 2562 5823 2591 5843
rect 2611 5823 2618 5843
rect 2562 5818 2618 5823
rect 2795 5846 2829 5853
rect 2795 5828 2803 5846
rect 2822 5828 2829 5846
rect 2795 5820 2829 5828
rect 3359 5840 3393 6046
rect 3599 6045 3638 6049
rect 3427 6019 4012 6025
rect 3427 5999 3443 6019
rect 3463 6018 4012 6019
rect 3463 5999 3983 6018
rect 3427 5998 3983 5999
rect 4003 5998 4012 6018
rect 3427 5990 4012 5998
rect 3359 5832 3394 5840
rect 2562 5612 2596 5818
rect 3359 5812 3367 5832
rect 3387 5812 3394 5832
rect 3359 5807 3394 5812
rect 3359 5806 3391 5807
rect 2630 5791 3215 5797
rect 2630 5771 2646 5791
rect 2666 5790 3215 5791
rect 2666 5771 3186 5790
rect 2630 5770 3186 5771
rect 3206 5770 3215 5790
rect 2630 5762 3215 5770
rect 3295 5761 3325 5762
rect 3295 5734 3631 5761
rect 3295 5733 3330 5734
rect 2562 5604 2597 5612
rect 2562 5584 2570 5604
rect 2590 5584 2597 5604
rect 2562 5579 2597 5584
rect 2562 5558 2596 5579
rect 3295 5558 3325 5733
rect 3381 5666 3416 5667
rect 2562 5532 3325 5558
rect 2563 5531 2596 5532
rect 3295 5530 3325 5532
rect 3360 5659 3416 5666
rect 3360 5639 3389 5659
rect 3409 5639 3416 5659
rect 3360 5634 3416 5639
rect 3595 5661 3630 5734
rect 3595 5641 3602 5661
rect 3622 5641 3630 5661
rect 3595 5634 3630 5641
rect 2390 5475 2729 5503
rect 2484 5440 2519 5441
rect 2463 5433 2519 5440
rect 2463 5413 2492 5433
rect 2512 5413 2519 5433
rect 2463 5408 2519 5413
rect 2698 5433 2729 5475
rect 2698 5414 2703 5433
rect 2724 5414 2729 5433
rect 2698 5408 2729 5414
rect 3360 5428 3394 5634
rect 3428 5607 4013 5613
rect 3428 5587 3444 5607
rect 3464 5606 4013 5607
rect 3464 5587 3984 5606
rect 3428 5586 3984 5587
rect 4004 5586 4013 5606
rect 3428 5578 4013 5586
rect 3360 5420 3395 5428
rect 2463 5202 2497 5408
rect 3360 5400 3368 5420
rect 3388 5400 3395 5420
rect 3360 5395 3395 5400
rect 3360 5394 3392 5395
rect 2531 5381 3116 5387
rect 2531 5361 2547 5381
rect 2567 5380 3116 5381
rect 2567 5361 3087 5380
rect 2531 5360 3087 5361
rect 3107 5360 3116 5380
rect 2531 5352 3116 5360
rect 2463 5194 2498 5202
rect 2463 5174 2471 5194
rect 2491 5186 2498 5194
rect 2491 5174 2502 5186
rect 2463 4937 2502 5174
rect 3333 5151 3619 5152
rect 2818 5143 3621 5151
rect 2818 5126 2829 5143
rect 2819 5121 2829 5126
rect 2853 5126 3621 5143
rect 2853 5121 2858 5126
rect 2819 5108 2858 5121
rect 3363 5060 3398 5061
rect 3342 5053 3398 5060
rect 3342 5033 3371 5053
rect 3391 5033 3398 5053
rect 3342 5028 3398 5033
rect 3582 5051 3621 5126
rect 3582 5031 3593 5051
rect 3613 5031 3621 5051
rect 2463 4903 2809 4937
rect 2780 4835 2809 4903
rect 2566 4832 2601 4833
rect 2545 4825 2601 4832
rect 2545 4805 2574 4825
rect 2594 4805 2601 4825
rect 2545 4800 2601 4805
rect 2778 4826 2813 4835
rect 2778 4807 2787 4826
rect 2808 4807 2813 4826
rect 2778 4801 2813 4807
rect 3342 4822 3376 5028
rect 3582 5027 3621 5031
rect 3410 5001 3995 5007
rect 3410 4981 3426 5001
rect 3446 5000 3995 5001
rect 3446 4981 3966 5000
rect 3410 4980 3966 4981
rect 3986 4980 3995 5000
rect 3410 4972 3995 4980
rect 3342 4814 3377 4822
rect 2545 4594 2579 4800
rect 3342 4794 3350 4814
rect 3370 4794 3377 4814
rect 3342 4789 3377 4794
rect 3342 4788 3374 4789
rect 2613 4773 3198 4779
rect 2613 4753 2629 4773
rect 2649 4772 3198 4773
rect 2649 4753 3169 4772
rect 2613 4752 3169 4753
rect 3189 4752 3198 4772
rect 2613 4744 3198 4752
rect 3278 4743 3308 4744
rect 3278 4716 3614 4743
rect 3278 4715 3313 4716
rect 2545 4586 2580 4594
rect 2545 4566 2553 4586
rect 2573 4566 2580 4586
rect 2545 4561 2580 4566
rect 2545 4540 2579 4561
rect 3278 4540 3308 4715
rect 3364 4648 3399 4649
rect 2545 4514 3308 4540
rect 2546 4513 2579 4514
rect 3278 4512 3308 4514
rect 3343 4641 3399 4648
rect 3343 4621 3372 4641
rect 3392 4621 3399 4641
rect 3343 4616 3399 4621
rect 3578 4643 3613 4716
rect 3578 4623 3585 4643
rect 3605 4623 3613 4643
rect 3578 4616 3613 4623
rect 2197 4493 2514 4496
rect 2197 4466 2200 4493
rect 2227 4466 2514 4493
rect 2197 4460 2514 4466
rect 2197 4457 2233 4460
rect 2478 4430 2514 4460
rect 2262 4426 2297 4427
rect 2241 4419 2297 4426
rect 2241 4399 2270 4419
rect 2290 4399 2297 4419
rect 2241 4394 2297 4399
rect 2476 4424 2514 4430
rect 2476 4398 2482 4424
rect 2508 4398 2514 4424
rect 2241 4195 2275 4394
rect 2476 4390 2514 4398
rect 3343 4410 3377 4616
rect 3411 4589 3996 4595
rect 3411 4569 3427 4589
rect 3447 4588 3996 4589
rect 3447 4569 3967 4588
rect 3411 4568 3967 4569
rect 3987 4568 3996 4588
rect 3411 4560 3996 4568
rect 3343 4402 3378 4410
rect 3343 4382 3351 4402
rect 3371 4382 3378 4402
rect 3343 4377 3378 4382
rect 3343 4376 3375 4377
rect 2309 4367 2894 4373
rect 2309 4347 2325 4367
rect 2345 4366 2894 4367
rect 2345 4347 2865 4366
rect 2309 4346 2865 4347
rect 2885 4346 2894 4366
rect 2309 4338 2894 4346
rect 2241 4180 2278 4195
rect 2241 4160 2249 4180
rect 2269 4160 2278 4180
rect 2241 4157 2278 4160
rect 2055 4046 2092 4049
rect 2055 4026 2064 4046
rect 2084 4026 2092 4046
rect 2055 4011 2092 4026
rect 1439 3860 2024 3868
rect 1439 3840 1448 3860
rect 1468 3859 2024 3860
rect 1468 3840 1988 3859
rect 1439 3839 1988 3840
rect 2008 3839 2024 3859
rect 1439 3833 2024 3839
rect 958 3829 990 3830
rect 955 3824 990 3829
rect 955 3804 962 3824
rect 982 3804 990 3824
rect 2058 3812 2092 4011
rect 2036 3807 2092 3812
rect 955 3796 990 3804
rect 337 3638 922 3646
rect 337 3618 346 3638
rect 366 3637 922 3638
rect 366 3618 886 3637
rect 337 3617 886 3618
rect 906 3617 922 3637
rect 337 3611 922 3617
rect 956 3590 990 3796
rect 1818 3805 1853 3807
rect 1818 3799 1856 3805
rect 1818 3776 1826 3799
rect 1849 3776 1856 3799
rect 2036 3787 2043 3807
rect 2063 3787 2092 3807
rect 2036 3780 2092 3787
rect 2036 3779 2071 3780
rect 1818 3770 1856 3776
rect 1818 3757 1853 3770
rect 1816 3699 1853 3757
rect 720 3583 755 3590
rect 720 3563 728 3583
rect 748 3563 755 3583
rect 720 3490 755 3563
rect 934 3585 990 3590
rect 934 3565 941 3585
rect 961 3565 990 3585
rect 934 3558 990 3565
rect 1025 3692 1055 3694
rect 1754 3692 1787 3693
rect 1025 3666 1788 3692
rect 934 3557 969 3558
rect 1025 3491 1055 3666
rect 1754 3645 1788 3666
rect 1816 3682 1851 3699
rect 1816 3681 2110 3682
rect 1816 3680 2153 3681
rect 1816 3673 2158 3680
rect 1816 3647 2118 3673
rect 2149 3647 2158 3673
rect 1753 3640 1788 3645
rect 2109 3644 2158 3647
rect 1753 3620 1760 3640
rect 1780 3620 1788 3640
rect 2115 3639 2158 3644
rect 1753 3612 1788 3620
rect 1020 3490 1055 3491
rect 719 3463 1055 3490
rect 1025 3462 1055 3463
rect 1135 3454 1720 3462
rect 1135 3434 1144 3454
rect 1164 3453 1720 3454
rect 1164 3434 1684 3453
rect 1135 3433 1684 3434
rect 1704 3433 1720 3453
rect 1135 3427 1720 3433
rect 959 3417 991 3418
rect 956 3412 991 3417
rect 956 3392 963 3412
rect 983 3392 991 3412
rect 1754 3406 1788 3612
rect 956 3384 991 3392
rect 338 3226 923 3234
rect 338 3206 347 3226
rect 367 3225 923 3226
rect 367 3206 887 3225
rect 338 3205 887 3206
rect 907 3205 923 3225
rect 338 3199 923 3205
rect 712 3175 751 3179
rect 957 3178 991 3384
rect 1520 3399 1555 3405
rect 1520 3380 1525 3399
rect 1546 3380 1555 3399
rect 1520 3371 1555 3380
rect 1732 3401 1788 3406
rect 1732 3381 1739 3401
rect 1759 3381 1788 3401
rect 1732 3374 1788 3381
rect 1732 3373 1767 3374
rect 1524 3303 1553 3371
rect 1524 3269 1870 3303
rect 712 3155 720 3175
rect 740 3155 751 3175
rect 712 3080 751 3155
rect 935 3173 991 3178
rect 935 3153 942 3173
rect 962 3153 991 3173
rect 935 3146 991 3153
rect 935 3145 970 3146
rect 1475 3085 1514 3098
rect 1475 3080 1480 3085
rect 712 3063 1480 3080
rect 1504 3080 1514 3085
rect 1504 3063 1515 3080
rect 712 3055 1515 3063
rect 714 3054 1000 3055
rect 1831 3032 1870 3269
rect 1831 3020 1842 3032
rect 1835 3012 1842 3020
rect 1862 3012 1870 3032
rect 1835 3004 1870 3012
rect 1217 2846 1802 2854
rect 1217 2826 1226 2846
rect 1246 2845 1802 2846
rect 1246 2826 1766 2845
rect 1217 2825 1766 2826
rect 1786 2825 1802 2845
rect 1217 2819 1802 2825
rect 941 2811 973 2812
rect 938 2806 973 2811
rect 938 2786 945 2806
rect 965 2786 973 2806
rect 1836 2798 1870 3004
rect 938 2778 973 2786
rect 320 2620 905 2628
rect 320 2600 329 2620
rect 349 2619 905 2620
rect 349 2600 869 2619
rect 320 2599 869 2600
rect 889 2599 905 2619
rect 320 2593 905 2599
rect 939 2572 973 2778
rect 1604 2792 1635 2798
rect 1604 2773 1609 2792
rect 1630 2773 1635 2792
rect 1604 2731 1635 2773
rect 1814 2793 1870 2798
rect 1814 2773 1821 2793
rect 1841 2773 1870 2793
rect 1814 2766 1870 2773
rect 1814 2765 1849 2766
rect 1604 2703 1943 2731
rect 703 2565 738 2572
rect 703 2545 711 2565
rect 731 2545 738 2565
rect 703 2472 738 2545
rect 917 2567 973 2572
rect 917 2547 924 2567
rect 944 2547 973 2567
rect 917 2540 973 2547
rect 1008 2674 1038 2676
rect 1737 2674 1770 2675
rect 1008 2648 1771 2674
rect 917 2539 952 2540
rect 1008 2473 1038 2648
rect 1737 2627 1771 2648
rect 1736 2622 1771 2627
rect 1736 2602 1743 2622
rect 1763 2602 1771 2622
rect 1736 2594 1771 2602
rect 1003 2472 1038 2473
rect 702 2445 1038 2472
rect 1008 2444 1038 2445
rect 1118 2436 1703 2444
rect 1118 2416 1127 2436
rect 1147 2435 1703 2436
rect 1147 2416 1667 2435
rect 1118 2415 1667 2416
rect 1687 2415 1703 2435
rect 1118 2409 1703 2415
rect 942 2399 974 2400
rect 939 2394 974 2399
rect 939 2374 946 2394
rect 966 2374 974 2394
rect 1737 2388 1771 2594
rect 939 2366 974 2374
rect 321 2208 906 2216
rect 321 2188 330 2208
rect 350 2207 906 2208
rect 350 2188 870 2207
rect 321 2187 870 2188
rect 890 2187 906 2207
rect 321 2181 906 2187
rect 695 2157 734 2161
rect 940 2160 974 2366
rect 1504 2378 1538 2386
rect 1504 2360 1511 2378
rect 1530 2360 1538 2378
rect 1504 2353 1538 2360
rect 1715 2383 1771 2388
rect 1715 2363 1722 2383
rect 1742 2363 1771 2383
rect 1715 2356 1771 2363
rect 1715 2355 1750 2356
rect 1508 2323 1537 2353
rect 1508 2315 1890 2323
rect 1508 2296 1861 2315
rect 1882 2296 1890 2315
rect 1508 2291 1890 2296
rect 695 2137 703 2157
rect 723 2137 734 2157
rect 695 2062 734 2137
rect 918 2155 974 2160
rect 918 2135 925 2155
rect 945 2135 974 2155
rect 918 2128 974 2135
rect 918 2127 953 2128
rect 1458 2067 1497 2080
rect 1458 2062 1463 2067
rect 695 2045 1463 2062
rect 1487 2062 1497 2067
rect 1487 2045 1498 2062
rect 695 2037 1498 2045
rect 697 2036 983 2037
rect 1914 2018 1943 2703
rect 2251 2457 2278 4157
rect 3314 4133 3600 4134
rect 2799 4125 3602 4133
rect 2799 4108 2810 4125
rect 2800 4103 2810 4108
rect 2834 4108 3602 4125
rect 2834 4103 2839 4108
rect 2800 4090 2839 4103
rect 3344 4042 3379 4043
rect 3323 4035 3379 4042
rect 3323 4015 3352 4035
rect 3372 4015 3379 4035
rect 3323 4010 3379 4015
rect 3563 4033 3602 4108
rect 3563 4013 3574 4033
rect 3594 4013 3602 4033
rect 2407 3874 2789 3879
rect 2407 3855 2415 3874
rect 2436 3855 2789 3874
rect 2407 3847 2789 3855
rect 2760 3817 2789 3847
rect 2547 3814 2582 3815
rect 2526 3807 2582 3814
rect 2526 3787 2555 3807
rect 2575 3787 2582 3807
rect 2526 3782 2582 3787
rect 2759 3810 2793 3817
rect 2759 3792 2767 3810
rect 2786 3792 2793 3810
rect 2759 3784 2793 3792
rect 3323 3804 3357 4010
rect 3563 4009 3602 4013
rect 3391 3983 3976 3989
rect 3391 3963 3407 3983
rect 3427 3982 3976 3983
rect 3427 3963 3947 3982
rect 3391 3962 3947 3963
rect 3967 3962 3976 3982
rect 3391 3954 3976 3962
rect 3323 3796 3358 3804
rect 2526 3576 2560 3782
rect 3323 3776 3331 3796
rect 3351 3776 3358 3796
rect 3323 3771 3358 3776
rect 3323 3770 3355 3771
rect 2594 3755 3179 3761
rect 2594 3735 2610 3755
rect 2630 3754 3179 3755
rect 2630 3735 3150 3754
rect 2594 3734 3150 3735
rect 3170 3734 3179 3754
rect 2594 3726 3179 3734
rect 3259 3725 3289 3726
rect 3259 3698 3595 3725
rect 3259 3697 3294 3698
rect 2526 3568 2561 3576
rect 2526 3548 2534 3568
rect 2554 3548 2561 3568
rect 2526 3543 2561 3548
rect 2526 3522 2560 3543
rect 3259 3522 3289 3697
rect 3345 3630 3380 3631
rect 2526 3496 3289 3522
rect 2527 3495 2560 3496
rect 3259 3494 3289 3496
rect 3324 3623 3380 3630
rect 3324 3603 3353 3623
rect 3373 3603 3380 3623
rect 3324 3598 3380 3603
rect 3559 3625 3594 3698
rect 3559 3605 3566 3625
rect 3586 3605 3594 3625
rect 3559 3598 3594 3605
rect 2349 3473 2381 3474
rect 2349 3468 2689 3473
rect 2349 3450 2352 3468
rect 2374 3450 2689 3468
rect 2349 3445 2689 3450
rect 2349 3444 2381 3445
rect 2663 3410 2689 3445
rect 2448 3404 2483 3405
rect 2427 3397 2483 3404
rect 2427 3377 2456 3397
rect 2476 3377 2483 3397
rect 2427 3372 2483 3377
rect 2659 3401 2695 3410
rect 2659 3384 2667 3401
rect 2686 3384 2695 3401
rect 2659 3375 2695 3384
rect 3324 3392 3358 3598
rect 3392 3571 3977 3577
rect 3392 3551 3408 3571
rect 3428 3570 3977 3571
rect 3428 3551 3948 3570
rect 3392 3550 3948 3551
rect 3968 3550 3977 3570
rect 3392 3542 3977 3550
rect 3324 3384 3359 3392
rect 2427 3166 2461 3372
rect 3324 3364 3332 3384
rect 3352 3364 3359 3384
rect 3324 3359 3359 3364
rect 3324 3358 3356 3359
rect 2495 3345 3080 3351
rect 2495 3325 2511 3345
rect 2531 3344 3080 3345
rect 2531 3325 3051 3344
rect 2495 3324 3051 3325
rect 3071 3324 3080 3344
rect 2495 3316 3080 3324
rect 2427 3158 2462 3166
rect 2427 3138 2435 3158
rect 2455 3150 2462 3158
rect 2455 3138 2466 3150
rect 2427 2901 2466 3138
rect 3297 3115 3583 3116
rect 2782 3107 3585 3115
rect 2782 3090 2793 3107
rect 2783 3085 2793 3090
rect 2817 3090 3585 3107
rect 2817 3085 2822 3090
rect 2783 3072 2822 3085
rect 3327 3024 3362 3025
rect 3306 3017 3362 3024
rect 3306 2997 3335 3017
rect 3355 2997 3362 3017
rect 3306 2992 3362 2997
rect 3546 3015 3585 3090
rect 3546 2995 3557 3015
rect 3577 2995 3585 3015
rect 2427 2867 2773 2901
rect 2744 2799 2773 2867
rect 2530 2796 2565 2797
rect 2509 2789 2565 2796
rect 2509 2769 2538 2789
rect 2558 2769 2565 2789
rect 2509 2764 2565 2769
rect 2742 2790 2777 2799
rect 2742 2771 2751 2790
rect 2772 2771 2777 2790
rect 2742 2765 2777 2771
rect 3306 2786 3340 2992
rect 3546 2991 3585 2995
rect 3374 2965 3959 2971
rect 3374 2945 3390 2965
rect 3410 2964 3959 2965
rect 3410 2945 3930 2964
rect 3374 2944 3930 2945
rect 3950 2944 3959 2964
rect 3374 2936 3959 2944
rect 3306 2778 3341 2786
rect 2509 2558 2543 2764
rect 3306 2758 3314 2778
rect 3334 2758 3341 2778
rect 3306 2753 3341 2758
rect 3306 2752 3338 2753
rect 2577 2737 3162 2743
rect 2577 2717 2593 2737
rect 2613 2736 3162 2737
rect 2613 2717 3133 2736
rect 2577 2716 3133 2717
rect 3153 2716 3162 2736
rect 2577 2708 3162 2716
rect 3242 2707 3272 2708
rect 3242 2680 3578 2707
rect 3242 2679 3277 2680
rect 2509 2550 2544 2558
rect 2509 2530 2517 2550
rect 2537 2530 2544 2550
rect 2509 2525 2544 2530
rect 2509 2504 2543 2525
rect 3242 2504 3272 2679
rect 3328 2612 3363 2613
rect 2509 2478 3272 2504
rect 2510 2477 2543 2478
rect 3242 2476 3272 2478
rect 3307 2605 3363 2612
rect 3307 2585 3336 2605
rect 3356 2585 3363 2605
rect 3307 2580 3363 2585
rect 3542 2607 3577 2680
rect 3542 2587 3549 2607
rect 3569 2587 3577 2607
rect 3542 2580 3577 2587
rect 2251 2421 2605 2457
rect 2267 2420 2605 2421
rect 2579 2390 2605 2420
rect 2365 2388 2400 2389
rect 2344 2381 2400 2388
rect 2344 2361 2373 2381
rect 2393 2361 2400 2381
rect 2344 2356 2400 2361
rect 2573 2382 2614 2390
rect 2573 2364 2586 2382
rect 2604 2364 2614 2382
rect 2344 2150 2378 2356
rect 2573 2353 2614 2364
rect 3307 2374 3341 2580
rect 3375 2553 3960 2559
rect 3375 2533 3391 2553
rect 3411 2552 3960 2553
rect 3411 2533 3931 2552
rect 3375 2532 3931 2533
rect 3951 2532 3960 2552
rect 3375 2524 3960 2532
rect 3307 2366 3342 2374
rect 3307 2346 3315 2366
rect 3335 2346 3342 2366
rect 3307 2341 3342 2346
rect 3307 2340 3339 2341
rect 2412 2329 2997 2335
rect 2412 2309 2428 2329
rect 2448 2328 2997 2329
rect 2448 2309 2968 2328
rect 2412 2308 2968 2309
rect 2988 2308 2997 2328
rect 2412 2300 2997 2308
rect 2344 2149 2379 2150
rect 2312 2142 2379 2149
rect 2312 2122 2352 2142
rect 2372 2122 2379 2142
rect 2312 2119 2379 2122
rect 2312 2116 2377 2119
rect 1883 2015 1948 2018
rect 1881 2012 1948 2015
rect 1881 1992 1888 2012
rect 1908 1992 1948 2012
rect 1881 1985 1948 1992
rect 1881 1984 1916 1985
rect 1263 1826 1848 1834
rect 1263 1806 1272 1826
rect 1292 1825 1848 1826
rect 1292 1806 1812 1825
rect 1263 1805 1812 1806
rect 1832 1805 1848 1825
rect 1263 1799 1848 1805
rect 921 1793 953 1794
rect 918 1788 953 1793
rect 918 1768 925 1788
rect 945 1768 953 1788
rect 918 1760 953 1768
rect 300 1602 885 1610
rect 300 1582 309 1602
rect 329 1601 885 1602
rect 329 1582 849 1601
rect 300 1581 849 1582
rect 869 1581 885 1601
rect 300 1575 885 1581
rect 919 1554 953 1760
rect 1648 1775 1681 1781
rect 1882 1778 1916 1984
rect 1648 1753 1653 1775
rect 1676 1753 1681 1775
rect 1648 1744 1681 1753
rect 1860 1773 1916 1778
rect 1860 1753 1867 1773
rect 1887 1753 1916 1773
rect 1860 1746 1916 1753
rect 1860 1745 1895 1746
rect 1650 1713 1677 1744
rect 2072 1713 2111 1725
rect 1650 1712 2113 1713
rect 1650 1690 2077 1712
rect 2101 1690 2113 1712
rect 1650 1682 2113 1690
rect 683 1547 718 1554
rect 683 1527 691 1547
rect 711 1527 718 1547
rect 683 1454 718 1527
rect 897 1549 953 1554
rect 897 1529 904 1549
rect 924 1529 953 1549
rect 897 1522 953 1529
rect 988 1656 1018 1658
rect 1717 1656 1750 1657
rect 988 1630 1751 1656
rect 897 1521 932 1522
rect 988 1455 1018 1630
rect 1717 1609 1751 1630
rect 1716 1604 1751 1609
rect 1716 1584 1723 1604
rect 1743 1584 1751 1604
rect 1716 1576 1751 1584
rect 983 1454 1018 1455
rect 682 1427 1018 1454
rect 988 1426 1018 1427
rect 1098 1418 1683 1426
rect 1098 1398 1107 1418
rect 1127 1417 1683 1418
rect 1127 1398 1647 1417
rect 1098 1397 1647 1398
rect 1667 1397 1683 1417
rect 1098 1391 1683 1397
rect 922 1381 954 1382
rect 919 1376 954 1381
rect 919 1356 926 1376
rect 946 1356 954 1376
rect 1717 1370 1751 1576
rect 919 1348 954 1356
rect 301 1190 886 1198
rect 301 1170 310 1190
rect 330 1189 886 1190
rect 330 1170 850 1189
rect 301 1169 850 1170
rect 870 1169 886 1189
rect 301 1163 886 1169
rect 675 1139 714 1143
rect 920 1142 954 1348
rect 1483 1363 1518 1369
rect 1483 1344 1488 1363
rect 1509 1344 1518 1363
rect 1483 1335 1518 1344
rect 1695 1365 1751 1370
rect 1695 1345 1702 1365
rect 1722 1345 1751 1365
rect 1695 1338 1751 1345
rect 1873 1516 1905 1528
rect 1873 1498 1880 1516
rect 1902 1498 1905 1516
rect 1695 1337 1730 1338
rect 1487 1267 1516 1335
rect 1487 1233 1833 1267
rect 675 1119 683 1139
rect 703 1119 714 1139
rect 675 1044 714 1119
rect 898 1137 954 1142
rect 898 1117 905 1137
rect 925 1117 954 1137
rect 898 1110 954 1117
rect 898 1109 933 1110
rect 1438 1049 1477 1062
rect 1438 1044 1443 1049
rect 675 1027 1443 1044
rect 1467 1044 1477 1049
rect 1467 1027 1478 1044
rect 675 1019 1478 1027
rect 677 1018 963 1019
rect 1794 996 1833 1233
rect 1794 984 1805 996
rect 1798 976 1805 984
rect 1825 976 1833 996
rect 1798 968 1833 976
rect 1180 810 1765 818
rect 1180 790 1189 810
rect 1209 809 1765 810
rect 1209 790 1729 809
rect 1180 789 1729 790
rect 1749 789 1765 809
rect 1180 783 1765 789
rect 904 775 936 776
rect 901 770 936 775
rect 901 750 908 770
rect 928 750 936 770
rect 1799 762 1833 968
rect 901 742 936 750
rect 283 584 868 592
rect 283 564 292 584
rect 312 583 868 584
rect 312 564 832 583
rect 283 563 832 564
rect 852 563 868 583
rect 283 557 868 563
rect 902 536 936 742
rect 1565 750 1601 759
rect 1565 733 1574 750
rect 1593 733 1601 750
rect 1565 724 1601 733
rect 1777 757 1833 762
rect 1777 737 1784 757
rect 1804 737 1833 757
rect 1777 730 1833 737
rect 1777 729 1812 730
rect 1571 689 1597 724
rect 1873 689 1905 1498
rect 2317 1431 2346 2116
rect 3277 2097 3563 2098
rect 2762 2089 3565 2097
rect 2762 2072 2773 2089
rect 2763 2067 2773 2072
rect 2797 2072 3565 2089
rect 2797 2067 2802 2072
rect 2763 2054 2802 2067
rect 3307 2006 3342 2007
rect 3286 1999 3342 2006
rect 3286 1979 3315 1999
rect 3335 1979 3342 1999
rect 3286 1974 3342 1979
rect 3526 1997 3565 2072
rect 3526 1977 3537 1997
rect 3557 1977 3565 1997
rect 2370 1838 2752 1843
rect 2370 1819 2378 1838
rect 2399 1819 2752 1838
rect 2370 1811 2752 1819
rect 2723 1781 2752 1811
rect 2510 1778 2545 1779
rect 2489 1771 2545 1778
rect 2489 1751 2518 1771
rect 2538 1751 2545 1771
rect 2489 1746 2545 1751
rect 2722 1774 2756 1781
rect 2722 1756 2730 1774
rect 2749 1756 2756 1774
rect 2722 1748 2756 1756
rect 3286 1768 3320 1974
rect 3526 1973 3565 1977
rect 3354 1947 3939 1953
rect 3354 1927 3370 1947
rect 3390 1946 3939 1947
rect 3390 1927 3910 1946
rect 3354 1926 3910 1927
rect 3930 1926 3939 1946
rect 3354 1918 3939 1926
rect 3286 1760 3321 1768
rect 2489 1540 2523 1746
rect 3286 1740 3294 1760
rect 3314 1740 3321 1760
rect 3286 1735 3321 1740
rect 3286 1734 3318 1735
rect 2557 1719 3142 1725
rect 2557 1699 2573 1719
rect 2593 1718 3142 1719
rect 2593 1699 3113 1718
rect 2557 1698 3113 1699
rect 3133 1698 3142 1718
rect 2557 1690 3142 1698
rect 3222 1689 3252 1690
rect 3222 1662 3558 1689
rect 3222 1661 3257 1662
rect 2489 1532 2524 1540
rect 2489 1512 2497 1532
rect 2517 1512 2524 1532
rect 2489 1507 2524 1512
rect 2489 1486 2523 1507
rect 3222 1486 3252 1661
rect 3308 1594 3343 1595
rect 2489 1460 3252 1486
rect 2490 1459 2523 1460
rect 3222 1458 3252 1460
rect 3287 1587 3343 1594
rect 3287 1567 3316 1587
rect 3336 1567 3343 1587
rect 3287 1562 3343 1567
rect 3522 1589 3557 1662
rect 3522 1569 3529 1589
rect 3549 1569 3557 1589
rect 3522 1562 3557 1569
rect 2317 1403 2656 1431
rect 2411 1368 2446 1369
rect 2390 1361 2446 1368
rect 2390 1341 2419 1361
rect 2439 1341 2446 1361
rect 2390 1336 2446 1341
rect 2625 1361 2656 1403
rect 2625 1342 2630 1361
rect 2651 1342 2656 1361
rect 2625 1336 2656 1342
rect 3287 1356 3321 1562
rect 3355 1535 3940 1541
rect 3355 1515 3371 1535
rect 3391 1534 3940 1535
rect 3391 1515 3911 1534
rect 3355 1514 3911 1515
rect 3931 1514 3940 1534
rect 3355 1506 3940 1514
rect 3287 1348 3322 1356
rect 2390 1130 2424 1336
rect 3287 1328 3295 1348
rect 3315 1328 3322 1348
rect 3287 1323 3322 1328
rect 3287 1322 3319 1323
rect 2458 1309 3043 1315
rect 2458 1289 2474 1309
rect 2494 1308 3043 1309
rect 2494 1289 3014 1308
rect 2458 1288 3014 1289
rect 3034 1288 3043 1308
rect 2458 1280 3043 1288
rect 2390 1122 2425 1130
rect 2390 1102 2398 1122
rect 2418 1114 2425 1122
rect 2418 1102 2429 1114
rect 2390 865 2429 1102
rect 3260 1079 3546 1080
rect 2745 1071 3548 1079
rect 2745 1054 2756 1071
rect 2746 1049 2756 1054
rect 2780 1054 3548 1071
rect 2780 1049 2785 1054
rect 2746 1036 2785 1049
rect 3290 988 3325 989
rect 3269 981 3325 988
rect 3269 961 3298 981
rect 3318 961 3325 981
rect 3269 956 3325 961
rect 3509 979 3548 1054
rect 3509 959 3520 979
rect 3540 959 3548 979
rect 2390 831 2736 865
rect 2707 763 2736 831
rect 2493 760 2528 761
rect 1571 661 1905 689
rect 2472 753 2528 760
rect 2472 733 2501 753
rect 2521 733 2528 753
rect 2472 728 2528 733
rect 2705 754 2740 763
rect 2705 735 2714 754
rect 2735 735 2740 754
rect 2705 729 2740 735
rect 3269 750 3303 956
rect 3509 955 3548 959
rect 3337 929 3922 935
rect 3337 909 3353 929
rect 3373 928 3922 929
rect 3373 909 3893 928
rect 3337 908 3893 909
rect 3913 908 3922 928
rect 3337 900 3922 908
rect 3269 742 3304 750
rect 666 529 701 536
rect 666 509 674 529
rect 694 509 701 529
rect 666 436 701 509
rect 880 531 936 536
rect 880 511 887 531
rect 907 511 936 531
rect 880 504 936 511
rect 971 638 1001 640
rect 1700 638 1733 639
rect 971 612 1734 638
rect 880 503 915 504
rect 971 437 1001 612
rect 1700 591 1734 612
rect 1699 586 1734 591
rect 1699 566 1706 586
rect 1726 566 1734 586
rect 1699 558 1734 566
rect 966 436 1001 437
rect 665 409 1001 436
rect 971 408 1001 409
rect 1081 400 1666 408
rect 1081 380 1090 400
rect 1110 399 1666 400
rect 1110 380 1630 399
rect 1081 379 1630 380
rect 1650 379 1666 399
rect 1081 373 1666 379
rect 905 363 937 364
rect 902 358 937 363
rect 902 338 909 358
rect 929 338 937 358
rect 1700 352 1734 558
rect 2472 522 2506 728
rect 3269 722 3277 742
rect 3297 722 3304 742
rect 3269 717 3304 722
rect 3269 716 3301 717
rect 2540 701 3125 707
rect 2540 681 2556 701
rect 2576 700 3125 701
rect 2576 681 3096 700
rect 2540 680 3096 681
rect 3116 680 3125 700
rect 2540 672 3125 680
rect 3205 671 3235 672
rect 3205 644 3541 671
rect 3205 643 3240 644
rect 2472 514 2507 522
rect 2472 494 2480 514
rect 2500 494 2507 514
rect 2472 489 2507 494
rect 2472 468 2506 489
rect 3205 468 3235 643
rect 3291 576 3326 577
rect 2472 442 3235 468
rect 2473 441 2506 442
rect 3205 440 3235 442
rect 3270 569 3326 576
rect 3270 549 3299 569
rect 3319 549 3326 569
rect 3270 544 3326 549
rect 3505 571 3540 644
rect 3505 551 3512 571
rect 3532 551 3540 571
rect 3505 544 3540 551
rect 902 330 937 338
rect 284 172 869 180
rect 284 152 293 172
rect 313 171 869 172
rect 313 152 833 171
rect 284 151 833 152
rect 853 151 869 171
rect 284 145 869 151
rect 658 121 697 125
rect 903 124 937 330
rect 1467 342 1501 350
rect 1467 324 1474 342
rect 1493 324 1501 342
rect 1467 317 1501 324
rect 1678 347 1734 352
rect 1678 327 1685 347
rect 1705 327 1734 347
rect 1678 320 1734 327
rect 3270 338 3304 544
rect 3338 517 3923 523
rect 3338 497 3354 517
rect 3374 516 3923 517
rect 3374 497 3894 516
rect 3338 496 3894 497
rect 3914 496 3923 516
rect 3338 488 3923 496
rect 3270 330 3305 338
rect 1678 319 1713 320
rect 1471 287 1500 317
rect 3270 310 3278 330
rect 3298 310 3305 330
rect 3270 305 3305 310
rect 3270 304 3302 305
rect 1471 279 1853 287
rect 1471 260 1824 279
rect 1845 260 1853 279
rect 1471 255 1853 260
rect 658 101 666 121
rect 686 101 697 121
rect 658 26 697 101
rect 881 119 937 124
rect 881 99 888 119
rect 908 99 937 119
rect 881 92 937 99
rect 881 91 916 92
rect 2116 44 2167 75
rect 1421 31 1460 44
rect 1421 26 1426 31
rect 658 9 1426 26
rect 1450 26 1460 31
rect 1450 9 1461 26
rect 658 1 1461 9
rect 2116 18 2133 44
rect 2161 18 2167 44
rect 660 0 946 1
rect 2116 -5 2167 18
rect 2196 50 2242 81
rect 4040 79 4083 87
rect 2196 19 2210 50
rect 2238 19 2242 50
rect 2196 12 2242 19
rect 4034 72 4089 79
rect 4034 47 4047 72
rect 4079 47 4089 72
rect 498 -16 559 -7
rect 498 -43 506 -16
rect 542 -22 559 -16
rect 600 -22 675 -18
rect 542 -24 675 -22
rect 542 -43 606 -24
rect 498 -60 606 -43
rect 651 -60 675 -24
rect 498 -62 675 -60
rect 600 -92 675 -62
rect 2129 -197 2160 -5
rect 2115 -218 2161 -197
rect 2115 -239 2122 -218
rect 2143 -239 2161 -218
rect 2115 -243 2161 -239
rect 2115 -246 2150 -243
rect 1497 -404 2082 -396
rect 1497 -424 1506 -404
rect 1526 -405 2082 -404
rect 1526 -424 2046 -405
rect 1497 -425 2046 -424
rect 2066 -425 2082 -405
rect 1497 -431 2082 -425
rect 2116 -452 2150 -246
rect 2198 -312 2232 12
rect 4034 -45 4089 47
rect 4034 -77 4045 -45
rect 4085 -77 4089 -45
rect 4034 -90 4089 -77
rect 2198 -332 2204 -312
rect 2224 -332 2232 -312
rect 2198 -338 2232 -332
rect 2094 -457 2150 -452
rect 2094 -477 2101 -457
rect 2121 -477 2150 -457
rect 2094 -484 2150 -477
rect 2094 -485 2129 -484
<< via1 >>
rect 2200 4466 2227 4493
rect 2118 3647 2149 3673
rect 2133 18 2161 44
rect 2210 19 2238 50
rect 606 -60 651 -24
rect 4045 -77 4085 -45
<< metal2 >>
rect 2195 4493 2232 4497
rect 2195 4466 2200 4493
rect 2227 4466 2232 4493
rect 2195 4456 2232 4466
rect 2110 3673 2158 3691
rect 2110 3647 2118 3673
rect 2149 3647 2158 3673
rect 2110 3615 2158 3647
rect 2118 69 2158 3615
rect 2199 1719 2225 4456
rect 2197 81 2225 1719
rect 2118 44 2164 69
rect 2118 18 2133 44
rect 2161 18 2164 44
rect 2118 -1 2164 18
rect 2196 50 2242 81
rect 2196 19 2210 50
rect 2238 19 2242 50
rect 2196 12 2242 19
rect 2122 -5 2164 -1
rect 592 -24 667 -12
rect 592 -60 606 -24
rect 651 -37 667 -24
rect 2109 -37 2203 -32
rect 651 -45 4089 -37
rect 651 -60 4045 -45
rect 592 -77 4045 -60
rect 4085 -77 4089 -45
rect 592 -86 4089 -77
rect 2109 -89 2203 -86
<< labels >>
rlabel locali 373 7692 395 7707 1 d0
rlabel locali 427 7880 456 7886 1 vdd
rlabel locali 424 7581 453 7587 1 gnd
rlabel space 530 7599 559 7608 1 gnd
rlabel nwell 562 7857 585 7860 1 vdd
rlabel locali 374 7280 396 7295 1 d0
rlabel locali 428 7468 457 7474 1 vdd
rlabel locali 425 7169 454 7175 1 gnd
rlabel space 531 7187 560 7196 1 gnd
rlabel nwell 563 7445 586 7448 1 vdd
rlabel locali 264 8125 288 8155 1 vref
rlabel locali 356 6674 378 6689 1 d0
rlabel locali 410 6862 439 6868 1 vdd
rlabel locali 407 6563 436 6569 1 gnd
rlabel space 513 6581 542 6590 1 gnd
rlabel nwell 545 6839 568 6842 1 vdd
rlabel locali 357 6262 379 6277 1 d0
rlabel locali 411 6450 440 6456 1 vdd
rlabel locali 408 6151 437 6157 1 gnd
rlabel space 514 6169 543 6178 1 gnd
rlabel nwell 546 6427 569 6430 1 vdd
rlabel locali 1225 7696 1254 7702 1 vdd
rlabel locali 1222 7397 1251 7403 1 gnd
rlabel space 1328 7415 1357 7424 1 gnd
rlabel nwell 1360 7673 1383 7676 1 vdd
rlabel locali 1165 7504 1187 7521 1 d1
rlabel locali 1208 6678 1237 6684 1 vdd
rlabel locali 1205 6379 1234 6385 1 gnd
rlabel space 1311 6397 1340 6406 1 gnd
rlabel nwell 1343 6655 1366 6658 1 vdd
rlabel locali 1148 6486 1170 6503 1 d1
rlabel locali 1307 7088 1336 7094 1 vdd
rlabel locali 1304 6789 1333 6795 1 gnd
rlabel space 1410 6807 1439 6816 1 gnd
rlabel nwell 1442 7065 1465 7068 1 vdd
rlabel locali 1249 6896 1269 6920 1 d2
rlabel locali 336 5656 358 5671 1 d0
rlabel locali 390 5844 419 5850 1 vdd
rlabel locali 387 5545 416 5551 1 gnd
rlabel space 493 5563 522 5572 1 gnd
rlabel nwell 525 5821 548 5824 1 vdd
rlabel locali 337 5244 359 5259 1 d0
rlabel locali 391 5432 420 5438 1 vdd
rlabel locali 388 5133 417 5139 1 gnd
rlabel space 494 5151 523 5160 1 gnd
rlabel nwell 526 5409 549 5412 1 vdd
rlabel locali 319 4638 341 4653 1 d0
rlabel locali 373 4826 402 4832 1 vdd
rlabel locali 370 4527 399 4533 1 gnd
rlabel space 476 4545 505 4554 1 gnd
rlabel nwell 508 4803 531 4806 1 vdd
rlabel locali 320 4226 342 4241 1 d0
rlabel locali 374 4414 403 4420 1 vdd
rlabel locali 371 4115 400 4121 1 gnd
rlabel space 477 4133 506 4142 1 gnd
rlabel nwell 509 4391 532 4394 1 vdd
rlabel locali 1188 5660 1217 5666 1 vdd
rlabel locali 1185 5361 1214 5367 1 gnd
rlabel space 1291 5379 1320 5388 1 gnd
rlabel nwell 1323 5637 1346 5640 1 vdd
rlabel locali 1128 5468 1150 5485 1 d1
rlabel locali 1171 4642 1200 4648 1 vdd
rlabel locali 1168 4343 1197 4349 1 gnd
rlabel space 1274 4361 1303 4370 1 gnd
rlabel nwell 1306 4619 1329 4622 1 vdd
rlabel locali 1111 4450 1133 4467 1 d1
rlabel locali 1270 5052 1299 5058 1 vdd
rlabel locali 1267 4753 1296 4759 1 gnd
rlabel space 1373 4771 1402 4780 1 gnd
rlabel nwell 1405 5029 1428 5032 1 vdd
rlabel locali 1212 4860 1232 4884 1 d2
rlabel locali 1353 6068 1382 6074 1 vdd
rlabel locali 1350 5769 1379 5775 1 gnd
rlabel space 1456 5787 1485 5796 1 gnd
rlabel nwell 1488 6045 1511 6048 1 vdd
rlabel locali 1297 5882 1317 5895 1 d3
rlabel locali 300 3620 322 3635 1 d0
rlabel locali 354 3808 383 3814 1 vdd
rlabel locali 351 3509 380 3515 1 gnd
rlabel space 457 3527 486 3536 1 gnd
rlabel nwell 489 3785 512 3788 1 vdd
rlabel locali 301 3208 323 3223 1 d0
rlabel locali 355 3396 384 3402 1 vdd
rlabel locali 352 3097 381 3103 1 gnd
rlabel space 458 3115 487 3124 1 gnd
rlabel nwell 490 3373 513 3376 1 vdd
rlabel locali 283 2602 305 2617 1 d0
rlabel locali 337 2790 366 2796 1 vdd
rlabel locali 334 2491 363 2497 1 gnd
rlabel space 440 2509 469 2518 1 gnd
rlabel nwell 472 2767 495 2770 1 vdd
rlabel locali 284 2190 306 2205 1 d0
rlabel locali 338 2378 367 2384 1 vdd
rlabel locali 335 2079 364 2085 1 gnd
rlabel space 441 2097 470 2106 1 gnd
rlabel nwell 473 2355 496 2358 1 vdd
rlabel locali 1152 3624 1181 3630 1 vdd
rlabel locali 1149 3325 1178 3331 1 gnd
rlabel space 1255 3343 1284 3352 1 gnd
rlabel nwell 1287 3601 1310 3604 1 vdd
rlabel locali 1092 3432 1114 3449 1 d1
rlabel locali 1135 2606 1164 2612 1 vdd
rlabel locali 1132 2307 1161 2313 1 gnd
rlabel space 1238 2325 1267 2334 1 gnd
rlabel nwell 1270 2583 1293 2586 1 vdd
rlabel locali 1075 2414 1097 2431 1 d1
rlabel locali 1234 3016 1263 3022 1 vdd
rlabel locali 1231 2717 1260 2723 1 gnd
rlabel space 1337 2735 1366 2744 1 gnd
rlabel nwell 1369 2993 1392 2996 1 vdd
rlabel locali 1176 2824 1196 2848 1 d2
rlabel locali 263 1584 285 1599 1 d0
rlabel locali 317 1772 346 1778 1 vdd
rlabel locali 314 1473 343 1479 1 gnd
rlabel space 420 1491 449 1500 1 gnd
rlabel nwell 452 1749 475 1752 1 vdd
rlabel locali 264 1172 286 1187 1 d0
rlabel locali 318 1360 347 1366 1 vdd
rlabel locali 315 1061 344 1067 1 gnd
rlabel space 421 1079 450 1088 1 gnd
rlabel nwell 453 1337 476 1340 1 vdd
rlabel locali 246 566 268 581 1 d0
rlabel locali 300 754 329 760 1 vdd
rlabel locali 297 455 326 461 1 gnd
rlabel space 403 473 432 482 1 gnd
rlabel nwell 435 731 458 734 1 vdd
rlabel locali 247 154 269 169 1 d0
rlabel locali 301 342 330 348 1 vdd
rlabel locali 298 43 327 49 1 gnd
rlabel space 404 61 433 70 1 gnd
rlabel nwell 436 319 459 322 1 vdd
rlabel locali 1115 1588 1144 1594 1 vdd
rlabel locali 1112 1289 1141 1295 1 gnd
rlabel space 1218 1307 1247 1316 1 gnd
rlabel nwell 1250 1565 1273 1568 1 vdd
rlabel locali 1055 1396 1077 1413 1 d1
rlabel locali 1098 570 1127 576 1 vdd
rlabel locali 1095 271 1124 277 1 gnd
rlabel space 1201 289 1230 298 1 gnd
rlabel nwell 1233 547 1256 550 1 vdd
rlabel locali 1038 378 1060 395 1 d1
rlabel locali 1197 980 1226 986 1 vdd
rlabel locali 1194 681 1223 687 1 gnd
rlabel space 1300 699 1329 708 1 gnd
rlabel nwell 1332 957 1355 960 1 vdd
rlabel locali 1139 788 1159 812 1 d2
rlabel locali 1280 1996 1309 2002 1 vdd
rlabel locali 1277 1697 1306 1703 1 gnd
rlabel space 1383 1715 1412 1724 1 gnd
rlabel nwell 1415 1973 1438 1976 1 vdd
rlabel locali 1224 1810 1244 1823 1 d3
rlabel locali 1456 4030 1485 4036 1 vdd
rlabel locali 1453 3731 1482 3737 1 gnd
rlabel space 1559 3749 1588 3758 1 gnd
rlabel nwell 1591 4007 1614 4010 1 vdd
rlabel locali 1402 3840 1421 3857 1 d4
rlabel locali 2912 4349 2931 4366 5 d4
rlabel nwell 2719 4196 2742 4199 5 vdd
rlabel space 2745 4448 2774 4457 5 gnd
rlabel locali 2851 4469 2880 4475 5 gnd
rlabel locali 2848 4170 2877 4176 5 vdd
rlabel locali 3089 6383 3109 6396 5 d3
rlabel nwell 2895 6230 2918 6233 5 vdd
rlabel space 2921 6482 2950 6491 5 gnd
rlabel locali 3027 6503 3056 6509 5 gnd
rlabel locali 3024 6204 3053 6210 5 vdd
rlabel locali 3174 7394 3194 7418 5 d2
rlabel nwell 2978 7246 3001 7249 5 vdd
rlabel space 3004 7498 3033 7507 5 gnd
rlabel locali 3110 7519 3139 7525 5 gnd
rlabel locali 3107 7220 3136 7226 5 vdd
rlabel locali 3273 7811 3295 7828 5 d1
rlabel nwell 3077 7656 3100 7659 5 vdd
rlabel space 3103 7908 3132 7917 5 gnd
rlabel locali 3209 7929 3238 7935 5 gnd
rlabel locali 3206 7630 3235 7636 5 vdd
rlabel locali 3256 6793 3278 6810 5 d1
rlabel nwell 3060 6638 3083 6641 5 vdd
rlabel space 3086 6890 3115 6899 5 gnd
rlabel locali 3192 6911 3221 6917 5 gnd
rlabel locali 3189 6612 3218 6618 5 vdd
rlabel locali 4192 8146 4220 8164 5 gnd
rlabel nwell 3874 7884 3897 7887 5 vdd
rlabel space 3900 8136 3929 8145 5 gnd
rlabel locali 4006 8157 4035 8163 5 gnd
rlabel locali 4003 7858 4032 7864 5 vdd
rlabel locali 4064 8037 4086 8052 5 d0
rlabel nwell 3875 7472 3898 7475 5 vdd
rlabel space 3901 7724 3930 7733 5 gnd
rlabel locali 4007 7745 4036 7751 5 gnd
rlabel locali 4004 7446 4033 7452 5 vdd
rlabel locali 4065 7625 4087 7640 5 d0
rlabel nwell 3857 6866 3880 6869 5 vdd
rlabel space 3883 7118 3912 7127 5 gnd
rlabel locali 3989 7139 4018 7145 5 gnd
rlabel locali 3986 6840 4015 6846 5 vdd
rlabel locali 4047 7019 4069 7034 5 d0
rlabel nwell 3858 6454 3881 6457 5 vdd
rlabel space 3884 6706 3913 6715 5 gnd
rlabel locali 3990 6727 4019 6733 5 gnd
rlabel locali 3987 6428 4016 6434 5 vdd
rlabel locali 4048 6607 4070 6622 5 d0
rlabel locali 3137 5358 3157 5382 5 d2
rlabel nwell 2941 5210 2964 5213 5 vdd
rlabel space 2967 5462 2996 5471 5 gnd
rlabel locali 3073 5483 3102 5489 5 gnd
rlabel locali 3070 5184 3099 5190 5 vdd
rlabel locali 3236 5775 3258 5792 5 d1
rlabel nwell 3040 5620 3063 5623 5 vdd
rlabel space 3066 5872 3095 5881 5 gnd
rlabel locali 3172 5893 3201 5899 5 gnd
rlabel locali 3169 5594 3198 5600 5 vdd
rlabel locali 3219 4757 3241 4774 5 d1
rlabel nwell 3023 4602 3046 4605 5 vdd
rlabel space 3049 4854 3078 4863 5 gnd
rlabel locali 3155 4875 3184 4881 5 gnd
rlabel locali 3152 4576 3181 4582 5 vdd
rlabel nwell 3837 5848 3860 5851 5 vdd
rlabel space 3863 6100 3892 6109 5 gnd
rlabel locali 3969 6121 3998 6127 5 gnd
rlabel locali 3966 5822 3995 5828 5 vdd
rlabel locali 4027 6001 4049 6016 5 d0
rlabel nwell 3838 5436 3861 5439 5 vdd
rlabel space 3864 5688 3893 5697 5 gnd
rlabel locali 3970 5709 3999 5715 5 gnd
rlabel locali 3967 5410 3996 5416 5 vdd
rlabel locali 4028 5589 4050 5604 5 d0
rlabel nwell 3820 4830 3843 4833 5 vdd
rlabel space 3846 5082 3875 5091 5 gnd
rlabel locali 3952 5103 3981 5109 5 gnd
rlabel locali 3949 4804 3978 4810 5 vdd
rlabel locali 4010 4983 4032 4998 5 d0
rlabel nwell 3821 4418 3844 4421 5 vdd
rlabel space 3847 4670 3876 4679 5 gnd
rlabel locali 3953 4691 3982 4697 5 gnd
rlabel locali 3950 4392 3979 4398 5 vdd
rlabel locali 4011 4571 4033 4586 5 d0
rlabel locali 3016 2311 3036 2324 5 d3
rlabel nwell 2822 2158 2845 2161 5 vdd
rlabel space 2848 2410 2877 2419 5 gnd
rlabel locali 2954 2431 2983 2437 5 gnd
rlabel locali 2951 2132 2980 2138 5 vdd
rlabel locali 3101 3322 3121 3346 5 d2
rlabel nwell 2905 3174 2928 3177 5 vdd
rlabel space 2931 3426 2960 3435 5 gnd
rlabel locali 3037 3447 3066 3453 5 gnd
rlabel locali 3034 3148 3063 3154 5 vdd
rlabel locali 3200 3739 3222 3756 5 d1
rlabel nwell 3004 3584 3027 3587 5 vdd
rlabel space 3030 3836 3059 3845 5 gnd
rlabel locali 3136 3857 3165 3863 5 gnd
rlabel locali 3133 3558 3162 3564 5 vdd
rlabel locali 3183 2721 3205 2738 5 d1
rlabel nwell 2987 2566 3010 2569 5 vdd
rlabel space 3013 2818 3042 2827 5 gnd
rlabel locali 3119 2839 3148 2845 5 gnd
rlabel locali 3116 2540 3145 2546 5 vdd
rlabel nwell 3801 3812 3824 3815 5 vdd
rlabel space 3827 4064 3856 4073 5 gnd
rlabel locali 3933 4085 3962 4091 5 gnd
rlabel locali 3930 3786 3959 3792 5 vdd
rlabel locali 3991 3965 4013 3980 5 d0
rlabel nwell 3802 3400 3825 3403 5 vdd
rlabel space 3828 3652 3857 3661 5 gnd
rlabel locali 3934 3673 3963 3679 5 gnd
rlabel locali 3931 3374 3960 3380 5 vdd
rlabel locali 3992 3553 4014 3568 5 d0
rlabel nwell 3784 2794 3807 2797 5 vdd
rlabel space 3810 3046 3839 3055 5 gnd
rlabel locali 3916 3067 3945 3073 5 gnd
rlabel locali 3913 2768 3942 2774 5 vdd
rlabel locali 3974 2947 3996 2962 5 d0
rlabel nwell 3785 2382 3808 2385 5 vdd
rlabel space 3811 2634 3840 2643 5 gnd
rlabel locali 3917 2655 3946 2661 5 gnd
rlabel locali 3914 2356 3943 2362 5 vdd
rlabel locali 3975 2535 3997 2550 5 d0
rlabel locali 3064 1286 3084 1310 5 d2
rlabel nwell 2868 1138 2891 1141 5 vdd
rlabel space 2894 1390 2923 1399 5 gnd
rlabel locali 3000 1411 3029 1417 5 gnd
rlabel locali 2997 1112 3026 1118 5 vdd
rlabel locali 3163 1703 3185 1720 5 d1
rlabel nwell 2967 1548 2990 1551 5 vdd
rlabel space 2993 1800 3022 1809 5 gnd
rlabel locali 3099 1821 3128 1827 5 gnd
rlabel locali 3096 1522 3125 1528 5 vdd
rlabel locali 3146 685 3168 702 5 d1
rlabel nwell 2950 530 2973 533 5 vdd
rlabel space 2976 782 3005 791 5 gnd
rlabel locali 3082 803 3111 809 5 gnd
rlabel locali 3079 504 3108 510 5 vdd
rlabel nwell 3764 1776 3787 1779 5 vdd
rlabel space 3790 2028 3819 2037 5 gnd
rlabel locali 3896 2049 3925 2055 5 gnd
rlabel locali 3893 1750 3922 1756 5 vdd
rlabel locali 3954 1929 3976 1944 5 d0
rlabel nwell 3765 1364 3788 1367 5 vdd
rlabel space 3791 1616 3820 1625 5 gnd
rlabel locali 3897 1637 3926 1643 5 gnd
rlabel locali 3894 1338 3923 1344 5 vdd
rlabel locali 3955 1517 3977 1532 5 d0
rlabel nwell 3747 758 3770 761 5 vdd
rlabel space 3773 1010 3802 1019 5 gnd
rlabel locali 3879 1031 3908 1037 5 gnd
rlabel locali 3876 732 3905 738 5 vdd
rlabel locali 3937 911 3959 926 5 d0
rlabel nwell 3748 346 3771 349 5 vdd
rlabel space 3774 598 3803 607 5 gnd
rlabel locali 3880 619 3909 625 5 gnd
rlabel locali 3877 320 3906 326 5 vdd
rlabel locali 3938 499 3960 514 5 d0
rlabel locali 1887 -387 1909 -372 1 vout
rlabel nwell 1649 -257 1672 -254 1 vdd
rlabel space 1617 -515 1646 -506 1 gnd
rlabel locali 1511 -533 1540 -527 1 gnd
rlabel locali 1514 -234 1543 -228 1 vdd
rlabel locali 1456 -421 1471 -408 1 d5
<< end >>

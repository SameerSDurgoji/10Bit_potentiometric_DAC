* SPICE3 file created from 9bit_DAC.ext - technology: sky130A

*.option scale=10000u

.lib "sky130_fd_pr/models/sky130.lib.spice" tt

X0 a_14463_5570# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1 a_26555_3913# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2 a_9220_5937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3 a_30648_4032# d0 a_31137_3926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X4 a_4769_2265# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X5 vdd d0 a_21008_3144# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X6 vdd d2 a_11534_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X7 vdd d0 a_34185_7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X8 a_30704_7086# d0 a_31193_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X9 a_9202_5331# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X10 a_23057_3521# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X11 a_9402_3901# a_9184_3901# a_8913_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X12 gnd d0 a_16722_2152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X13 a_30711_7304# d0 a_31192_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X14 a_6986_5378# d0 a_7783_5606# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X15 vdd d4 a_33047_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X16 a_31119_3320# d1 a_31917_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X17 a_1514_7158# d2 a_1565_6667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X18 a_33062_3379# d0 a_33859_3607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X19 a_26284_4019# a_26291_4237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X20 a_2545_1470# d0 a_3347_1109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X21 a_17496_1158# d0 a_17977_1246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X22 a_12101_2329# a_12358_2139# a_11303_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X23 a_17597_6755# a_17599_7048# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X24 gnd d0 a_29784_5617# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X25 gnd d0 a_29712_1133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X26 a_19838_1913# a_20091_1900# a_19788_3110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X27 a_4609_8067# a_4616_8285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X28 a_4987_2265# a_4769_2265# a_4512_2360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X29 a_11327_3354# a_11580_3341# a_11241_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X30 a_10182_6573# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X31 a_1482_5651# a_1276_6140# a_696_6324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X32 a_14551_3653# a_14345_4142# a_13765_4326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X33 a_12174_6401# a_12431_6211# a_11376_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X34 vdd d0 a_29728_2563# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X35 a_4988_1853# d1 a_5773_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X36 a_11158_3123# d2 a_11204_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X37 a_3379_3734# a_3636_3544# a_2586_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X38 a_3456_7629# a_3470_8412# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X39 a_28784_8633# d0 a_29586_8272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X40 a_6023_6561# a_5805_6561# a_5924_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X41 a_27553_3123# a_27335_3123# a_26755_3307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X42 a_28657_1507# a_28914_1317# a_28575_2115# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X43 a_30684_6068# a_30691_6286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X44 a_25191_7654# a_25205_8437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X45 a_21926_5025# a_21933_5243# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X46 a_26265_2708# a_26267_3001# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X47 a_24156_2946# d2 a_24239_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X48 a_13331_6781# a_13333_7074# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X49 a_15568_2116# d1 a_15654_1331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X50 gnd d0 a_16741_3582# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X51 a_26735_2289# a_26517_2289# a_26254_2201# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X52 a_15641_6188# a_15898_5998# a_15595_7208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X53 a_2603_4347# d0 a_3396_4752# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X54 a_24202_1926# a_24455_1913# a_24152_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X55 a_29531_5630# a_29545_6413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X56 a_26735_2289# d1 a_27521_1616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X57 a_26809_5949# a_26591_5949# a_26318_5956# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X58 a_15641_6188# d1 a_15727_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X59 a_22124_847# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X60 a_25078_1311# a_25082_1134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X61 a_20730_2728# a_20734_2551# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X62 a_14291_1088# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X63 a_14587_5689# a_14381_6178# a_13802_5950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X64 vdd d0 a_16722_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X65 a_28533_2958# a_28786_2945# a_28426_5173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X66 a_20754_3569# a_21007_3556# a_19957_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X67 gnd d0 a_8090_8647# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X68 a_27388_6177# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X69 a_22938_2093# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X70 a_18957_2488# a_18739_2488# a_18863_2607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X71 a_27589_5159# a_27371_5159# a_26792_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X72 vdd d0 a_29712_1133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X73 a_7711_1122# a_7706_1711# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X74 a_4506_2177# a_4512_2360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X75 a_23011_6165# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X76 a_12141_4600# a_12157_5383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X77 a_11323_3531# a_11580_3341# a_11241_4139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X78 a_25204_8849# a_25208_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X79 a_14831_403# a_14649_4548# a_14764_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X80 a_21993_8480# a_20844_8659# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X81 a_17850_5924# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X82 a_23254_7712# a_23048_8201# a_22469_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X83 a_5759_7581# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X84 a_21941_5944# d0 a_22432_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X85 a_185_4383# d0 a_660_4288# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X86 a_7711_1122# a_7964_1109# a_6909_1483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X87 a_2494_6993# d2 a_2573_8186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X88 a_31735_5172# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X89 a_6090_378# a_5908_4523# a_6023_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X90 a_7784_5194# a_7779_5783# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X91 a_13785_4932# a_13567_4932# a_13296_5038# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X92 gnd d0 a_8001_3145# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X93 gnd d1 a_15961_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X94 a_27932_283# d6 a_26029_208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X95 a_10150_1604# a_9944_2093# a_9364_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X96 vdd d0 a_16741_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X97 a_228_7036# d0 a_717_6930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X98 a_18812_3098# d2 a_18863_2607# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X99 vdd d0 a_21061_6198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X100 a_2603_4347# d0 a_3400_4575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X101 gnd d1 a_20300_8418# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X102 a_515_8360# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X103 a_17487_841# a_17489_940# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X104 a_22358_2277# a_22140_2277# a_21883_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X105 gnd d1 a_28951_3353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X106 gnd d1 a_16034_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X107 a_14826_284# d5 a_12951_197# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X108 a_16525_5219# a_16778_5206# a_15723_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X109 gnd d0 a_12340_1533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X110 a_22359_1865# d1 a_23144_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X111 a_17869_7354# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X112 gnd d1 a_29024_7425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X113 a_2536_6150# d1 a_2618_5542# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X114 a_20750_3746# a_21007_3556# a_19957_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X115 a_4609_8067# d0 a_5098_7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X116 a_23394_6573# a_23176_6573# a_23295_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X117 vdd d0 a_8073_7629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X118 a_9183_4313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X119 a_26610_7379# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X120 a_1240_4104# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X121 a_6678_5149# d3 a_6785_2934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X122 a_28602_7207# d2 a_28652_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X123 a_10223_5676# d2 a_10301_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X124 a_20717_1533# a_20970_1520# a_19920_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X125 a_3379_3734# a_3383_3557# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X126 a_16468_2577# a_16721_2564# a_15671_2349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X127 a_11417_8444# d0 a_12214_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X128 vdd d0 a_34149_5218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X129 a_5080_7355# d1 a_5878_7171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X130 a_3432_6788# a_3689_6598# a_2639_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X131 a_32135_6598# a_31917_6598# a_32041_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X132 gnd d1 a_33388_7438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X133 a_30711_7304# a_30717_7487# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X134 a_29458_1558# a_29711_1545# a_28661_1330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X135 a_29454_1735# a_29458_1558# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X136 a_15654_1331# d0 a_16447_1736# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X137 gnd d1 a_2802_1280# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X138 a_31958_5701# a_31752_6190# a_31173_5962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X139 a_13258_2709# d0 a_13749_2896# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X140 vdd d0 a_8001_3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X141 vdd d1 a_15961_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X142 a_18885_7170# a_18667_7170# a_18087_7354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X143 a_1358_5532# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X144 vdd d1 a_16034_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X145 a_9219_6349# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X146 vdd d1 a_28951_3353# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X147 vdd d2 a_7121_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X148 a_24334_4549# a_24591_4359# a_24239_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X149 vdd d0 a_12340_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X150 vdd d1 a_29024_7425# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X151 a_2536_6150# d1 a_2622_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X152 a_6831_1914# a_7084_1901# a_6781_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X153 a_2586_3329# a_2839_3316# a_2500_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X154 a_11396_7603# d0 a_12198_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X155 a_18031_4300# a_17813_4300# a_17550_4212# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X156 a_17148_133# a_25910_208# a_21680_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X157 a_1186_1050# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X158 a_1560_6548# a_1358_5532# a_1482_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X159 vdd d0 a_12413_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X160 gnd d4 a_2571_4946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X161 a_20713_1710# a_20970_1520# a_19920_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X162 a_19937_2323# a_20190_2310# a_19838_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X163 a_16464_2754# a_16721_2564# a_15671_2349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X164 a_4752_1247# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X165 a_228_7036# a_235_7254# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X166 a_9437_6349# a_9219_6349# a_8962_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X167 a_21868_1872# a_21870_1971# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X168 a_4579_6249# a_4585_6432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X169 a_2314_5136# a_2571_4946# a_1721_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X170 a_25188_7419# a_25445_7229# a_24390_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X171 a_29454_1735# a_29711_1545# a_28661_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X172 a_5851_2489# a_5649_1473# a_5768_1063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X173 a_21956_6444# a_21961_6768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X174 a_28730_5579# d0 a_29528_5395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X175 a_20768_4352# a_20772_4175# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X176 a_17759_1246# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X177 a_33895_5643# a_34148_5630# a_33098_5415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X178 a_15654_1331# d0 a_16451_1559# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X179 vdd d1 a_2802_1280# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X180 a_19907_6162# d1 a_19989_5554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X181 a_21866_1354# d0 a_22341_1259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X182 gnd d0 a_25351_2551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X183 a_25115_3347# a_25119_3170# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X184 a_33873_4390# a_33877_4213# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X185 a_18105_7960# a_17887_7960# a_17616_8066# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X186 a_26333_6456# d0 a_26808_6361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X187 a_28678_2348# d0 a_29471_2753# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X188 a_24049_5161# d3 a_24156_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X189 a_31716_4154# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X190 gnd d0 a_25424_6623# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X191 a_13566_5344# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X192 a_162_3182# a_168_3365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X193 a_22178_3901# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X194 a_13766_3914# a_13548_3914# a_13277_4020# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X195 a_31917_3136# a_31699_3136# a_31120_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X196 a_13729_1878# a_13511_1878# a_13240_1984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X197 a_17977_1246# a_17759_1246# a_17502_1341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X198 gnd d1 a_2929_8406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X199 a_8930_4926# a_8932_5025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X200 a_1820_246# a_1602_246# a_1721_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X201 a_27599_2513# d3 a_27698_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X202 a_26756_2895# a_26538_2895# a_26267_3001# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X203 a_2582_3506# a_2839_3316# a_2500_4114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X204 a_25188_7419# a_25192_7242# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X205 a_18574_2080# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X206 a_31990_7208# a_31772_7208# a_31193_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X207 a_9421_4919# a_9203_4919# a_8932_5025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X208 a_3396_4752# a_3400_4575# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X209 a_19933_2500# a_20190_2310# a_19838_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X210 gnd d0 a_12451_7229# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X211 a_643_3270# d1 a_1441_3086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X212 a_16506_4201# a_16759_4188# a_15704_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X213 gnd d2 a_24528_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X214 a_2504_3937# d1 a_2599_4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X215 a_30728_8322# a_30734_8505# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X216 a_7821_7230# a_7816_7819# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X217 a_4532_3378# a_4534_3896# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X218 gnd d0 a_25335_1121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X219 a_27714_283# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X220 a_8976_7279# d0 a_9457_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X221 a_716_7342# d1 a_1514_7158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X222 a_29496_3182# a_29749_3169# a_28694_3543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X223 a_14582_5160# a_14364_5160# a_13784_5344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X224 a_22921_1075# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X225 a_15522_3136# d2 a_15572_1939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X226 a_31834_5582# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X227 vdd d4 a_15676_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X228 a_10260_7712# d2 a_10306_6692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X229 a_19907_6162# d1 a_19993_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X230 a_33891_5820# a_34148_5630# a_33098_5415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X231 vdd d0 a_25351_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X232 a_33877_4213# a_33872_4802# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X233 vdd d0 a_34130_4200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X234 a_24407_8621# d0 a_25209_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X235 a_18067_6336# d1 a_18853_5663# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X236 a_28678_2348# d0 a_29475_2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X237 a_23176_3111# a_22958_3111# a_22378_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X238 a_7816_7819# a_7820_7642# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X239 a_7838_8248# a_8091_8235# a_7036_8609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X240 a_4605_7450# a_4607_7968# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X241 a_8926_4408# a_8930_4926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X242 vdd d0 a_25424_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X243 a_5686_3509# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X244 a_2318_4959# d3 a_2494_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X245 vdd d2 a_2757_3924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X246 a_162_3182# d0 a_643_3270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X247 a_15691_3367# d0 a_16484_3772# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X248 a_13346_7475# d0 a_13821_7380# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X249 a_30691_6286# d0 a_31172_6374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X250 a_33872_4802# a_33876_4625# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X251 gnd d2 a_11498_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X252 a_30938_4944# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X253 a_7710_1534# a_7963_1521# a_6913_1306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X254 a_22431_6349# a_22213_6349# a_21950_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X255 a_30882_1890# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X256 a_6085_259# d4 a_6682_4972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X257 a_26501_859# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X258 a_13247_2202# a_13253_2385# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X259 a_3347_1109# a_3600_1096# a_2545_1470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X260 a_17797_2870# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X261 a_9256_8385# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X262 a_2504_3937# d1 a_2603_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X263 a_30881_2302# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X264 a_4517_2684# d0 a_5008_2871# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X265 a_31173_5962# d1 a_31958_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X266 vdd d0 a_25335_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X267 a_8876_1971# a_8883_2189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X268 a_2577_8009# d1 a_2676_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X269 a_8658_196# d7 a_8757_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X270 a_20731_2316# a_20735_2139# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X271 a_33152_8469# d0 a_33945_8874# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X272 a_12105_2152# a_12358_2139# a_11303_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X273 a_17539_3377# d0 a_18014_3282# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X274 vdd d1 a_7276_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X275 a_28612_4151# a_28869_3961# a_28533_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X276 a_1519_7687# a_1313_8176# a_734_7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X277 a_7834_8425# a_8091_8235# a_7036_8609# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X278 a_12161_5206# a_12414_5193# a_11359_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X279 a_20043_8608# d0 a_20841_8424# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X280 a_28711_4561# d0 a_29509_4377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X281 a_17599_7048# d0 a_18088_6942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X282 a_17579_6030# a_17586_6248# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X283 a_15671_2349# a_15924_2336# a_15572_1939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X284 a_9384_3295# d1 a_10182_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X285 a_12832_197# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X286 a_7820_7642# a_7834_8425# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X287 a_19875_3949# d1 a_19970_4536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X288 a_33876_4625# a_34129_4612# a_33079_4397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X289 a_28784_8633# d0 a_29582_8449# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X290 a_8872_1354# d0 a_9347_1259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X291 a_15691_3367# d0 a_16488_3595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X292 a_28661_1330# a_28914_1317# a_28575_2115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X293 a_125_1146# a_131_1329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X294 a_12101_2329# a_12105_2152# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X295 a_21903_3390# d0 a_22378_3295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X296 a_4210_172# a_5966_259# a_6090_378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X297 a_7706_1711# a_7963_1521# a_6913_1306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X298 a_6930_2324# a_7183_2311# a_6831_1914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X299 a_11059_4984# d3 a_11235_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X300 a_20786_5782# a_20790_5605# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X301 a_15568_2116# d1 a_15650_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X302 a_9129_1259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X303 a_258_8455# vref SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X304 a_5878_7171# a_5660_7171# a_5081_6943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X305 a_3437_6199# a_3432_6788# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X306 a_11290_1318# d0 a_12083_1723# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X307 a_32062_2526# a_31844_2526# a_31963_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X308 a_30638_3232# d0 a_31119_3320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X309 a_22233_7367# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X310 a_24225_7195# a_24482_7005# a_24053_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X311 a_8883_2189# a_8889_2372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X312 a_23300_6692# a_23130_7593# a_23249_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X313 a_4826_4907# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X314 a_32976_4164# d1 a_33058_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X315 vdd d2 a_20128_3936# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X316 a_33152_8469# d0 gnd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X317 a_33053_8059# a_33306_8046# a_32970_7043# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X318 a_16520_5808# a_16777_5618# a_15727_5403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X319 a_16465_2342# a_16469_2165# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X320 vdd d2 a_15862_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X321 a_25081_1546# a_25334_1533# a_24284_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X322 a_30902_2908# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X323 vdd d0 a_16759_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X324 a_32893_3148# a_33150_2958# a_32790_5186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X325 a_33840_2177# a_33835_2766# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X326 a_20043_8608# d0 a_20845_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X327 gnd d3 a_33223_7030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X328 gnd d1 a_20263_6382# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X329 a_4971_835# d1 a_5768_1063# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X330 a_15667_2526# a_15924_2336# a_15572_1939# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X331 a_29568_7666# a_29582_8449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X332 a_215_6236# d0 a_696_6324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X333 a_9438_5937# d1 a_10223_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X334 a_4568_5414# a_4570_5932# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X335 a_6781_3111# d2 a_6827_2091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X336 a_23048_8201# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X337 a_19875_3949# d1 a_19974_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X338 a_33872_4802# a_34129_4612# a_33079_4397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X339 a_26247_1983# d0 a_26736_1877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X340 a_3380_3322# a_3384_3145# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X341 gnd d1 a_29004_6407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X342 a_26237_1183# d0 a_26718_1271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X343 a_10343_271# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X344 a_33912_6661# a_33929_7444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X345 a_26230_965# a_26237_1183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X346 a_18656_1472# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X347 a_6926_2501# a_7183_2311# a_6831_1914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X348 a_18105_7960# a_17887_7960# a_17614_7967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X349 a_30702_6793# a_30704_7086# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X350 a_26254_2201# d0 a_26735_2289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X351 a_27677_6704# d3 a_27771_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X352 a_19689_4971# a_19942_4958# a_19092_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X353 a_26718_1271# d1 a_27516_1087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X354 a_9364_2277# a_9146_2277# a_8883_2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X355 a_11290_1318# d0 a_12087_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X356 a_28579_1938# d1 a_28674_2525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X357 a_12177_6636# a_12194_7419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X358 a_14592_2514# a_14390_1498# a_14514_1617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X359 a_6930_2324# d0 a_7727_2552# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X360 a_30919_3926# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X361 a_26303_5037# a_26310_5255# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X362 a_22469_7973# a_22251_7973# a_21978_7980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X363 a_10109_2501# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X364 a_1721_246# d4 a_2314_5136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X365 a_30992_7998# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X366 a_32976_4164# d1 a_33062_3379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X367 a_1477_5122# a_1259_5122# a_680_4894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X368 a_23020_1485# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X369 a_1602_246# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X370 a_33049_8236# a_33306_8046# a_32970_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X371 gnd d0 a_8073_7629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X372 a_25077_1723# a_25334_1533# a_24284_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X373 a_5567_2081# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X374 a_31210_7998# a_30992_7998# a_30719_8005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X375 a_21851_854# d0 a_22342_847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X376 a_17504_1859# d0 a_17995_1852# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X377 a_31136_4338# a_30918_4338# a_30661_4433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X378 a_22468_8385# a_22250_8385# a_21993_8480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X379 a_11417_8444# d0 a_12210_8849# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X380 vdd d3 a_33223_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X381 vdd d1 a_20263_6382# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X382 gnd d0 a_34149_5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X383 a_30717_7487# a_30719_8005# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X384 a_26029_208# a_30203_209# a_30322_209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X385 gnd d2 a_20091_1900# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X386 a_24301_2336# d0 a_25094_2741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X387 a_22123_1259# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X388 a_10327_2501# a_10109_2501# a_10233_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X389 a_2566_2311# a_2819_2298# a_2467_1901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X390 a_26590_6361# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X391 gnd d0 a_3727_8222# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X392 a_28734_5402# d0 a_29531_5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X393 a_19030_6560# d4 a_19097_377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X394 a_21868_1872# d0 a_22359_1865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X395 a_12193_7831# a_12197_7654# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X396 a_22197_4919# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X397 a_10467_390# a_10285_4535# a_10327_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X398 a_12174_6401# a_12178_6224# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X399 a_31958_5701# d2 a_32036_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X400 gnd d2 a_28832_1925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X401 vdd d4 a_11312_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X402 a_9130_847# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X403 a_23222_2501# d3 a_23321_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X404 a_22379_2883# a_22161_2883# a_21890_2989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X405 vdd d1 a_24610_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X406 a_28579_1938# d1 a_28678_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X407 a_27480_2513# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X408 vdd d0 a_20987_2538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X409 a_14691_2514# a_14473_2514# a_14592_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X410 a_13333_7074# d0 a_13822_6968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X411 a_24338_4372# a_24591_4359# a_24239_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X412 a_22341_1259# a_22123_1259# a_21866_1354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X413 vdd d1 a_24627_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X414 a_30954_6374# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X415 a_31120_2908# a_30902_2908# a_30631_3014# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X416 a_23394_6573# d4 a_23461_390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X417 a_31761_1510# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X418 a_25135_4600# a_25151_5383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X419 a_21890_2989# a_21897_3207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X420 a_11396_7603# d0 a_12194_7419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X421 a_18853_5663# a_18647_6152# a_18068_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X422 gnd d4 a_28683_4983# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X423 a_1223_3086# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X424 a_15605_4152# d1 a_15687_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X425 a_13258_2709# a_13260_3002# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X426 a_7036_8609# d0 a_7834_8425# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X427 a_15682_8047# a_15935_8034# a_15599_7031# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X428 gnd d2 a_33196_1938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X429 a_4599_7267# d0 a_5080_7355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X430 a_24225_7195# d2 a_24271_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X431 a_607_822# a_389_822# a_116_829# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X432 a_13236_1367# a_13238_1885# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X433 a_27626_7195# d2 a_27677_6704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X434 a_25192_7242# a_25445_7229# a_24390_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X435 a_16501_4790# a_16758_4600# a_15708_4385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X436 a_24301_2336# d0 a_25098_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X437 a_4789_3283# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X438 a_4863_6943# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X439 a_17760_834# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X440 a_19792_2933# a_20045_2920# a_19685_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X441 vdd d0 a_3727_8222# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X442 a_30719_8005# a_30721_8104# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X443 a_498_7342# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X444 a_8757_196# a_8539_196# a_8658_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X445 a_30665_4951# a_30667_5050# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X446 a_8920_4225# a_8926_4408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X447 a_13547_4326# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X448 a_5008_2871# a_4790_2871# a_4519_2977# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X449 a_12197_7654# a_12211_8437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X450 a_26338_6780# d0 a_26829_6967# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X451 a_13603_7380# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X452 a_31082_1284# a_30864_1284# a_30601_1196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X453 a_3342_1698# a_3346_1521# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X454 a_26537_3307# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X455 a_30721_8104# a_30728_8322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X456 a_7817_7407# a_7821_7230# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X457 vdd d1 a_2912_7388# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X458 a_31156_4944# a_30938_4944# a_30665_4951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X459 a_6963_4537# a_7220_4347# a_6868_3950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X460 a_734_7948# a_516_7948# a_243_7955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X461 a_26291_4237# d0 a_26772_4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X462 a_26230_965# d0 a_26719_859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X463 a_18014_3282# a_17796_3282# a_17533_3194# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X464 a_15605_4152# d1 a_15691_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X465 a_8993_8297# a_8999_8480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X466 a_7036_8609# d0 a_7838_8248# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X467 gnd d0 a_21098_8234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X468 a_716_7342# a_498_7342# a_241_7437# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X469 a_5805_3099# a_5587_3099# a_5007_3283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X470 a_15678_8224# a_15935_8034# a_15599_7031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X471 gnd d1 a_7256_6383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X472 a_19920_1305# a_20173_1292# a_19834_2090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X473 gnd d0 a_16832_8260# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X474 a_16575_8450# a_16579_8273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X475 gnd d1 a_33332_4384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X476 a_20845_8247# a_20840_8836# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X477 a_29582_8449# a_29839_8259# a_28784_8633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X478 a_12142_4188# a_12137_4777# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X479 a_9402_3901# a_9184_3901# a_8911_3908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X480 a_1446_3615# a_1240_4104# a_661_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X481 a_6937_8199# a_7194_8009# a_6858_7006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X482 a_26260_2384# a_26265_2708# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X483 a_5097_8373# a_4879_8373# a_4622_8468# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X484 a_30661_4433# a_30665_4951# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X485 a_6831_1914# d1 a_6926_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X486 a_18684_8188# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X487 a_28606_7030# d2 a_28685_8223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X488 a_133_1847# d0 a_624_1840# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X489 a_14619_7196# a_14401_7196# a_13821_7380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X490 a_24407_8621# d0 a_25205_8437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X491 a_26340_7073# a_26347_7291# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X492 a_4495_1342# d0 a_4970_1247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X493 gnd d0 a_25407_5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X494 a_3473_8647# a_3726_8634# a_2676_8419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X495 gnd d0 a_34186_7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X496 a_17487_841# d0 a_17978_834# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X497 a_22160_3295# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X498 a_25172_6224# a_25167_6813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X499 a_17575_5413# a_17577_5931# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X500 a_28715_4384# d0 a_29512_4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X501 a_23031_7183# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X502 a_4568_5414# d0 a_5043_5319# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X503 a_21581_184# a_23337_271# a_23461_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X504 a_1586_2476# a_1368_2476# a_1487_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X505 a_18812_6560# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X506 vdd d1 a_24591_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X507 a_25081_1546# a_25095_2329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X508 a_32790_5186# d3 a_32897_2971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X509 vdd d0 a_21098_8234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X510 a_1659_6548# d4 a_1726_365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X511 vdd d1 a_7256_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X512 vdd d0 a_16832_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X513 a_5081_6943# a_4863_6943# a_4592_7049# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X514 a_5924_6561# d3 a_6023_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X515 a_25167_6813# a_25171_6636# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X516 vdd d1 a_33332_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X517 a_16579_8273# a_16574_8862# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X518 gnd d0 a_29801_6635# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X519 gnd d0 a_29729_2151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X520 a_9364_2277# d1 a_10150_1604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X521 a_4770_1853# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X522 a_2618_5542# d0 a_3420_5181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X523 vdd d0 a_16778_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X524 a_3384_3145# a_3637_3132# a_2582_3506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X525 a_31209_8410# d1 a_31995_7737# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X526 a_2573_8186# d1 a_2655_7578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X527 a_11204_2103# d1 a_11290_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X528 gnd d1 a_20190_2310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X529 a_6831_1914# d1 a_6930_2324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X530 gnd d3 a_2747_6980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X531 a_17586_6248# d0 a_18067_6336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X532 a_15704_4562# d0 a_16506_4201# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X533 a_405_2252# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X534 a_26355_7992# d0 a_26846_7985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X535 a_18936_6679# d3 a_19030_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X536 a_17777_1852# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X537 a_11417_8444# a_11670_8431# a_11318_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X538 a_28606_7030# d2 a_28689_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X539 a_5550_1063# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X540 a_10145_1075# a_9927_1075# a_9348_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X541 a_606_1234# a_388_1234# a_125_1146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X542 a_26347_7291# a_26353_7474# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X543 a_24280_1495# a_24537_1305# a_24198_2103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X544 a_3469_8824# a_3726_8634# a_2676_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X545 vdd d0 a_34186_7254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X546 a_17850_5924# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X547 a_13711_1272# a_13493_1272# a_13230_1184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X548 a_26500_1271# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X549 a_21943_6043# d0 a_22432_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X550 a_18557_1062# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X551 a_21933_5243# d0 a_22414_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X552 a_30203_209# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X553 a_22341_1259# d1 a_23139_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X554 a_22342_847# a_22124_847# a_21853_953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X555 a_15645_6011# d1 a_15744_6421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X556 a_27553_6585# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X557 a_13785_4932# a_13567_4932# a_13294_4939# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X558 a_32041_6717# d3 a_32135_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X559 a_17995_1852# a_17777_1852# a_17506_1958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X560 a_24202_1926# d1 a_24297_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X561 a_14308_2106# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X562 a_22414_5331# d1 a_23212_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X563 a_21860_1171# a_21866_1354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X564 a_28648_6187# d1 a_28734_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X565 a_5060_6337# a_4842_6337# a_4579_6249# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X566 a_27298_1087# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X567 vdd d0 a_29801_6635# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X568 vdd d0 a_29729_2151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X569 a_31844_2526# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X570 a_18775_1062# a_18557_1062# a_17977_1246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X571 a_6785_2934# a_7038_2921# a_6678_5149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X572 a_3380_3322# a_3637_3132# a_2582_3506# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X573 a_11340_4549# a_11597_4359# a_11245_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X574 a_26245_1884# a_26247_1983# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X575 vdd d1 a_20190_2310# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X576 a_1721_246# d5 a_1820_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X577 a_3453_7394# a_3710_7204# a_2655_7578# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X578 a_11413_8621# a_11670_8431# a_11318_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X579 a_16524_5631# a_16777_5618# a_15727_5403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X580 a_14707_284# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X581 a_1492_2595# a_1322_3496# a_1446_3615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X582 a_2599_4524# d0 a_3397_4340# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X583 vdd d2 a_24455_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X584 vdd d1 a_28914_1317# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X585 a_389_822# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X586 a_30624_2397# d0 a_31099_2302# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X587 a_4309_172# a_4091_172# a_4210_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X588 gnd d0 a_3616_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X589 a_426_2858# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X590 a_258_8455# d0 a_733_8360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X591 a_5024_4301# d1 a_5810_3628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X592 a_20755_3157# a_21008_3144# a_19953_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X593 gnd d0 a_8091_8235# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X594 a_6913_1306# a_7166_1293# a_6827_2091# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X595 gnd d0 a_25388_4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X596 a_24202_1926# d1 a_24301_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X597 a_13531_2896# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X598 a_9964_3111# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X599 gnd d3 a_20118_6992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X600 a_23103_2501# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X601 a_24271_6175# d1 a_24357_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X602 vdd d0 a_29785_5205# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X603 gnd d1 a_29041_8443# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X604 a_5966_259# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X605 a_27558_3652# d2 a_27604_2632# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X606 a_13530_3308# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X607 a_11055_5161# d3 a_11162_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X608 a_13838_8398# a_13620_8398# a_13357_8310# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X609 gnd d4 a_24306_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X610 a_644_2858# a_426_2858# a_155_2964# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X611 gnd d0 a_12430_6623# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X612 gnd d2 a_2720_1888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X613 a_14597_2633# a_14427_3534# a_14546_3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X614 a_6930_2324# d0 a_7723_2729# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X615 a_27434_3533# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X616 a_13838_8398# d1 a_14624_7725# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X617 a_20823_7818# a_21080_7628# a_20030_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X618 a_16542_6237# a_16537_6826# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X619 a_26828_7379# a_26610_7379# a_26347_7291# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X620 a_21943_6043# a_21950_6261# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X621 a_6854_7183# a_7111_6993# a_6682_4972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X622 a_29475_2576# a_29728_2563# a_28678_2348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X623 a_24152_3123# a_24409_2933# a_24049_5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X624 gnd d3 a_33150_2958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X625 a_24053_4984# d3 a_24225_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X626 a_2599_4524# d0 a_3401_4163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X627 gnd d0 a_7964_1109# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X628 a_19792_2933# d2 a_19871_4126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X629 a_31798_3546# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X630 a_516_7948# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X631 a_29548_6648# a_29801_6635# a_28751_6420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X632 a_13223_966# d0 a_13712_860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X633 a_31880_1100# a_31662_1100# a_31083_872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X634 vdd d0 a_3616_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X635 gnd d1 a_2892_6370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X636 a_15744_6421# d0 a_16537_6826# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X637 gnd d0 a_12341_1121# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X638 a_21905_3908# a_21907_4007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X639 a_31871_7618# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X640 a_8930_4926# d0 a_9421_4919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X641 a_20751_3334# a_21008_3144# a_19953_3518# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X642 vdd d0 a_8091_8235# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X643 a_11277_6175# a_11534_5985# a_11231_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X644 a_8876_1971# d0 a_9365_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X645 vdd d0 a_8074_7217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X646 a_9184_3901# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X647 a_26611_6967# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X648 a_28734_5402# d0 a_29527_5807# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X649 a_606_1234# d1 a_1404_1050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X650 vdd d1 a_29041_8443# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X651 a_9147_1865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X652 a_16469_2165# a_16722_2152# a_15667_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X653 a_32790_5186# a_33047_4996# a_32197_296# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X654 a_5768_1063# d2 a_5851_2489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X655 a_18087_7354# a_17869_7354# a_17612_7449# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X656 a_21914_4225# d0 a_22395_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X657 a_6858_7006# d2 a_6941_8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X658 a_28652_6010# a_28905_5997# a_28602_7207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X659 gnd d1 a_24610_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X660 a_12141_4600# a_12394_4587# a_11344_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X661 a_13766_3914# a_13548_3914# a_13275_3921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X662 vdd d0 a_12430_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X663 a_29459_1146# a_29712_1133# a_28657_1507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X664 a_20730_2728# a_20987_2538# a_19937_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X665 gnd d0 a_20987_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X666 a_4519_2977# a_4526_3195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X667 a_16484_3772# a_16488_3595# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X668 a_10255_7183# a_10037_7183# a_9457_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X669 a_4769_2265# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X670 a_7723_2729# a_7727_2552# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X671 a_1276_6140# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X672 a_22395_4313# d1 a_23181_3640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X673 a_30975_6980# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X674 a_15650_1508# d0 a_16448_1324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X675 a_9421_4919# a_9203_4919# a_8930_4926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X676 a_29471_2753# a_29728_2563# a_28678_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X677 a_5805_6561# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X678 a_18853_5663# d2 a_18931_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X679 a_16524_5631# a_16538_6414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X680 a_135_1946# a_142_2164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X681 a_31120_2908# d1 a_31917_3136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X682 a_4592_7049# a_4599_7267# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X683 a_22452_6955# d1 a_23249_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X684 a_29544_6825# a_29801_6635# a_28751_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X685 a_8913_4007# a_8920_4225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X686 a_24229_7018# d2 a_24308_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X687 a_26517_2289# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X688 a_27631_7724# a_27425_8213# a_26846_7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X689 vdd d1 a_2892_6370# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X690 a_15744_6421# d0 a_16541_6649# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X691 vdd d0 a_12341_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X692 gnd d0 a_3710_7204# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X693 a_21956_6444# d0 a_22431_6349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X694 a_16561_7667# a_16814_7654# a_15764_7439# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X695 a_3436_6611# a_3453_7394# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X696 vdd d2 a_24492_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X697 a_6023_6561# a_5805_6561# a_5929_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X698 a_17994_2264# d1 a_18780_1591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X699 vdd d0 a_12414_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X700 a_20714_1298# a_20971_1108# a_19916_1482# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X701 a_16465_2342# a_16722_2152# a_15667_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X702 a_2467_1901# d1 a_2566_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X703 a_19834_2090# d1 a_19920_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X704 vdd d2 a_20201_8008# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X705 a_9438_5937# a_9220_5937# a_8949_6043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X706 gnd d1 a_2839_3316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X707 a_31995_7737# a_31789_8226# a_31210_7998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X708 a_2672_8596# a_2929_8406# a_2577_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X709 a_29455_1323# a_29712_1133# a_28657_1507# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X710 a_20713_1710# a_20717_1533# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X711 a_26736_1877# d1 a_27521_1616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X712 a_30938_4944# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X713 a_31119_3320# a_30901_3320# a_30638_3232# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X714 a_6967_4360# a_7220_4347# a_6868_3950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X715 a_15650_1508# d0 a_16452_1147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X716 a_27932_283# a_27714_283# a_27838_402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X717 a_33839_2589# a_33856_3372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X718 a_733_8360# d1 a_1519_7687# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X719 a_189_4901# a_191_5000# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X720 a_33928_7856# a_33932_7679# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X721 a_14587_5689# a_14381_6178# a_13801_6362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X722 a_28674_2525# d0 a_29472_2341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X723 gnd d3 a_15779_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X724 a_1565_6667# a_1395_7568# a_1514_7158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X725 a_15723_5580# d0 a_16525_5219# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X726 gnd d0 a_25425_6211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X727 a_13567_4932# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X728 a_21462_184# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X729 a_29586_8272# a_29839_8259# a_28784_8633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X730 a_24229_7018# d2 a_24312_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X731 a_27589_5159# a_27371_5159# a_26791_5343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X732 a_23011_6165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X733 gnd d3 a_7111_6993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X734 a_25168_6401# a_25172_6224# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X735 a_11231_7195# a_11488_7005# a_11059_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X736 a_18050_5318# a_17832_5318# a_17569_5230# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X737 a_13221_867# a_13223_966# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X738 a_22141_1865# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X739 a_16557_7844# a_16814_7654# a_15764_7439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X740 a_33038_2538# a_33295_2348# a_32943_1951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X741 a_15781_8457# a_16034_8444# a_15682_8047# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X742 a_23254_7712# a_23048_8201# a_22468_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X743 a_4482_941# d0 a_4971_835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X744 a_28771_7438# a_29024_7425# a_28685_8223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X745 a_23176_6573# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X746 a_30601_1196# d0 a_31082_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X747 vdd d1 a_2839_3316# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X748 a_7816_7819# a_8073_7629# a_7023_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X749 a_1404_1050# d2 a_1487_2476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X750 a_15781_8457# d0 a_16574_8862# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X751 a_30322_209# d6 a_26029_208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X752 a_8967_6768# d0 a_9458_6955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X753 a_26338_6780# a_26340_7073# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X754 a_16447_1736# a_16451_1559# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X755 a_7710_1534# a_7724_2317# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X756 a_28771_7438# d0 a_29564_7843# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X757 a_33892_5408# a_34149_5218# a_33094_5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X758 gnd d1 a_24591_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X759 a_28674_2525# d0 a_29476_2164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X760 a_23394_6573# a_23176_6573# a_23300_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X761 gnd d1 a_24574_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X762 vdd d0 a_25425_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X763 a_9385_2883# a_9167_2883# a_8894_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X764 a_13821_7380# a_13603_7380# a_13346_7475# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X765 a_31752_6190# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X766 a_10218_5147# d2 a_10301_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X767 a_1240_4104# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X768 a_4555_5013# a_4562_5231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X769 a_6827_2091# d1 a_6909_1483# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X770 a_18667_7170# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X771 a_2618_5542# d0 a_3416_5358# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X772 a_15687_3544# d0 a_16485_3360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X773 a_9384_3295# a_9166_3295# a_8909_3390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X774 a_30682_5969# d0 a_31173_5962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X775 a_17629_8467# d0 a_18104_8372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X776 a_5081_6943# d1 a_5878_7171# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X777 a_32202_415# a_32020_4560# a_32135_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X778 a_15777_8634# a_16034_8444# a_15682_8047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X779 a_20026_7590# a_20283_7400# a_19944_8198# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X780 a_14514_1617# d2 a_14592_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X781 gnd d0 a_16704_1546# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X782 a_5098_7961# d1 a_5883_7700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X783 a_3383_3557# a_3397_4340# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X784 a_19685_5148# d3 a_19792_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X785 a_10233_2620# a_10063_3521# a_10182_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X786 a_9474_8385# d1 a_10260_7712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X787 a_252_8272# a_258_8455# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X788 a_28767_7615# a_29024_7425# a_28685_8223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X789 a_3469_8824# a_3473_8647# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X790 a_4549_4396# a_4553_4914# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X791 a_17813_4300# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X792 a_20030_7413# d0 a_20827_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X793 gnd d0 a_7963_1521# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X794 a_15781_8457# d0 a_16578_8685# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X795 a_31100_1890# a_30882_1890# a_30609_1897# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X796 a_21993_8480# d0 a_22468_8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X797 a_12156_5795# a_12413_5605# a_11363_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X798 a_26280_3402# a_26282_3920# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X799 a_1358_5532# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X800 a_6682_4972# d3 a_6858_7006# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X801 a_29458_1558# a_29472_2341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X802 a_23181_3640# d2 a_23227_2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X803 a_11307_2336# d0 a_12100_2741# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X804 a_30721_8104# d0 a_31210_7998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X805 a_28771_7438# d0 a_29568_7666# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X806 a_9219_6349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X807 a_14345_4142# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X808 a_33148_8646# d0 a_33946_8462# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X809 a_29544_6825# a_29548_6648# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X810 a_25136_4188# a_25131_4777# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X811 a_30624_2397# a_30629_2721# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X812 a_11380_6408# d0 a_12173_6813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X813 a_12161_5206# a_12156_5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X814 a_2417_3098# d2 a_2463_2078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X815 a_9475_7973# a_9257_7973# a_8986_8079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X816 vdd d1 a_24574_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X817 a_30728_8322# d0 a_31209_8410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X818 a_4842_6337# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X819 a_27335_3123# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X820 a_23130_7593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X821 a_30680_5451# a_30682_5969# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X822 a_30919_3926# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X823 a_25192_7242# a_25187_7831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X824 a_1544_4510# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X825 a_17526_2976# a_17533_3194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X826 a_30975_6980# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X827 a_15687_3544# d0 a_16489_3183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X828 a_11344_4372# a_11597_4359# a_11245_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X829 a_33839_2589# a_34092_2576# a_33042_2361# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X830 vdd d2 a_28869_3961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X831 a_25171_6636# a_25424_6623# a_24374_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X832 a_7707_1299# a_7964_1109# a_6909_1483# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X833 vdd d0 a_16704_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X834 gnd d1 a_15924_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X835 a_5732_2489# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X836 a_30974_7392# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X837 a_32197_296# d4 a_32794_5009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X838 a_5851_2489# a_5649_1473# a_5773_1592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X839 a_2490_7170# d2 a_2540_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X840 a_31699_3136# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X841 a_32078_296# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X842 a_11231_7195# d2 a_11277_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X843 a_17759_1246# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X844 a_14597_2633# d3 a_14691_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X845 gnd d1 a_28914_1317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X846 a_4499_1959# d0 a_4988_1853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X847 a_11286_1495# d0 a_12084_1311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X848 a_21860_1171# d0 a_22341_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X849 a_19948_8021# d1 a_20047_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X850 a_31772_7208# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X851 a_9203_4919# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X852 vdd d0 a_7963_1521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X853 a_30629_2721# d0 a_31120_2908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X854 a_22234_6955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X855 a_26327_6273# d0 a_26808_6361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X856 a_24198_2103# d1 a_24280_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X857 a_27599_2513# a_27397_1497# a_27516_1087# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X858 a_11307_2336# d0 a_12104_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X859 a_24275_5998# a_24528_5985# a_24225_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X860 a_33148_8646# d0 a_33950_8285# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X861 a_14649_4548# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X862 a_31917_3136# a_31699_3136# a_31119_3320# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X863 a_14546_6586# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X864 a_26808_6361# d1 a_27594_5688# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X865 a_25082_1134# a_25335_1121# a_24280_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X866 a_24271_6175# d1 a_24353_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X867 a_11380_6408# d0 a_12177_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X868 a_14364_5160# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X869 a_1820_246# a_1602_246# a_1726_365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X870 a_13333_7074# a_13340_7292# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X871 a_15419_5174# a_15676_4984# a_14826_284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X872 a_31990_7208# a_31772_7208# a_31192_7392# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X873 a_206_5919# d0 a_697_5912# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X874 a_31120_2908# a_30902_2908# a_30629_2721# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X875 a_20827_7641# a_21080_7628# a_20030_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X876 a_33049_8236# d1 a_33135_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X877 a_33835_2766# a_34092_2576# a_33042_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X878 a_25167_6813# a_25424_6623# a_24374_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X879 vdd d1 a_20173_1292# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X880 vdd d1 a_15924_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X881 a_717_6930# d1 a_1514_7158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X882 a_26301_4938# d0 a_26792_4931# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X883 a_2500_4114# a_2757_3924# a_2421_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X884 a_4480_842# a_4482_941# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X885 a_624_1840# a_406_1840# a_133_1847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X886 gnd d0 a_3599_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X887 a_4534_3896# a_4536_3995# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X888 a_11286_1495# d0 a_12088_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X889 vdd d2 a_7084_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X890 a_2655_7578# d0 a_3453_7394# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X891 a_22213_6349# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X892 a_24357_5390# d0 a_25154_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X893 a_6926_2501# d0 a_7728_2140# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X894 vdd d3 a_2674_2908# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X895 a_5007_3283# d1 a_5805_3099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X896 a_18068_5924# d1 a_18853_5663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X897 a_30680_5451# d0 a_31155_5356# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X898 a_4622_8468# a_3473_8647# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X899 gnd d3 a_11415_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X900 a_2639_6383# a_2892_6370# a_2540_5973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X901 a_13350_8092# d0 a_13839_7986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X902 gnd d0 a_8074_7217# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X903 a_25078_1311# a_25335_1121# a_24280_1495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X904 a_31137_3926# a_30919_3926# a_30648_4032# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X905 a_27698_2513# a_27480_2513# a_27599_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X906 a_13357_8310# d0 a_13838_8398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X907 a_26340_7073# d0 a_26829_6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X908 a_22431_6349# a_22213_6349# a_21956_6444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X909 a_3397_4340# a_3401_4163# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X910 a_20827_7641# a_20841_8424# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X911 a_31210_7998# a_30992_7998# a_30721_8104# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X912 a_26501_859# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X913 a_7019_7591# a_7276_7401# a_6937_8199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X914 a_13821_7380# d1 a_14619_7196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X915 a_15682_8047# d1 a_15777_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X916 a_20734_2551# a_20987_2538# a_19937_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X917 a_1313_8176# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X918 a_29455_1323# a_29459_1146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X919 a_26247_1983# a_26254_2201# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X920 a_30648_4032# a_30655_4250# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X921 a_15419_5174# d3 a_15522_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X922 a_21961_6768# a_21963_7061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X923 gnd d1 a_11543_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X924 a_5878_7171# d2 a_5929_6680# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X925 a_9457_7367# a_9239_7367# a_8976_7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X926 a_28685_8223# d1 a_28767_7615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X927 a_7023_7414# d0 a_7820_7642# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X928 a_32020_4560# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X929 a_21581_184# d6 a_21680_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X930 a_27833_283# d4 a_28430_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X931 a_17543_3994# d0 a_18032_3888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X932 gnd d1 a_2819_2298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X933 a_33929_7444# a_33933_7267# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X934 a_17562_5012# a_17569_5230# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X935 a_1519_7687# a_1313_8176# a_733_8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X936 a_2635_6560# a_2892_6370# a_2540_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X937 a_9385_2883# d1 a_10182_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X938 a_1565_6667# d3 a_1659_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X939 a_8909_3390# a_8911_3908# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X940 a_4590_6756# d0 a_5081_6943# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X941 a_8866_1171# d0 a_9347_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X942 a_31172_6374# a_30954_6374# a_30691_6286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X943 a_19871_4126# a_20128_3936# a_19792_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X944 a_24394_7426# d0 a_25187_7831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X945 a_17556_4395# a_17560_4913# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X946 a_10150_1604# d2 a_10228_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X947 a_16561_7667# a_16575_8450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X948 a_16502_4378# a_16759_4188# a_15704_4562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X949 gnd d2 a_15935_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X950 a_5878_7171# a_5660_7171# a_5080_7355# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X951 a_31995_7737# d2 a_32041_6717# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X952 a_24297_2513# d0 a_25099_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X953 a_15682_8047# d1 a_15781_8457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X954 vdd d3 a_20045_2920# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X955 a_5883_7700# a_5677_8189# a_5097_8373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X956 a_26846_7985# a_26628_7985# a_26355_7992# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X957 a_17612_7449# a_17614_7967# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X958 a_32970_7043# a_33223_7030# a_32794_5009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X959 a_20010_6395# a_20263_6382# a_19911_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X960 a_26254_2201# a_26260_2384# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X961 a_32062_2526# a_31844_2526# a_31968_2645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X962 a_7748_3158# a_7743_3747# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X963 a_30655_4250# a_30661_4433# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X964 a_20790_5605# a_20804_6388# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X965 a_28685_8223# d1 a_28771_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X966 vdd d3 a_28786_2945# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X967 a_9944_2093# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X968 a_6941_8022# d1 a_7040_8432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X969 a_5081_6943# a_4863_6943# a_4590_6756# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X970 a_16448_1324# a_16452_1147# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X971 a_13236_1367# d0 a_13711_1272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X972 a_26845_8397# a_26627_8397# a_26370_8492# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X973 a_28751_6420# a_29004_6407# a_28652_6010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X974 a_204_5401# d0 a_679_5306# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X975 a_9420_5331# d1 a_10218_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X976 a_27626_7195# a_27408_7195# a_26829_6967# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X977 a_5924_6561# a_5722_5545# a_5841_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X978 a_14390_1498# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X979 a_13309_5439# d0 a_13784_5344# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X980 a_26282_3920# d0 a_26773_3913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X981 a_17832_5318# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X982 a_33042_2361# a_33295_2348# a_32943_1951# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X983 a_23048_8201# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X984 a_4585_6432# d0 a_5060_6337# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X985 a_26245_1884# d0 a_26736_1877# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X986 a_13363_8493# a_12214_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X987 a_33098_5415# a_33351_5402# a_33012_6200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X988 a_10343_271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X989 vdd d2 a_11461_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X990 a_22250_8385# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X991 a_24394_7426# d0 a_25191_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X992 a_7820_7642# a_8073_7629# a_7023_7414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X993 a_1259_5122# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X994 a_33042_2361# d0 a_33835_2766# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X995 a_5098_7961# a_4880_7961# a_4609_8067# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X996 vdd d2 a_15935_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X997 vdd d1 a_7166_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X998 a_5851_2489# d3 a_5950_2489# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X999 a_3470_8412# a_3474_8235# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1000 a_9364_2277# a_9146_2277# a_8889_2372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1001 a_19933_2500# d0 a_20731_2316# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1002 a_1409_1579# a_1203_2068# a_624_1840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1003 a_1441_3086# d2 a_1492_2595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1004 a_32966_7220# a_33223_7030# a_32794_5009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1005 a_20006_6572# a_20263_6382# a_19911_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1006 a_19861_7182# d2 a_19907_6162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1007 a_33896_5231# a_34149_5218# a_33094_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1008 a_26320_6055# a_26327_6273# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1009 a_28575_2115# a_28832_1925# a_28529_3135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1010 a_4988_1853# a_4770_1853# a_4497_1860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1011 a_11277_6175# d1 a_11363_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1012 a_8932_5025# a_8939_5243# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1013 a_10109_2501# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1014 a_2314_5136# d3 a_2417_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1015 gnd d0 a_25408_5193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1016 a_4480_842# a_7707_1299# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1017 a_3474_8235# a_3727_8222# a_2672_8596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1018 a_1477_5122# a_1259_5122# a_679_5306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1019 a_11281_5998# d1 a_11380_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1020 a_10285_4535# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1021 a_28711_4561# d0 a_29513_4200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1022 vdd d1 a_15980_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1023 a_5768_1063# a_5550_1063# a_4971_835# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1024 a_11055_5161# a_11312_4971# a_10462_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1025 a_13728_2290# a_13510_2290# a_13247_2202# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1026 a_696_6324# a_478_6324# a_215_6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1027 a_10223_5676# a_10017_6165# a_9438_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1028 a_26029_208# a_30203_209# a_27932_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1029 a_14473_2514# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1030 a_24370_6585# a_24627_6395# a_24275_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1031 a_22123_1259# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1032 a_19957_3341# d0 a_20750_3746# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1033 a_13801_6362# a_13583_6362# a_13320_6274# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1034 a_26718_1271# a_26500_1271# a_26237_1183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1035 a_32897_2971# d2 a_32980_3987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1036 a_26590_6361# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1037 a_8872_1354# a_8874_1872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1038 a_18957_2488# d4 a_19097_377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1039 a_23222_2501# a_23020_1485# a_23139_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1040 a_10467_390# a_10285_4535# a_10400_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1041 a_17541_3895# a_17543_3994# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1042 a_20030_7413# d0 a_20823_7818# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1043 a_22431_6349# d1 a_23217_5676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1044 a_26791_5343# a_26573_5343# a_26310_5255# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1045 a_33042_2361# d0 a_33839_2589# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1046 a_14624_7725# d2 a_14670_6705# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1047 a_17577_5931# d0 a_18068_5924# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1048 a_23295_6573# a_23093_5557# a_23212_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1049 a_14826_284# d4 a_15419_5174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1050 a_13311_5957# a_13313_6056# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1051 a_31083_872# a_30865_872# a_30592_879# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1052 a_19933_2500# d0 a_20735_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1053 a_14691_2514# a_14473_2514# a_14597_2633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1054 gnd d2 a_2830_7996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1055 a_30954_6374# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1056 a_23321_2501# d4 a_23461_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1057 vdd d0 a_12377_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1058 a_12951_197# a_14707_284# a_14826_284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1059 a_3470_8412# a_3727_8222# a_2672_8596# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1060 a_18853_5663# a_18647_6152# a_18067_6336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1061 a_607_822# a_389_822# a_118_928# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1062 a_2421_2921# d2 a_2500_4114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1063 a_9401_4313# d1 a_10187_3640# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1064 a_442_4288# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1065 a_21980_8079# a_21987_8297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1066 vdd d1 a_29004_6407# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1067 a_17487_841# a_20714_1298# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1068 a_9457_7367# d1 a_10255_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1069 a_17760_834# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1070 a_21851_854# a_21853_953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1071 a_19957_3341# d0 a_20754_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1072 a_15727_5403# a_15980_5390# a_15641_6188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1073 a_13290_4421# d0 a_13765_4326# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1074 a_516_7948# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1075 a_13326_6457# a_13331_6781# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1076 a_22359_1865# a_22141_1865# a_21868_1872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1077 a_17796_3282# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1078 a_19944_8198# d1 a_20026_7590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1079 vdd d3 a_7038_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1080 a_30882_1890# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1081 a_498_7342# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1082 a_26538_2895# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1083 a_5587_3099# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1084 a_19948_8021# d1 a_20043_8608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1085 a_13621_7986# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1086 a_7003_6396# a_7256_6383# a_6904_5986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1087 a_13547_4326# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1088 a_26280_3402# d0 a_26755_3307# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1089 a_8932_5025# d0 a_9421_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1090 a_4549_4396# d0 a_5024_4301# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1091 a_5929_6680# a_5759_7581# a_5883_7700# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1092 a_33079_4397# a_33332_4384# a_32980_3987# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1093 a_13748_3308# a_13530_3308# a_13267_3220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1094 a_15595_7208# a_15852_7018# a_15423_4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1095 a_26611_6967# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1096 a_26537_3307# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1097 a_9184_3901# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1098 a_13620_8398# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1099 a_18032_3888# a_17814_3888# a_17541_3895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1100 a_11363_5390# d0 a_12156_5795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1101 vdd d2 a_11498_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1102 a_29569_7254# a_29564_7843# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1103 a_14401_7196# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1104 a_26228_866# d0 a_26719_859# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1105 a_18031_4300# a_17813_4300# a_17556_4395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1106 gnd d0 a_3617_2114# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1107 vdd d1 a_7203_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1108 a_24308_8211# d1 a_24390_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1109 a_21680_184# d7 a_17148_133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1110 a_3432_6788# a_3436_6611# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1111 a_12125_3170# a_12120_3759# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1112 a_27677_6704# a_27507_7605# a_27626_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1113 a_18812_3098# a_18594_3098# a_18015_2870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1114 a_25154_5618# a_25407_5605# a_24357_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1115 a_23456_271# d4 a_24053_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1116 a_33049_8236# d1 a_33131_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1117 a_7800_6624# a_7817_7407# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1118 gnd d0 a_25389_4175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1119 a_26243_1366# a_26245_1884# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1120 a_30644_3415# a_30646_3933# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1121 a_2494_6993# d2 a_2577_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1122 gnd d0 a_8054_6199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1123 a_7760_4765# a_7764_4588# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1124 a_1446_3615# a_1240_4104# a_660_4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1125 a_2562_2488# a_2819_2298# a_2467_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1126 a_13531_2896# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1127 a_15526_2959# d2 a_15609_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1128 a_1368_2476# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1129 gnd d0 a_12431_6211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1130 a_15572_1939# a_15825_1926# a_15522_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1131 a_6926_2501# d0 a_7724_2317# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1132 a_6999_6573# a_7256_6383# a_6904_5986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1133 a_4489_1159# d0 a_4970_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1134 a_33835_2766# a_33839_2589# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1135 a_1487_2476# a_1285_1460# a_1404_1050# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1136 a_25155_5206# a_25150_5795# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1137 a_27516_1087# d2 a_27599_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1138 a_23337_271# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1139 a_33075_4574# a_33332_4384# a_32980_3987# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1140 a_696_6324# d1 a_1482_5651# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1141 a_29476_2164# a_29729_2151# a_28674_2525# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1142 gnd d0 a_3709_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1143 a_4562_5231# d0 a_5043_5319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1144 a_16521_5396# a_16778_5206# a_15723_5580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1145 a_26772_4325# a_26554_4325# a_26291_4237# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1146 a_2494_6993# a_2747_6980# a_2318_4959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1147 a_9438_5937# a_9220_5937# a_8947_5944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1148 a_1586_2476# a_1368_2476# a_1492_2595# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1149 a_30704_7086# a_30711_7304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1150 a_29549_6236# a_29802_6223# a_28747_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1151 vdd d0 a_3617_2114# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1152 a_24308_8211# d1 a_24394_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1153 a_17575_5413# d0 a_18050_5318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1154 a_388_1234# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1155 a_15740_6598# d0 a_16538_6414# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1156 a_28430_4996# d3 a_28606_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1157 vdd d0 a_25389_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1158 a_13311_5957# d0 a_13802_5950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1159 a_13493_1272# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1160 a_31210_7998# d1 a_31995_7737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1161 a_23249_7183# a_23031_7183# a_22452_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1162 a_461_5306# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1163 vdd d0 a_25372_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1164 a_20750_3746# a_20754_3569# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1165 a_5640_6153# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1166 a_5950_2489# a_5732_2489# a_5851_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1167 a_7023_7414# d0 a_7816_7819# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1168 a_18088_6942# a_17870_6942# a_17599_7048# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1169 a_13567_4932# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1170 gnd d1 a_11580_3341# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1171 a_30646_3933# a_30648_4032# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1172 a_21905_3908# d0 a_22396_3901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1173 a_17777_1852# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1174 a_12142_4188# a_12395_4175# a_11340_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1175 a_10145_1075# a_9927_1075# a_9347_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1176 vdd d0 a_12431_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1177 gnd d2 a_20164_5972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1178 a_680_4894# a_462_4894# a_189_4901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1179 a_606_1234# a_388_1234# a_131_1329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1180 gnd d0 a_20988_2126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1181 gnd d1 a_11653_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1182 a_15708_4385# a_15961_4372# a_15609_3975# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1183 a_13711_1272# a_13493_1272# a_13236_1367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1184 a_25095_2329# a_25099_2152# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1185 gnd d2 a_28905_5997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1186 gnd d0 a_29765_4599# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1187 a_29472_2341# a_29729_2151# a_28674_2525# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1188 a_11158_3123# d2 a_11208_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1189 a_18557_1062# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1190 vdd d0 a_3709_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1191 a_22342_847# d1 a_23139_1075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1192 a_14764_6586# a_14546_6586# a_14665_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1193 a_18915_4522# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1194 a_28698_3366# a_28951_3353# a_28612_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1195 a_8909_3390# d0 a_9384_3295# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1196 a_13340_7292# d0 a_13821_7380# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1197 a_31193_6980# a_30975_6980# a_30704_7086# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1198 a_29545_6413# a_29802_6223# a_28747_6597# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1199 a_19685_5148# a_19942_4958# a_19092_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1200 a_31209_8410# a_30991_8410# a_30728_8322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1201 a_8969_7061# d0 a_9458_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1202 a_22415_4919# d1 a_23212_5147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1203 a_28529_3135# d2 a_28575_2115# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1204 a_1322_3496# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1205 a_5060_6337# a_4842_6337# a_4585_6432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1206 a_21680_184# a_21462_184# a_19191_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1207 a_24198_2103# a_24455_1913# a_24152_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1208 a_3419_5593# a_3433_6376# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1209 a_15740_6598# d0 a_16542_6237# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1210 a_14509_1088# a_14291_1088# a_13711_1272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1211 a_24297_2513# d0 a_25095_2329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1212 a_16562_7255# a_16815_7242# a_15760_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1213 a_10187_3640# d2 a_10233_2620# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1214 a_24353_5567# d0 a_25151_5383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1215 a_31844_2526# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1216 a_3363_2539# a_3616_2526# a_2566_2311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1217 a_28730_5579# d0 a_29532_5218# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1218 a_6937_8199# d1 a_7019_7591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1219 a_28529_3135# a_28786_2945# a_28426_5173# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1220 a_18067_6336# a_17849_6336# a_17586_6248# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1221 a_26316_5438# a_26318_5956# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1222 a_4553_4914# a_4555_5013# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1223 a_6941_8022# d1 a_7036_8609# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1224 a_10462_271# d4 a_11055_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1225 a_30611_1996# d0 a_31100_1890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1226 a_4512_2360# a_4517_2684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1227 a_21950_6261# a_21956_6444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1228 a_3343_1286# a_3347_1109# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1229 vdd d1 a_11580_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1230 gnd d0 a_16814_7654# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1231 vdd d0 a_34075_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1232 a_19865_7005# a_20118_6992# a_19689_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1233 a_12138_4365# a_12395_4175# a_11340_4549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1234 vdd d0 a_20988_2126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1235 a_155_2964# d0 a_644_2858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1236 a_10136_7593# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1237 a_30684_6068# d0 a_31173_5962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1238 a_30618_2214# d0 a_31099_2302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1239 vdd d1 a_11653_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1240 a_4309_172# a_4091_172# a_1820_246# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1241 a_15704_4562# a_15961_4372# a_15609_3975# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1242 a_24053_4984# a_24306_4971# a_23456_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1243 a_426_2858# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1244 a_8984_7980# a_8986_8079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1245 a_5025_3889# d1 a_5810_3628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1246 a_25099_2152# a_25094_2741# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1247 a_14427_3534# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1248 a_22414_5331# a_22196_5331# a_21933_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1249 a_11162_2946# d2 a_11241_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1250 vdd d1 a_2929_8406# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1251 a_31099_2302# d1 a_31885_1629# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1252 a_28694_3543# a_28951_3353# a_28612_4151# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1253 a_31155_5356# d1 a_31953_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1254 a_6963_4537# d0 a_7761_4353# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1255 a_14500_7606# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1256 a_30667_5050# a_30674_5268# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1257 a_6090_378# d5 a_4210_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1258 a_25171_6636# a_25188_7419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1259 a_208_6018# a_215_6236# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1260 a_11307_2336# a_11560_2323# a_11208_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1261 a_27553_3123# d2 a_27604_2632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1262 a_18031_4300# d1 a_18817_3627# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1263 a_24239_3962# a_24492_3949# a_24156_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1264 a_28616_3974# d1 a_28711_4561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1265 a_18863_2607# a_18693_3508# a_18812_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1266 a_16558_7432# a_16815_7242# a_15760_7616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1267 a_2573_8186# d1 a_2659_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1268 a_31662_1100# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1269 a_3359_2716# a_3616_2526# a_2566_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1270 a_14597_2633# a_14427_3534# a_14551_3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1271 gnd d1 a_24664_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1272 a_29495_3594# a_29509_4377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1273 a_13839_7986# d1 a_14624_7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1274 a_9475_7973# a_9257_7973# a_8984_7980# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1275 a_26828_7379# a_26610_7379# a_26353_7474# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1276 gnd d3 a_24482_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1277 a_11277_6175# d1 a_11359_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1278 vdd d2 a_33196_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1279 gnd d0 a_16721_2564# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1280 a_7817_7407# a_8074_7217# a_7019_7591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1281 a_15777_8634# d0 a_16575_8450# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1282 vdd d0 a_16814_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1283 a_26829_6967# d1 a_27626_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1284 a_9474_8385# a_9256_8385# a_8999_8480# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1285 a_4543_4213# a_4549_4396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1286 a_5024_4301# a_4806_4301# a_4543_4213# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1287 a_25114_3759# a_25371_3569# a_24321_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1288 gnd d0 a_29711_1545# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1289 a_12137_4777# a_12141_4600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1290 a_32202_415# d5 a_30322_209# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1291 a_28767_7615# d0 a_29565_7431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1292 a_21888_2696# a_21890_2989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1293 a_27594_5688# d2 a_27672_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1294 a_717_6930# a_499_6930# a_228_7036# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1295 a_21976_7462# a_21978_7980# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1296 a_661_3876# a_443_3876# a_170_3883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1297 gnd d0 a_8053_6611# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1298 a_8874_1872# d0 a_9365_1865# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1299 a_13822_6968# a_13604_6968# a_13333_7074# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1300 a_9203_4919# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1301 a_6963_4537# d0 a_7765_4176# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1302 a_30631_3014# d0 a_31120_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1303 a_22234_6955# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1304 a_3343_1286# a_3600_1096# a_2545_1470# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1305 a_33131_7628# a_33388_7438# a_33049_8236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1306 a_660_4288# a_442_4288# a_185_4383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1307 a_11303_2513# a_11560_2323# a_11208_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1308 a_19916_1482# d0 a_20714_1298# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1309 a_9385_2883# a_9167_2883# a_8896_2989# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1310 a_28616_3974# d1 a_28715_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1311 gnd d0 a_16705_1134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1312 a_2463_2078# a_2720_1888# a_2417_3098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1313 vdd d1 a_24664_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1314 a_148_2347# d0 a_623_2252# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1315 a_27425_8213# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1316 gnd d0 a_12377_3569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1317 a_22396_3901# d1 a_23181_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1318 gnd d2 a_7157_5973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1319 vdd d0 a_16721_2564# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1320 a_208_6018# d0 a_697_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1321 a_15777_8634# d0 a_16579_8273# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1322 a_30322_209# a_32078_296# a_32202_415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1323 a_13260_3002# a_13267_3220# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1324 gnd d2 a_33233_3974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1325 a_16488_3595# a_16502_4378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1326 a_5805_6561# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1327 a_12157_5383# a_12414_5193# a_11359_5567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1328 vdd d4 a_2571_4946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1329 a_15650_1508# a_15907_1318# a_15568_2116# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1330 a_18848_5134# d2 a_18931_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1331 a_10228_2501# a_10026_1485# a_10150_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1332 vdd d0 a_29711_1545# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1333 gnd d1 a_28931_2335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1334 a_16574_8862# a_16578_8685# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1335 a_13313_6056# d0 a_13802_5950# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1336 a_31789_8226# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1337 a_28767_7615# d0 a_29569_7254# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1338 vdd d0 a_7980_2539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1339 a_4753_835# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1340 a_27631_7724# a_27425_8213# a_26845_8397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1341 a_26303_5037# d0 a_26792_4931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1342 a_10561_271# d6 a_8658_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1343 a_11376_6585# d0 a_12174_6401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1344 a_21950_6261# d0 a_22431_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1345 vdd d0 a_25388_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1346 vdd d0 a_8053_6611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1347 a_13728_2290# d1 a_14514_1617# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1348 a_30719_8005# d0 a_31210_7998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1349 a_23139_1075# d2 a_23222_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1350 a_13784_5344# d1 a_14582_5160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1351 a_7761_4353# a_7765_4176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1352 a_2586_3329# d0 a_3379_3734# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1353 a_24275_5998# d1 a_24370_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1354 gnd d1 a_33278_1330# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1355 a_15526_2959# a_15779_2946# a_15419_5174# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1356 a_18630_5134# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1357 a_22395_4313# a_22177_4313# a_21914_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1358 a_33840_2177# a_34093_2164# a_33038_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1359 a_31995_7737# a_31789_8226# a_31209_8410# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1360 a_2659_7401# d0 a_3452_7806# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1361 a_1395_7568# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1362 a_5060_6337# d1 a_5846_5664# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1363 a_25172_6224# a_25425_6211# a_24370_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1364 vdd d0 a_16705_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1365 a_15599_7031# a_15852_7018# a_15423_4997# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1366 a_31137_3926# a_30919_3926# a_30646_3933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1367 a_33836_2354# a_33840_2177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1368 a_20844_8659# a_21097_8646# a_20047_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1369 a_31193_6980# a_30975_6980# a_30702_6793# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1370 a_31917_6598# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1371 a_30865_872# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1372 a_31761_1510# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1373 a_22994_5147# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1374 a_734_7948# d1 a_1519_7687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1375 vdd d0 a_7964_1109# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1376 gnd d1 a_7203_3329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1377 a_31192_7392# a_30974_7392# a_30717_7487# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1378 a_19788_3110# d2 a_19838_1913# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1379 a_13267_3220# a_13273_3403# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1380 a_1565_6667# a_1395_7568# a_1519_7687# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1381 a_21924_4926# d0 a_22415_4919# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1382 vdd d1 a_28931_2335# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1383 vdd d2 a_24528_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1384 a_12124_3582# a_12138_4365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1385 a_12100_2741# a_12104_2564# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1386 a_11241_4139# d1 a_11323_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1387 gnd d0 a_3689_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1388 a_31885_1629# d2 a_31963_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1389 a_8896_2989# a_8903_3207# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1390 a_11318_8034# a_11571_8021# a_11235_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1391 a_11376_6585# d0 a_12178_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1392 gnd d0 a_3672_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1393 a_17560_4913# a_17562_5012# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1394 a_27771_6585# d4 a_27838_402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1395 a_22141_1865# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1396 a_18050_5318# a_17832_5318# a_17575_5413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1397 a_5773_1592# a_5567_2081# a_4987_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1398 a_33932_7679# a_34185_7666# a_33135_7451# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1399 a_21939_5426# a_21941_5944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1400 a_2586_3329# d0 a_3383_3557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1401 a_28575_2115# d1 a_28661_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1402 a_20751_3334# a_20755_3157# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1403 a_4480_842# d0 a_4971_835# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1404 gnd d1 a_16017_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1405 a_28648_6187# a_28905_5997# a_28602_7207# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1406 vdd d1 a_33278_1330# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1407 a_4532_3378# d0 a_5007_3283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1408 a_23176_6573# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1409 a_24321_3354# a_24574_3341# a_24235_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1410 a_20828_7229# a_21081_7216# a_20026_7590# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1411 a_12137_4777# a_12394_4587# a_11344_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1412 a_33836_2354# a_34093_2164# a_33038_2538# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1413 a_2659_7401# d0 a_3456_7629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1414 a_25168_6401# a_25425_6211# a_24370_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1415 a_9167_2883# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1416 a_13603_7380# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1417 a_17599_7048# a_17606_7266# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1418 a_4592_7049# d0 a_5081_6943# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1419 a_24152_3123# d2 a_24198_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1420 a_27521_1616# a_27315_2105# a_26736_1877# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1421 a_20840_8836# a_21097_8646# a_20047_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1422 a_10026_1485# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1423 a_9166_3295# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1424 gnd d0 a_3600_1096# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1425 a_16451_1559# a_16704_1546# a_15654_1331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1426 a_28426_5173# d3 a_28529_3135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1427 a_18015_2870# d1 a_18812_3098# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1428 a_10063_3521# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1429 a_16451_1559# a_16465_2342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1430 gnd d1 a_11633_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1431 gnd d0 a_29838_8671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1432 a_3457_7217# a_3452_7806# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1433 a_31885_1629# a_31679_2118# a_31100_1890# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1434 a_28430_4996# d3 a_28602_7207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1435 a_16537_6826# a_16541_6649# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1436 gnd d0 a_25372_3157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1437 a_11241_4139# d1 a_11327_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1438 a_31953_5172# a_31735_5172# a_31156_4944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1439 a_17623_8284# d0 a_18104_8372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1440 a_11314_8211# a_11571_8021# a_11235_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1441 vdd d0 a_3672_5580# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1442 a_1441_3086# a_1223_3086# a_643_3270# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1443 a_13348_7993# d0 a_13839_7986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1444 a_22432_5937# a_22214_5937# a_21943_6043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1445 a_33928_7856# a_34185_7666# a_33135_7451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1446 a_6909_1483# d0 a_7707_1299# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1447 a_10233_2620# a_10063_3521# a_10187_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1448 a_3452_7806# a_3456_7629# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1449 a_623_2252# d1 a_1409_1579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1450 a_7724_2317# a_7728_2140# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1451 a_643_3270# a_425_3270# a_162_3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1452 a_9475_7973# d1 a_10260_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1453 a_9257_7973# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1454 a_18104_8372# d1 a_18890_7699# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1455 vdd d1 a_16017_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1456 a_20735_2139# a_20988_2126# a_19933_2500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1457 a_21941_5944# a_21943_6043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1458 a_24317_3531# a_24574_3341# a_24235_4139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1459 a_26284_4019# d0 a_26773_3913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1460 a_20824_7406# a_21081_7216# a_20026_7590# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1461 a_17496_1158# a_17502_1341# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1462 a_33860_3195# a_33855_3784# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1463 a_717_6930# a_499_6930# a_226_6743# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1464 a_131_1329# a_133_1847# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1465 a_13765_4326# d1 a_14551_3653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1466 a_23176_3111# d2 a_23227_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1467 a_7019_7591# d0 a_7821_7230# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1468 a_18611_4116# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1469 gnd d0 a_21043_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1470 a_14345_4142# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1471 a_26755_3307# d1 a_27553_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1472 gnd d0 a_29822_7241# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1473 a_23461_390# d5 a_21581_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1474 a_16447_1736# a_16704_1546# a_15654_1331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1475 a_23144_1604# a_22938_2093# a_22358_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1476 a_1586_2476# d4 a_1726_365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1477 a_33877_4213# a_34130_4200# a_33075_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1478 a_17541_3895# d0 a_18032_3888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1479 a_5098_7961# a_4880_7961# a_4607_7968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1480 a_4842_6337# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1481 a_14546_3124# a_14328_3124# a_13749_2896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1482 a_204_5401# a_206_5919# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1483 a_7779_5783# a_7783_5606# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1484 a_27335_3123# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1485 a_13230_1184# a_13236_1367# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1486 vdd d0 a_29838_8671# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1487 a_10301_6573# a_10099_5557# a_10218_5147# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1488 a_6682_4972# a_6935_4959# a_6085_259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1489 a_19920_1305# d0 a_20713_1710# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1490 a_13326_6457# d0 a_13801_6362# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1491 a_5043_5319# a_4825_5319# a_4562_5231# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1492 a_15671_2349# d0 a_16464_2754# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1493 a_22975_4129# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1494 a_17849_6336# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1495 a_18931_6560# d3 a_19030_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1496 a_28661_1330# d0 a_29454_1735# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1497 a_8859_953# a_8866_1171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1498 a_27397_1497# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1499 vdd d3 a_33150_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1500 a_26316_5438# d0 a_26791_5343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1501 gnd d0 a_34075_1558# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1502 a_31699_3136# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1503 a_23217_5676# d2 a_23295_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1504 a_21961_6768# d0 a_22452_6955# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1505 a_13303_5256# a_13309_5439# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1506 a_20714_1298# a_20718_1121# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1507 a_20731_2316# a_20988_2126# a_19933_2500# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1508 a_14592_2514# d3 a_14691_2514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1509 a_17616_8066# a_17623_8284# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1510 a_27470_5569# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1511 a_4497_1860# d0 a_4988_1853# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1512 gnd d2 a_2793_5960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1513 gnd d0 a_3653_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1514 a_31772_7208# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1515 a_18739_2488# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1516 a_14665_6586# d3 a_14764_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1517 a_12138_4365# a_12142_4188# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1518 a_26846_7985# a_26628_7985# a_26357_8091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1519 a_24239_3962# d1 a_24338_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1520 a_17519_2359# d0 a_17994_2264# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1521 a_26809_5949# d1 a_27594_5688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1522 a_14649_4548# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1523 a_19916_1482# a_20173_1292# a_19834_2090# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1524 vdd d0 a_29822_7241# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1525 a_6023_6561# d4 a_6090_378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1526 a_17579_6030# d0 a_18068_5924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1527 a_406_1840# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1528 a_241_7437# a_243_7955# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1529 a_3401_4163# a_3396_4752# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1530 a_19920_1305# d0 a_20717_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1531 a_15671_2349# d0 a_16468_2577# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1532 a_2417_3098# a_2674_2908# a_2314_5136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1533 a_27558_3652# a_27352_4141# a_26773_3913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1534 a_21883_2372# d0 a_22358_2277# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1535 a_11162_2946# a_11415_2933# a_11055_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1536 a_1721_246# d4 a_2318_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1537 a_27833_283# d5 a_27932_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1538 a_24390_7603# d0 a_25192_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1539 a_18050_5318# d1 a_18848_5134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1540 a_28661_1330# d0 a_29458_1558# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1541 a_7821_7230# a_8074_7217# a_7019_7591# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1542 a_8866_1171# a_8872_1354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1543 a_33038_2538# d0 a_33836_2354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1544 a_5846_5664# a_5640_6153# a_5061_5925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1545 vdd d0 a_25407_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1546 a_25118_3582# a_25371_3569# a_24321_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1547 a_29476_2164# a_29471_2753# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1548 a_4517_2684# a_4519_2977# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1549 a_17513_2176# a_17519_2359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1550 a_10037_7183# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1551 a_22213_6349# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1552 vdd d0 a_3653_4562# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1553 a_20047_8431# d0 a_20840_8836# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1554 a_26808_6361# a_26590_6361# a_26327_6273# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1555 a_30674_5268# d0 a_31155_5356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1556 a_33823_1159# a_33818_1748# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1557 a_252_8272# d0 a_733_8360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1558 a_29548_6648# a_29565_7431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1559 a_32939_2128# d1 a_33021_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1560 a_13275_3921# a_13277_4020# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1561 a_11290_1318# a_11543_1305# a_11204_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1562 a_30864_1284# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1563 a_3437_6199# a_3690_6186# a_2635_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1564 a_12088_1134# a_12083_1723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1565 a_33135_7451# a_33388_7438# a_33049_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1566 vdd d2 a_28832_1925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1567 a_27698_2513# a_27480_2513# a_27604_2632# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1568 a_31963_2526# a_31761_1510# a_31880_1100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1569 vdd d0 a_12467_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1570 a_27838_402# a_27656_4547# a_27698_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1571 a_27771_6585# a_27553_6585# a_27677_6704# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1572 gnd d0 a_21024_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1573 a_6868_3950# a_7121_3937# a_6785_2934# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1574 a_1313_8176# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1575 a_33135_7451# d0 a_33928_7856# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1576 a_243_7955# a_245_8054# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1577 vdd d4 a_28683_4983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1578 a_9457_7367# a_9239_7367# a_8982_7462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1579 a_5007_3283# a_4789_3283# a_4526_3195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1580 a_1514_7158# a_1296_7158# a_717_6930# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1581 a_24225_7195# d2 a_24275_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1582 a_20026_7590# d0 a_20824_7406# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1583 a_33038_2538# d0 a_33840_2177# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1584 a_18890_7699# d2 a_18936_6679# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1585 a_15654_1331# a_15907_1318# a_15568_2116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1586 a_10306_6692# a_10136_7593# a_10255_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1587 a_7743_3747# a_8000_3557# a_6950_3342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1588 a_29545_6413# a_29549_6236# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1589 a_1482_5651# d2 a_1560_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1590 a_31880_1100# a_31662_1100# a_31082_1284# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1591 gnd d0 a_7980_2539# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1592 a_20047_8431# d0 a_20844_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1593 a_13221_867# d0 a_13712_860# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1594 a_17886_8372# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1595 a_30955_5962# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1596 a_8962_6444# d0 a_9437_6349# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1597 gnd d0 a_8036_5593# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1598 a_8859_953# d0 a_9348_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1599 a_19788_3110# a_20045_2920# a_19685_5148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1600 vdd d0 a_12378_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1601 a_24338_4372# d0 a_25131_4777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1602 a_32939_2128# d1 a_33025_1343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1603 gnd d0 a_34112_3594# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1604 a_5677_8189# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1605 a_26628_7985# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1606 a_23254_7712# d2 a_23300_6692# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1607 a_1560_6548# d3 a_1659_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1608 a_3433_6376# a_3690_6186# a_2635_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1609 a_31172_6374# a_30954_6374# a_30697_6469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1610 a_607_822# d1 a_1404_1050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1611 a_28602_7207# a_28859_7017# a_28430_4996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1612 a_5649_1473# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1613 a_6913_1306# d0 a_7706_1711# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1614 a_26627_8397# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1615 vdd d1 a_7220_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1616 a_27408_7195# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1617 vdd d0 a_21024_4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1618 a_8911_3908# a_8913_4007# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1619 a_31990_7208# d2 a_32041_6717# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1620 a_5722_5545# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1621 a_8999_8480# a_7837_8660# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1622 a_33053_8059# d1 a_33148_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1623 a_33135_7451# d0 a_33932_7679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1624 a_19953_3518# a_20210_3328# a_19871_4126# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1625 vdd d1 a_7293_8419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1626 a_4562_5231# a_4568_5414# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1627 a_26228_866# a_26230_965# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1628 a_191_5000# d0 a_680_4894# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1629 a_18890_7699# a_18684_8188# a_18105_7960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1630 a_13240_1984# d0 a_13729_1878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1631 a_20026_7590# d0 a_20828_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1632 a_12156_5795# a_12160_5618# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1633 a_8658_196# a_12832_197# a_12951_197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1634 vdd d0 a_3599_1508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1635 gnd d1 a_20246_5364# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1636 a_13548_3914# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1637 gnd d1 a_15997_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1638 a_9421_4919# d1 a_10218_5147# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1639 a_13230_1184# d0 a_13711_1272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1640 a_20808_6211# a_21061_6198# a_20006_6572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1641 a_198_5218# d0 a_679_5306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1642 a_13247_2202# d0 a_13728_2290# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1643 a_26538_2895# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1644 a_13621_7986# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1645 a_5924_6561# a_5722_5545# a_5846_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1646 a_13303_5256# d0 a_13784_5344# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1647 gnd d1 a_28987_5389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1648 a_31100_1890# a_30882_1890# a_30611_1996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1649 a_7838_8248# a_7833_8837# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1650 a_11359_5567# d0 a_12157_5383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1651 a_13711_1272# d1 a_14509_1088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1652 a_8757_196# d8 vout SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1653 a_6909_1483# a_7166_1293# a_6827_2091# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1654 a_18088_6942# a_17870_6942# a_17597_6755# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1655 a_1203_2068# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1656 a_15572_1939# d1 a_15667_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1657 a_10182_3111# a_9964_3111# a_9385_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1658 a_21907_4007# d0 a_22396_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1659 vdd d3 a_20118_6992# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1660 a_17832_5318# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1661 a_33075_4574# d0 a_33873_4390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1662 a_16538_6414# a_16542_6237# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1663 a_18032_3888# a_17814_3888# a_17543_3994# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1664 a_4579_6249# d0 a_5060_6337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1665 a_12105_2152# a_12100_2741# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1666 vdd d3 a_15852_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1667 a_28575_2115# d1 a_28657_1507# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1668 a_18931_6560# a_18729_5544# a_18848_5134# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1669 a_17995_1852# d1 a_18780_1591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1670 a_22378_3295# a_22160_3295# a_21897_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1671 a_6913_1306# d0 a_7710_1534# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1672 a_25155_5206# a_25408_5193# a_24353_5567# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1673 a_20804_6388# a_20808_6211# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1674 a_1259_5122# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1675 a_22378_3295# d1 a_23176_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1676 a_12197_7654# a_12450_7641# a_11400_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1677 a_22451_7367# a_22233_7367# a_21970_7279# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1678 a_1409_1579# a_1203_2068# a_623_2252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1679 a_33053_8059# d1 a_33152_8469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1680 a_29513_4200# a_29508_4789# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1681 a_18863_2607# d3 a_18957_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1682 a_31119_3320# a_30901_3320# a_30644_3415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1683 a_4499_1959# a_4506_2177# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1684 a_478_6324# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1685 a_24053_4984# d3 a_24229_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1686 a_4988_1853# a_4770_1853# a_4499_1959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1687 vdd d1 a_2819_2298# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1688 vdd d1 a_20246_5364# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1689 a_13583_6362# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1690 a_26318_5956# d0 a_26809_5949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1691 a_198_5218# a_204_5401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1692 vdd d0 a_25462_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1693 a_15727_5403# d0 a_16524_5631# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1694 a_24284_1318# d0 a_25077_1723# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1695 a_10285_4535# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1696 a_11245_3962# a_11498_3949# a_11162_2946# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1697 a_3346_1521# a_3360_2304# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1698 a_4553_4914# d0 a_5044_4907# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1699 a_26573_5343# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1700 gnd d1 a_11670_8431# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1701 a_215_6236# a_221_6419# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1702 a_7780_5371# a_7784_5194# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1703 gnd d2 a_15825_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1704 a_17994_2264# a_17776_2264# a_17513_2176# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1705 vdd d3 a_2747_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1706 a_5768_1063# a_5550_1063# a_4970_1247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1707 a_10223_5676# a_10017_6165# a_9437_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1708 a_23093_5557# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1709 a_15572_1939# d1 a_15671_2349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1710 gnd d3 a_11488_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1711 a_696_6324# a_478_6324# a_221_6419# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1712 a_14473_2514# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1713 a_26736_1877# a_26518_1877# a_26245_1884# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1714 a_28715_4384# a_28968_4371# a_28616_3974# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1715 a_26718_1271# a_26500_1271# a_26243_1366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1716 a_13801_6362# a_13583_6362# a_13326_6457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1717 a_12120_3759# a_12377_3569# a_11327_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1718 gnd d0 a_8017_4575# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1719 a_26735_2289# a_26517_2289# a_26260_2384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1720 a_8999_8480# d0 a_9474_8385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1721 a_22432_5937# d1 a_23217_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1722 a_26791_5343# a_26573_5343# a_26316_5438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1723 a_27516_1087# a_27298_1087# a_26719_859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1724 a_12193_7831# a_12450_7641# a_11400_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1725 a_19092_258# d4 a_19685_5148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1726 a_14619_7196# d2 a_14670_6705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1727 a_7019_7591# d0 a_7817_7407# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1728 a_23295_6573# a_23093_5557# a_23217_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1729 a_8874_1872# a_8876_1971# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1730 a_31083_872# a_30865_872# a_30594_978# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1731 a_25910_208# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1732 a_8962_6444# a_8967_6768# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1733 a_25118_3582# a_25132_4365# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1734 a_28747_6597# a_29004_6407# a_28652_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1735 a_22938_2093# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1736 a_25094_2741# a_25098_2564# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1737 a_21883_2372# a_21888_2696# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1738 gnd d0 a_16831_8672# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1739 a_24284_1318# d0 a_25081_1546# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1740 a_6781_3111# a_7038_2921# a_6678_5149# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1741 a_680_4894# a_462_4894# a_191_5000# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1742 a_172_3982# d0 a_661_3876# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1743 gnd d0 a_29766_4187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1744 vdd d0 a_3710_7204# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1745 vdd d1 a_11670_8431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1746 a_16562_7255# a_16557_7844# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1747 vdd d0 a_34165_6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1748 gnd d2 a_7194_8009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1749 a_21963_7061# a_21970_7279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1750 gnd d1 a_20227_4346# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1751 a_5759_7581# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1752 a_9402_3901# d1 a_10187_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1753 a_179_4200# d0 a_660_4288# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1754 gnd d1 a_20283_7400# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1755 a_8539_196# d7 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1756 a_17814_3888# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1757 a_5061_5925# a_4843_5925# a_4572_6031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1758 a_26267_3001# d0 a_26756_2895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1759 a_28711_4561# a_28968_4371# a_28616_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1760 a_13284_4238# d0 a_13765_4326# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1761 a_2463_2078# d1 a_2545_1470# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1762 a_22359_1865# a_22141_1865# a_21870_1971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1763 a_31172_6374# d1 a_31958_5701# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1764 vdd d0 a_8017_4575# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1765 a_19097_377# a_18915_4522# a_18957_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1766 a_6785_2934# d2 a_6864_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1767 a_9240_6955# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1768 a_2540_5973# a_2793_5960# a_2490_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1769 a_17813_4300# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1770 a_3364_2127# a_3617_2114# a_2562_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1771 a_32036_6598# a_31834_5582# a_31953_5172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1772 a_13749_2896# a_13531_2896# a_13258_2709# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1773 a_6946_3519# a_7203_3329# a_6864_4127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1774 a_26274_3219# d0 a_26755_3307# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1775 a_8857_854# a_8859_953# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1776 a_18594_3098# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1777 a_27507_7605# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1778 a_4543_4213# d0 a_5024_4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1779 a_13822_6968# a_13604_6968# a_13331_6781# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1780 gnd d1 a_7239_5365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1781 a_13748_3308# a_13530_3308# a_13273_3403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1782 a_18936_6679# a_18766_7580# a_18885_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1783 gnd d0 a_16815_7242# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1784 a_24239_3962# d1 a_24334_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1785 a_7801_6212# a_8054_6199# a_6999_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1786 a_23461_390# a_23279_4535# a_23321_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1787 gnd d1 a_33315_3366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1788 a_9348_847# a_9130_847# a_8857_854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1789 vdd d0 a_21080_7628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1790 a_17556_4395# d0 a_18031_4300# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1791 vdd d0 a_16831_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1792 a_15599_7031# d2 a_15678_8224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1793 vdd d4 a_24306_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1794 a_30601_1196# a_30607_1379# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1795 a_26029_208# d7 a_17148_133# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1796 a_27677_6704# a_27507_7605# a_27631_7724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1797 vdd d3 a_7111_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1798 a_26370_8492# d0 a_26845_8397# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1799 a_1285_1460# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1800 a_7743_3747# a_7747_3570# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1801 a_25204_8849# a_25461_8659# a_24411_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1802 vdd d1 a_20227_4346# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1803 a_24390_7603# d0 a_25188_7419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1804 a_9146_2277# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1805 a_3456_7629# a_3709_7616# a_2659_7401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1806 a_19792_2933# d2 a_19875_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1807 a_2463_2078# d1 a_2549_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1808 a_26554_4325# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1809 a_1368_2476# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1810 a_155_2964# a_162_3182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1811 a_30661_4433# d0 a_31136_4338# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1812 a_12215_8260# a_12210_8849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1813 a_11323_3531# d0 a_12125_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1814 a_3360_2304# a_3617_2114# a_2562_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1815 a_30717_7487# d0 a_31192_7392# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1816 a_20807_6623# a_21060_6610# a_20010_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1817 a_26333_6456# a_26338_6780# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1818 a_30734_8505# a_29585_8684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1819 a_26829_6967# a_26611_6967# a_26340_7073# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1820 a_23337_271# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1821 vdd d1 a_7239_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1822 vdd d0 a_16815_7242# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1823 a_10233_2620# d3 a_10327_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1824 a_20006_6572# d0 a_20804_6388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1825 vdd d1 a_33315_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1826 a_25115_3347# a_25372_3157# a_24317_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1827 a_6868_3950# d1 a_6967_4360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1828 a_9347_1259# d1 a_10145_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1829 a_30901_3320# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1830 a_26772_4325# a_26554_4325# a_26297_4420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1831 a_4987_2265# d1 a_5773_1592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1832 a_31192_7392# d1 a_31990_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1833 vout a_17029_133# a_17148_133# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1834 a_15599_7031# d2 a_15682_8047# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1835 a_6827_2091# d1 a_6913_1306# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1836 gnd d0 a_12467_8659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1837 a_19911_5985# a_20164_5972# a_19861_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1838 a_17569_5230# d0 a_18050_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1839 a_462_4894# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1840 a_388_1234# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1841 a_13511_1878# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1842 a_11400_7426# a_11653_7413# a_11314_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1843 a_4971_835# a_4753_835# a_4480_842# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1844 a_13493_1272# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1845 a_17506_1958# a_17513_2176# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1846 a_5640_6153# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1847 a_461_5306# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1848 a_29512_4612# a_29765_4599# a_28715_4384# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1849 a_21907_4007# a_21914_4225# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1850 a_13510_2290# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1851 a_3452_7806# a_3709_7616# a_2659_7401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1852 a_21926_5025# d0 a_22415_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1853 a_5841_5135# a_5623_5135# a_5044_4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1854 a_14291_1088# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1855 a_624_1840# a_406_1840# a_135_1946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1856 a_7747_3570# a_8000_3557# a_6950_3342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1857 a_12157_5383# a_12161_5206# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1858 a_20754_3569# a_20768_4352# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1859 a_20803_6800# a_21060_6610# a_20010_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1860 a_18647_6152# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1861 a_14665_6586# a_14463_5570# a_14582_5160# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1862 a_28430_4996# a_28683_4983# a_27833_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1863 a_18957_2488# a_18739_2488# a_18858_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1864 a_32943_1951# a_33196_1938# a_32893_3148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1865 a_2676_8419# d0 a_3469_8824# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1866 gnd d0 a_12378_3157# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1867 a_20840_8836# a_20844_8659# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1868 a_13240_1984# a_13247_2202# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1869 a_3364_2127# a_3359_2716# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1870 gnd d1 a_33368_6420# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1871 a_18915_4522# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1872 a_30618_2214# a_30624_2397# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1873 a_28606_7030# a_28859_7017# a_28430_4996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1874 a_1726_365# a_1544_4510# a_1586_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1875 a_33818_1748# a_34075_1558# a_33025_1343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1876 vdd d0 a_7981_2127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1877 a_13221_867# a_16448_1324# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1878 gnd d1 a_7220_4347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1879 a_644_2858# d1 a_1441_3086# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1880 vdd d1 a_15907_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1881 vdd d0 a_8054_6199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1882 a_10150_1604# a_9944_2093# a_9365_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1883 a_11396_7603# a_11653_7413# a_11314_8211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1884 a_7727_2552# a_7744_3335# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1885 a_10182_3111# d2 a_10233_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1886 gnd d1 a_7293_8419# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1887 a_26591_5949# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1888 a_19957_3341# a_20210_3328# a_19871_4126# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1889 a_2582_3506# d0 a_3380_3322# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1890 a_7706_1711# a_7710_1534# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1891 a_4495_1342# a_4497_1860# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1892 vdd d3 a_15779_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1893 a_21933_5243# a_21939_5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1894 a_22196_5331# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1895 a_2549_1293# d0 a_3342_1698# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1896 a_10255_7183# d2 a_10306_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1897 a_18067_6336# a_17849_6336# a_17592_6431# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1898 a_32020_4560# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1899 a_15744_6421# a_15997_6408# a_15645_6011# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1900 gnd d4 a_19942_4958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1901 a_14831_403# d5 a_12951_197# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1902 a_241_7437# d0 a_716_7342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1903 a_19097_377# d5 a_19191_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1904 a_11318_8034# d1 a_11413_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1905 a_22358_2277# d1 a_23144_1604# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1906 a_153_2671# d0 a_644_2858# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1907 a_28734_5402# a_28987_5389# a_28648_6187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1908 a_24198_2103# d1 a_24284_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1909 a_14551_3653# d2 a_14597_2633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1910 a_20845_8247# a_21098_8234# a_20043_8608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1911 a_26355_7992# a_26357_8091# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1912 a_2676_8419# d0 a_3473_8647# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1913 a_8967_6768# a_8969_7061# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1914 a_22432_5937# a_22214_5937# a_21941_5944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1915 a_18693_3508# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1916 a_4622_8468# d0 a_5097_8373# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1917 vdd d1 a_33368_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1918 a_14427_3534# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1919 a_24411_8444# a_24664_8431# a_24312_8034# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1920 a_22414_5331# a_22196_5331# a_21939_5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1921 a_32135_6598# d4 a_32202_415# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1922 a_23139_1075# a_22921_1075# a_22342_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1923 gnd d3 a_15852_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1924 a_3433_6376# a_3437_6199# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1925 a_31100_1890# d1 a_31885_1629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1926 a_9257_7973# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1927 a_32135_6598# a_31917_6598# a_32036_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1928 a_31156_4944# d1 a_31953_5172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1929 a_14500_7606# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1930 a_6085_259# d5 a_4210_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1931 a_23212_5147# a_22994_5147# a_22415_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1932 a_18032_3888# d1 a_18817_3627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1933 a_9256_8385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1934 a_4806_4301# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1935 gnd d0 a_3690_6186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1936 a_18051_4906# a_17833_4906# a_17562_5012# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1937 a_29475_2576# a_29492_3359# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1938 a_18863_2607# a_18693_3508# a_18817_3627# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1939 a_30592_879# a_33819_1336# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1940 a_33933_7267# a_34186_7254# a_33131_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1941 a_17526_2976# d0 a_18015_2870# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1942 a_2582_3506# d0 a_3384_3145# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1943 a_11245_3962# d1 a_11344_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1944 a_29564_7843# a_29568_7666# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1945 a_499_6930# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1946 a_185_4383# a_189_4901# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1947 a_7800_6624# a_8053_6611# a_7003_6396# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1948 a_17533_3194# d0 a_18014_3282# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1949 a_2655_7578# d0 a_3457_7217# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1950 a_11318_8034# d1 a_11417_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1951 gnd d0 a_25462_8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1952 a_13604_6968# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1953 a_15727_5403# d0 a_16520_5808# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1954 a_5024_4301# a_4806_4301# a_4549_4396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1955 a_31099_2302# a_30881_2302# a_30618_2214# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1956 a_21890_2989# d0 a_22379_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1957 a_20841_8424# a_21098_8234# a_20043_8608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1958 vdd d2 a_28905_5997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1959 a_9167_2883# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1960 a_6999_6573# d0 a_7797_6389# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1961 vdd d0 a_29765_4599# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1962 a_12832_197# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1963 a_733_8360# a_515_8360# a_252_8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1964 a_1441_6548# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1965 a_5810_3628# a_5604_4117# a_5025_3889# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1966 a_16452_1147# a_16705_1134# a_15650_1508# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1967 a_27589_5159# d2 a_27672_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1968 a_13284_4238# a_13290_4421# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X1969 a_24407_8621# a_24664_8431# a_24312_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1970 a_21963_7061# d0 a_22452_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1971 a_21897_3207# d0 a_22378_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1972 a_28652_6010# d1 a_28747_6597# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1973 a_661_3876# a_443_3876# a_172_3982# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1974 a_12124_3582# a_12377_3569# a_11327_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1975 a_6904_5986# a_7157_5973# a_6854_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1976 a_26772_4325# d1 a_27558_3652# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1977 a_6900_6163# d1 a_6982_5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1978 a_27604_2632# a_27434_3533# a_27553_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1979 a_32980_3987# a_33233_3974# a_32897_2971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1980 vdd d0 a_3690_6186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1981 a_13494_860# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1982 a_26845_8397# d1 a_27631_7724# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1983 vdd d0 a_3673_5168# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1984 vdd d1 a_11543_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1985 a_33929_7444# a_34186_7254# a_33131_7628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1986 a_14624_7725# a_14418_8214# a_13839_7986# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1987 a_142_2164# d0 a_623_2252# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1988 a_27425_8213# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1989 a_23300_6692# a_23130_7593# a_23254_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1990 a_7796_6801# a_8053_6611# a_7003_6396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1991 a_20010_6395# d0 a_20803_6800# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1992 a_21978_7980# d0 a_22469_7973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1993 a_33025_1343# a_33278_1330# a_32939_2128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1994 a_22177_4313# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1995 a_31789_8226# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1996 gnd d0 a_34165_6648# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1997 a_4753_835# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X1998 a_17977_1246# d1 a_18775_1062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X1999 gnd d0 a_21044_5180# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2000 a_16448_1324# a_16705_1134# a_15650_1508# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2001 a_4091_172# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2002 gnd d1 a_24554_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2003 a_13729_1878# d1 a_14514_1617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2004 a_4843_5925# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2005 a_11231_7195# d2 a_11281_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2006 a_9365_1865# a_9147_1865# a_8874_1872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2007 a_13350_8092# a_13357_8310# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2008 a_27672_6585# d3 a_27771_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2009 a_27714_283# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2010 a_3363_2539# a_3380_3322# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2011 vdd d0 a_29839_8259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2012 a_1404_1050# a_1186_1050# a_607_822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2013 a_26719_859# d1 a_27516_1087# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2014 a_235_7254# a_241_7437# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2015 a_6900_6163# d1 a_6986_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2016 a_33098_5415# d0 a_33891_5820# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2017 a_29532_5218# a_29527_5807# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2018 a_18630_5134# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2019 a_31834_5582# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2020 a_17550_4212# a_17556_4395# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2021 a_15667_2526# d0 a_16465_2342# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2022 a_6950_3342# a_7203_3329# a_6864_4127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2023 a_22395_4313# a_22177_4313# a_21920_4408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2024 a_5061_5925# d1 a_5846_5664# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2025 a_1395_7568# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2026 a_24271_6175# a_24528_5985# a_24225_7195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2027 a_11344_4372# d0 a_12137_4777# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2028 a_28657_1507# d0 a_29455_1323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2029 gnd d4 a_6935_4959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2030 a_16502_4378# a_16506_4201# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2031 a_19937_2323# d0 a_20734_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2032 gnd d0 a_34076_1146# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2033 a_30865_872# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2034 a_30629_2721# a_30631_3014# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2035 a_23181_3640# a_22975_4129# a_22396_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2036 a_3419_5593# a_3672_5580# a_2622_5365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2037 a_170_3883# a_172_3982# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2038 a_20010_6395# d0 a_20807_6623# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2039 a_29527_5807# a_29531_5630# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2040 a_5567_2081# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2041 a_25119_3170# a_25114_3759# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2042 a_22994_5147# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2043 gnd d0 a_3654_4150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2044 a_148_2347# a_153_2671# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2045 gnd d0 a_21080_7628# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2046 a_32893_3148# d2 a_32939_2128# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2047 a_25135_4600# a_25388_4587# a_24338_4372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2048 a_12104_2564# a_12121_3347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2049 a_15764_7439# a_16017_7426# a_15678_8224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2050 a_118_928# d0 a_607_822# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2051 a_33021_1520# a_33278_1330# a_32939_2128# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2052 a_26267_3001# a_26274_3219# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2053 a_25208_8672# a_25461_8659# a_24411_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2054 vdd d0 a_21044_5180# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2055 a_33094_5592# a_33351_5402# a_33012_6200# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2056 vdd d1 a_24554_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2057 a_27698_2513# d4 a_27838_402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2058 a_33025_1343# d0 a_33822_1571# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2059 a_27315_2105# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2060 a_15764_7439# d0 a_16557_7844# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2061 a_221_6419# a_226_6743# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2062 a_13357_8310# a_13363_8493# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2063 a_31953_5172# d2 a_32036_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2064 a_18780_1591# a_18574_2080# a_17995_1852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2065 a_11323_3531# d0 a_12121_3347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2066 a_4536_3995# d0 a_5025_3889# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2067 a_30955_5962# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2068 a_19916_1482# d0 a_20718_1121# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2069 a_15667_2526# d0 a_16469_2165# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2070 a_15609_3975# a_15862_3962# a_15526_2959# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2071 a_33016_6023# d1 a_33111_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2072 a_33098_5415# d0 a_33895_5643# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2073 vdd d3 a_11415_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2074 a_4309_172# d7 a_8757_196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2075 a_11380_6408# a_11633_6395# a_11281_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2076 a_8986_8079# a_8993_8297# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2077 a_28657_1507# d0 a_29459_1146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2078 a_31679_2118# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2079 a_16525_5219# a_16520_5808# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2080 vdd d0 a_34076_1146# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2081 vdd d0 a_25408_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2082 a_27521_1616# a_27315_2105# a_26735_2289# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2083 a_25119_3170# a_25372_3157# a_24317_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2084 a_20841_8424# a_20845_8247# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2085 a_6868_3950# d1 a_6963_4537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2086 a_4790_2871# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2087 a_19689_4971# d3 a_19861_7182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2088 a_3415_5770# a_3672_5580# a_2622_5365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2089 a_1223_3086# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2090 a_30609_1897# d0 a_31100_1890# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2091 a_22214_5937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2092 vdd d0 a_3654_4150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2093 a_10063_3521# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2094 a_17612_7449# d0 a_18087_7354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2095 a_30665_4951# d0 a_31156_4944# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2096 a_425_3270# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2097 a_243_7955# d0 a_734_7948# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2098 a_15760_7616# a_16017_7426# a_15678_8224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2099 a_4607_7968# a_4609_8067# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2100 a_15419_5174# d3 a_15526_2959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2101 a_31885_1629# a_31679_2118# a_31099_2302# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2102 a_26274_3219# a_26280_3402# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2103 a_499_6930# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2104 a_31953_5172# a_31735_5172# a_31155_5356# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2105 a_13548_3914# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2106 a_32943_1951# d1 a_33042_2361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2107 a_8911_3908# d0 a_9402_3901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2108 a_15764_7439# d0 a_16561_7667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2109 a_31958_5701# a_31752_6190# a_31172_6374# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2110 a_21976_7462# d0 a_22451_7367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2111 a_7707_1299# a_7711_1122# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2112 a_20790_5605# a_21043_5592# a_19993_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2113 a_8757_196# a_8539_196# a_4309_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2114 vdd d0 a_12468_8247# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2115 gnd d0 a_21025_4162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2116 a_624_1840# d1 a_1409_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2117 gnd d0 a_34202_8684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2118 a_33016_6023# d1 a_33115_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2119 a_31082_1284# a_30864_1284# a_30607_1379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2120 a_18015_2870# a_17797_2870# a_17524_2683# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2121 a_33131_7628# d0 a_33929_7444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2122 a_14328_3124# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2123 a_1487_2476# a_1285_1460# a_1409_1579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2124 vdd d2 a_2830_7996# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2125 a_9458_6955# a_9240_6955# a_8969_7061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2126 a_697_5912# d1 a_1482_5651# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2127 a_10099_5557# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2128 a_11162_2946# d2 a_11245_3962# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2129 a_7003_6396# d0 a_7796_6801# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2130 a_13766_3914# d1 a_14551_3653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2131 a_4880_7961# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2132 a_4825_5319# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2133 a_18014_3282# a_17796_3282# a_17539_3377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2134 a_20735_2139# a_20730_2728# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2135 a_33079_4397# d0 a_33872_4802# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2136 a_18611_4116# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2137 a_11208_1926# a_11461_1913# a_11158_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2138 a_23456_271# d5 a_21581_184# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2139 a_133_1847# a_135_1946# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2140 a_26756_2895# d1 a_27553_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2141 gnd d0 a_7981_2127# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2142 a_33822_1571# a_34075_1558# a_33025_1343# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2143 a_28533_2958# d2 a_28612_4151# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2144 a_33950_8285# a_33945_8874# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2145 a_20043_8608# a_20300_8418# a_19948_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2146 a_17586_6248# a_17592_6431# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2147 a_24235_4139# a_24492_3949# a_24156_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2148 gnd d0 a_8037_5181# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2149 a_17029_133# d8 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2150 a_14546_3124# a_14328_3124# a_13748_3308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2151 gnd d2 a_24565_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2152 a_24334_4549# d0 a_25132_4365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2153 gnd d1 a_15907_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2154 a_26260_2384# d0 a_26735_2289# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2155 gnd d0 a_34113_3182# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2156 vdd d0 a_3689_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2157 a_10301_6573# a_10099_5557# a_10223_5676# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2158 a_3400_4575# a_3653_4562# a_2603_4347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2159 a_5043_5319# a_4825_5319# a_4568_5414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2160 a_13320_6274# d0 a_13801_6362# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2161 a_22975_4129# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2162 a_6854_7183# d2 a_6900_6163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2163 a_31173_5962# a_30955_5962# a_30684_6068# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2164 a_15723_5580# a_15980_5390# a_15641_6188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2165 a_18104_8372# a_17886_8372# a_17623_8284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2166 a_26320_6055# d0 a_26809_5949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2167 a_19944_8198# d1 a_20030_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2168 a_17849_6336# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2169 a_7783_5606# a_7797_6389# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2170 a_14592_2514# a_14390_1498# a_14509_1088# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2171 a_26628_7985# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2172 a_26310_5255# d0 a_26791_5343# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2173 a_22161_2883# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2174 a_13801_6362# d1 a_14587_5689# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2175 a_13320_6274# a_13326_6457# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2176 a_23212_5147# d2 a_23295_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2177 a_4555_5013# d0 a_5044_4907# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2178 vdd d0 a_21025_4162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2179 a_10260_7712# a_10054_8201# a_9475_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2180 vdd d0 a_34202_8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2181 a_33131_7628# d0 a_33933_7267# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2182 a_27470_5569# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2183 a_26791_5343# d1 a_27589_5159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2184 a_23020_1485# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2185 a_22160_3295# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2186 vdd d3 a_28859_7017# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2187 gnd d1 a_33351_5402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2188 a_22468_8385# a_22250_8385# a_21987_8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2189 a_11363_5390# d0 a_12160_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2190 a_9420_5331# a_9202_5331# a_8939_5243# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2191 a_7003_6396# d0 a_7800_6624# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2192 a_23227_2620# a_23057_3521# a_23176_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2193 a_27352_4141# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2194 a_8949_6043# a_8956_6261# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2195 a_31136_4338# d1 a_31922_3665# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2196 gnd d2 a_7084_1901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2197 a_16469_2165# a_16464_2754# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2198 a_22468_8385# d1 a_23254_7712# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2199 a_189_4901# d0 a_680_4894# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2200 a_33079_4397# d0 a_33876_4625# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2201 a_2577_8009# a_2830_7996# a_2494_6993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2202 a_17513_2176# d0 a_17994_2264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2203 a_5950_2489# d4 a_6090_378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2204 a_13294_4939# d0 a_13785_4932# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2205 a_31209_8410# a_30991_8410# a_30734_8505# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2206 a_25150_5795# a_25407_5605# a_24357_5390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2207 vdd d0 a_8037_5181# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2208 a_17539_3377# a_17541_3895# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2209 a_9365_1865# d1 a_10150_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2210 a_24334_4549# d0 a_25136_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2211 vdd d2 a_24565_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2212 a_16541_6649# a_16558_7432# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2213 a_19191_258# a_18973_258# a_19092_258# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2214 a_3384_3145# a_3379_3734# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2215 a_10400_6573# a_10182_6573# a_10301_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2216 a_19861_7182# d2 a_19911_5985# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2217 a_17833_4906# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2218 vdd d0 a_34113_3182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2219 a_3396_4752# a_3653_4562# a_2603_4347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2220 a_27558_3652# a_27352_4141# a_26772_4325# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2221 a_4570_5932# a_4572_6031# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2222 a_4570_5932# d0 a_5061_5925# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2223 a_20803_6800# a_20807_6623# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2224 a_11245_3962# d1 a_11340_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2225 a_21877_2189# d0 a_22358_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2226 a_26237_1183# a_26243_1366# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2227 a_22251_7973# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2228 a_24374_6408# d0 a_25167_6813# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2229 a_6909_1483# d0 a_7711_1122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2230 a_20771_4587# a_20787_5370# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2231 gnd d0 a_16758_4600# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2232 a_19834_2090# a_20091_1900# a_19788_3110# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2233 a_18051_4906# d1 a_18848_5134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2234 a_2622_5365# a_2875_5352# a_2536_6150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2235 a_25131_4777# a_25135_4600# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2236 a_5846_5664# a_5640_6153# a_5060_6337# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2237 a_23300_6692# d3 a_23394_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2238 a_10467_390# d5 a_10561_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2239 gnd d0 a_29748_3581# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2240 a_1820_246# d6 a_4309_172# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2241 a_26808_6361# a_26590_6361# a_26333_6456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2242 a_12210_8849# a_12467_8659# a_11417_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2243 a_27656_4547# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2244 a_27553_6585# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2245 a_5061_5925# a_4843_5925# a_4570_5932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2246 a_20771_4587# a_21024_4574# a_19974_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2247 a_8956_6261# a_8962_6444# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2248 a_32036_6598# d3 a_32135_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2249 a_5810_3628# d2 a_5856_2608# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2250 a_9240_6955# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2251 a_27594_5688# a_27388_6177# a_26809_5949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2252 a_24280_1495# d0 a_25078_1311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2253 a_13346_7475# a_13348_7993# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2254 a_15678_8224# d1 a_15760_7616# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2255 a_4789_3283# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2256 a_1296_7158# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2257 a_14826_284# d4 a_15423_4997# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2258 a_33913_6249# a_33908_6838# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2259 gnd d0 a_3673_5168# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2260 a_4862_7355# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2261 a_697_5912# a_479_5912# a_208_6018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2262 gnd d0 a_16742_3170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2263 a_27838_402# a_27656_4547# a_27771_6585# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2264 a_31662_1100# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2265 a_19865_7005# d2 a_19944_8198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2266 a_3453_7394# a_3457_7217# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2267 a_226_6743# a_228_7036# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2268 a_7783_5606# a_8036_5593# a_6986_5378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2269 a_12121_3347# a_12378_3157# a_11323_3531# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2270 a_5025_3889# a_4807_3889# a_4534_3896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2271 a_24374_6408# d0 a_25171_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2272 gnd d0 a_8018_4163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2273 a_14707_284# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2274 a_33859_3607# a_34112_3594# a_33062_3379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2275 a_1514_7158# a_1296_7158# a_716_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2276 a_2618_5542# a_2875_5352# a_2536_6150# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2277 a_2421_2921# d2 a_2504_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2278 a_19948_8021# a_20201_8008# a_19865_7005# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2279 a_26792_4931# a_26574_4931# a_26303_5037# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2280 a_12194_7419# a_12451_7229# a_11396_7603# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2281 a_29528_5395# a_29532_5218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2282 gnd d1 a_28968_4371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2283 vdd d0 a_29748_3581# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2284 a_31082_1284# d1 a_31880_1100# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2285 a_5805_3099# a_5587_3099# a_5008_2871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2286 a_1477_5122# d2 a_1560_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2287 a_31155_5356# a_30937_5356# a_30674_5268# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2288 gnd d0 a_12357_2551# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2289 a_17886_8372# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2290 a_2540_5973# d1 a_2635_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2291 a_20767_4764# a_21024_4574# a_19974_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2292 a_8857_854# d0 a_9348_847# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2293 a_21897_3207# a_21903_3390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2294 a_8956_6261# d0 a_9437_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2295 a_13839_7986# a_13621_7986# a_13348_7993# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2296 a_29532_5218# a_29785_5205# a_28730_5579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2297 a_24280_1495# d0 a_25082_1134# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2298 gnd d0 a_29839_8259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2299 a_18684_8188# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2300 a_15678_8224# d1 a_15764_7439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2301 a_7797_6389# a_7801_6212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2302 a_26829_6967# a_26611_6967# a_26338_6780# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2303 a_19993_5377# a_20246_5364# a_19907_6162# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2304 a_9401_4313# a_9183_4313# a_8920_4225# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2305 a_5649_1473# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2306 a_26282_3920# a_26284_4019# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2307 a_13838_8398# a_13620_8398# a_13363_8493# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2308 gnd d3 a_24409_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2309 a_17524_2683# a_17526_2976# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2310 a_33855_3784# a_33859_3607# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2311 a_13348_7993# a_13350_8092# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2312 gnd d1 a_33405_8456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2313 a_17614_7967# d0 a_18105_7960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2314 a_24353_5567# d0 a_25155_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2315 a_26370_8492# a_25208_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2316 a_14619_7196# a_14401_7196# a_13822_6968# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2317 a_9927_1075# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2318 vdd d0 a_16742_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2319 a_6937_8199# d1 a_7023_7414# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2320 a_19937_2323# d0 a_20730_2728# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2321 a_5722_5545# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2322 a_5043_5319# d1 a_5841_5135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2323 a_13294_4939# a_13296_5038# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2324 a_19993_5377# d0 a_20786_5782# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2325 a_13275_3921# d0 a_13766_3914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2326 a_10000_5147# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2327 vdd d0 a_8018_4163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2328 a_23031_7183# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2329 a_19861_7182# a_20118_6992# a_19689_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2330 a_14587_5689# d2 a_14665_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2331 a_26719_859# a_26501_859# a_26228_866# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2332 a_13238_1885# d0 a_13729_1878# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2333 a_17814_3888# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2334 gnd d2 a_11534_5985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2335 a_18729_5544# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2336 gnd d0 a_20971_1108# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2337 a_26265_2708# d0 a_26756_2895# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2338 a_17870_6942# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2339 vdd d1 a_28968_4371# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2340 a_13749_2896# a_13531_2896# a_13260_3002# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2341 gnd d1 a_24537_1305# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2342 a_12160_5618# a_12174_6401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2343 vdd d0 a_12357_2551# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2344 a_2540_5973# d1 a_2639_6383# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2345 a_2603_4347# a_2856_4334# a_2504_3937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2346 a_11413_8621# d0 a_12215_8260# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2347 a_17148_133# d8 vout vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2348 a_10182_3111# a_9964_3111# a_9384_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2349 a_1203_2068# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2350 a_33025_1343# d0 a_33818_1748# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2351 gnd d1 a_7183_2311# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2352 a_1659_6548# a_1441_6548# a_1560_6548# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2353 a_13785_4932# d1 a_14582_5160# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2354 a_18931_6560# a_18729_5544# a_18853_5663# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2355 a_15568_2116# a_15825_1926# a_15522_3136# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2356 a_20787_5370# a_20791_5193# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2357 a_13290_4421# a_13294_4939# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2358 a_15595_7208# d2 a_15641_6188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2359 a_19989_5554# a_20246_5364# a_19907_6162# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2360 a_18780_1591# d2 a_18858_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2361 a_25205_8437# a_25462_8247# a_24407_8621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2362 a_22379_2883# d1 a_23176_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2363 vdd d1 a_33405_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2364 a_4970_1247# a_4752_1247# a_4489_1159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2365 a_30991_8410# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2366 a_22451_7367# a_22233_7367# a_21976_7462# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2367 a_3346_1521# a_3599_1508# a_2549_1293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2368 a_32041_6717# a_31871_7618# a_31990_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2369 a_6827_2091# a_7084_1901# a_6781_3111# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2370 vdd d3 a_24482_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2371 a_4482_941# a_4489_1159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2372 a_17776_2264# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2373 a_2490_7170# a_2747_6980# a_2318_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2374 a_32794_5009# d3 a_32966_7220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2375 a_19911_5985# d1 a_20006_6572# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2376 a_5908_4523# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2377 a_478_6324# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2378 a_118_928# a_125_1146# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2379 a_16488_3595# a_16741_3582# a_15691_3367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2380 a_26518_1877# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2381 a_10218_5147# a_10000_5147# a_9421_4919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2382 a_13583_6362# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2383 a_679_5306# a_461_5306# a_198_5218# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2384 a_6678_5149# a_6935_4959# a_6085_259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2385 a_7764_4588# a_8017_4575# a_6967_4360# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2386 a_26591_5949# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2387 a_26517_2289# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2388 a_3415_5770# a_3419_5593# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2389 a_20718_1121# a_20713_1710# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2390 a_31922_3665# a_31716_4154# a_31137_3926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2391 a_13784_5344# a_13566_5344# a_13303_5256# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2392 a_24338_4372# d0 a_25135_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2393 a_21914_4225# a_21920_4408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2394 a_17577_5931# a_17579_6030# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2395 a_26573_5343# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2396 a_27298_1087# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2397 a_17994_2264# a_17776_2264# a_17519_2359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2398 a_14381_6178# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2399 a_2599_4524# a_2856_4334# a_2504_3937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2400 a_31880_1100# d2 a_31963_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2401 a_23093_5557# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2402 a_26228_866# a_29455_1323# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2403 a_26773_3913# a_26555_3913# a_26284_4019# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2404 a_17569_5230# a_17575_5413# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2405 a_26736_1877# a_26518_1877# a_26247_1983# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2406 a_32943_1951# d1 a_33038_2538# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2407 vdd d1 a_7183_2311# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2408 a_21970_7279# a_21976_7462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2409 vdd d2 a_20164_5972# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2410 a_33012_6200# d1 a_33094_5592# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2411 a_27371_5159# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2412 gnd d0 a_12468_8247# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2413 a_19030_6560# a_18812_6560# a_18931_6560# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2414 a_17560_4913# d0 a_18051_4906# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2415 a_9239_7367# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2416 a_1492_2595# a_1322_3496# a_1441_3086# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2417 a_33818_1748# a_33822_1571# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2418 a_462_4894# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2419 a_29513_4200# a_29766_4187# a_28711_4561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2420 a_30607_1379# a_30609_1897# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2421 a_33908_6838# a_34165_6648# a_33115_6433# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2422 a_8945_5426# a_8947_5944# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2423 a_172_3982# a_179_4200# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2424 a_32794_5009# d3 a_32970_7043# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2425 a_19911_5985# d1 a_20010_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2426 a_19974_4359# a_20227_4346# a_19875_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2427 a_25910_208# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2428 a_7748_3158# a_8001_3145# a_6946_3519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2429 vdd d1 a_15997_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2430 a_28529_3135# d2 a_28579_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2431 a_16484_3772# a_16741_3582# a_15691_3367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2432 a_12083_1723# a_12087_1546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2433 a_20804_6388# a_21061_6198# a_20006_6572# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2434 a_20047_8431# a_20300_8418# a_19948_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2435 a_2672_8596# d0 a_3470_8412# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2436 a_18051_4906# a_17833_4906# a_17560_4913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2437 vdd d1 a_28987_5389# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2438 a_7760_4765# a_8017_4575# a_6967_4360# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2439 a_19974_4359# d0 a_20767_4764# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2440 a_2639_6383# d0 a_3432_6788# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2441 a_170_3883# d0 a_661_3876# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2442 a_9981_4129# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2443 a_15708_4385# d0 a_16501_4790# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2444 a_13273_3403# d0 a_13748_3308# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2445 a_5856_2608# a_5686_3509# a_5805_3099# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2446 a_245_8054# a_252_8272# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2447 a_12087_1546# a_12340_1533# a_11290_1318# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2448 a_31968_2645# d3 a_32062_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2449 a_10462_271# d4 a_11059_4984# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2450 a_6678_5149# d3 a_6781_3111# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2451 a_29491_3771# a_29495_3594# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2452 a_28698_3366# d0 a_29491_3771# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2453 a_13604_6968# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2454 a_6986_5378# a_7239_5365# a_6900_6163# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2455 a_18766_7580# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2456 a_24275_5998# d1 a_24374_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2457 gnd d0 a_25444_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2458 a_23279_4535# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2459 a_33062_3379# a_33315_3366# a_32976_4164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2460 a_643_3270# a_425_3270# a_168_3365# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2461 a_19097_377# a_18915_4522# a_19030_6560# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2462 a_25132_4365# a_25136_4188# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2463 gnd d3 a_28859_7017# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2464 a_23217_5676# a_23011_6165# a_22432_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2465 a_6986_5378# d0 a_7779_5783# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2466 a_24049_5161# a_24306_4971# a_23456_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2467 gnd d4 a_33047_4996# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2468 vdd d0 a_25352_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2469 a_14670_6705# a_14500_7606# a_14619_7196# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2470 a_27507_7605# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2471 a_2545_1470# d0 a_3343_1286# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2472 a_33062_3379# d0 a_33855_3784# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2473 a_18068_5924# a_17850_5924# a_17579_6030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2474 gnd d1 a_11560_2323# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2475 a_19970_4536# a_20227_4346# a_19875_3949# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2476 a_19953_3518# d0 a_20751_3334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2477 a_7744_3335# a_8001_3145# a_6946_3519# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2478 a_23461_390# a_23279_4535# a_23394_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2479 a_8947_5944# a_8949_6043# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2480 a_17616_8066# d0 a_18105_7960# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2481 a_9348_847# a_9130_847# a_8859_953# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2482 a_2672_8596# d0 a_3474_8235# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2483 a_19974_4359# d0 a_20771_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2484 a_6864_4127# a_7121_3937# a_6785_2934# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2485 a_3400_4575# a_3416_5358# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2486 a_28678_2348# a_28931_2335# a_28579_1938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2487 a_8889_2372# d0 a_9364_2277# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2488 a_12083_1723# a_12340_1533# a_11290_1318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2489 a_3359_2716# a_3363_2539# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2490 a_14509_1088# d2 a_14592_2514# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2491 a_7723_2729# a_7980_2539# a_6930_2324# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2492 vdd d0 a_25371_3569# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2493 a_10187_3640# a_9981_4129# a_9402_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2494 a_18087_7354# d1 a_18885_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2495 a_28698_3366# d0 a_29495_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2496 a_6982_5555# a_7239_5365# a_6900_6163# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2497 a_9146_2277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2498 a_21980_8079# d0 a_22469_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2499 a_10255_7183# a_10037_7183# a_9458_6955# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2500 vdd d0 a_25444_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2501 a_30691_6286# a_30697_6469# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2502 a_15641_6188# d1 a_15723_5580# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2503 a_2318_4959# a_2571_4946# a_1721_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2504 a_33058_3556# a_33315_3366# a_32976_4164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2505 a_679_5306# d1 a_1477_5122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2506 a_13765_4326# a_13547_4326# a_13284_4238# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2507 a_26554_4325# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2508 a_7747_3570# a_7761_4353# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2509 a_9347_1259# a_9129_1259# a_8866_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2510 a_30655_4250# d0 a_31136_4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2511 a_21987_8297# d0 a_22468_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2512 gnd d0 a_20970_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2513 a_7833_8837# a_7837_8660# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2514 a_6904_5986# d1 a_6999_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2515 a_13712_860# a_13494_860# a_13221_867# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2516 a_26755_3307# a_26537_3307# a_26274_3219# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2517 a_12214_8672# a_12467_8659# a_11417_8444# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2518 a_17978_834# a_17760_834# a_17487_841# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2519 a_22451_7367# d1 a_23249_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2520 a_32980_3987# d1 a_33075_4574# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2521 vdd d0 a_3600_1096# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2522 a_4843_5925# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2523 vdd d1 a_11560_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2524 a_15423_4997# d3 a_15599_7031# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2525 gnd d0 a_16794_6636# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2526 a_25082_1134# a_25077_1723# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2527 a_25098_2564# a_25351_2551# a_24301_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2528 a_10228_2501# d3 a_10327_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2529 a_24049_5161# d3 a_24152_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2530 vdd d1 a_11616_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2531 a_19953_3518# d0 a_20755_3157# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2532 gnd d3 a_2674_2908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2533 a_9348_847# d1 a_10145_1075# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2534 vdd d1 a_11633_6395# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2535 a_29527_5807# a_29784_5617# a_28734_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2536 vdd d2 a_2720_1888# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2537 a_10400_6573# d4 a_10467_390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2538 vout a_17029_133# a_8757_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2539 a_22958_3111# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2540 a_31193_6980# d1 a_31990_7208# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2541 a_5623_5135# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2542 a_406_1840# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2543 vdd d0 a_29766_4187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2544 vdd d2 a_7194_8009# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2545 a_32970_7043# d2 a_33049_8236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2546 a_10561_271# a_10343_271# a_10462_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2547 a_14463_5570# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2548 a_18973_258# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2549 a_13511_1878# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2550 a_28674_2525# a_28931_2335# a_28579_1938# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2551 a_21888_2696# d0 a_22379_2883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2552 a_29508_4789# a_29512_4612# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2553 a_4971_835# a_4753_835# a_4482_941# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2554 a_33856_3372# a_33860_3195# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2555 vdd d2 a_7157_5973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2556 a_12125_3170# a_12378_3157# a_11323_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2557 a_20828_7229# a_20823_7818# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2558 gnd d2 a_15898_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2559 vdd d2 a_33233_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2560 a_33115_6433# a_33368_6420# a_33016_6023# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2561 a_18858_2488# a_18656_1472# a_18775_1062# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2562 a_27932_283# a_27714_283# a_27833_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2563 a_15691_3367# a_15944_3354# a_15605_4152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2564 a_12198_7242# a_12451_7229# a_11396_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2565 a_5841_5135# a_5623_5135# a_5043_5319# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2566 a_20734_2551# a_20751_3334# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2567 a_6781_3111# d2 a_6831_1914# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2568 a_4526_3195# a_4532_3378# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2569 vdd d0 a_20970_1520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2570 a_6904_5986# d1 a_7003_6396# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2571 a_18647_6152# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2572 gnd d4 a_15676_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2573 a_30937_5356# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2574 a_15522_3136# d2 a_15568_2116# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2575 a_20823_7818# a_20827_7641# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2576 a_12120_3759# a_12124_3582# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2577 a_13223_966# a_13230_1184# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2578 a_21462_184# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2579 a_27599_2513# a_27397_1497# a_27521_1616# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2580 a_32980_3987# d1 a_33079_4397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2581 a_1482_5651# a_1276_6140# a_697_5912# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2582 a_7797_6389# a_8054_6199# a_6999_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2583 vdd d0 a_21043_5592# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2584 vdd d0 a_16794_6636# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2585 a_18848_5134# a_18630_5134# a_18051_4906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2586 a_25094_2741# a_25351_2551# a_24301_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2587 a_33873_4390# a_34130_4200# a_33075_4574# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2588 a_6967_4360# d0 a_7760_4765# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2589 a_142_2164# a_148_2347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2590 a_15522_3136# a_15779_2946# a_15419_5174# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2591 a_2318_4959# d3 a_2490_7170# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2592 gnd d2 a_2757_3924# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2593 gnd d0 a_34166_6236# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2594 a_31963_2526# a_31761_1510# a_31885_1629# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2595 a_32970_7043# d2 a_33053_8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2596 a_116_829# a_3343_1286# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2597 a_22140_2277# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2598 a_30607_1379# d0 a_31082_1284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2599 a_25150_5795# a_25154_5618# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2600 a_13802_5950# a_13584_5950# a_13313_6056# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2601 a_22214_5937# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2602 a_33111_6610# a_33368_6420# a_33016_6023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2603 a_30667_5050# d0 a_31156_4944# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2604 a_245_8054# d0 a_734_7948# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2605 a_22196_5331# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2606 a_15687_3544# a_15944_3354# a_15605_4152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2607 a_22396_3901# a_22178_3901# a_21907_4007# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2608 a_235_7254# d0 a_716_7342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2609 a_18885_7170# d2 a_18936_6679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2610 a_19092_258# d5 a_19191_258# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2611 a_11241_4139# a_11498_3949# a_11162_2946# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2612 vdd d2 a_20091_1900# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2613 a_16468_2577# a_16485_3360# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2614 a_5008_2871# d1 a_5805_3099# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2615 gnd d2 a_11571_8021# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2616 a_11340_4549# d0 a_12138_4365# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2617 a_33115_6433# d0 a_33912_6661# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2618 a_4497_1860# a_4499_1959# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2619 a_14546_3124# d2 a_14597_2633# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2620 a_16557_7844# a_16561_7667# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2621 a_8913_4007# d0 a_9402_3901# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2622 a_15609_3975# d1 a_15704_4562# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2623 a_11413_8621# d0 a_12211_8437# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2624 a_4585_6432# a_4590_6756# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2625 a_20006_6572# d0 a_20808_6211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2626 gnd d0 a_12413_5605# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2627 a_660_4288# d1 a_1446_3615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2628 a_18693_3508# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2629 a_28616_3974# a_28869_3961# a_28533_2958# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2630 a_3416_5358# a_3420_5181# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2631 a_4616_8285# d0 a_5097_8373# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2632 gnd d0 a_21081_7216# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2633 a_25136_4188# a_25389_4175# a_24334_4549# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2634 a_23139_1075# a_22921_1075# a_22341_1259# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2635 a_9384_3295# a_9166_3295# a_8903_3207# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2636 a_6967_4360# d0 a_7764_4588# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2637 a_28612_4151# d1 a_28694_3543# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2638 a_33932_7679# a_33946_8462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2639 a_7744_3335# a_7748_3158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2640 a_28689_8046# a_28942_8033# a_28606_7030# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2641 a_6950_3342# d0 a_7747_3570# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2642 gnd d1 a_24647_7413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2643 vdd d0 a_34166_6236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2644 a_5097_8373# d1 a_5883_7700# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2645 a_13822_6968# d1 a_14619_7196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2646 a_9458_6955# a_9240_6955# a_8967_6768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2647 a_19092_258# d4 a_19689_4971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2648 a_25209_8260# a_25462_8247# a_24407_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2649 a_23212_5147# a_22994_5147# a_22414_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2650 a_24152_3123# d2 a_24202_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2651 a_4880_7961# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2652 a_4806_4301# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2653 vdd d1 a_11597_4359# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2654 a_15760_7616# d0 a_16558_7432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2655 a_29508_4789# a_29765_4599# a_28715_4384# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2656 a_2566_2311# d0 a_3359_2716# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2657 a_515_8360# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2658 a_33819_1336# a_33823_1159# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2659 a_20772_4175# a_20767_4764# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2660 a_5604_4117# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2661 a_28426_5173# d3 a_28533_2958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2662 a_33094_5592# d0 a_33896_5231# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2663 a_1492_2595# d3 a_1586_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2664 a_5660_7171# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2665 a_8945_5426# d0 a_9420_5331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2666 a_4534_3896# d0 a_5025_3889# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2667 vdd d2 a_11571_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2668 a_11340_4549# d0 a_12142_4188# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2669 a_5846_5664# d2 a_5924_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2670 gnd d2 a_20128_3936# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2671 a_31173_5962# a_30955_5962# a_30682_5969# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2672 a_31099_2302# a_30881_2302# a_30624_2397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2673 gnd d2 a_15862_3962# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2674 a_31922_3665# d2 a_31968_2645# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2675 a_23130_7593# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2676 a_3416_5358# a_3673_5168# a_2618_5542# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2677 a_15609_3975# d1 a_15708_4385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2678 a_1441_6548# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2679 a_11286_1495# a_11543_1305# a_11204_2103# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2680 a_2659_7401# a_2912_7388# a_2573_8186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2681 a_5810_3628# a_5604_4117# a_5024_4301# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2682 vdd d0 a_21081_7216# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2683 a_14418_8214# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2684 a_28612_4151# d1 a_28698_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2685 a_25132_4365# a_25389_4175# a_24334_4549# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2686 a_17502_1341# a_17504_1859# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2687 a_30918_4338# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2688 a_6785_2934# d2 a_6868_3950# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2689 a_10306_6692# d3 a_10400_6573# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2690 a_29492_3359# a_29496_3182# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2691 a_28685_8223# a_28942_8033# a_28606_7030# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2692 vdd d1 a_24647_7413# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2693 a_10145_1075# d2 a_10228_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2694 a_5732_2489# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2695 a_26773_3913# d1 a_27558_3652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2696 a_30974_7392# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2697 a_131_1329# d0 a_606_1234# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2698 a_11208_1926# d1 a_11303_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2699 a_18817_3627# a_18611_4116# a_18032_3888# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2700 a_32078_296# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2701 a_27604_2632# a_27434_3533# a_27558_3652# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2702 a_26846_7985# d1 a_27631_7724# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2703 a_18885_7170# a_18667_7170# a_18088_6942# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2704 a_24156_2946# d2 a_24235_4139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2705 gnd d0 a_34130_4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2706 a_15760_7616# d0 a_16562_7255# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2707 a_2566_2311# d0 a_3363_2539# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2708 a_33912_6661# a_34165_6648# a_33115_6433# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2709 a_20791_5193# a_21044_5180# a_19989_5554# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2710 a_2549_1293# d0 a_3346_1521# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2711 a_9944_2093# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2712 a_14624_7725# a_14418_8214# a_13838_8398# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2713 a_15740_6598# a_15997_6408# a_15645_6011# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2714 a_13296_5038# d0 a_13785_4932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2715 a_4512_2360# d0 a_4987_2265# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2716 a_24301_2336# a_24554_2323# a_24202_1926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2717 gnd d0 a_34203_8272# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2718 a_27626_7195# a_27408_7195# a_26828_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2719 a_17833_4906# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2720 a_14546_6586# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2721 a_28730_5579# a_28987_5389# a_28648_6187# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2722 a_24321_3354# d0 a_25118_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2723 a_4572_6031# d0 a_5061_5925# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2724 a_1186_1050# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2725 a_14390_1498# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2726 a_13253_2385# a_13258_2709# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2727 vdd d0 a_8036_5593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2728 a_22251_7973# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2729 a_22177_4313# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2730 a_17978_834# d1 a_18775_1062# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2731 vdd d0 a_34112_3594# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2732 a_16520_5808# a_16524_5631# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2733 a_13309_5439# a_13311_5957# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2734 a_27672_6585# a_27470_5569# a_27589_5159# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2735 a_19788_3110# d2 a_19834_2090# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2736 a_33823_1159# a_34076_1146# a_33021_1520# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2737 a_4091_172# d6 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2738 a_3360_2304# a_3364_2127# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2739 a_22250_8385# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2740 a_9365_1865# a_9147_1865# a_8876_1971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2741 vdd d2 a_2793_5960# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2742 a_29496_3182# a_29491_3771# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2743 a_17533_3194# a_17539_3377# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2744 a_3401_4163# a_3654_4150# a_2599_4524# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2745 a_5044_4907# a_4826_4907# a_4555_5013# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2746 gnd d0 a_12394_4587# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2747 gnd d0 a_25352_2139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2748 a_11208_1926# d1 a_11307_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2749 a_2577_8009# d1 a_2672_8596# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2750 a_30682_5969# a_30684_6068# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2751 a_21924_4926# a_21926_5025# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2752 gnd d1 a_7276_7401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2753 a_2417_3098# d2 a_2467_1901# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2754 a_30594_978# d0 a_31083_872# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2755 a_20787_5370# a_21044_5180# a_19989_5554# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2756 a_623_2252# a_405_2252# a_142_2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2757 gnd d4 a_11312_4971# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2758 a_23181_3640# a_22975_4129# a_22395_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2759 a_14764_6586# d4 a_14831_403# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2760 a_24297_2513# a_24554_2323# a_24202_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2761 vdd d0 a_34203_8272# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2762 a_22161_2883# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2763 a_697_5912# a_479_5912# a_206_5919# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2764 a_24353_5567# a_24610_5377# a_24271_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2765 a_18574_2080# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2766 a_11359_5567# d0 a_12161_5206# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2767 a_6999_6573# d0 a_7801_6212# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2768 a_116_829# d0 a_607_822# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2769 a_13363_8493# d0 a_13838_8398# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2770 a_13802_5950# a_13584_5950# a_13311_5957# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2771 a_11158_3123# a_11415_2933# a_11055_5161# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2772 a_11059_4984# d3 a_11231_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2773 a_7727_2552# a_7980_2539# a_6930_2324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2774 gnd d0 a_25371_3569# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2775 a_33075_4574# d0 a_33877_4213# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2776 gnd d0 a_29802_6223# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2777 a_8926_4408# d0 a_9401_4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2778 a_26353_7474# d0 a_26828_7379# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2779 a_28652_6010# d1 a_28751_6420# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2780 a_26792_4931# a_26574_4931# a_26301_4938# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2781 a_17519_2359# a_17524_2683# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2782 a_25209_8260# a_25204_8849# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2783 a_21920_4408# a_21924_4926# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2784 a_33819_1336# a_34076_1146# a_33021_1520# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2785 a_14514_1617# a_14308_2106# a_13729_1878# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2786 a_29509_4377# a_29513_4200# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2787 a_25151_5383# a_25408_5193# a_24353_5567# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2788 a_27315_2105# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2789 a_23222_2501# a_23020_1485# a_23144_1604# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2790 a_14582_5160# a_14364_5160# a_13785_4932# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2791 a_5883_7700# d2 a_5929_6680# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2792 a_24229_7018# a_24482_7005# a_24053_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2793 a_3397_4340# a_3654_4150# a_2599_4524# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2794 a_19191_258# d6 a_21680_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2795 a_26357_8091# a_26364_8309# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2796 a_29565_7431# a_29569_7254# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2797 a_191_5000# a_198_5218# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2798 a_32939_2128# a_33196_1938# a_32893_3148# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2799 gnd d2 a_33269_6010# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2800 a_24370_6585# d0 a_25168_6401# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2801 a_4879_8373# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2802 a_16541_6649# a_16794_6636# a_15744_6421# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2803 a_31679_2118# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2804 a_15423_4997# d3 a_15595_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2805 a_12121_3347# a_12125_3170# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2806 a_18936_6679# a_18766_7580# a_18890_7699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2807 gnd d1 a_11616_5377# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2808 gnd d0 a_29821_7653# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2809 a_12951_197# a_14707_284# a_14831_403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2810 a_4790_2871# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2811 a_168_3365# d0 a_643_3270# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2812 a_29531_5630# a_29784_5617# a_28734_5402# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2813 gnd d2 a_7121_3937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2814 a_31752_6190# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2815 a_17550_4212# d0 a_18031_4300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2816 a_21870_1971# a_21877_2189# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2817 a_443_3876# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2818 a_6864_4127# d1 a_6950_3342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2819 a_12211_8437# a_12468_8247# a_11413_8621# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2820 a_17606_7266# d0 a_18087_7354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2821 gnd d1 a_2875_5352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2822 a_20772_4175# a_21025_4162# a_19970_4536# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2823 a_13238_1885# a_13240_1984# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2824 gnd a_34202_8684# a_33152_8469# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2825 a_22415_4919# a_22197_4919# a_21926_5025# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2826 a_17797_2870# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2827 a_13277_4020# d0 a_13766_3914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2828 vdd d3 a_11488_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2829 a_442_4288# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2830 a_1285_1460# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2831 vdd d1 a_33295_2348# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2832 a_9458_6955# d1 a_10255_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2833 vdd d0 a_29802_6223# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2834 a_15645_6011# a_15898_5998# a_15595_7208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2835 vdd d0 a_8000_3557# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2836 vdd d4 a_19942_4958# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2837 a_11235_7018# d2 a_11314_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2838 a_17870_6942# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2839 a_25151_5383# a_25155_5206# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2840 a_17796_3282# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2841 a_5883_7700# a_5677_8189# a_5098_7961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2842 a_13277_4020# a_13284_4238# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2843 a_23321_2501# a_23103_2501# a_23222_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2844 a_21970_7279# d0 a_22451_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2845 a_13748_3308# d1 a_14546_3124# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2846 a_29459_1146# a_29454_1735# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2847 a_26364_8309# a_26370_8492# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2848 a_26845_8397# a_26627_8397# a_26364_8309# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2849 a_11344_4372# d0 a_12141_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2850 a_24235_4139# d1 a_24317_3531# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2851 vdd d2 a_33269_6010# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2852 a_7784_5194# a_8037_5181# a_6982_5555# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2853 a_14328_3124# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2854 a_24312_8034# a_24565_8021# a_24229_7018# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2855 a_24370_6585# d0 a_25172_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2856 a_33860_3195# a_34113_3182# a_33058_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2857 a_16537_6826# a_16794_6636# a_15744_6421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2858 a_10099_5557# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2859 a_5080_7355# a_4862_7355# a_4599_7267# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2860 a_16558_7432# a_16562_7255# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2861 a_4825_5319# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2862 a_26310_5255# a_26316_5438# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2863 a_14401_7196# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2864 a_5025_3889# a_4807_3889# a_4536_3995# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2865 vdd d0 a_29821_7653# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2866 vdd d0 a_29749_3169# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2867 a_30901_3320# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2868 a_10017_6165# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2869 a_25131_4777# a_25388_4587# a_24338_4372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2870 a_21877_2189# a_21883_2372# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2871 vdd d1 a_20210_3328# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2872 a_31968_2645# a_31798_3546# a_31917_3136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2873 a_18812_3098# a_18594_3098# a_18014_3282# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2874 a_10054_8201# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2875 vdd d1 a_2875_5352# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2876 a_17029_133# d8 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2877 a_20768_4352# a_21025_4162# a_19970_4536# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2878 a_8947_5944# d0 a_9438_5937# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2879 a_33945_8874# a_34202_8684# a_33152_8469# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2880 vdd d1 a_20283_7400# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2881 a_28751_6420# d0 a_29544_6825# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2882 gnd d0 a_21061_6198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2883 a_9202_5331# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2884 a_5856_2608# d3 a_5950_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2885 a_30644_3415# d0 a_31119_3320# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2886 a_19838_1913# d1 a_19933_2500# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2887 a_23057_3521# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2888 a_18104_8372# a_17886_8372# a_17629_8467# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2889 a_11235_7018# d2 a_11318_8034# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2890 a_1446_3615# d2 a_1492_2595# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2891 gnd d0 a_3636_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2892 a_13839_7986# a_13621_7986# a_13350_8092# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2893 gnd d1 a_24627_6395# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2894 a_13802_5950# d1 a_14587_5689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2895 a_10260_7712# a_10054_8201# a_9474_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2896 a_1519_7687# d2 a_1565_6667# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2897 a_33115_6433# d0 a_33908_6838# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2898 a_24235_4139# d1 a_24321_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2899 a_14665_6586# a_14463_5570# a_14587_5689# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2900 a_7780_5371# a_8037_5181# a_6982_5555# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2901 a_17502_1341# d0 a_17977_1246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2902 a_30594_978# a_30601_1196# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2903 a_26773_3913# a_26555_3913# a_26282_3920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2904 a_19989_5554# d0 a_20787_5370# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2905 a_26792_4931# d1 a_27589_5159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2906 a_24308_8211# a_24565_8021# a_24229_7018# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2907 a_4987_2265# a_4769_2265# a_4506_2177# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2908 a_17614_7967# a_17616_8066# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2909 a_10182_6573# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2910 a_33856_3372# a_34113_3182# a_33058_3556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2911 a_28602_7207# d2 a_28648_6187# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2912 a_9420_5331# a_9202_5331# a_8945_5426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2913 a_27352_4141# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2914 a_14551_3653# a_14345_4142# a_13766_3914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2915 a_17562_5012# d0 a_18051_4906# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2916 a_23227_2620# a_23057_3521# a_23181_3640# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2917 a_31137_3926# d1 a_31922_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2918 a_22469_7973# d1 a_23254_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2919 gnd d0 a_12450_7641# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2920 a_3436_6611# a_3689_6598# a_2639_6383# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2921 a_27553_3123# a_27335_3123# a_26756_2895# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2922 a_16505_4613# a_16758_4600# a_15708_4385# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2923 a_6950_3342# d0 a_7743_3747# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2924 a_1726_365# a_1544_4510# a_1659_6548# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2925 vdd d0 a_12358_2139# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2926 gnd d1 a_11597_4359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2927 gnd d0 a_34092_2576# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2928 a_29495_3594# a_29748_3581# a_28698_3366# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2929 a_16578_8685# a_16831_8672# a_15781_8457# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2930 a_6085_259# d4 a_6678_5149# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2931 a_19191_258# a_18973_258# a_19097_377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2932 a_23249_7183# a_23031_7183# a_22451_7367# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2933 a_10400_6573# a_10182_6573# a_10306_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2934 a_33021_1520# d0 a_33819_1336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2935 a_8894_2696# a_8896_2989# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2936 a_28751_6420# d0 a_29548_6648# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2937 a_5950_2489# a_5732_2489# a_5856_2608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2938 a_8982_7462# a_8984_7980# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2939 a_29568_7666# a_29821_7653# a_28771_7438# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2940 a_22124_847# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2941 a_19838_1913# d1 a_19937_2323# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2942 a_33094_5592# d0 a_33892_5408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2943 gnd d1 a_2856_4334# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2944 a_25114_3759# a_25118_3582# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2945 vdd d0 a_3636_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2946 a_21903_3390# a_21905_3908# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2947 a_17629_8467# a_16578_8685# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2948 a_27388_6177# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2949 a_22452_6955# a_22234_6955# a_21963_7061# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2950 a_23295_6573# d3 a_23394_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2951 a_10462_271# d5 a_10561_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2952 a_3474_8235# a_3469_8824# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2953 a_8896_2989# d0 a_9385_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2954 vdd d2 a_15825_1926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2955 a_19989_5554# d0 a_20791_5193# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2956 gnd d2 a_24455_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2957 a_26327_6273# a_26333_6456# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2958 a_3420_5181# a_3673_5168# a_2618_5542# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2959 a_4210_172# d6 a_4309_172# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2960 a_479_5912# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2961 a_14831_403# a_14649_4548# a_14691_2514# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2962 a_16489_3183# a_16742_3170# a_15687_3544# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2963 a_14764_6586# a_14546_6586# a_14670_6705# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2964 a_27656_4547# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2965 a_8903_3207# d0 a_9384_3295# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2966 a_32062_2526# d4 a_32202_415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2967 a_16521_5396# a_16525_5219# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2968 a_5805_3099# d2 a_5856_2608# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2969 a_4807_3889# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2970 vdd d0 a_12450_7641# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2971 a_31735_5172# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2972 a_7765_4176# a_8018_4163# a_6963_4537# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2973 gnd d0 a_21007_3556# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2974 a_27594_5688# a_27388_6177# a_26808_6361# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2975 a_6090_378# a_5908_4523# a_5950_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2976 a_1296_7158# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2977 a_26574_4931# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2978 a_18068_5924# a_17850_5924# a_17577_5931# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2979 a_16574_8862# a_16831_8672# a_15781_8457# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2980 a_7801_6212# a_7796_6801# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2981 vdd d0 a_34092_2576# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2982 a_29491_3771# a_29748_3581# a_28698_3366# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2983 a_18817_3627# d2 a_18863_2607# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2984 vdd d4 a_6935_4959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2985 a_33021_1520# d0 a_33823_1159# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2986 a_4862_7355# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2987 a_4536_3995# a_4543_4213# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X2988 a_2314_5136# d3 a_2421_2921# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2989 a_5587_3099# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2990 a_17524_2683# d0 a_18015_2870# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2991 a_22358_2277# a_22140_2277# a_21877_2189# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2992 a_12104_2564# a_12357_2551# a_11307_2336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2993 a_29564_7843# a_29821_7653# a_28771_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2994 a_11055_5161# d3 a_11158_3123# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2995 a_28788_8456# a_29041_8443# a_28689_8046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2996 a_5929_6680# a_5759_7581# a_5878_7171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X2997 a_7833_8837# a_8090_8647# a_7040_8432# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2998 vdd d1 a_2856_4334# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X2999 a_32893_3148# d2 a_32943_1951# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3000 a_13620_8398# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3001 a_17869_7354# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3002 a_8984_7980# d0 a_9475_7973# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3003 a_12177_6636# a_12430_6623# a_11380_6408# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3004 a_2467_1901# a_2720_1888# a_2417_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3005 a_24321_3354# d0 a_25114_3759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3006 a_30611_1996# a_30618_2214# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3007 a_28788_8456# d0 a_29581_8861# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3008 a_26610_7379# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3009 a_9183_4313# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3010 a_24156_2946# a_24409_2933# a_24049_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3011 a_33152_8469# a_33405_8456# a_33053_8059# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3012 a_31155_5356# a_30937_5356# a_30680_5451# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3013 a_733_8360# a_515_8360# a_258_8455# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3014 a_16485_3360# a_16742_3170# a_15687_3544# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3015 a_32897_2971# a_33150_2958# a_32790_5186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3016 a_2536_6150# a_2793_5960# a_2490_7170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3017 a_32966_7220# d2 a_33012_6200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3018 gnd d0 a_16778_5206# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3019 a_7761_4353# a_8018_4163# a_6963_4537# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3020 a_19970_4536# d0 a_20768_4352# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3021 a_11204_2103# d1 a_11286_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3022 vdd d0 a_21007_3556# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3023 a_2635_6560# d0 a_3433_6376# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3024 a_11281_5998# a_11534_5985# a_11231_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3025 a_29512_4612# a_29528_5395# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3026 a_9401_4313# a_9183_4313# a_8926_4408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3027 a_12088_1134# a_12341_1121# a_11286_1495# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3028 a_29471_2753# a_29475_2576# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3029 a_26353_7474# a_26355_7992# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3030 a_20791_5193# a_20786_5782# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3031 a_13494_860# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3032 a_21987_8297# a_21993_8480# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3033 a_9927_1075# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3034 a_24284_1318# a_24537_1305# a_24198_2103# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3035 a_5044_4907# d1 a_5841_5135# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3036 a_12100_2741# a_12357_2551# a_11307_2336# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3037 a_28784_8633# a_29041_8443# a_28689_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3038 a_27521_1616# d2 a_27599_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3039 a_33859_3607# a_33873_4390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3040 a_10000_5147# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3041 a_26719_859# a_26501_859# a_26230_965# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3042 a_4489_1159# a_4495_1342# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3043 a_25098_2564# a_25115_3347# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3044 a_206_5919# a_208_6018# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3045 a_6982_5555# d0 a_7780_5371# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3046 a_24357_5390# a_24610_5377# a_24271_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3047 vdd d0 a_25461_8659# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3048 a_33945_8874# gnd SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3049 a_12173_6813# a_12430_6623# a_11380_6408# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3050 a_21866_1354# a_21868_1872# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3051 a_18729_5544# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3052 a_32197_296# d5 a_30322_209# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3053 a_17148_133# a_25910_208# a_26029_208# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3054 a_33058_3556# d0 a_33856_3372# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3055 a_28788_8456# d0 a_29585_8684# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3056 a_33891_5820# a_33895_5643# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3057 a_1560_6548# a_1358_5532# a_1477_5122# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3058 a_33148_8646# a_33405_8456# a_33053_8059# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3059 a_4752_1247# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3060 a_9437_6349# a_9219_6349# a_8956_6261# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3061 gnd d0 a_21060_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3062 a_1659_6548# a_1441_6548# a_1565_6667# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3063 a_32966_7220# d2 a_33016_6023# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3064 a_13273_3403# a_13275_3921# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3065 a_19970_4536# d0 a_20772_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3066 a_2635_6560# d0 a_3437_6199# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3067 a_1404_1050# a_1186_1050# a_606_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3068 a_135_1946# d0 a_624_1840# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3069 a_12084_1311# a_12341_1121# a_11286_1495# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3070 a_18775_1062# d2 a_18858_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3071 a_3457_7217# a_3710_7204# a_2655_7578# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3072 a_7724_2317# a_7981_2127# a_6926_2501# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3073 a_19865_7005# d2 a_19948_8021# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3074 a_4970_1247# a_4752_1247# a_4495_1342# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3075 a_28694_3543# d0 a_29496_3182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3076 a_31716_4154# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3077 a_32041_6717# a_31871_7618# a_31995_7737# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3078 a_13566_5344# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3079 a_16505_4613# a_16521_5396# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3080 vdd d0 a_25445_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3081 a_17776_2264# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3082 a_16464_2754# a_16468_2577# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3083 a_19871_4126# d1 a_19957_3341# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3084 a_26555_3913# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3085 a_19944_8198# a_20201_8008# a_19865_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3086 a_9220_5937# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3087 a_5908_4523# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3088 a_30638_3232# a_30644_3415# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3089 a_30646_3933# d0 a_31137_3926# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3090 a_26301_4938# a_26303_5037# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3091 a_179_4200# a_185_4383# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3092 a_26518_1877# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3093 a_13729_1878# a_13511_1878# a_13238_1885# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3094 gnd d0 a_34148_5630# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3095 a_6982_5555# d0 a_7784_5194# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3096 a_17977_1246# a_17759_1246# a_17496_1158# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3097 a_27604_2632# d3 a_27698_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3098 a_18812_6560# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3099 a_19907_6162# a_20164_5972# a_19861_7182# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3100 a_6864_4127# d1 a_6946_3519# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3101 a_12215_8260# a_12468_8247# a_11413_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3102 a_10218_5147# a_10000_5147# a_9420_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3103 a_679_5306# a_461_5306# a_204_5401# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3104 a_33058_3556# d0 a_33860_3195# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3105 a_25205_8437# a_25209_8260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3106 gnd d0 a_29785_5205# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3107 a_13728_2290# a_13510_2290# a_13253_2385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3108 gnd d0 a_16795_6224# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3109 a_1322_3496# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3110 a_4572_6031# a_4579_6249# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3111 a_12951_197# d6 a_8658_196# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3112 a_31922_3665# a_31716_4154# a_31136_4338# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3113 a_13784_5344# a_13566_5344# a_13309_5439# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3114 a_14509_1088# a_14291_1088# a_13712_860# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3115 a_21680_184# a_21462_184# a_21581_184# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3116 gnd d1 a_33295_2348# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3117 gnd d0 a_8000_3557# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3118 a_14381_6178# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3119 a_33895_5643# a_33909_6426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3120 a_22396_3901# a_22178_3901# a_21905_3908# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3121 a_8982_7462# d0 a_9457_7367# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3122 vdd d0 a_21060_6610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3123 a_27371_5159# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3124 a_22921_1075# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3125 a_18780_1591# a_18574_2080# a_17994_2264# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3126 a_28426_5173# a_28683_4983# a_27833_283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3127 a_9239_7367# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3128 a_6858_7006# a_7111_6993# a_6682_4972# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3129 a_20808_6211# a_20803_6800# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3130 a_23176_3111# a_22958_3111# a_22379_2883# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3131 a_11400_7426# d0 a_12193_7831# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3132 a_10136_7593# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3133 a_26297_4420# a_26301_4938# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3134 gnd d0 a_16759_4188# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3135 a_31917_6598# d3 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3136 a_21851_854# a_25078_1311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3137 a_5686_3509# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3138 a_20717_1533# a_20731_2316# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3139 a_11303_2513# d0 a_12105_2152# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3140 gnd d0 a_29749_3169# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3141 a_2549_1293# a_2802_1280# a_2463_2078# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3142 a_30697_6469# d0 a_31172_6374# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3143 vdd d0 a_20971_1108# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3144 a_33822_1571# a_33836_2354# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3145 a_12178_6224# a_12173_6813# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3146 vdd d0 a_34148_5630# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3147 a_30609_1897# a_30611_1996# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3148 a_25191_7654# a_25444_7641# a_24394_7426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3149 a_26809_5949# a_26591_5949# a_26320_6055# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3150 a_13260_3002# d0 a_13749_2896# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3151 gnd d1 a_20210_3328# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3152 a_425_3270# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3153 a_33908_6838# a_33912_6661# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3154 gnd d1 a_15944_3354# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3155 a_30697_6469# a_30702_6793# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3156 vdd d0 a_16795_6224# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3157 a_32794_5009# a_33047_4996# a_32197_296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3158 a_9981_4129# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3159 a_17543_3994# a_17550_4212# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3160 a_25095_2329# a_25352_2139# a_24297_2513# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3161 a_12087_1546# a_12101_2329# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3162 a_5856_2608# a_5686_3509# a_5810_3628# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3163 a_30881_2302# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3164 a_13267_3220# d0 a_13748_3308# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3165 a_31963_2526# d3 a_32062_2526# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3166 a_4519_2977# d0 a_5008_2871# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3167 a_12173_6813# a_12177_6636# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3168 a_17489_940# a_17496_1158# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3169 a_15595_7208# d2 a_15645_6011# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3170 a_7036_8609# a_7293_8419# a_6941_8022# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3171 a_23279_4535# d4 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3172 a_4526_3195# d0 a_5007_3283# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3173 a_11327_3354# d0 a_12124_3582# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3174 a_3342_1698# a_3599_1508# a_2549_1293# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3175 a_18015_2870# a_17797_2870# a_17526_2976# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3176 a_19685_5148# d3 a_19788_3110# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3177 a_26828_7379# d1 a_27626_7195# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3178 a_28689_8046# d1 a_28784_8633# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3179 a_9474_8385# a_9256_8385# a_8993_8297# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3180 a_23217_5676# a_23011_6165# a_22431_6349# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3181 a_11400_7426# d0 a_12197_7654# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3182 a_7040_8432# d0 a_7837_8660# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3183 a_29581_8861# a_29585_8684# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3184 a_14670_6705# a_14500_7606# a_14624_7725# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3185 a_10026_1485# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3186 a_3347_1109# a_3342_1698# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3187 a_26318_5956# a_26320_6055# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3188 a_2545_1470# a_2802_1280# a_2463_2078# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3189 a_4210_172# a_5966_259# a_6085_259# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3190 a_25187_7831# a_25444_7641# a_24394_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3191 gnd d0 a_12358_2139# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3192 a_17887_7960# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3193 a_4599_7267# a_4605_7450# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3194 a_9129_1259# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3195 vdd d1 a_15944_3354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3196 gnd d0 a_12414_5193# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3197 a_32790_5186# d3 a_32893_3148# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3198 a_660_4288# a_442_4288# a_179_4200# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3199 a_4607_7968# d0 a_5098_7961# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3200 a_8883_2189# d0 a_9364_2277# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3201 a_13296_5038# a_13303_5256# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3202 a_19834_2090# d1 a_19916_1482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3203 gnd d0 a_34129_4612# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3204 a_22233_7367# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3205 a_10187_3640# a_9981_4129# a_9401_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3206 a_2676_8419# a_2929_8406# a_2577_8009# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3207 a_30674_5268# a_30680_5451# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3208 gnd d2 a_28869_3961# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3209 a_11359_5567# a_11616_5377# a_11277_6175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3210 a_2421_2921# a_2674_2908# a_2314_5136# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3211 a_18105_7960# d1 a_18890_7699# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3212 a_26756_2895# a_26538_2895# a_26265_2708# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3213 a_680_4894# d1 a_1477_5122# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3214 a_13765_4326# a_13547_4326# a_13290_4421# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3215 a_9347_1259# a_9129_1259# a_8872_1354# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3216 a_11376_6585# a_11633_6395# a_11281_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3217 a_16501_4790# a_16505_4613# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3218 a_2490_7170# d2 a_2536_6150# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3219 a_2562_2488# d0 a_3360_2304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3220 a_29509_4377# a_29766_4187# a_28711_4561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3221 gnd d2 a_28942_8033# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3222 a_30322_209# a_32078_296# a_32197_296# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3223 a_28689_8046# d1 a_28788_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3224 a_26755_3307# a_26537_3307# a_26280_3402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3225 a_15723_5580# d0 a_16521_5396# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3226 a_4970_1247# d1 a_5768_1063# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3227 a_17978_834# a_17760_834# a_17489_940# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3228 a_10228_2501# a_10026_1485# a_10145_1075# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3229 a_13253_2385# d0 a_13728_2290# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3230 a_19689_4971# d3 a_19865_7005# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3231 a_9437_6349# d1 a_10223_5676# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3232 a_221_6419# d0 a_696_6324# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3233 a_6900_6163# a_7157_5973# a_6854_7183# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3234 a_5044_4907# a_4826_4907# a_4553_4914# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3235 a_26243_1366# d0 a_26718_1271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3236 a_32976_4164# a_33233_3974# a_32897_2971# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3237 a_18656_1472# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3238 gnd d2 a_33306_8046# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3239 a_11235_7018# a_11488_7005# a_11059_4984# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3240 vdd d0 a_16777_5618# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3241 a_23144_1604# d2 a_23222_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3242 gnd d0 a_25334_1533# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3243 a_22958_3111# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3244 a_2639_6383# d0 a_3436_6611# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3245 a_10327_2501# d4 a_10467_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3246 a_5623_5135# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3247 a_15423_4997# a_15676_4984# a_14826_284# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3248 a_10561_271# a_10343_271# a_10467_390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3249 a_18973_258# d5 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3250 a_29472_2341# a_29476_2164# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3251 vdd d0 a_34129_4612# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3252 a_24411_8444# d0 a_25208_8672# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3253 a_21978_7980# a_21980_8079# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3254 a_27397_1497# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3255 a_1276_6140# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3256 a_20786_5782# a_21043_5592# a_19993_5377# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3257 a_7837_8660# a_8090_8647# a_7040_8432# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3258 a_30592_879# a_30594_978# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3259 a_18858_2488# a_18656_1472# a_18780_1591# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3260 a_168_3365# a_170_3883# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3261 gnd d1 a_2912_7388# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3262 a_1602_246# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3263 a_21853_953# d0 a_22342_847# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3264 a_31136_4338# a_30918_4338# a_30655_4250# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3265 a_2504_3937# a_2757_3924# a_2421_2921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3266 a_17506_1958# d0 a_17995_1852# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3267 a_2562_2488# d0 a_3364_2127# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3268 a_33946_8462# a_33950_8285# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3269 vdd d2 a_28942_8033# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3270 a_33913_6249# a_34166_6236# a_33111_6610# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3271 a_31192_7392# a_30974_7392# a_30711_7304# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3272 a_30937_5356# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3273 a_12084_1311# a_12088_1134# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3274 a_2500_4114# d1 a_2582_3506# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3275 a_18848_5134# a_18630_5134# a_18050_5318# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3276 a_33892_5408# a_33896_5231# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3277 a_13584_5950# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3278 a_10327_2501# a_10109_2501# a_10228_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3279 a_6941_8022# a_7194_8009# a_6858_7006# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3280 a_24317_3531# d0 a_25119_3170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3281 a_4616_8285# a_4622_8468# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3282 a_3420_5181# a_3415_5770# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3283 a_21870_1971# d0 a_22359_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3284 vdd d2 a_33306_8046# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3285 a_20030_7413# a_20283_7400# a_19944_8198# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3286 a_5773_1592# a_5567_2081# a_4988_1853# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3287 vdd d0 a_25334_1533# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3288 a_22178_3901# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3289 a_12210_8849# a_12214_8672# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3290 a_13313_6056# a_13320_6274# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3291 a_22140_2277# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3292 a_23227_2620# d3 a_23321_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3293 a_9130_847# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3294 a_11314_8211# d1 a_11396_7603# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3295 a_7765_4176# a_7760_4765# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3296 a_27480_2513# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3297 a_22341_1259# a_22123_1259# a_21860_1171# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3298 a_12160_5618# a_12413_5605# a_11363_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3299 a_28715_4384# d0 a_29508_4789# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3300 a_6682_4972# d3 a_6854_7183# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3301 gnd d0 a_12395_4175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3302 a_9166_3295# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3303 gnd d0 a_25461_8659# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3304 a_22415_4919# a_22197_4919# a_21924_4926# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3305 a_10037_7183# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3306 a_25154_5618# a_25168_6401# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3307 vdd d1 a_33351_5402# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3308 a_4605_7450# d0 a_5080_7355# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3309 a_24394_7426# a_24647_7413# a_24308_8211# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3310 a_33909_6426# a_34166_6236# a_33111_6610# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3311 a_31083_872# d1 a_31880_1100# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3312 a_27631_7724# d2 a_27677_6704# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3313 a_18014_3282# d1 a_18812_3098# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3314 a_27833_283# d4 a_28426_5173# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3315 vdd d0 a_29784_5617# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3316 a_2500_4114# d1 a_2586_3329# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3317 a_2573_8186# a_2830_7996# a_2494_6993# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3318 a_661_3876# d1 a_1446_3615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3319 a_33896_5231# a_33891_5820# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3320 a_30631_3014# a_30638_3232# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3321 a_15605_4152# a_15862_3962# a_15526_2959# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3322 a_1441_3086# a_1223_3086# a_644_2858# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3323 a_15704_4562# d0 a_16502_4378# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3324 a_32197_296# d4 a_32790_5186# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3325 a_7728_2140# a_7981_2127# a_6926_2501# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3326 a_26291_4237# a_26297_4420# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3327 a_5008_2871# a_4790_2871# a_4517_2684# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3328 a_8903_3207# a_8909_3390# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3329 a_1409_1579# d2 a_1487_2476# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3330 a_28694_3543# d0 a_29492_3359# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3331 a_19875_3949# a_20128_3936# a_19792_2933# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3332 a_11314_8211# d1 a_11400_7426# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3333 vdd d2 a_15898_5998# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3334 gnd d0 a_25445_7229# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3335 vdd d0 a_16758_4600# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3336 a_16485_3360# a_16489_3183# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3337 a_20755_3157# a_20750_3746# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3338 a_19871_4126# d1 a_19953_3518# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3339 a_5007_3283# a_4789_3283# a_4532_3378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3340 gnd d3 a_20045_2920# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3341 a_7834_8425# a_7838_8248# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3342 a_14582_5160# d2 a_14665_6586# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3343 a_5604_4117# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3344 a_26297_4420# d0 a_26772_4325# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3345 a_17887_7960# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3346 vdd d0 a_12395_4175# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3347 a_1487_2476# d3 a_1586_2476# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3348 a_153_2671# a_155_2964# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3349 a_10306_6692# a_10136_7593# a_10260_7712# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3350 a_5660_7171# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3351 a_15645_6011# d1 a_15740_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3352 a_8949_6043# d0 a_9438_5937# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3353 a_716_7342# a_498_7342# a_235_7254# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3354 a_17606_7266# a_17612_7449# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3355 a_8939_5243# d0 a_9420_5331# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3356 gnd d3 a_28786_2945# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3357 vdd d0 a_8090_8647# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3358 a_24390_7603# a_24647_7413# a_24308_8211# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3359 a_23144_1604# a_22938_2093# a_22359_1865# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3360 a_16542_6237# a_16795_6224# a_15740_6598# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3361 a_13821_7380# a_13603_7380# a_13340_7292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3362 a_5841_5135# d2 a_5924_6561# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3363 a_28648_6187# d1 a_28730_5579# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3364 a_33909_6426# a_33913_6249# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3365 a_18667_7170# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3366 a_31917_3136# d2 a_31968_2645# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3367 a_23249_7183# d2 a_23300_6692# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3368 a_5097_8373# a_4879_8373# a_4616_8285# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3369 a_24312_8034# d1 a_24407_8621# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3370 a_32202_415# a_32020_4560# a_32062_2526# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3371 a_14418_8214# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3372 a_17597_6755# d0 a_18088_6942# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3373 a_30992_7998# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3374 a_10301_6573# d3 a_10400_6573# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3375 a_8889_2372# a_8894_2696# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3376 a_30918_4338# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3377 a_33950_8285# a_34203_8272# a_33148_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3378 a_13340_7292# a_13346_7475# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3379 gnd d1 a_20173_1292# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3380 gnd d2 a_24492_3949# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3381 a_27408_7195# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3382 a_125_1146# d0 a_606_1234# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3383 a_18817_3627# a_18611_4116# a_18031_4300# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3384 a_30991_8410# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3385 a_33876_4625# a_33892_5408# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3386 a_17489_940# d0 a_17978_834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3387 gnd d2 a_11461_1913# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3388 a_7779_5783# a_8036_5593# a_6986_5378# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3389 a_17504_1859# a_17506_1958# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3390 a_8969_7061# a_8976_7279# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3391 a_25077_1723# a_25081_1546# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3392 a_11204_2103# a_11461_1913# a_11158_3123# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3393 vdd d1 a_20300_8418# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3394 a_24357_5390# d0 a_25150_5795# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3395 a_18739_2488# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3396 a_33855_3784# a_34112_3594# a_33062_3379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3397 a_18890_7699# a_18684_8188# a_18104_8372# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3398 a_17592_6431# a_17597_6755# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3399 a_11303_2513# d0 a_12101_2329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3400 a_16489_3183# a_16484_3772# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3401 a_29582_8449# a_29586_8272# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3402 a_14670_6705# d3 a_14764_6586# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3403 a_8658_196# a_12832_197# a_10561_271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3404 a_7728_2140# a_7723_2729# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3405 a_20824_7406# a_20828_7229# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3406 a_4506_2177# d0 a_4987_2265# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3407 a_28533_2958# d2 a_28616_3974# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3408 a_21581_184# a_23337_271# a_23456_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3409 a_30702_6793# d0 a_31193_6980# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3410 a_28579_1938# a_28832_1925# a_28529_3135# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3411 a_30734_8505# d0 a_31209_8410# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3412 a_5929_6680# d3 a_6023_6561# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3413 a_16538_6414# a_16795_6224# a_15740_6598# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3414 a_13712_860# d1 a_14509_1088# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3415 gnd d0 a_3726_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3416 a_4826_4907# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3417 a_25099_2152# a_25352_2139# a_24297_2513# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3418 a_4590_6756# a_4592_7049# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3419 a_6854_7183# d2 a_6904_5986# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3420 a_1544_4510# d4 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3421 a_4770_1853# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3422 a_22379_2883# a_22161_2883# a_21888_2696# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3423 a_30902_2908# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3424 a_29528_5395# a_29785_5205# a_28730_5579# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3425 a_7023_7414# a_7276_7401# a_6937_8199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3426 a_12194_7419# a_12198_7242# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3427 a_24312_8034# d1 a_24411_8444# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3428 a_22452_6955# a_22234_6955# a_21961_6768# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3429 a_17592_6431# d0 a_18067_6336# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3430 a_27672_6585# a_27470_5569# a_27594_5688# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3431 a_22378_3295# a_22160_3295# a_21903_3390# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3432 a_405_2252# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3433 a_7040_8432# a_7293_8419# a_6941_8022# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3434 vdd d1 a_33388_7438# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3435 a_19030_6560# a_18812_6560# a_18936_6679# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3436 a_11059_4984# a_11312_4971# a_10462_271# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3437 a_27838_402# d5 a_27932_283# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3438 a_11327_3354# d0 a_12120_3759# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3439 a_33946_8462# a_34203_8272# a_33148_8646# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3440 a_5550_1063# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3441 a_13510_2290# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3442 a_479_5912# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3443 a_28747_6597# d0 a_29545_6413# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3444 a_32897_2971# d2 a_32976_4164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3445 a_116_829# a_118_928# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3446 a_19993_5377# d0 a_20790_5605# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3447 a_7040_8432# d0 a_7833_8837# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3448 a_13584_5950# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3449 a_26500_1271# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3450 a_18858_2488# d3 a_18957_2488# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3451 gnd d0 a_3637_3132# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3452 a_8976_7279# a_8982_7462# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3453 a_30203_209# d6 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3454 a_21939_5426# d0 a_22414_5331# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3455 a_22342_847# a_22124_847# a_21851_854# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3456 a_30592_879# d0 a_31083_872# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3457 a_623_2252# a_405_2252# a_148_2347# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3458 a_29585_8684# a_29838_8671# a_28788_8456# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3459 a_29586_8272# a_29581_8861# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3460 a_26574_4931# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3461 a_17623_8284# a_17629_8467# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3462 a_33111_6610# d0 a_33909_6426# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3463 a_14691_2514# d4 a_14831_403# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3464 a_17995_1852# a_17777_1852# a_17504_1859# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3465 a_14308_2106# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3466 a_14364_5160# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3467 a_22469_7973# a_22251_7973# a_21980_8079# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3468 a_33933_7267# a_33928_7856# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3469 vdd d1 a_24537_1305# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3470 a_30864_1284# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3471 vdd d0 a_3726_8634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3472 a_6858_7006# d2 a_6937_8199# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3473 a_2655_7578# a_2912_7388# a_2573_8186# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3474 a_33016_6023# a_33269_6010# a_32966_7220# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3475 a_18775_1062# a_18557_1062# a_17978_834# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3476 a_7796_6801# a_7800_6624# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3477 a_6946_3519# d0 a_7744_3335# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3478 a_8986_8079# d0 a_9475_7973# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3479 a_26347_7291# d0 a_26828_7379# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3480 a_27771_6585# a_27553_6585# a_27672_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3481 a_8920_4225# d0 a_9401_4313# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3482 a_12198_7242# a_12193_7831# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3483 a_1726_365# d5 a_1820_246# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3484 a_18766_7580# d2 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3485 a_11363_5390# a_11616_5377# a_11277_6175# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3486 a_7764_4588# a_7780_5371# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3487 a_14514_1617# a_14308_2106# a_13728_2290# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3488 gnd d0 a_34093_2164# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3489 a_16579_8273# a_16832_8260# a_15777_8634# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3490 a_8993_8297# d0 a_9474_8385# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3491 a_28747_6597# d0 a_29549_6236# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3492 a_389_822# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3493 a_27516_1087# a_27298_1087# a_26718_1271# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3494 a_29569_7254# a_29822_7241# a_28767_7615# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3495 gnd d0 a_21097_8646# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3496 gnd d3 a_7038_2921# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3497 a_22197_4919# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3498 a_16506_4201# a_16501_4790# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3499 vdd d0 a_3637_3132# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3500 a_4879_8373# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3501 a_226_6743# d0 a_717_6930# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3502 a_29581_8861# a_29838_8671# a_28788_8456# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3503 a_16452_1147# a_16447_1736# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3504 a_33111_6610# d0 a_33913_6249# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3505 a_2622_5365# d0 a_3415_5770# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3506 gnd d0 a_16777_5618# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3507 a_21853_953# a_21860_1171# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3508 a_9964_3111# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3509 a_5677_8189# d1 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3510 a_13331_6781# d0 a_13822_6968# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3511 a_23103_2501# d3 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3512 a_443_3876# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3513 a_5966_259# d5 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3514 a_13530_3308# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3515 a_20718_1121# a_20971_1108# a_19916_1482# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3516 a_8894_2696# d0 a_9385_2883# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3517 a_26627_8397# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3518 a_2467_1901# d1 a_2562_2488# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3519 a_644_2858# a_426_2858# a_153_2671# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3520 a_12211_8437# a_12215_8260# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3521 gnd d2 a_20201_8008# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3522 a_20807_6623# a_20824_7406# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3523 a_33012_6200# a_33269_6010# a_32966_7220# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3524 a_27434_3533# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3525 a_24411_8444# d0 a_25204_8849# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3526 vdd d0 a_12451_7229# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3527 a_8539_196# d7 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3528 gnd d0 a_21008_3144# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3529 a_20767_4764# a_20771_4587# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3530 gnd d1 a_7166_1293# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3531 a_6946_3519# d0 a_7748_3158# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3532 gnd d0 a_34185_7666# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3533 a_18088_6942# d1 a_18885_7170# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3534 a_33012_6200# d1 a_33098_5415# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3535 a_23456_271# d4 a_24049_5161# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3536 a_23321_2501# a_23103_2501# a_23227_2620# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3537 a_4807_3889# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3538 a_16575_8450# a_16832_8260# a_15777_8634# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3539 vdd d0 a_12394_4587# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3540 vdd d0 a_34093_2164# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3541 a_29492_3359# a_29749_3169# a_28694_3543# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3542 a_4863_6943# d0 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3543 a_32036_6598# a_31834_5582# a_31958_5701# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3544 a_13749_2896# d1 a_14546_3124# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3545 a_15526_2959# d2 a_15605_4152# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3546 a_31798_3546# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3547 a_18594_3098# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3548 a_29565_7431# a_29822_7241# a_28767_7615# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3549 a_13712_860# a_13494_860# a_13223_966# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3550 vdd d0 a_21097_8646# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3551 a_11281_5998# d1 a_11376_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3552 a_5080_7355# a_4862_7355# a_4605_7450# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3553 a_31871_7618# d2 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3554 a_12178_6224# a_12431_6211# a_11376_6585# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3555 gnd d1 a_15980_5390# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3556 a_24317_3531# d0 a_25115_3347# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3557 a_25187_7831# a_25191_7654# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3558 a_8939_5243# a_8945_5426# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3559 gnd d0 a_29728_2563# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3560 a_26357_8091# d0 a_26846_7985# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3561 vdd d3 a_24409_2933# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3562 a_10017_6165# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3563 a_2622_5365# d0 a_3419_5593# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3564 a_8857_854# a_12084_1311# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3565 a_3383_3557# a_3636_3544# a_2586_3329# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3566 a_29549_6236# a_29544_6825# SUB sky130_fd_pr__res_generic_nd w=0.17 l=0.81
X3567 a_24374_6408# a_24627_6395# a_24275_5998# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3568 a_31156_4944# a_30938_4944# a_30667_5050# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3569 a_15708_4385# d0 a_16505_4613# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3570 a_5773_1592# d2 a_5851_2489# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3571 a_9147_1865# d0 gnd SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3572 a_31968_2645# a_31798_3546# a_31922_3665# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3573 a_734_7948# a_516_7948# a_245_8054# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3574 a_26364_8309# d0 a_26845_8397# vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
X3575 a_18087_7354# a_17869_7354# a_17606_7266# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3576 a_21920_4408# d0 a_22395_4313# SUB sky130_fd_pr__nfet_01v8 w=0.42 l=0.5
X3577 a_10054_8201# d1 vdd vdd sky130_fd_pr__pfet_01v8 w=1.0 l=0.5
C0 a_19092_258# a_19097_377# 5.60fF
C1 d1 vdd 4.27fF
C2 a_1721_246# a_1726_365# 5.60fF
C3 a_10462_271# a_10467_390# 5.60fF
C4 d2 vdd 3.73fF
C5 a_23456_271# a_23461_390# 5.60fF
C6 a_32197_296# a_32202_415# 5.60fF
C7 d0 gnd 19.14fF
C8 a_14826_284# a_14831_403# 5.60fF
C9 a_6085_259# a_6090_378# 5.60fF
C10 d1 gnd 10.12fF
C11 vdd gnd 9.71fF
C12 d3 gnd 2.53fF
C13 d2 gnd 5.06fF
C14 d0 vdd 7.22fF
C15 a_27833_283# a_27838_402# 5.60fF
C16 gnd SUB 109.45fF
C17 a_30322_209# SUB 3.15fF
C18 vdd SUB 481.72fF
C19 a_27932_283# SUB 3.77fF
C20 a_26029_208# SUB 5.68fF
C21 a_21581_184# SUB 3.15fF
C22 a_21680_184# SUB 5.69fF
C23 a_19191_258# SUB 3.77fF
C24 d5 SUB 3.90fF
C25 a_12951_197# SUB 3.15fF
C26 a_10561_271# SUB 3.77fF
C27 a_8658_196# SUB 5.73fF
C28 a_8757_196# SUB 9.23fF
C29 a_4210_172# SUB 3.15fF
C30 a_4309_172# SUB 5.69fF
C31 a_1820_246# SUB 3.77fF
C32 a_30592_879# SUB 5.34fF
C33 d0 SUB 157.68fF
C34 a_26228_866# SUB 5.34fF
C35 a_21851_854# SUB 5.34fF
C36 a_17487_841# SUB 5.34fF
C37 a_13221_867# SUB 5.34fF
C38 a_31083_872# SUB 2.21fF
C39 d1 SUB 81.44fF
C40 a_26719_859# SUB 2.21fF
C41 a_31082_1284# SUB 2.30fF
C42 a_22342_847# SUB 2.21fF
C43 a_8857_854# SUB 5.34fF
C44 a_4480_842# SUB 5.34fF
C45 a_116_829# SUB 5.34fF
C46 a_33021_1520# SUB 2.30fF
C47 a_26718_1271# SUB 2.30fF
C48 a_17978_834# SUB 2.21fF
C49 a_28657_1507# SUB 2.30fF
C50 a_22341_1259# SUB 2.30fF
C51 a_13712_860# SUB 2.21fF
C52 a_24280_1495# SUB 2.30fF
C53 a_17977_1246# SUB 2.30fF
C54 d2 SUB 37.77fF
C55 a_33025_1343# SUB 2.21fF
C56 a_19916_1482# SUB 2.30fF
C57 a_13711_1272# SUB 2.30fF
C58 a_4971_835# SUB 2.21fF
C59 a_28661_1330# SUB 2.21fF
C60 a_15650_1508# SUB 2.30fF
C61 a_9347_1259# SUB 2.30fF
C62 a_607_822# SUB 2.21fF
C63 a_24284_1318# SUB 2.21fF
C64 a_11286_1495# SUB 2.30fF
C65 a_4970_1247# SUB 2.30fF
C66 a_19920_1305# SUB 2.21fF
C67 a_6909_1483# SUB 2.30fF
C68 a_606_1234# SUB 2.30fF
C69 a_15654_1331# SUB 2.21fF
C70 a_2545_1470# SUB 2.30fF
C71 a_11290_1318# SUB 2.21fF
C72 a_6913_1306# SUB 2.21fF
C73 a_2549_1293# SUB 2.21fF
C74 a_31100_1890# SUB 2.21fF
C75 a_26736_1877# SUB 2.21fF
C76 a_31099_2302# SUB 2.30fF
C77 a_22359_1865# SUB 2.21fF
C78 a_26735_2289# SUB 2.30fF
C79 a_17995_1852# SUB 2.21fF
C80 a_33038_2538# SUB 2.30fF
C81 a_22358_2277# SUB 2.30fF
C82 a_13729_1878# SUB 2.21fF
C83 a_28674_2525# SUB 2.30fF
C84 a_31963_2526# SUB 2.37fF
C85 a_17994_2264# SUB 2.30fF
C86 a_9365_1865# SUB 2.21fF
C87 a_24297_2513# SUB 2.30fF
C88 d3 SUB 22.79fF
C89 a_33042_2361# SUB 2.21fF
C90 a_27599_2513# SUB 2.37fF
C91 a_13728_2290# SUB 2.30fF
C92 a_4988_1853# SUB 2.21fF
C93 a_19933_2500# SUB 2.30fF
C94 a_28678_2348# SUB 2.21fF
C95 a_23222_2501# SUB 2.37fF
C96 a_624_1840# SUB 2.21fF
C97 a_15667_2526# SUB 2.30fF
C98 a_24301_2336# SUB 2.21fF
C99 a_18858_2488# SUB 2.37fF
C100 a_4987_2265# SUB 2.30fF
C101 a_11303_2513# SUB 2.30fF
C102 a_19937_2323# SUB 2.21fF
C103 a_14592_2514# SUB 2.37fF
C104 a_623_2252# SUB 2.30fF
C105 a_6926_2501# SUB 2.30fF
C106 a_15671_2349# SUB 2.21fF
C107 a_10228_2501# SUB 2.37fF
C108 a_2562_2488# SUB 2.30fF
C109 a_11307_2336# SUB 2.21fF
C110 a_5851_2489# SUB 2.37fF
C111 a_6930_2324# SUB 2.21fF
C112 a_1487_2476# SUB 2.37fF
C113 a_2566_2311# SUB 2.21fF
C114 a_31120_2908# SUB 2.21fF
C115 a_26756_2895# SUB 2.21fF
C116 a_31119_3320# SUB 2.30fF
C117 a_22379_2883# SUB 2.21fF
C118 a_33058_3556# SUB 2.30fF
C119 a_18015_2870# SUB 2.21fF
C120 a_28694_3543# SUB 2.30fF
C121 a_22378_3295# SUB 2.30fF
C122 a_13749_2896# SUB 2.21fF
C123 a_24317_3531# SUB 2.30fF
C124 a_18014_3282# SUB 2.30fF
C125 a_9385_2883# SUB 2.21fF
C126 a_33062_3379# SUB 2.21fF
C127 a_19953_3518# SUB 2.30fF
C128 a_13748_3308# SUB 2.30fF
C129 a_5008_2871# SUB 2.21fF
C130 a_28698_3366# SUB 2.21fF
C131 a_15687_3544# SUB 2.30fF
C132 a_9384_3295# SUB 2.30fF
C133 a_644_2858# SUB 2.21fF
C134 a_24321_3354# SUB 2.21fF
C135 a_11323_3531# SUB 2.30fF
C136 a_5007_3283# SUB 2.30fF
C137 a_19957_3341# SUB 2.21fF
C138 a_6946_3519# SUB 2.30fF
C139 a_643_3270# SUB 2.30fF
C140 a_15691_3367# SUB 2.21fF
C141 a_2582_3506# SUB 2.30fF
C142 a_11327_3354# SUB 2.21fF
C143 a_6950_3342# SUB 2.21fF
C144 a_2586_3329# SUB 2.21fF
C145 a_32897_2971# SUB 2.63fF
C146 a_28533_2958# SUB 2.63fF
C147 a_31137_3926# SUB 2.21fF
C148 a_24156_2946# SUB 2.63fF
C149 a_19792_2933# SUB 2.63fF
C150 a_31136_4338# SUB 2.30fF
C151 a_22396_3901# SUB 2.21fF
C152 a_15526_2959# SUB 2.63fF
C153 a_18032_3888# SUB 2.21fF
C154 a_11162_2946# SUB 2.63fF
C155 a_33075_4574# SUB 2.30fF
C156 a_22395_4313# SUB 2.30fF
C157 a_13766_3914# SUB 2.21fF
C158 a_6785_2934# SUB 2.63fF
C159 a_28711_4561# SUB 2.30fF
C160 a_32062_2526# SUB 4.04fF
C161 a_32202_415# SUB 5.00fF
C162 a_18031_4300# SUB 2.30fF
C163 a_9402_3901# SUB 2.21fF
C164 a_2421_2921# SUB 2.63fF
C165 a_24334_4549# SUB 2.30fF
C166 d4 SUB 11.46fF
C167 a_33079_4397# SUB 2.21fF
C168 a_27698_2513# SUB 4.04fF
C169 a_27838_402# SUB 5.00fF
C170 a_19970_4536# SUB 2.30fF
C171 a_28715_4384# SUB 2.21fF
C172 a_23321_2501# SUB 4.04fF
C173 a_23461_390# SUB 5.00fF
C174 a_13765_4326# SUB 2.30fF
C175 a_5025_3889# SUB 2.21fF
C176 a_9401_4313# SUB 2.30fF
C177 a_661_3876# SUB 2.21fF
C178 a_15704_4562# SUB 2.30fF
C179 a_24338_4372# SUB 2.21fF
C180 a_18957_2488# SUB 4.04fF
C181 a_19097_377# SUB 5.00fF
C182 a_5024_4301# SUB 2.30fF
C183 a_11340_4549# SUB 2.30fF
C184 a_19974_4359# SUB 2.21fF
C185 a_14691_2514# SUB 4.04fF
C186 a_14831_403# SUB 5.00fF
C187 a_660_4288# SUB 2.30fF
C188 a_6963_4537# SUB 2.30fF
C189 a_15708_4385# SUB 2.21fF
C190 a_10327_2501# SUB 4.04fF
C191 a_10467_390# SUB 5.00fF
C192 a_2599_4524# SUB 2.30fF
C193 a_11344_4372# SUB 2.21fF
C194 a_5950_2489# SUB 4.04fF
C195 a_6090_378# SUB 5.00fF
C196 a_6967_4360# SUB 2.21fF
C197 a_1586_2476# SUB 4.04fF
C198 a_1726_365# SUB 5.00fF
C199 a_2603_4347# SUB 2.21fF
C200 a_32197_296# SUB 5.75fF
C201 a_32790_5186# SUB 2.94fF
C202 a_27833_283# SUB 5.75fF
C203 a_28426_5173# SUB 2.94fF
C204 a_31156_4944# SUB 2.21fF
C205 a_23456_271# SUB 5.75fF
C206 a_24049_5161# SUB 2.94fF
C207 a_19092_258# SUB 5.75fF
C208 a_19685_5148# SUB 2.94fF
C209 a_31155_5356# SUB 2.30fF
C210 a_22415_4919# SUB 2.21fF
C211 a_14826_284# SUB 5.75fF
C212 a_15419_5174# SUB 2.94fF
C213 a_33094_5592# SUB 2.30fF
C214 a_18051_4906# SUB 2.21fF
C215 a_10462_271# SUB 5.75fF
C216 a_11055_5161# SUB 2.94fF
C217 a_28730_5579# SUB 2.30fF
C218 a_22414_5331# SUB 2.30fF
C219 a_13785_4932# SUB 2.21fF
C220 a_6085_259# SUB 5.75fF
C221 a_6678_5149# SUB 2.94fF
C222 a_24353_5567# SUB 2.30fF
C223 a_18050_5318# SUB 2.30fF
C224 a_9421_4919# SUB 2.21fF
C225 a_1721_246# SUB 5.75fF
C226 a_2314_5136# SUB 2.94fF
C227 a_33098_5415# SUB 2.21fF
C228 a_19989_5554# SUB 2.30fF
C229 a_13784_5344# SUB 2.30fF
C230 a_5044_4907# SUB 2.21fF
C231 a_28734_5402# SUB 2.21fF
C232 a_15723_5580# SUB 2.30fF
C233 a_9420_5331# SUB 2.30fF
C234 a_680_4894# SUB 2.21fF
C235 a_24357_5390# SUB 2.21fF
C236 a_11359_5567# SUB 2.30fF
C237 a_5043_5319# SUB 2.30fF
C238 a_19993_5377# SUB 2.21fF
C239 a_6982_5555# SUB 2.30fF
C240 a_679_5306# SUB 2.30fF
C241 a_15727_5403# SUB 2.21fF
C242 a_2618_5542# SUB 2.30fF
C243 a_11363_5390# SUB 2.21fF
C244 a_6986_5378# SUB 2.21fF
C245 a_2622_5365# SUB 2.21fF
C246 a_31173_5962# SUB 2.21fF
C247 a_31172_6374# SUB 2.30fF
C248 a_22432_5937# SUB 2.21fF
C249 a_18068_5924# SUB 2.21fF
C250 a_33111_6610# SUB 2.30fF
C251 a_22431_6349# SUB 2.30fF
C252 a_13802_5950# SUB 2.21fF
C253 a_28747_6597# SUB 2.30fF
C254 a_32036_6598# SUB 2.63fF
C255 a_32135_6598# SUB 2.94fF
C256 a_18067_6336# SUB 2.30fF
C257 a_9438_5937# SUB 2.21fF
C258 a_24370_6585# SUB 2.30fF
C259 a_33115_6433# SUB 2.21fF
C260 a_27672_6585# SUB 2.63fF
C261 a_27771_6585# SUB 2.94fF
C262 a_13801_6362# SUB 2.30fF
C263 a_20006_6572# SUB 2.30fF
C264 a_28751_6420# SUB 2.21fF
C265 a_23295_6573# SUB 2.63fF
C266 a_23394_6573# SUB 2.94fF
C267 a_9437_6349# SUB 2.30fF
C268 a_697_5912# SUB 2.21fF
C269 a_15740_6598# SUB 2.30fF
C270 a_24374_6408# SUB 2.21fF
C271 a_18931_6560# SUB 2.63fF
C272 a_19030_6560# SUB 2.94fF
C273 a_5060_6337# SUB 2.30fF
C274 a_11376_6585# SUB 2.30fF
C275 a_20010_6395# SUB 2.21fF
C276 a_14665_6586# SUB 2.63fF
C277 a_14764_6586# SUB 2.94fF
C278 a_696_6324# SUB 2.30fF
C279 a_6999_6573# SUB 2.30fF
C280 a_15744_6421# SUB 2.21fF
C281 a_10301_6573# SUB 2.63fF
C282 a_10400_6573# SUB 2.94fF
C283 a_2635_6560# SUB 2.30fF
C284 a_11380_6408# SUB 2.21fF
C285 a_5924_6561# SUB 2.63fF
C286 a_6023_6561# SUB 2.94fF
C287 a_7003_6396# SUB 2.21fF
C288 a_1560_6548# SUB 2.63fF
C289 a_1659_6548# SUB 2.94fF
C290 a_2639_6383# SUB 2.21fF
C291 a_32794_5009# SUB 4.03fF
C292 a_28430_4996# SUB 4.03fF
C293 a_31193_6980# SUB 2.21fF
C294 a_24053_4984# SUB 4.03fF
C295 a_26829_6967# SUB 2.21fF
C296 a_19689_4971# SUB 4.03fF
C297 a_31192_7392# SUB 2.30fF
C298 a_22452_6955# SUB 2.21fF
C299 a_15423_4997# SUB 4.03fF
C300 a_33131_7628# SUB 2.30fF
C301 a_18088_6942# SUB 2.21fF
C302 a_11059_4984# SUB 4.03fF
C303 a_28767_7615# SUB 2.30fF
C304 a_22451_7367# SUB 2.30fF
C305 a_13822_6968# SUB 2.21fF
C306 a_6682_4972# SUB 4.03fF
C307 a_24390_7603# SUB 2.30fF
C308 a_18087_7354# SUB 2.30fF
C309 a_9458_6955# SUB 2.21fF
C310 a_2318_4959# SUB 4.03fF
C311 a_33135_7451# SUB 2.21fF
C312 a_20026_7590# SUB 2.30fF
C313 a_13821_7380# SUB 2.30fF
C314 a_5081_6943# SUB 2.21fF
C315 a_28771_7438# SUB 2.21fF
C316 a_15760_7616# SUB 2.30fF
C317 a_9457_7367# SUB 2.30fF
C318 a_717_6930# SUB 2.21fF
C319 a_24394_7426# SUB 2.21fF
C320 a_11396_7603# SUB 2.30fF
C321 a_20030_7413# SUB 2.21fF
C322 a_7019_7591# SUB 2.30fF
C323 a_716_7342# SUB 2.30fF
C324 a_15764_7439# SUB 2.21fF
C325 a_2655_7578# SUB 2.30fF
C326 a_11400_7426# SUB 2.21fF
C327 a_7023_7414# SUB 2.21fF
C328 a_2659_7401# SUB 2.21fF
C329 a_32970_7043# SUB 2.37fF
C330 a_28606_7030# SUB 2.37fF
C331 a_31210_7998# SUB 2.21fF
C332 a_24229_7018# SUB 2.37fF
C333 a_19865_7005# SUB 2.37fF
C334 a_31209_8410# SUB 2.30fF
C335 a_22469_7973# SUB 2.21fF
C336 a_15599_7031# SUB 2.37fF
C337 a_26845_8397# SUB 2.30fF
C338 a_18105_7960# SUB 2.21fF
C339 a_11235_7018# SUB 2.37fF
C340 a_22468_8385# SUB 2.30fF
C341 a_13839_7986# SUB 2.21fF
C342 a_6858_7006# SUB 2.37fF
C343 a_18104_8372# SUB 2.30fF
C344 a_9475_7973# SUB 2.21fF
C345 a_2494_6993# SUB 2.37fF
C346 a_33148_8646# SUB 2.30fF
C347 a_28784_8633# SUB 2.30fF
C348 a_24407_8621# SUB 2.30fF
C349 a_33152_8469# SUB 2.21fF
C350 a_20043_8608# SUB 2.30fF
C351 a_13838_8398# SUB 2.30fF
C352 a_9474_8385# SUB 2.30fF
C353 a_734_7948# SUB 2.21fF
C354 a_5097_8373# SUB 2.30fF
C355 a_733_8360# SUB 2.30fF
C356 a_28788_8456# SUB 2.21fF
C357 a_15777_8634# SUB 2.30fF
C358 a_25208_8672# SUB 2.54fF
C359 a_24411_8444# SUB 2.21fF
C360 a_11413_8621# SUB 2.30fF
C361 a_20844_8659# SUB 2.31fF
C362 a_20047_8431# SUB 2.21fF
C363 a_7036_8609# SUB 2.30fF
C364 a_16578_8685# SUB 2.37fF
C365 a_15781_8457# SUB 2.21fF
C366 a_2672_8596# SUB 2.30fF
C367 a_12214_8672# SUB 2.31fF
C368 a_11417_8444# SUB 2.21fF
C369 a_7837_8660# SUB 2.54fF
C370 a_7040_8432# SUB 2.21fF
C371 a_3473_8647# SUB 2.31fF
C372 a_2676_8419# SUB 2.21fF

Vdd vdd 0 dc 1.8
Vsub SUB 0 dc 0
Vin1 vref 0 dc 3.3
Vd0 d0 0 pulse(0 1.8 0ns 0.1ns 0.1ns 5ns 10ns)
Vd1 d1 0 pulse(0 1.8 0ns 0.1ns 0.1ns 10ns 20ns)
Vd2 d2 0 pulse(0 1.8 0ns 0.1ns 0.1ns 20ns 40ns)
Vd3 d3 0 pulse(0 1.8 0ns 0.1ns 0.1ns 40ns 80ns)
Vd4 d4 0 pulse(0 1.8 0ns 0.1ns 0.1ns 80ns 160ns)
Vd5 d5 0 pulse(0 1.8 0ns 0.1ns 0.1ns 160ns 320ns)
Vd6 d6 0 pulse(0 1.8 0ns 0.1ns 0.1ns 320ns 640ns)
Vd7 d7 0 pulse(0 1.8 0ns 0.1ns 0.1ns 640ns 1280ns)
Vd8 d8 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1280ns 2560ns)


.tran 5ns 2560ns
.control
run
plot V(vout) 
.endc
.end

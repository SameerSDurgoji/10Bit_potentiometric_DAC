magic
tech sky130A
timestamp 1616086883
<< nwell >>
rect 1047 -185 1655 -35
<< nmos >>
rect 1111 -286 1161 -244
rect 1329 -286 1379 -244
rect 1537 -286 1587 -244
<< pmos >>
rect 1111 -167 1161 -67
rect 1329 -167 1379 -67
rect 1537 -167 1587 -67
<< ndiff >>
rect 1062 -254 1111 -244
rect 1062 -274 1073 -254
rect 1093 -274 1111 -254
rect 1062 -286 1111 -274
rect 1161 -250 1205 -244
rect 1161 -270 1176 -250
rect 1196 -270 1205 -250
rect 1161 -286 1205 -270
rect 1280 -254 1329 -244
rect 1280 -274 1291 -254
rect 1311 -274 1329 -254
rect 1280 -286 1329 -274
rect 1379 -250 1423 -244
rect 1379 -270 1394 -250
rect 1414 -270 1423 -250
rect 1379 -286 1423 -270
rect 1493 -250 1537 -244
rect 1493 -270 1502 -250
rect 1522 -270 1537 -250
rect 1493 -286 1537 -270
rect 1587 -254 1636 -244
rect 1587 -274 1605 -254
rect 1625 -274 1636 -254
rect 1587 -286 1636 -274
<< pdiff >>
rect 1067 -105 1111 -67
rect 1067 -125 1079 -105
rect 1099 -125 1111 -105
rect 1067 -167 1111 -125
rect 1161 -105 1203 -67
rect 1161 -125 1175 -105
rect 1195 -125 1203 -105
rect 1161 -167 1203 -125
rect 1285 -105 1329 -67
rect 1285 -125 1297 -105
rect 1317 -125 1329 -105
rect 1285 -167 1329 -125
rect 1379 -105 1421 -67
rect 1379 -125 1393 -105
rect 1413 -125 1421 -105
rect 1379 -167 1421 -125
rect 1495 -105 1537 -67
rect 1495 -125 1503 -105
rect 1523 -125 1537 -105
rect 1495 -167 1537 -125
rect 1587 -98 1632 -67
rect 1587 -105 1631 -98
rect 1587 -125 1599 -105
rect 1619 -125 1631 -105
rect 1587 -167 1631 -125
<< ndiffc >>
rect 1073 -274 1093 -254
rect 1176 -270 1196 -250
rect 1291 -274 1311 -254
rect 1394 -270 1414 -250
rect 1502 -270 1522 -250
rect 1605 -274 1625 -254
<< pdiffc >>
rect 1079 -125 1099 -105
rect 1175 -125 1195 -105
rect 1297 -125 1317 -105
rect 1393 -125 1413 -105
rect 1503 -125 1523 -105
rect 1599 -125 1619 -105
<< poly >>
rect 1111 -67 1161 -54
rect 1329 -67 1379 -54
rect 1537 -67 1587 -54
rect 1111 -195 1161 -167
rect 1111 -215 1124 -195
rect 1144 -215 1161 -195
rect 1111 -244 1161 -215
rect 1329 -192 1379 -167
rect 1329 -212 1342 -192
rect 1362 -212 1379 -192
rect 1329 -244 1379 -212
rect 1537 -194 1587 -167
rect 1537 -214 1560 -194
rect 1580 -214 1587 -194
rect 1537 -244 1587 -214
rect 1111 -302 1161 -286
rect 1329 -302 1379 -286
rect 1537 -302 1587 -286
<< polycont >>
rect 1124 -215 1144 -195
rect 1342 -212 1362 -192
rect 1560 -214 1580 -194
<< locali >>
rect 1419 -9 1484 -8
rect 1070 -34 1257 -10
rect 1288 -29 1681 -9
rect 1701 -29 1704 -9
rect 1288 -34 1704 -29
rect 1070 -105 1107 -34
rect 1288 -35 1629 -34
rect 1222 -95 1253 -94
rect 1070 -125 1079 -105
rect 1099 -125 1107 -105
rect 1070 -135 1107 -125
rect 1166 -105 1253 -95
rect 1166 -125 1175 -105
rect 1195 -125 1253 -105
rect 1166 -134 1253 -125
rect 1166 -135 1203 -134
rect 1222 -185 1253 -134
rect 1288 -105 1325 -35
rect 1591 -36 1628 -35
rect 1440 -95 1476 -94
rect 1288 -125 1297 -105
rect 1317 -125 1325 -105
rect 1288 -135 1325 -125
rect 1384 -105 1532 -95
rect 1632 -98 1728 -96
rect 1384 -125 1393 -105
rect 1413 -125 1503 -105
rect 1523 -125 1532 -105
rect 1384 -134 1532 -125
rect 1590 -105 1728 -98
rect 1590 -125 1599 -105
rect 1619 -125 1728 -105
rect 1590 -134 1728 -125
rect 1384 -135 1421 -134
rect 1114 -188 1155 -187
rect 1006 -195 1155 -188
rect 1006 -215 1065 -195
rect 1085 -215 1124 -195
rect 1144 -215 1155 -195
rect 1006 -223 1155 -215
rect 1222 -192 1379 -185
rect 1222 -212 1342 -192
rect 1362 -212 1379 -192
rect 1222 -222 1379 -212
rect 1222 -223 1257 -222
rect 1222 -244 1253 -223
rect 1440 -244 1476 -134
rect 1495 -135 1532 -134
rect 1591 -135 1628 -134
rect 1551 -194 1641 -188
rect 1551 -214 1560 -194
rect 1580 -196 1641 -194
rect 1580 -214 1605 -196
rect 1551 -216 1605 -214
rect 1625 -216 1641 -196
rect 1551 -222 1641 -216
rect 1065 -245 1102 -244
rect 1064 -254 1102 -245
rect 1064 -274 1073 -254
rect 1093 -274 1102 -254
rect 1064 -282 1102 -274
rect 1168 -250 1253 -244
rect 1283 -245 1320 -244
rect 1168 -270 1176 -250
rect 1196 -270 1253 -250
rect 1168 -278 1253 -270
rect 1282 -254 1320 -245
rect 1282 -274 1291 -254
rect 1311 -274 1320 -254
rect 1168 -279 1204 -278
rect 1282 -282 1320 -274
rect 1386 -250 1530 -244
rect 1386 -270 1394 -250
rect 1414 -270 1502 -250
rect 1522 -270 1530 -250
rect 1386 -278 1530 -270
rect 1386 -279 1422 -278
rect 1494 -279 1530 -278
rect 1596 -245 1633 -244
rect 1596 -246 1634 -245
rect 1596 -254 1660 -246
rect 1596 -274 1605 -254
rect 1625 -268 1660 -254
rect 1680 -268 1683 -248
rect 1625 -273 1683 -268
rect 1625 -274 1660 -273
rect 1065 -311 1102 -282
rect 1066 -313 1102 -311
rect 1066 -335 1257 -313
rect 1283 -314 1320 -282
rect 1596 -286 1660 -274
rect 1700 -312 1727 -134
rect 1559 -314 1727 -312
rect 1283 -340 1727 -314
rect 1393 -564 1433 -340
rect 1559 -341 1727 -340
rect 1393 -586 1401 -564
rect 1425 -586 1433 -564
rect 1393 -594 1433 -586
<< viali >>
rect 1681 -29 1701 -9
rect 1065 -215 1085 -195
rect 1605 -216 1625 -196
rect 1660 -268 1680 -248
rect 1401 -586 1425 -564
<< metal1 >>
rect 1674 -9 1709 -6
rect 1674 -29 1681 -9
rect 1701 -29 1709 -9
rect 1674 -37 1709 -29
rect 1056 -195 1641 -187
rect 1056 -215 1065 -195
rect 1085 -196 1641 -195
rect 1085 -215 1605 -196
rect 1056 -216 1605 -215
rect 1625 -216 1641 -196
rect 1056 -222 1641 -216
rect 1675 -243 1709 -37
rect 1653 -248 1709 -243
rect 1653 -268 1660 -248
rect 1680 -268 1709 -248
rect 1653 -275 1709 -268
rect 1653 -276 1688 -275
rect 1396 -564 1435 -551
rect 1396 -569 1401 -564
rect 988 -586 1401 -569
rect 1425 -569 1435 -564
rect 1425 -586 1436 -569
rect 988 -594 1436 -586
<< labels >>
rlabel locali 1073 -25 1102 -19 1 vdd
rlabel locali 1070 -324 1099 -318 1 gnd
rlabel space 1176 -306 1205 -297 1 gnd
rlabel nwell 1208 -48 1231 -45 1 vdd
rlabel locali 1446 -178 1468 -163 1 vout
rlabel locali 1013 -217 1035 -200 1 d1
<< end >>
